module fake_ariane_516_n_17181 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_17181);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_17181;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_9872;
wire n_14741;
wire n_16050;
wire n_9604;
wire n_10943;
wire n_10453;
wire n_12407;
wire n_15048;
wire n_7329;
wire n_4030;
wire n_12343;
wire n_13909;
wire n_7029;
wire n_6790;
wire n_4770;
wire n_14469;
wire n_11913;
wire n_8165;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_12760;
wire n_11172;
wire n_12018;
wire n_14470;
wire n_3056;
wire n_3500;
wire n_15304;
wire n_6603;
wire n_2679;
wire n_6557;
wire n_17159;
wire n_10678;
wire n_5402;
wire n_11190;
wire n_13957;
wire n_6581;
wire n_15154;
wire n_16227;
wire n_2182;
wire n_5553;
wire n_6002;
wire n_7277;
wire n_2680;
wire n_11458;
wire n_16683;
wire n_11999;
wire n_3264;
wire n_16580;
wire n_1250;
wire n_5717;
wire n_10649;
wire n_13176;
wire n_10794;
wire n_12945;
wire n_2993;
wire n_17013;
wire n_17081;
wire n_4283;
wire n_9297;
wire n_11627;
wire n_2879;
wire n_4403;
wire n_10557;
wire n_13125;
wire n_8139;
wire n_15369;
wire n_11453;
wire n_416;
wire n_4962;
wire n_1430;
wire n_14456;
wire n_7832;
wire n_16166;
wire n_8438;
wire n_2002;
wire n_12806;
wire n_12244;
wire n_11135;
wire n_1238;
wire n_11306;
wire n_15390;
wire n_15157;
wire n_2729;
wire n_4302;
wire n_14658;
wire n_12589;
wire n_5791;
wire n_7127;
wire n_13109;
wire n_4547;
wire n_14209;
wire n_13718;
wire n_5090;
wire n_3765;
wire n_8321;
wire n_864;
wire n_5302;
wire n_15105;
wire n_1096;
wire n_1379;
wire n_10000;
wire n_2376;
wire n_12103;
wire n_7922;
wire n_7805;
wire n_9807;
wire n_2790;
wire n_7542;
wire n_12354;
wire n_2207;
wire n_11783;
wire n_7053;
wire n_16181;
wire n_11614;
wire n_9892;
wire n_5712;
wire n_14807;
wire n_11143;
wire n_3954;
wire n_6297;
wire n_4982;
wire n_2042;
wire n_10704;
wire n_14334;
wire n_16576;
wire n_11431;
wire n_11799;
wire n_462;
wire n_16966;
wire n_8699;
wire n_9263;
wire n_9734;
wire n_1131;
wire n_8037;
wire n_5479;
wire n_2646;
wire n_8257;
wire n_737;
wire n_2653;
wire n_4610;
wire n_16300;
wire n_6058;
wire n_11246;
wire n_11377;
wire n_10213;
wire n_232;
wire n_13029;
wire n_3115;
wire n_9886;
wire n_15093;
wire n_4028;
wire n_5263;
wire n_10904;
wire n_15293;
wire n_5565;
wire n_9096;
wire n_6358;
wire n_8546;
wire n_6293;
wire n_8997;
wire n_13215;
wire n_14066;
wire n_2482;
wire n_9985;
wire n_15841;
wire n_9665;
wire n_16698;
wire n_1682;
wire n_14300;
wire n_12233;
wire n_11349;
wire n_7001;
wire n_10169;
wire n_10903;
wire n_13875;
wire n_16759;
wire n_11906;
wire n_958;
wire n_6129;
wire n_13755;
wire n_14335;
wire n_2554;
wire n_14473;
wire n_13910;
wire n_15347;
wire n_4321;
wire n_15801;
wire n_10574;
wire n_13066;
wire n_1985;
wire n_5590;
wire n_10468;
wire n_2621;
wire n_14226;
wire n_9241;
wire n_146;
wire n_6524;
wire n_16188;
wire n_16032;
wire n_9286;
wire n_16284;
wire n_4853;
wire n_9592;
wire n_338;
wire n_8744;
wire n_1909;
wire n_5229;
wire n_15921;
wire n_12574;
wire n_6313;
wire n_12260;
wire n_7464;
wire n_8449;
wire n_15404;
wire n_9683;
wire n_10380;
wire n_10968;
wire n_14979;
wire n_4260;
wire n_13491;
wire n_903;
wire n_7626;
wire n_9939;
wire n_3348;
wire n_239;
wire n_15874;
wire n_12315;
wire n_10688;
wire n_3261;
wire n_9358;
wire n_1761;
wire n_16157;
wire n_9466;
wire n_8953;
wire n_11756;
wire n_7965;
wire n_16817;
wire n_13636;
wire n_7368;
wire n_9787;
wire n_1690;
wire n_8399;
wire n_16825;
wire n_2807;
wire n_6664;
wire n_8598;
wire n_10276;
wire n_15671;
wire n_7562;
wire n_11604;
wire n_9997;
wire n_7534;
wire n_13196;
wire n_1018;
wire n_12581;
wire n_7428;
wire n_4512;
wire n_17012;
wire n_6190;
wire n_8460;
wire n_12085;
wire n_14960;
wire n_4132;
wire n_16108;
wire n_13980;
wire n_14861;
wire n_16646;
wire n_1364;
wire n_8068;
wire n_2390;
wire n_7373;
wire n_6891;
wire n_4500;
wire n_9318;
wire n_10281;
wire n_16224;
wire n_13715;
wire n_12089;
wire n_625;
wire n_2322;
wire n_8734;
wire n_12671;
wire n_16798;
wire n_1107;
wire n_14592;
wire n_15750;
wire n_8720;
wire n_331;
wire n_559;
wire n_2663;
wire n_10528;
wire n_8097;
wire n_5481;
wire n_6539;
wire n_13120;
wire n_12993;
wire n_495;
wire n_8422;
wire n_4824;
wire n_8114;
wire n_12728;
wire n_7467;
wire n_16641;
wire n_14572;
wire n_350;
wire n_16657;
wire n_8126;
wire n_381;
wire n_5340;
wire n_3545;
wire n_6797;
wire n_16841;
wire n_7392;
wire n_9714;
wire n_14598;
wire n_14405;
wire n_16147;
wire n_15441;
wire n_10399;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_8664;
wire n_10131;
wire n_14378;
wire n_11721;
wire n_7526;
wire n_561;
wire n_11736;
wire n_4143;
wire n_14430;
wire n_10634;
wire n_4273;
wire n_507;
wire n_11444;
wire n_901;
wire n_11891;
wire n_13058;
wire n_4136;
wire n_14094;
wire n_9809;
wire n_11492;
wire n_3144;
wire n_14636;
wire n_2359;
wire n_9613;
wire n_9354;
wire n_17139;
wire n_1519;
wire n_5896;
wire n_7338;
wire n_4567;
wire n_12647;
wire n_9897;
wire n_786;
wire n_9295;
wire n_5833;
wire n_6249;
wire n_15363;
wire n_6887;
wire n_15602;
wire n_10595;
wire n_11767;
wire n_13180;
wire n_6253;
wire n_15577;
wire n_9119;
wire n_6128;
wire n_3552;
wire n_2950;
wire n_9058;
wire n_17000;
wire n_8326;
wire n_7200;
wire n_6197;
wire n_11807;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_11944;
wire n_2301;
wire n_13090;
wire n_3121;
wire n_15161;
wire n_2847;
wire n_5589;
wire n_11474;
wire n_11819;
wire n_15423;
wire n_16768;
wire n_8504;
wire n_3015;
wire n_5744;
wire n_8920;
wire n_3870;
wire n_12080;
wire n_6808;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_277;
wire n_5691;
wire n_7937;
wire n_16257;
wire n_8985;
wire n_3482;
wire n_7490;
wire n_13069;
wire n_6295;
wire n_11409;
wire n_5403;
wire n_823;
wire n_11692;
wire n_1900;
wire n_620;
wire n_13138;
wire n_12599;
wire n_6096;
wire n_4268;
wire n_6338;
wire n_587;
wire n_863;
wire n_6992;
wire n_303;
wire n_3960;
wire n_10644;
wire n_12863;
wire n_16369;
wire n_2433;
wire n_352;
wire n_899;
wire n_3975;
wire n_8035;
wire n_11856;
wire n_16652;
wire n_5830;
wire n_9516;
wire n_15063;
wire n_365;
wire n_2004;
wire n_13996;
wire n_13064;
wire n_4018;
wire n_1495;
wire n_8660;
wire n_334;
wire n_192;
wire n_15593;
wire n_3325;
wire n_6681;
wire n_661;
wire n_4227;
wire n_15788;
wire n_5158;
wire n_9917;
wire n_12185;
wire n_5152;
wire n_8939;
wire n_11737;
wire n_533;
wire n_11652;
wire n_16701;
wire n_15326;
wire n_11038;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_13991;
wire n_1924;
wire n_6542;
wire n_13466;
wire n_9202;
wire n_13689;
wire n_13896;
wire n_11925;
wire n_1811;
wire n_16277;
wire n_14115;
wire n_6161;
wire n_16705;
wire n_15930;
wire n_3612;
wire n_273;
wire n_4505;
wire n_11974;
wire n_12457;
wire n_6452;
wire n_10426;
wire n_1840;
wire n_5247;
wire n_9923;
wire n_9512;
wire n_8469;
wire n_8715;
wire n_5464;
wire n_7306;
wire n_10070;
wire n_4476;
wire n_6740;
wire n_16368;
wire n_6978;
wire n_12792;
wire n_579;
wire n_7507;
wire n_13458;
wire n_844;
wire n_1267;
wire n_8176;
wire n_9677;
wire n_2956;
wire n_5210;
wire n_7379;
wire n_149;
wire n_1213;
wire n_2382;
wire n_7441;
wire n_7215;
wire n_237;
wire n_15481;
wire n_780;
wire n_5292;
wire n_1918;
wire n_8327;
wire n_12556;
wire n_8991;
wire n_7438;
wire n_11200;
wire n_8855;
wire n_4119;
wire n_4443;
wire n_9811;
wire n_4000;
wire n_13762;
wire n_9508;
wire n_13441;
wire n_13532;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_6136;
wire n_1140;
wire n_14236;
wire n_3458;
wire n_570;
wire n_11597;
wire n_5843;
wire n_7874;
wire n_11309;
wire n_14156;
wire n_15702;
wire n_8539;
wire n_13118;
wire n_8630;
wire n_9308;
wire n_14587;
wire n_15566;
wire n_8533;
wire n_13830;
wire n_11233;
wire n_7108;
wire n_3511;
wire n_2077;
wire n_9638;
wire n_1121;
wire n_11047;
wire n_15665;
wire n_11068;
wire n_490;
wire n_17144;
wire n_3012;
wire n_13912;
wire n_15057;
wire n_15429;
wire n_1947;
wire n_13768;
wire n_4529;
wire n_3850;
wire n_575;
wire n_11476;
wire n_8435;
wire n_7695;
wire n_10245;
wire n_6156;
wire n_11611;
wire n_13111;
wire n_1216;
wire n_4908;
wire n_8098;
wire n_3754;
wire n_8204;
wire n_11957;
wire n_5060;
wire n_13290;
wire n_12509;
wire n_12663;
wire n_9199;
wire n_12155;
wire n_15221;
wire n_13379;
wire n_15828;
wire n_11210;
wire n_4432;
wire n_7162;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_9808;
wire n_7331;
wire n_10457;
wire n_5913;
wire n_8958;
wire n_13838;
wire n_4530;
wire n_11333;
wire n_11682;
wire n_9821;
wire n_1432;
wire n_2245;
wire n_5614;
wire n_13692;
wire n_16187;
wire n_16483;
wire n_5391;
wire n_5452;
wire n_10715;
wire n_11381;
wire n_3359;
wire n_7944;
wire n_3841;
wire n_11922;
wire n_5249;
wire n_13126;
wire n_249;
wire n_14762;
wire n_851;
wire n_12068;
wire n_444;
wire n_10579;
wire n_3900;
wire n_3413;
wire n_7850;
wire n_5076;
wire n_10707;
wire n_3539;
wire n_5757;
wire n_15682;
wire n_9265;
wire n_6872;
wire n_15357;
wire n_15098;
wire n_12332;
wire n_12858;
wire n_17042;
wire n_6644;
wire n_11352;
wire n_9143;
wire n_5062;
wire n_2134;
wire n_16387;
wire n_3862;
wire n_12641;
wire n_930;
wire n_4912;
wire n_12140;
wire n_9845;
wire n_4226;
wire n_10112;
wire n_14505;
wire n_10556;
wire n_14150;
wire n_4311;
wire n_3284;
wire n_8542;
wire n_8572;
wire n_5046;
wire n_14292;
wire n_7607;
wire n_13330;
wire n_7642;
wire n_8373;
wire n_16075;
wire n_8424;
wire n_13417;
wire n_8442;
wire n_1386;
wire n_9304;
wire n_14492;
wire n_7104;
wire n_6236;
wire n_8147;
wire n_3506;
wire n_15909;
wire n_4827;
wire n_6801;
wire n_11152;
wire n_13505;
wire n_1842;
wire n_4993;
wire n_7397;
wire n_16950;
wire n_3678;
wire n_7205;
wire n_10080;
wire n_366;
wire n_2791;
wire n_14951;
wire n_1661;
wire n_555;
wire n_3212;
wire n_11022;
wire n_4871;
wire n_11025;
wire n_12517;
wire n_16321;
wire n_3529;
wire n_4405;
wire n_16228;
wire n_6563;
wire n_5968;
wire n_11251;
wire n_992;
wire n_966;
wire n_3549;
wire n_13821;
wire n_3914;
wire n_10766;
wire n_13787;
wire n_6398;
wire n_11222;
wire n_5586;
wire n_14065;
wire n_7461;
wire n_8519;
wire n_1692;
wire n_11650;
wire n_14310;
wire n_2611;
wire n_15420;
wire n_14958;
wire n_17115;
wire n_15690;
wire n_8075;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_7638;
wire n_10781;
wire n_2398;
wire n_11091;
wire n_13243;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_8642;
wire n_15565;
wire n_6319;
wire n_11713;
wire n_8648;
wire n_10217;
wire n_16666;
wire n_7224;
wire n_6966;
wire n_9791;
wire n_5056;
wire n_9449;
wire n_16346;
wire n_9934;
wire n_9149;
wire n_9686;
wire n_13063;
wire n_1178;
wire n_2015;
wire n_13186;
wire n_14639;
wire n_15101;
wire n_13463;
wire n_15748;
wire n_7259;
wire n_7838;
wire n_8556;
wire n_5984;
wire n_12961;
wire n_14039;
wire n_11398;
wire n_9844;
wire n_5204;
wire n_6705;
wire n_6724;
wire n_12389;
wire n_2877;
wire n_7307;
wire n_6776;
wire n_15472;
wire n_11208;
wire n_203;
wire n_9458;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_150;
wire n_2930;
wire n_8585;
wire n_7840;
wire n_15994;
wire n_16404;
wire n_9717;
wire n_12595;
wire n_11858;
wire n_16283;
wire n_11487;
wire n_14194;
wire n_2745;
wire n_8455;
wire n_16418;
wire n_2087;
wire n_8444;
wire n_16831;
wire n_13237;
wire n_619;
wire n_9128;
wire n_14788;
wire n_10638;
wire n_14559;
wire n_14255;
wire n_2161;
wire n_11745;
wire n_10239;
wire n_746;
wire n_12368;
wire n_13353;
wire n_6624;
wire n_1357;
wire n_7888;
wire n_8560;
wire n_292;
wire n_15360;
wire n_12816;
wire n_14730;
wire n_11525;
wire n_6710;
wire n_1787;
wire n_6883;
wire n_9558;
wire n_8108;
wire n_16633;
wire n_1389;
wire n_8158;
wire n_3172;
wire n_14990;
wire n_16076;
wire n_2659;
wire n_4033;
wire n_10464;
wire n_13054;
wire n_15923;
wire n_3747;
wire n_10446;
wire n_15010;
wire n_15957;
wire n_14166;
wire n_9715;
wire n_6553;
wire n_4905;
wire n_10219;
wire n_9016;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_6261;
wire n_3651;
wire n_1812;
wire n_9399;
wire n_15615;
wire n_6659;
wire n_16735;
wire n_4894;
wire n_15215;
wire n_16402;
wire n_428;
wire n_7351;
wire n_16803;
wire n_3614;
wire n_7256;
wire n_959;
wire n_12967;
wire n_2257;
wire n_14458;
wire n_1101;
wire n_1343;
wire n_12907;
wire n_14353;
wire n_3116;
wire n_12020;
wire n_4141;
wire n_13877;
wire n_15368;
wire n_3784;
wire n_16211;
wire n_6893;
wire n_12377;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_12007;
wire n_13272;
wire n_11087;
wire n_8814;
wire n_5778;
wire n_7021;
wire n_15779;
wire n_5179;
wire n_2435;
wire n_10394;
wire n_15700;
wire n_6337;
wire n_5680;
wire n_1932;
wire n_7583;
wire n_6210;
wire n_1780;
wire n_14368;
wire n_2825;
wire n_5685;
wire n_13394;
wire n_15240;
wire n_16431;
wire n_5974;
wire n_10776;
wire n_14032;
wire n_14375;
wire n_10917;
wire n_5723;
wire n_14914;
wire n_15815;
wire n_15085;
wire n_542;
wire n_5922;
wire n_6378;
wire n_14822;
wire n_5549;
wire n_1087;
wire n_13536;
wire n_632;
wire n_9094;
wire n_2388;
wire n_13524;
wire n_2273;
wire n_8130;
wire n_15212;
wire n_1911;
wire n_11483;
wire n_14075;
wire n_3496;
wire n_14093;
wire n_4364;
wire n_3493;
wire n_12944;
wire n_14705;
wire n_9510;
wire n_11049;
wire n_7488;
wire n_16101;
wire n_3700;
wire n_7690;
wire n_12706;
wire n_14817;
wire n_12973;
wire n_12319;
wire n_4307;
wire n_14178;
wire n_2795;
wire n_14053;
wire n_6044;
wire n_1841;
wire n_1680;
wire n_15825;
wire n_16567;
wire n_16138;
wire n_12388;
wire n_6206;
wire n_7893;
wire n_2954;
wire n_16807;
wire n_11031;
wire n_382;
wire n_9429;
wire n_14929;
wire n_489;
wire n_11599;
wire n_4438;
wire n_11292;
wire n_15740;
wire n_6538;
wire n_11568;
wire n_15016;
wire n_7966;
wire n_251;
wire n_974;
wire n_506;
wire n_3814;
wire n_6996;
wire n_5831;
wire n_9653;
wire n_4367;
wire n_5134;
wire n_11468;
wire n_13815;
wire n_2467;
wire n_7599;
wire n_9648;
wire n_7231;
wire n_14626;
wire n_10240;
wire n_4195;
wire n_7007;
wire n_7717;
wire n_6579;
wire n_12470;
wire n_12711;
wire n_5091;
wire n_16651;
wire n_4866;
wire n_7230;
wire n_15483;
wire n_1447;
wire n_8675;
wire n_1220;
wire n_12216;
wire n_9095;
wire n_7900;
wire n_11203;
wire n_2019;
wire n_5708;
wire n_8123;
wire n_698;
wire n_9003;
wire n_9048;
wire n_16080;
wire n_12879;
wire n_14228;
wire n_13801;
wire n_16879;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_5454;
wire n_14472;
wire n_13659;
wire n_17015;
wire n_307;
wire n_1209;
wire n_4254;
wire n_10578;
wire n_14946;
wire n_11206;
wire n_646;
wire n_12649;
wire n_12093;
wire n_13473;
wire n_8913;
wire n_9932;
wire n_15247;
wire n_3438;
wire n_16815;
wire n_8220;
wire n_12165;
wire n_15170;
wire n_404;
wire n_2625;
wire n_11779;
wire n_13497;
wire n_16262;
wire n_9309;
wire n_8355;
wire n_12724;
wire n_9661;
wire n_14557;
wire n_9799;
wire n_12447;
wire n_5373;
wire n_7403;
wire n_1578;
wire n_6665;
wire n_8883;
wire n_15480;
wire n_15910;
wire n_3147;
wire n_13822;
wire n_17096;
wire n_299;
wire n_3661;
wire n_7168;
wire n_10427;
wire n_15514;
wire n_15527;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_16975;
wire n_11927;
wire n_11609;
wire n_10626;
wire n_11676;
wire n_16793;
wire n_17143;
wire n_1029;
wire n_2649;
wire n_6033;
wire n_6461;
wire n_10138;
wire n_15556;
wire n_1247;
wire n_6860;
wire n_9063;
wire n_522;
wire n_1568;
wire n_2919;
wire n_7322;
wire n_10364;
wire n_6060;
wire n_10532;
wire n_3108;
wire n_5983;
wire n_5788;
wire n_15734;
wire n_15719;
wire n_9895;
wire n_10288;
wire n_367;
wire n_6709;
wire n_11602;
wire n_15601;
wire n_13843;
wire n_2632;
wire n_11865;
wire n_15263;
wire n_12566;
wire n_5557;
wire n_12383;
wire n_6914;
wire n_8816;
wire n_15873;
wire n_4314;
wire n_8418;
wire n_14943;
wire n_2980;
wire n_5951;
wire n_1728;
wire n_4315;
wire n_5647;
wire n_16145;
wire n_6117;
wire n_7287;
wire n_12035;
wire n_7789;
wire n_15684;
wire n_3239;
wire n_2631;
wire n_12212;
wire n_9110;
wire n_3311;
wire n_11427;
wire n_3516;
wire n_11613;
wire n_15739;
wire n_4442;
wire n_424;
wire n_10668;
wire n_4857;
wire n_8739;
wire n_9969;
wire n_11375;
wire n_8927;
wire n_10398;
wire n_15749;
wire n_1651;
wire n_3087;
wire n_6009;
wire n_11870;
wire n_5523;
wire n_4637;
wire n_12053;
wire n_2697;
wire n_13250;
wire n_7221;
wire n_15004;
wire n_1263;
wire n_1817;
wire n_8243;
wire n_3704;
wire n_8798;
wire n_13228;
wire n_7963;
wire n_13893;
wire n_6382;
wire n_8423;
wire n_13869;
wire n_15278;
wire n_14326;
wire n_9028;
wire n_15335;
wire n_670;
wire n_2677;
wire n_4296;
wire n_14699;
wire n_379;
wire n_138;
wire n_162;
wire n_16539;
wire n_13100;
wire n_9654;
wire n_10683;
wire n_14232;
wire n_16926;
wire n_2483;
wire n_10249;
wire n_7938;
wire n_5088;
wire n_6615;
wire n_17132;
wire n_9810;
wire n_441;
wire n_7294;
wire n_7414;
wire n_5773;
wire n_6192;
wire n_1032;
wire n_12852;
wire n_16907;
wire n_12123;
wire n_1592;
wire n_9701;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_9270;
wire n_11373;
wire n_11878;
wire n_16738;
wire n_3589;
wire n_6418;
wire n_1743;
wire n_8548;
wire n_9437;
wire n_8996;
wire n_13185;
wire n_207;
wire n_9483;
wire n_720;
wire n_6263;
wire n_1943;
wire n_14593;
wire n_8156;
wire n_6731;
wire n_15774;
wire n_5138;
wire n_8845;
wire n_4588;
wire n_16151;
wire n_6048;
wire n_13738;
wire n_7185;
wire n_10229;
wire n_194;
wire n_12268;
wire n_5149;
wire n_9256;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_10889;
wire n_16625;
wire n_11070;
wire n_6234;
wire n_16046;
wire n_4153;
wire n_14966;
wire n_8992;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_7141;
wire n_11107;
wire n_15459;
wire n_2373;
wire n_14116;
wire n_3881;
wire n_13195;
wire n_12298;
wire n_6224;
wire n_12930;
wire n_8510;
wire n_5089;
wire n_11394;
wire n_17005;
wire n_5775;
wire n_9854;
wire n_2099;
wire n_16630;
wire n_3759;
wire n_15190;
wire n_9737;
wire n_8961;
wire n_12890;
wire n_14551;
wire n_9964;
wire n_11154;
wire n_3323;
wire n_16870;
wire n_14940;
wire n_4643;
wire n_9719;
wire n_16822;
wire n_10826;
wire n_6142;
wire n_2617;
wire n_6119;
wire n_10358;
wire n_12301;
wire n_15086;
wire n_13886;
wire n_6619;
wire n_808;
wire n_2476;
wire n_11973;
wire n_13200;
wire n_2814;
wire n_4133;
wire n_11073;
wire n_13876;
wire n_2636;
wire n_1439;
wire n_6759;
wire n_6903;
wire n_3466;
wire n_7416;
wire n_15466;
wire n_2074;
wire n_5031;
wire n_6768;
wire n_1665;
wire n_7092;
wire n_7233;
wire n_2122;
wire n_4543;
wire n_14442;
wire n_4337;
wire n_9679;
wire n_9669;
wire n_11186;
wire n_12382;
wire n_5082;
wire n_4788;
wire n_10835;
wire n_13095;
wire n_12996;
wire n_1414;
wire n_2067;
wire n_16757;
wire n_15947;
wire n_17129;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_10416;
wire n_3465;
wire n_12661;
wire n_8402;
wire n_8978;
wire n_14097;
wire n_15125;
wire n_2117;
wire n_7191;
wire n_14279;
wire n_6189;
wire n_1053;
wire n_5796;
wire n_15339;
wire n_13907;
wire n_9105;
wire n_13085;
wire n_14411;
wire n_7173;
wire n_9699;
wire n_11360;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_6761;
wire n_14304;
wire n_16686;
wire n_9673;
wire n_15313;
wire n_2194;
wire n_10860;
wire n_11823;
wire n_16672;
wire n_4780;
wire n_4640;
wire n_16549;
wire n_8685;
wire n_1828;
wire n_10997;
wire n_16688;
wire n_9240;
wire n_15162;
wire n_1304;
wire n_7202;
wire n_14033;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_2267;
wire n_9212;
wire n_5858;
wire n_13889;
wire n_7445;
wire n_5985;
wire n_8595;
wire n_16778;
wire n_10602;
wire n_15327;
wire n_604;
wire n_12088;
wire n_478;
wire n_11181;
wire n_9040;
wire n_1349;
wire n_9478;
wire n_10261;
wire n_10817;
wire n_12277;
wire n_12062;
wire n_14045;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_9742;
wire n_11806;
wire n_3477;
wire n_7868;
wire n_10124;
wire n_13386;
wire n_16405;
wire n_16999;
wire n_3370;
wire n_874;
wire n_16238;
wire n_7654;
wire n_16604;
wire n_3949;
wire n_2286;
wire n_8779;
wire n_5192;
wire n_15844;
wire n_4247;
wire n_707;
wire n_5051;
wire n_10132;
wire n_15034;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_8520;
wire n_4583;
wire n_17055;
wire n_14305;
wire n_8555;
wire n_12421;
wire n_10730;
wire n_9456;
wire n_6366;
wire n_16742;
wire n_1015;
wire n_11321;
wire n_1162;
wire n_6304;
wire n_4292;
wire n_2118;
wire n_9146;
wire n_11702;
wire n_688;
wire n_7176;
wire n_14233;
wire n_14835;
wire n_636;
wire n_8565;
wire n_8334;
wire n_13605;
wire n_1490;
wire n_6074;
wire n_5552;
wire n_7547;
wire n_12133;
wire n_442;
wire n_11970;
wire n_15167;
wire n_3764;
wire n_1553;
wire n_10111;
wire n_15083;
wire n_13283;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_13596;
wire n_15912;
wire n_3025;
wire n_9573;
wire n_14983;
wire n_15257;
wire n_3051;
wire n_11286;
wire n_986;
wire n_1104;
wire n_2802;
wire n_8030;
wire n_16671;
wire n_8513;
wire n_14511;
wire n_887;
wire n_13746;
wire n_13327;
wire n_14550;
wire n_16921;
wire n_9379;
wire n_10948;
wire n_13534;
wire n_9219;
wire n_16186;
wire n_2125;
wire n_14056;
wire n_10927;
wire n_11496;
wire n_15356;
wire n_1156;
wire n_14151;
wire n_13149;
wire n_4974;
wire n_5123;
wire n_6689;
wire n_2861;
wire n_8245;
wire n_13727;
wire n_13992;
wire n_14846;
wire n_7942;
wire n_4344;
wire n_17178;
wire n_5242;
wire n_12186;
wire n_3130;
wire n_8753;
wire n_1188;
wire n_1498;
wire n_15230;
wire n_7527;
wire n_16487;
wire n_9706;
wire n_4856;
wire n_2618;
wire n_7948;
wire n_7096;
wire n_11863;
wire n_15776;
wire n_4216;
wire n_957;
wire n_1242;
wire n_9206;
wire n_2707;
wire n_14139;
wire n_15002;
wire n_8485;
wire n_5596;
wire n_6482;
wire n_10118;
wire n_8106;
wire n_2849;
wire n_15585;
wire n_1489;
wire n_15847;
wire n_8325;
wire n_2756;
wire n_15329;
wire n_3781;
wire n_14619;
wire n_2217;
wire n_17031;
wire n_10875;
wire n_4864;
wire n_11225;
wire n_15018;
wire n_2226;
wire n_6335;
wire n_5742;
wire n_5127;
wire n_15239;
wire n_10731;
wire n_4313;
wire n_14071;
wire n_15169;
wire n_11355;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_9434;
wire n_3713;
wire n_6229;
wire n_1863;
wire n_5933;
wire n_13113;
wire n_5536;
wire n_13097;
wire n_13198;
wire n_15256;
wire n_15928;
wire n_4798;
wire n_10350;
wire n_10654;
wire n_1500;
wire n_616;
wire n_7293;
wire n_9874;
wire n_11261;
wire n_11862;
wire n_13369;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_12579;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_5810;
wire n_3750;
wire n_10564;
wire n_3424;
wire n_12342;
wire n_13653;
wire n_3356;
wire n_14832;
wire n_14691;
wire n_11584;
wire n_9082;
wire n_7144;
wire n_12877;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_16612;
wire n_12256;
wire n_2516;
wire n_4991;
wire n_11893;
wire n_10262;
wire n_13360;
wire n_11500;
wire n_11044;
wire n_7316;
wire n_7508;
wire n_13785;
wire n_9596;
wire n_15861;
wire n_3070;
wire n_1005;
wire n_8677;
wire n_15065;
wire n_16986;
wire n_16741;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_11109;
wire n_12909;
wire n_13044;
wire n_3245;
wire n_12859;
wire n_16025;
wire n_10729;
wire n_2894;
wire n_9559;
wire n_15463;
wire n_9709;
wire n_10973;
wire n_15525;
wire n_2452;
wire n_4182;
wire n_8626;
wire n_16318;
wire n_12822;
wire n_2827;
wire n_7869;
wire n_13217;
wire n_3214;
wire n_13943;
wire n_10069;
wire n_10810;
wire n_16001;
wire n_12468;
wire n_9356;
wire n_8166;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_14948;
wire n_5009;
wire n_12267;
wire n_15515;
wire n_3710;
wire n_12170;
wire n_12426;
wire n_15689;
wire n_1844;
wire n_15876;
wire n_6943;
wire n_10791;
wire n_1957;
wire n_1953;
wire n_12900;
wire n_10553;
wire n_16532;
wire n_1219;
wire n_14555;
wire n_710;
wire n_16833;
wire n_6631;
wire n_5889;
wire n_12846;
wire n_8602;
wire n_9609;
wire n_15467;
wire n_10284;
wire n_3944;
wire n_7151;
wire n_16736;
wire n_7762;
wire n_13469;
wire n_15346;
wire n_13836;
wire n_13840;
wire n_16343;
wire n_5632;
wire n_17060;
wire n_16970;
wire n_12855;
wire n_11501;
wire n_4729;
wire n_8002;
wire n_6728;
wire n_16260;
wire n_13569;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_7472;
wire n_9342;
wire n_14229;
wire n_4800;
wire n_14425;
wire n_1373;
wire n_15324;
wire n_7075;
wire n_13076;
wire n_1540;
wire n_14917;
wire n_5427;
wire n_12234;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_6770;
wire n_14317;
wire n_5450;
wire n_7611;
wire n_11437;
wire n_7796;
wire n_6508;
wire n_16663;
wire n_14682;
wire n_832;
wire n_13320;
wire n_13082;
wire n_8047;
wire n_12120;
wire n_16598;
wire n_7989;
wire n_15863;
wire n_15064;
wire n_744;
wire n_2821;
wire n_3696;
wire n_9233;
wire n_10474;
wire n_7936;
wire n_10694;
wire n_215;
wire n_10529;
wire n_13117;
wire n_15622;
wire n_16863;
wire n_1331;
wire n_4781;
wire n_12042;
wire n_6031;
wire n_1529;
wire n_3531;
wire n_14328;
wire n_15457;
wire n_5124;
wire n_655;
wire n_16084;
wire n_4237;
wire n_8751;
wire n_5297;
wire n_11722;
wire n_4828;
wire n_3333;
wire n_12568;
wire n_12149;
wire n_14444;
wire n_15138;
wire n_8800;
wire n_4652;
wire n_12278;
wire n_4114;
wire n_7105;
wire n_7013;
wire n_7655;
wire n_10622;
wire n_1007;
wire n_9435;
wire n_1580;
wire n_3135;
wire n_13318;
wire n_4925;
wire n_5719;
wire n_7254;
wire n_2448;
wire n_9557;
wire n_11639;
wire n_2211;
wire n_8955;
wire n_9551;
wire n_16991;
wire n_951;
wire n_8039;
wire n_12231;
wire n_12116;
wire n_13677;
wire n_9073;
wire n_8193;
wire n_7546;
wire n_8432;
wire n_15343;
wire n_17128;
wire n_14422;
wire n_5904;
wire n_11997;
wire n_14876;
wire n_16088;
wire n_6628;
wire n_5318;
wire n_5374;
wire n_8684;
wire n_2424;
wire n_10270;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_6456;
wire n_722;
wire n_16069;
wire n_13158;
wire n_7407;
wire n_12014;
wire n_13230;
wire n_9388;
wire n_3277;
wire n_10463;
wire n_9721;
wire n_11731;
wire n_14061;
wire n_4863;
wire n_10880;
wire n_11610;
wire n_12097;
wire n_14612;
wire n_12363;
wire n_13115;
wire n_16579;
wire n_15599;
wire n_13427;
wire n_16307;
wire n_1766;
wire n_5463;
wire n_16339;
wire n_1338;
wire n_2978;
wire n_6328;
wire n_11498;
wire n_16499;
wire n_12008;
wire n_6929;
wire n_11509;
wire n_4859;
wire n_4568;
wire n_8628;
wire n_15097;
wire n_14401;
wire n_14034;
wire n_15518;
wire n_15820;
wire n_13559;
wire n_15400;
wire n_3617;
wire n_6012;
wire n_704;
wire n_2958;
wire n_15723;
wire n_7481;
wire n_11447;
wire n_1044;
wire n_1714;
wire n_6484;
wire n_5435;
wire n_4429;
wire n_11706;
wire n_3340;
wire n_5053;
wire n_7182;
wire n_11055;
wire n_14498;
wire n_10689;
wire n_9507;
wire n_5476;
wire n_5483;
wire n_12534;
wire n_9539;
wire n_8617;
wire n_14517;
wire n_14297;
wire n_7605;
wire n_8591;
wire n_16362;
wire n_8090;
wire n_1243;
wire n_15513;
wire n_9268;
wire n_5511;
wire n_9718;
wire n_8661;
wire n_13512;
wire n_10068;
wire n_15330;
wire n_16595;
wire n_3486;
wire n_11258;
wire n_6639;
wire n_358;
wire n_608;
wire n_9672;
wire n_12748;
wire n_11168;
wire n_9890;
wire n_12272;
wire n_9187;
wire n_2457;
wire n_9572;
wire n_16272;
wire n_12148;
wire n_2992;
wire n_10363;
wire n_6124;
wire n_16130;
wire n_12142;
wire n_12615;
wire n_16164;
wire n_13201;
wire n_9527;
wire n_317;
wire n_3197;
wire n_11234;
wire n_15375;
wire n_16771;
wire n_9949;
wire n_13388;
wire n_14484;
wire n_7423;
wire n_13674;
wire n_3256;
wire n_1878;
wire n_16308;
wire n_15115;
wire n_7375;
wire n_7076;
wire n_16269;
wire n_7689;
wire n_8189;
wire n_13858;
wire n_8811;
wire n_6344;
wire n_266;
wire n_9952;
wire n_11612;
wire n_7736;
wire n_6435;
wire n_13949;
wire n_10888;
wire n_12714;
wire n_13782;
wire n_14486;
wire n_3646;
wire n_14759;
wire n_5829;
wire n_2520;
wire n_14580;
wire n_7419;
wire n_811;
wire n_13612;
wire n_6600;
wire n_14087;
wire n_13681;
wire n_7010;
wire n_13700;
wire n_14421;
wire n_16095;
wire n_14193;
wire n_791;
wire n_17172;
wire n_10277;
wire n_15242;
wire n_5881;
wire n_9798;
wire n_17041;
wire n_3864;
wire n_4694;
wire n_11895;
wire n_8192;
wire n_9251;
wire n_16972;
wire n_1025;
wire n_4664;
wire n_6201;
wire n_17162;
wire n_10537;
wire n_14703;
wire n_3450;
wire n_14653;
wire n_8573;
wire n_14684;
wire n_687;
wire n_4633;
wire n_13770;
wire n_2026;
wire n_10807;
wire n_4050;
wire n_3173;
wire n_480;
wire n_14048;
wire n_13920;
wire n_7918;
wire n_642;
wire n_9546;
wire n_10331;
wire n_1406;
wire n_5073;
wire n_6555;
wire n_16495;
wire n_4306;
wire n_6360;
wire n_13130;
wire n_6735;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_9181;
wire n_9602;
wire n_12812;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_13377;
wire n_15846;
wire n_11455;
wire n_6803;
wire n_4288;
wire n_3452;
wire n_14816;
wire n_474;
wire n_4098;
wire n_2691;
wire n_10981;
wire n_5894;
wire n_13750;
wire n_9635;
wire n_11868;
wire n_4511;
wire n_3422;
wire n_12639;
wire n_12189;
wire n_14063;
wire n_15542;
wire n_14521;
wire n_4675;
wire n_13701;
wire n_695;
wire n_11934;
wire n_13518;
wire n_2991;
wire n_16571;
wire n_5419;
wire n_8339;
wire n_16506;
wire n_14737;
wire n_386;
wire n_1596;
wire n_11969;
wire n_13668;
wire n_4289;
wire n_4972;
wire n_11571;
wire n_197;
wire n_2723;
wire n_1476;
wire n_6036;
wire n_9405;
wire n_7346;
wire n_2016;
wire n_16561;
wire n_15255;
wire n_3925;
wire n_17007;
wire n_12428;
wire n_12069;
wire n_14384;
wire n_4689;
wire n_5165;
wire n_8775;
wire n_678;
wire n_10780;
wire n_10158;
wire n_11481;
wire n_651;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_6102;
wire n_16173;
wire n_16948;
wire n_14276;
wire n_12057;
wire n_3780;
wire n_12050;
wire n_1657;
wire n_13587;
wire n_9726;
wire n_13488;
wire n_15852;
wire n_8804;
wire n_16559;
wire n_9577;
wire n_6650;
wire n_10024;
wire n_6573;
wire n_11774;
wire n_15271;
wire n_6904;
wire n_12214;
wire n_3753;
wire n_6329;
wire n_13805;
wire n_7385;
wire n_15425;
wire n_9802;
wire n_1488;
wire n_6244;
wire n_4846;
wire n_9250;
wire n_1330;
wire n_906;
wire n_6204;
wire n_9540;
wire n_13365;
wire n_13767;
wire n_13972;
wire n_12381;
wire n_10191;
wire n_2295;
wire n_5225;
wire n_16627;
wire n_283;
wire n_7295;
wire n_4076;
wire n_7824;
wire n_12157;
wire n_7148;
wire n_13938;
wire n_3142;
wire n_9171;
wire n_7169;
wire n_3129;
wire n_16054;
wire n_13443;
wire n_15297;
wire n_9350;
wire n_374;
wire n_3843;
wire n_3495;
wire n_11257;
wire n_12330;
wire n_16909;
wire n_6756;
wire n_17046;
wire n_4805;
wire n_2606;
wire n_9441;
wire n_7600;
wire n_15268;
wire n_15814;
wire n_15838;
wire n_9124;
wire n_10675;
wire n_2386;
wire n_5826;
wire n_8697;
wire n_11598;
wire n_9626;
wire n_14011;
wire n_14645;
wire n_4822;
wire n_11327;
wire n_6946;
wire n_12926;
wire n_7947;
wire n_8645;
wire n_5931;
wire n_8820;
wire n_9408;
wire n_14712;
wire n_1829;
wire n_8146;
wire n_4635;
wire n_8154;
wire n_7847;
wire n_1450;
wire n_12824;
wire n_12392;
wire n_13094;
wire n_5532;
wire n_14545;
wire n_7311;
wire n_3740;
wire n_6804;
wire n_16189;
wire n_5441;
wire n_14103;
wire n_2417;
wire n_6179;
wire n_6059;
wire n_1815;
wire n_16858;
wire n_7039;
wire n_8027;
wire n_7807;
wire n_1493;
wire n_2911;
wire n_14976;
wire n_515;
wire n_8063;
wire n_3313;
wire n_13798;
wire n_14677;
wire n_8406;
wire n_15580;
wire n_2354;
wire n_6427;
wire n_17100;
wire n_14474;
wire n_14459;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_12070;
wire n_3726;
wire n_8480;
wire n_11265;
wire n_14037;
wire n_11788;
wire n_14112;
wire n_14811;
wire n_16696;
wire n_9754;
wire n_10477;
wire n_4419;
wire n_14296;
wire n_11904;
wire n_8849;
wire n_17078;
wire n_13071;
wire n_17063;
wire n_5405;
wire n_9750;
wire n_10296;
wire n_7660;
wire n_13676;
wire n_13735;
wire n_14127;
wire n_1256;
wire n_5365;
wire n_9566;
wire n_3560;
wire n_3345;
wire n_5772;
wire n_9529;
wire n_10339;
wire n_11901;
wire n_12848;
wire n_15528;
wire n_16357;
wire n_6442;
wire n_10307;
wire n_8241;
wire n_140;
wire n_10606;
wire n_6188;
wire n_12161;
wire n_16249;
wire n_3421;
wire n_1448;
wire n_10066;
wire n_11755;
wire n_1009;
wire n_230;
wire n_3548;
wire n_4906;
wire n_11754;
wire n_15610;
wire n_13825;
wire n_6846;
wire n_10054;
wire n_4630;
wire n_8261;
wire n_10343;
wire n_6840;
wire n_142;
wire n_6645;
wire n_16616;
wire n_15020;
wire n_8535;
wire n_8348;
wire n_4829;
wire n_13985;
wire n_16916;
wire n_6749;
wire n_12238;
wire n_6915;
wire n_12956;
wire n_12320;
wire n_7831;
wire n_13342;
wire n_8138;
wire n_2612;
wire n_11413;
wire n_13953;
wire n_10652;
wire n_13040;
wire n_5259;
wire n_15735;
wire n_3236;
wire n_8702;
wire n_11601;
wire n_1995;
wire n_7455;
wire n_8273;
wire n_14250;
wire n_10944;
wire n_16479;
wire n_1397;
wire n_5921;
wire n_6247;
wire n_10367;
wire n_15365;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_11129;
wire n_11710;
wire n_833;
wire n_4966;
wire n_14602;
wire n_2250;
wire n_8235;
wire n_15510;
wire n_17035;
wire n_13685;
wire n_1117;
wire n_6104;
wire n_15476;
wire n_3321;
wire n_9940;
wire n_15444;
wire n_8294;
wire n_1303;
wire n_12476;
wire n_4188;
wire n_10016;
wire n_2001;
wire n_15273;
wire n_9036;
wire n_9165;
wire n_7509;
wire n_9283;
wire n_6205;
wire n_2506;
wire n_11010;
wire n_8349;
wire n_15901;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_9822;
wire n_10036;
wire n_15199;
wire n_2626;
wire n_9607;
wire n_9443;
wire n_7497;
wire n_16201;
wire n_10749;
wire n_17092;
wire n_7315;
wire n_10166;
wire n_8429;
wire n_13765;
wire n_2892;
wire n_6939;
wire n_16214;
wire n_2605;
wire n_7887;
wire n_10419;
wire n_2804;
wire n_15726;
wire n_9298;
wire n_5884;
wire n_16312;
wire n_15470;
wire n_5006;
wire n_14200;
wire n_4882;
wire n_3206;
wire n_10006;
wire n_5728;
wire n_1035;
wire n_13334;
wire n_3475;
wire n_14902;
wire n_4878;
wire n_8486;
wire n_11240;
wire n_9052;
wire n_2070;
wire n_426;
wire n_6706;
wire n_13123;
wire n_12154;
wire n_16149;
wire n_7431;
wire n_8140;
wire n_398;
wire n_11734;
wire n_14450;
wire n_3842;
wire n_12645;
wire n_15276;
wire n_1367;
wire n_14477;
wire n_4202;
wire n_6909;
wire n_13933;
wire n_2044;
wire n_5679;
wire n_6487;
wire n_166;
wire n_12668;
wire n_8117;
wire n_15143;
wire n_15633;
wire n_3886;
wire n_10348;
wire n_13884;
wire n_825;
wire n_732;
wire n_2619;
wire n_7521;
wire n_10058;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_6627;
wire n_4503;
wire n_15975;
wire n_8129;
wire n_1291;
wire n_11156;
wire n_10355;
wire n_7253;
wire n_5208;
wire n_9535;
wire n_16933;
wire n_13511;
wire n_5113;
wire n_10304;
wire n_12928;
wire n_3987;
wire n_11955;
wire n_5205;
wire n_4249;
wire n_15110;
wire n_9943;
wire n_7569;
wire n_12538;
wire n_13745;
wire n_12151;
wire n_16202;
wire n_3160;
wire n_10966;
wire n_14697;
wire n_13112;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_13646;
wire n_12130;
wire n_14608;
wire n_15049;
wire n_2711;
wire n_3223;
wire n_7452;
wire n_12409;
wire n_13031;
wire n_6551;
wire n_3386;
wire n_12350;
wire n_400;
wire n_15767;
wire n_7972;
wire n_8672;
wire n_13455;
wire n_15411;
wire n_7505;
wire n_13993;
wire n_17073;
wire n_3921;
wire n_282;
wire n_14280;
wire n_16545;
wire n_467;
wire n_2177;
wire n_13946;
wire n_16884;
wire n_6516;
wire n_14567;
wire n_2766;
wire n_10060;
wire n_7524;
wire n_16668;
wire n_16600;
wire n_15763;
wire n_13931;
wire n_4196;
wire n_1197;
wire n_11270;
wire n_8934;
wire n_14961;
wire n_11020;
wire n_7318;
wire n_2613;
wire n_9977;
wire n_10722;
wire n_13314;
wire n_7411;
wire n_13378;
wire n_7326;
wire n_5667;
wire n_168;
wire n_9555;
wire n_15980;
wire n_1517;
wire n_13618;
wire n_10957;
wire n_2647;
wire n_14277;
wire n_8847;
wire n_16524;
wire n_8005;
wire n_5508;
wire n_16659;
wire n_5105;
wire n_3920;
wire n_11344;
wire n_15446;
wire n_3444;
wire n_14952;
wire n_3851;
wire n_16624;
wire n_5879;
wire n_1671;
wire n_6500;
wire n_11303;
wire n_5027;
wire n_1048;
wire n_2343;
wire n_775;
wire n_12847;
wire n_667;
wire n_3380;
wire n_14340;
wire n_16891;
wire n_16995;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_9030;
wire n_869;
wire n_11216;
wire n_15652;
wire n_846;
wire n_1398;
wire n_1921;
wire n_8221;
wire n_13638;
wire n_7573;
wire n_6630;
wire n_14886;
wire n_5629;
wire n_5759;
wire n_10409;
wire n_2411;
wire n_13167;
wire n_4631;
wire n_8191;
wire n_6798;
wire n_13758;
wire n_5999;
wire n_1504;
wire n_9590;
wire n_2110;
wire n_14646;
wire n_11511;
wire n_7498;
wire n_7895;
wire n_6421;
wire n_10322;
wire n_16655;
wire n_11339;
wire n_11346;
wire n_11829;
wire n_12680;
wire n_5377;
wire n_6180;
wire n_12530;
wire n_17002;
wire n_11581;
wire n_8225;
wire n_16721;
wire n_3822;
wire n_889;
wire n_4355;
wire n_7453;
wire n_3818;
wire n_12163;
wire n_16184;
wire n_14131;
wire n_7932;
wire n_9651;
wire n_7890;
wire n_5599;
wire n_10825;
wire n_16199;
wire n_3587;
wire n_16129;
wire n_2608;
wire n_15575;
wire n_6004;
wire n_9583;
wire n_16347;
wire n_9763;
wire n_10349;
wire n_9944;
wire n_13709;
wire n_13035;
wire n_1948;
wire n_6652;
wire n_9888;
wire n_7183;
wire n_4155;
wire n_810;
wire n_10040;
wire n_10844;
wire n_10636;
wire n_4710;
wire n_12738;
wire n_4278;
wire n_1959;
wire n_6275;
wire n_6403;
wire n_3497;
wire n_6395;
wire n_9862;
wire n_14622;
wire n_4542;
wire n_5451;
wire n_6578;
wire n_3243;
wire n_15267;
wire n_4326;
wire n_9966;
wire n_2121;
wire n_15455;
wire n_10242;
wire n_3865;
wire n_6350;
wire n_16115;
wire n_5460;
wire n_4685;
wire n_16023;
wire n_9936;
wire n_565;
wire n_3927;
wire n_6141;
wire n_8559;
wire n_11165;
wire n_2068;
wire n_3595;
wire n_7189;
wire n_6875;
wire n_1194;
wire n_9617;
wire n_10727;
wire n_4060;
wire n_1647;
wire n_9341;
wire n_6194;
wire n_14984;
wire n_1454;
wire n_14864;
wire n_2459;
wire n_15000;
wire n_941;
wire n_8689;
wire n_11231;
wire n_3396;
wire n_9749;
wire n_5517;
wire n_9629;
wire n_13654;
wire n_5807;
wire n_14985;
wire n_15944;
wire n_11448;
wire n_12227;
wire n_5426;
wire n_6475;
wire n_12525;
wire n_10679;
wire n_4093;
wire n_11132;
wire n_452;
wire n_10524;
wire n_12282;
wire n_5693;
wire n_13426;
wire n_5695;
wire n_12932;
wire n_14849;
wire n_4123;
wire n_13799;
wire n_14207;
wire n_16064;
wire n_16407;
wire n_4294;
wire n_8330;
wire n_10011;
wire n_1521;
wire n_12037;
wire n_1940;
wire n_3683;
wire n_6502;
wire n_11410;
wire n_6944;
wire n_10030;
wire n_14365;
wire n_4452;
wire n_15147;
wire n_284;
wire n_3887;
wire n_16288;
wire n_3195;
wire n_8304;
wire n_9349;
wire n_13480;
wire n_15658;
wire n_5587;
wire n_4722;
wire n_11267;
wire n_16929;
wire n_13780;
wire n_6318;
wire n_10119;
wire n_11348;
wire n_11940;
wire n_16726;
wire n_13613;
wire n_10845;
wire n_8163;
wire n_6805;
wire n_11947;
wire n_3048;
wire n_3339;
wire n_16914;
wire n_4126;
wire n_5030;
wire n_4164;
wire n_7240;
wire n_15630;
wire n_8907;
wire n_409;
wire n_2963;
wire n_14227;
wire n_5674;
wire n_2561;
wire n_7499;
wire n_9423;
wire n_1056;
wire n_526;
wire n_5584;
wire n_674;
wire n_12424;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_15227;
wire n_1653;
wire n_6075;
wire n_10063;
wire n_12942;
wire n_6559;
wire n_4088;
wire n_9038;
wire n_8777;
wire n_11149;
wire n_2669;
wire n_8698;
wire n_10709;
wire n_3911;
wire n_6068;
wire n_3802;
wire n_12236;
wire n_4366;
wire n_1584;
wire n_6541;
wire n_11436;
wire n_13326;
wire n_9034;
wire n_848;
wire n_5125;
wire n_4922;
wire n_11909;
wire n_12547;
wire n_13554;
wire n_6066;
wire n_14372;
wire n_6080;
wire n_629;
wire n_13421;
wire n_4733;
wire n_7927;
wire n_161;
wire n_8928;
wire n_13967;
wire n_1814;
wire n_13150;
wire n_13014;
wire n_7219;
wire n_2441;
wire n_10526;
wire n_11439;
wire n_8081;
wire n_12192;
wire n_4041;
wire n_12747;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_216;
wire n_6150;
wire n_11462;
wire n_14564;
wire n_6638;
wire n_16155;
wire n_7063;
wire n_7402;
wire n_9676;
wire n_6351;
wire n_4509;
wire n_4935;
wire n_2073;
wire n_7382;
wire n_8384;
wire n_10861;
wire n_4004;
wire n_5238;
wire n_750;
wire n_13795;
wire n_834;
wire n_8650;
wire n_14729;
wire n_14992;
wire n_3630;
wire n_1612;
wire n_11272;
wire n_800;
wire n_14044;
wire n_12989;
wire n_16415;
wire n_1910;
wire n_5906;
wire n_16005;
wire n_16792;
wire n_7767;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2672;
wire n_2018;
wire n_11759;
wire n_10494;
wire n_14431;
wire n_2602;
wire n_16908;
wire n_17001;
wire n_16258;
wire n_5780;
wire n_10478;
wire n_11061;
wire n_724;
wire n_11653;
wire n_2931;
wire n_3433;
wire n_8284;
wire n_10534;
wire n_8374;
wire n_5556;
wire n_16702;
wire n_6006;
wire n_3597;
wire n_6474;
wire n_13662;
wire n_13864;
wire n_16677;
wire n_5743;
wire n_6481;
wire n_10078;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_5633;
wire n_11478;
wire n_12273;
wire n_7510;
wire n_15475;
wire n_9041;
wire n_3786;
wire n_875;
wire n_15809;
wire n_9995;
wire n_12200;
wire n_6022;
wire n_10629;
wire n_13863;
wire n_2828;
wire n_6991;
wire n_7434;
wire n_1626;
wire n_5950;
wire n_1335;
wire n_9035;
wire n_13926;
wire n_16320;
wire n_9011;
wire n_1715;
wire n_14240;
wire n_4204;
wire n_7691;
wire n_296;
wire n_3553;
wire n_5323;
wire n_7745;
wire n_11748;
wire n_14165;
wire n_17110;
wire n_9135;
wire n_9776;
wire n_3645;
wire n_6744;
wire n_793;
wire n_15055;
wire n_5705;
wire n_12660;
wire n_11867;
wire n_14192;
wire n_15673;
wire n_14678;
wire n_6927;
wire n_7335;
wire n_12400;
wire n_13072;
wire n_14708;
wire n_10695;
wire n_10472;
wire n_17099;
wire n_10286;
wire n_9413;
wire n_4996;
wire n_9107;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_16718;
wire n_17068;
wire n_15823;
wire n_4317;
wire n_7735;
wire n_8531;
wire n_15713;
wire n_6116;
wire n_9548;
wire n_8074;
wire n_15117;
wire n_15479;
wire n_14246;
wire n_494;
wire n_3550;
wire n_8780;
wire n_7956;
wire n_5510;
wire n_15536;
wire n_7651;
wire n_7495;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_9775;
wire n_13857;
wire n_16143;
wire n_16867;
wire n_13033;
wire n_1805;
wire n_12922;
wire n_8580;
wire n_4068;
wire n_15736;
wire n_5440;
wire n_12193;
wire n_9288;
wire n_2270;
wire n_4163;
wire n_15594;
wire n_16036;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_185;
wire n_5011;
wire n_6757;
wire n_7536;
wire n_1554;
wire n_3279;
wire n_15047;
wire n_12243;
wire n_5513;
wire n_10218;
wire n_5875;
wire n_14671;
wire n_16855;
wire n_8358;
wire n_972;
wire n_7734;
wire n_4262;
wire n_2923;
wire n_10441;
wire n_164;
wire n_2843;
wire n_3714;
wire n_9305;
wire n_9093;
wire n_184;
wire n_11764;
wire n_13696;
wire n_15200;
wire n_7671;
wire n_15924;
wire n_16045;
wire n_12950;
wire n_10043;
wire n_4832;
wire n_8033;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_6485;
wire n_13041;
wire n_15021;
wire n_5848;
wire n_1679;
wire n_5834;
wire n_14269;
wire n_7926;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_11882;
wire n_5784;
wire n_13418;
wire n_14820;
wire n_3125;
wire n_12250;
wire n_5128;
wire n_10628;
wire n_13498;
wire n_14290;
wire n_15806;
wire n_16358;
wire n_8643;
wire n_15715;
wire n_2356;
wire n_14792;
wire n_11787;
wire n_12403;
wire n_5618;
wire n_11539;
wire n_15760;
wire n_15099;
wire n_10440;
wire n_15618;
wire n_10134;
wire n_12904;
wire n_6495;
wire n_7528;
wire n_14669;
wire n_12444;
wire n_11163;
wire n_6209;
wire n_16107;
wire n_4672;
wire n_8094;
wire n_2564;
wire n_3558;
wire n_11695;
wire n_13489;
wire n_14520;
wire n_9425;
wire n_15225;
wire n_13373;
wire n_3034;
wire n_10317;
wire n_13739;
wire n_11730;
wire n_13101;
wire n_11916;
wire n_13723;
wire n_3502;
wire n_783;
wire n_13000;
wire n_13556;
wire n_15238;
wire n_4053;
wire n_16713;
wire n_14821;
wire n_11311;
wire n_1127;
wire n_14525;
wire n_7413;
wire n_14435;
wire n_7993;
wire n_11980;
wire n_7821;
wire n_160;
wire n_11151;
wire n_14238;
wire n_7620;
wire n_15520;
wire n_1008;
wire n_3963;
wire n_13153;
wire n_12837;
wire n_12356;
wire n_581;
wire n_15195;
wire n_3091;
wire n_13091;
wire n_13937;
wire n_13032;
wire n_16442;
wire n_6274;
wire n_1024;
wire n_176;
wire n_5157;
wire n_12764;
wire n_14654;
wire n_4496;
wire n_9347;
wire n_12269;
wire n_16962;
wire n_14556;
wire n_2518;
wire n_12079;
wire n_14687;
wire n_936;
wire n_13508;
wire n_10706;
wire n_4596;
wire n_5178;
wire n_9420;
wire n_13350;
wire n_13901;
wire n_12972;
wire n_3105;
wire n_6237;
wire n_13635;
wire n_1525;
wire n_4628;
wire n_6802;
wire n_13224;
wire n_7343;
wire n_16163;
wire n_5982;
wire n_8477;
wire n_16548;
wire n_1775;
wire n_908;
wire n_13306;
wire n_1036;
wire n_9344;
wire n_14657;
wire n_12438;
wire n_7109;
wire n_8028;
wire n_15435;
wire n_16082;
wire n_14245;
wire n_14254;
wire n_12125;
wire n_341;
wire n_4083;
wire n_14993;
wire n_1270;
wire n_12554;
wire n_10297;
wire n_1272;
wire n_549;
wire n_15608;
wire n_2794;
wire n_6155;
wire n_2901;
wire n_7506;
wire n_3940;
wire n_9530;
wire n_6809;
wire n_10160;
wire n_6099;
wire n_10849;
wire n_3225;
wire n_10605;
wire n_11296;
wire n_13259;
wire n_8530;
wire n_14343;
wire n_15165;
wire n_10379;
wire n_9446;
wire n_15434;
wire n_3621;
wire n_5529;
wire n_15094;
wire n_244;
wire n_16234;
wire n_7561;
wire n_3473;
wire n_6349;
wire n_3680;
wire n_11081;
wire n_8500;
wire n_13278;
wire n_8713;
wire n_6716;
wire n_12860;
wire n_3565;
wire n_7885;
wire n_14554;
wire n_8297;
wire n_14100;
wire n_15410;
wire n_6905;
wire n_15519;
wire n_15616;
wire n_8926;
wire n_9865;
wire n_14974;
wire n_8456;
wire n_7722;
wire n_5388;
wire n_7470;
wire n_11230;
wire n_5824;
wire n_8025;
wire n_10282;
wire n_5354;
wire n_15498;
wire n_2453;
wire n_7898;
wire n_11357;
wire n_3331;
wire n_11027;
wire n_13179;
wire n_1788;
wire n_10458;
wire n_12206;
wire n_11393;
wire n_6203;
wire n_12947;
wire n_2138;
wire n_6407;
wire n_14468;
wire n_3040;
wire n_4230;
wire n_11892;
wire n_6899;
wire n_7980;
wire n_7817;
wire n_6413;
wire n_445;
wire n_3360;
wire n_1930;
wire n_17111;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_7070;
wire n_9025;
wire n_17097;
wire n_2000;
wire n_5276;
wire n_11105;
wire n_4037;
wire n_9713;
wire n_11160;
wire n_13043;
wire n_3804;
wire n_14675;
wire n_4659;
wire n_8293;
wire n_13962;
wire n_3211;
wire n_7299;
wire n_917;
wire n_5196;
wire n_2440;
wire n_2096;
wire n_2556;
wire n_10382;
wire n_8029;
wire n_14892;
wire n_2215;
wire n_13468;
wire n_9314;
wire n_3847;
wire n_12270;
wire n_15830;
wire n_15325;
wire n_6960;
wire n_4073;
wire n_14235;
wire n_8880;
wire n_1261;
wire n_7249;
wire n_16715;
wire n_9660;
wire n_16675;
wire n_5763;
wire n_3633;
wire n_15062;
wire n_857;
wire n_13018;
wire n_363;
wire n_12739;
wire n_6061;
wire n_1235;
wire n_13831;
wire n_16105;
wire n_9769;
wire n_2584;
wire n_4001;
wire n_8471;
wire n_1462;
wire n_15031;
wire n_5701;
wire n_7002;
wire n_14529;
wire n_15940;
wire n_1064;
wire n_633;
wire n_16758;
wire n_1446;
wire n_15688;
wire n_12906;
wire n_16436;
wire n_12490;
wire n_9902;
wire n_1701;
wire n_6273;
wire n_14424;
wire n_7094;
wire n_7396;
wire n_3111;
wire n_12751;
wire n_11397;
wire n_16601;
wire n_8726;
wire n_10640;
wire n_731;
wire n_8977;
wire n_1813;
wire n_315;
wire n_2997;
wire n_7018;
wire n_16783;
wire n_11897;
wire n_14949;
wire n_10522;
wire n_1573;
wire n_6746;
wire n_15248;
wire n_3258;
wire n_10691;
wire n_758;
wire n_12650;
wire n_10914;
wire n_10244;
wire n_10764;
wire n_13348;
wire n_7175;
wire n_3691;
wire n_2252;
wire n_8316;
wire n_6174;
wire n_10272;
wire n_15070;
wire n_6545;
wire n_14690;
wire n_6763;
wire n_7773;
wire n_15116;
wire n_1996;
wire n_1106;
wire n_13415;
wire n_2009;
wire n_5907;
wire n_784;
wire n_4339;
wire n_7297;
wire n_7730;
wire n_10980;
wire n_12279;
wire n_13265;
wire n_8134;
wire n_17027;
wire n_6013;
wire n_6182;
wire n_6754;
wire n_4690;
wire n_14916;
wire n_2987;
wire n_6279;
wire n_1473;
wire n_16315;
wire n_1076;
wire n_1348;
wire n_5895;
wire n_9588;
wire n_2651;
wire n_753;
wire n_12242;
wire n_9410;
wire n_2445;
wire n_2733;
wire n_16285;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_10071;
wire n_4023;
wire n_8610;
wire n_4253;
wire n_7637;
wire n_2522;
wire n_3632;
wire n_12588;
wire n_309;
wire n_1344;
wire n_485;
wire n_16241;
wire n_4064;
wire n_16296;
wire n_3351;
wire n_5478;
wire n_13382;
wire n_6131;
wire n_16703;
wire n_10176;
wire n_435;
wire n_6113;
wire n_1141;
wire n_3457;
wire n_9740;
wire n_14767;
wire n_5384;
wire n_6477;
wire n_7486;
wire n_840;
wire n_2324;
wire n_11719;
wire n_6575;
wire n_5283;
wire n_9910;
wire n_3454;
wire n_5961;
wire n_7544;
wire n_2139;
wire n_7613;
wire n_9061;
wire n_15178;
wire n_15810;
wire n_7995;
wire n_9941;
wire n_14794;
wire n_8113;
wire n_9579;
wire n_2521;
wire n_5686;
wire n_6391;
wire n_10254;
wire n_2740;
wire n_14446;
wire n_1991;
wire n_8724;
wire n_14121;
wire n_10332;
wire n_14955;
wire n_15877;
wire n_15769;
wire n_16117;
wire n_7140;
wire n_12775;
wire n_614;
wire n_12173;
wire n_4066;
wire n_10938;
wire n_10257;
wire n_9668;
wire n_6252;
wire n_6426;
wire n_14031;
wire n_4681;
wire n_11956;
wire n_8253;
wire n_12167;
wire n_15091;
wire n_9258;
wire n_15033;
wire n_9228;
wire n_3303;
wire n_13461;
wire n_17056;
wire n_7910;
wire n_6592;
wire n_4414;
wire n_10214;
wire n_11874;
wire n_2541;
wire n_16626;
wire n_5094;
wire n_10195;
wire n_14918;
wire n_16096;
wire n_3232;
wire n_13979;
wire n_1113;
wire n_9598;
wire n_10354;
wire n_248;
wire n_7741;
wire n_12060;
wire n_3768;
wire n_4295;
wire n_10436;
wire n_1615;
wire n_11450;
wire n_4100;
wire n_228;
wire n_11723;
wire n_6668;
wire n_9311;
wire n_11982;
wire n_1265;
wire n_14062;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_11822;
wire n_12179;
wire n_14448;
wire n_11522;
wire n_4087;
wire n_8232;
wire n_12842;
wire n_1409;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_8803;
wire n_10866;
wire n_1673;
wire n_4473;
wire n_14715;
wire n_4619;
wire n_12499;
wire n_6670;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_17043;
wire n_5026;
wire n_16316;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_7679;
wire n_3018;
wire n_8818;
wire n_16525;
wire n_12693;
wire n_14906;
wire n_16764;
wire n_10811;
wire n_7698;
wire n_1875;
wire n_10073;
wire n_14873;
wire n_6962;
wire n_14187;
wire n_16927;
wire n_2429;
wire n_6779;
wire n_10164;
wire n_5286;
wire n_9608;
wire n_4449;
wire n_14779;
wire n_13172;
wire n_3285;
wire n_4607;
wire n_10205;
wire n_1039;
wire n_16800;
wire n_5676;
wire n_16065;
wire n_14716;
wire n_5949;
wire n_5040;
wire n_10515;
wire n_12326;
wire n_1150;
wire n_7800;
wire n_15438;
wire n_6901;
wire n_4266;
wire n_6336;
wire n_13713;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_15384;
wire n_4695;
wire n_6503;
wire n_15362;
wire n_7835;
wire n_1136;
wire n_12542;
wire n_16040;
wire n_15080;
wire n_13650;
wire n_458;
wire n_15187;
wire n_1190;
wire n_16276;
wire n_6049;
wire n_5885;
wire n_11499;
wire n_3628;
wire n_14390;
wire n_9818;
wire n_7100;
wire n_4777;
wire n_7243;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_11034;
wire n_7415;
wire n_14747;
wire n_8823;
wire n_5399;
wire n_8536;
wire n_14004;
wire n_9433;
wire n_16563;
wire n_11746;
wire n_658;
wire n_11698;
wire n_15462;
wire n_362;
wire n_8795;
wire n_2846;
wire n_16526;
wire n_3371;
wire n_10430;
wire n_12934;
wire n_11560;
wire n_10338;
wire n_9599;
wire n_8674;
wire n_9186;
wire n_14054;
wire n_4918;
wire n_5856;
wire n_8016;
wire n_13941;
wire n_15805;
wire n_3872;
wire n_5760;
wire n_12483;
wire n_7747;
wire n_9935;
wire n_14263;
wire n_17107;
wire n_12404;
wire n_12258;
wire n_4415;
wire n_16449;
wire n_5110;
wire n_8966;
wire n_11871;
wire n_14694;
wire n_1964;
wire n_3659;
wire n_14872;
wire n_3928;
wire n_14826;
wire n_16291;
wire n_7552;
wire n_10018;
wire n_9537;
wire n_10500;
wire n_1777;
wire n_9552;
wire n_9421;
wire n_3366;
wire n_15537;
wire n_6998;
wire n_7395;
wire n_16537;
wire n_13209;
wire n_15888;
wire n_5844;
wire n_10359;
wire n_6298;
wire n_8132;
wire n_7650;
wire n_3441;
wire n_199;
wire n_3020;
wire n_12823;
wire n_4146;
wire n_4947;
wire n_7535;
wire n_14775;
wire n_15795;
wire n_708;
wire n_6609;
wire n_10548;
wire n_2545;
wire n_2513;
wire n_7635;
wire n_4408;
wire n_12905;
wire n_10291;
wire n_2115;
wire n_15124;
wire n_8567;
wire n_8259;
wire n_15638;
wire n_2017;
wire n_10667;
wire n_1810;
wire n_12274;
wire n_12849;
wire n_1347;
wire n_11167;
wire n_11297;
wire n_4976;
wire n_9473;
wire n_860;
wire n_6525;
wire n_10208;
wire n_11183;
wire n_3555;
wire n_9469;
wire n_11285;
wire n_5938;
wire n_14270;
wire n_7274;
wire n_3534;
wire n_450;
wire n_11740;
wire n_8578;
wire n_14859;
wire n_10757;
wire n_4548;
wire n_7819;
wire n_8495;
wire n_15428;
wire n_14679;
wire n_2670;
wire n_13975;
wire n_6494;
wire n_15680;
wire n_3556;
wire n_896;
wire n_4574;
wire n_15624;
wire n_8160;
wire n_8980;
wire n_2644;
wire n_6132;
wire n_10631;
wire n_10864;
wire n_11136;
wire n_4557;
wire n_3071;
wire n_11434;
wire n_16480;
wire n_8336;
wire n_11133;
wire n_1698;
wire n_14710;
wire n_14781;
wire n_13711;
wire n_1337;
wire n_774;
wire n_2148;
wire n_5548;
wire n_7788;
wire n_16903;
wire n_16261;
wire n_6974;
wire n_13477;
wire n_1168;
wire n_10748;
wire n_14783;
wire n_4663;
wire n_219;
wire n_5840;
wire n_6882;
wire n_3296;
wire n_9909;
wire n_15087;
wire n_3794;
wire n_3762;
wire n_15718;
wire n_4624;
wire n_16024;
wire n_16877;
wire n_656;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_6498;
wire n_12303;
wire n_6562;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_12002;
wire n_15512;
wire n_8600;
wire n_8229;
wire n_12442;
wire n_415;
wire n_4686;
wire n_9236;
wire n_9751;
wire n_2384;
wire n_10751;
wire n_14649;
wire n_7794;
wire n_17131;
wire n_1705;
wire n_13579;
wire n_768;
wire n_3707;
wire n_1091;
wire n_3895;
wire n_10434;
wire n_16079;
wire n_16311;
wire n_9369;
wire n_3149;
wire n_3934;
wire n_13634;
wire n_14844;
wire n_16846;
wire n_4338;
wire n_13987;
wire n_12597;
wire n_5917;
wire n_15853;
wire n_9757;
wire n_12419;
wire n_6965;
wire n_16399;
wire n_11886;
wire n_2058;
wire n_3231;
wire n_14804;
wire n_14210;
wire n_8761;
wire n_15732;
wire n_1846;
wire n_14316;
wire n_7630;
wire n_15607;
wire n_11804;
wire n_16731;
wire n_13262;
wire n_4161;
wire n_304;
wire n_14673;
wire n_9076;
wire n_17036;
wire n_6168;
wire n_17049;
wire n_5304;
wire n_15943;
wire n_5437;
wire n_6951;
wire n_6963;
wire n_16416;
wire n_1581;
wire n_946;
wire n_757;
wire n_2047;
wire n_3058;
wire n_375;
wire n_1655;
wire n_3709;
wire n_3398;
wire n_1146;
wire n_5355;
wire n_9729;
wire n_11531;
wire n_12943;
wire n_13543;
wire n_6284;
wire n_998;
wire n_3592;
wire n_12039;
wire n_15024;
wire n_16203;
wire n_10663;
wire n_14393;
wire n_5321;
wire n_14144;
wire n_7454;
wire n_2536;
wire n_10263;
wire n_12295;
wire n_1604;
wire n_3399;
wire n_8473;
wire n_9366;
wire n_4772;
wire n_11883;
wire n_6931;
wire n_8351;
wire n_6521;
wire n_5915;
wire n_7276;
wire n_174;
wire n_11792;
wire n_6379;
wire n_16059;
wire n_9647;
wire n_12410;
wire n_1368;
wire n_963;
wire n_7085;
wire n_6306;
wire n_12938;
wire n_4120;
wire n_925;
wire n_7753;
wire n_12891;
wire n_13493;
wire n_12304;
wire n_6834;
wire n_2880;
wire n_1313;
wire n_1001;
wire n_3722;
wire n_4716;
wire n_4654;
wire n_1115;
wire n_8948;
wire n_13166;
wire n_14760;
wire n_13541;
wire n_15412;
wire n_15695;
wire n_1339;
wire n_12572;
wire n_10318;
wire n_13551;
wire n_1051;
wire n_14356;
wire n_5116;
wire n_3771;
wire n_10740;
wire n_7225;
wire n_15131;
wire n_719;
wire n_11634;
wire n_15535;
wire n_7541;
wire n_3158;
wire n_11039;
wire n_3221;
wire n_10062;
wire n_2316;
wire n_7913;
wire n_10128;
wire n_8020;
wire n_7946;
wire n_8944;
wire n_1010;
wire n_2830;
wire n_10717;
wire n_11965;
wire n_5500;
wire n_13890;
wire n_9275;
wire n_4622;
wire n_15158;
wire n_15265;
wire n_4757;
wire n_15955;
wire n_803;
wire n_1871;
wire n_9520;
wire n_6471;
wire n_6949;
wire n_11477;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_9493;
wire n_6760;
wire n_14852;
wire n_2940;
wire n_15006;
wire n_548;
wire n_3427;
wire n_8875;
wire n_3162;
wire n_5966;
wire n_4591;
wire n_5569;
wire n_9102;
wire n_14128;
wire n_5515;
wire n_11588;
wire n_11818;
wire n_6589;
wire n_11592;
wire n_3083;
wire n_4570;
wire n_10721;
wire n_7014;
wire n_10945;
wire n_12290;
wire n_9801;
wire n_11742;
wire n_2491;
wire n_13902;
wire n_12718;
wire n_7920;
wire n_16452;
wire n_11312;
wire n_1931;
wire n_5559;
wire n_8649;
wire n_2259;
wire n_5337;
wire n_849;
wire n_11235;
wire n_5059;
wire n_4655;
wire n_7459;
wire n_14185;
wire n_1820;
wire n_7841;
wire n_10013;
wire n_9424;
wire n_7324;
wire n_7160;
wire n_9333;
wire n_16099;
wire n_8205;
wire n_11505;
wire n_12469;
wire n_15387;
wire n_15986;
wire n_6046;
wire n_11673;
wire n_7054;
wire n_1233;
wire n_4493;
wire n_8975;
wire n_16896;
wire n_6055;
wire n_7161;
wire n_9004;
wire n_1808;
wire n_6364;
wire n_8919;
wire n_6091;
wire n_6348;
wire n_9987;
wire n_1635;
wire n_8440;
wire n_11555;
wire n_1704;
wire n_13917;
wire n_15102;
wire n_15663;
wire n_4896;
wire n_8041;
wire n_16388;
wire n_4851;
wire n_16920;
wire n_9860;
wire n_2479;
wire n_10565;
wire n_6848;
wire n_886;
wire n_14327;
wire n_7837;
wire n_359;
wire n_13548;
wire n_9670;
wire n_6788;
wire n_1308;
wire n_13903;
wire n_11241;
wire n_6144;
wire n_15730;
wire n_15868;
wire n_10389;
wire n_1451;
wire n_16810;
wire n_1487;
wire n_675;
wire n_9200;
wire n_5528;
wire n_15035;
wire n_7806;
wire n_5605;
wire n_15905;
wire n_17108;
wire n_3432;
wire n_2163;
wire n_12336;
wire n_1938;
wire n_13080;
wire n_11059;
wire n_9417;
wire n_6896;
wire n_15534;
wire n_2484;
wire n_16729;
wire n_5753;
wire n_15681;
wire n_5358;
wire n_8076;
wire n_12248;
wire n_12931;
wire n_1469;
wire n_14047;
wire n_11066;
wire n_16200;
wire n_4901;
wire n_3480;
wire n_8757;
wire n_1355;
wire n_10020;
wire n_7201;
wire n_16669;
wire n_13408;
wire n_4213;
wire n_4127;
wire n_6221;
wire n_2500;
wire n_9386;
wire n_12713;
wire n_8897;
wire n_12810;
wire n_7676;
wire n_8177;
wire n_11683;
wire n_13733;
wire n_2334;
wire n_14311;
wire n_5467;
wire n_7241;
wire n_15612;
wire n_1169;
wire n_789;
wire n_3181;
wire n_14147;
wire n_5493;
wire n_9207;
wire n_13592;
wire n_1916;
wire n_6285;
wire n_12717;
wire n_10356;
wire n_610;
wire n_13915;
wire n_16645;
wire n_7644;
wire n_9276;
wire n_4602;
wire n_1713;
wire n_14186;
wire n_8829;
wire n_12119;
wire n_7816;
wire n_1436;
wire n_2818;
wire n_14149;
wire n_4900;
wire n_10110;
wire n_17038;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_6748;
wire n_11275;
wire n_7430;
wire n_14540;
wire n_13589;
wire n_3487;
wire n_16267;
wire n_16618;
wire n_3668;
wire n_11329;
wire n_17091;
wire n_2011;
wire n_8638;
wire n_1515;
wire n_817;
wire n_14272;
wire n_13189;
wire n_13260;
wire n_5901;
wire n_9980;
wire n_1566;
wire n_2837;
wire n_11923;
wire n_717;
wire n_952;
wire n_11718;
wire n_16310;
wire n_2446;
wire n_6582;
wire n_4116;
wire n_7724;
wire n_5360;
wire n_10501;
wire n_7269;
wire n_15160;
wire n_16058;
wire n_12003;
wire n_7047;
wire n_2671;
wire n_12292;
wire n_16348;
wire n_2702;
wire n_16113;
wire n_10908;
wire n_9176;
wire n_6937;
wire n_4363;
wire n_16365;
wire n_12405;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_214;
wire n_9728;
wire n_11809;
wire n_4103;
wire n_10777;
wire n_2529;
wire n_8101;
wire n_2374;
wire n_13712;
wire n_15549;
wire n_5439;
wire n_8687;
wire n_6115;
wire n_1225;
wire n_3154;
wire n_9866;
wire n_137;
wire n_14685;
wire n_8721;
wire n_1366;
wire n_8749;
wire n_12780;
wire n_13349;
wire n_9465;
wire n_13277;
wire n_3938;
wire n_11975;
wire n_8937;
wire n_2278;
wire n_6272;
wire n_12087;
wire n_13233;
wire n_13808;
wire n_7067;
wire n_16331;
wire n_14478;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_12662;
wire n_10965;
wire n_4416;
wire n_7879;
wire n_8730;
wire n_11441;
wire n_12416;
wire n_14895;
wire n_15555;
wire n_9702;
wire n_16323;
wire n_10998;
wire n_13503;
wire n_6607;
wire n_12854;
wire n_4439;
wire n_520;
wire n_870;
wire n_4985;
wire n_13056;
wire n_9000;
wire n_12936;
wire n_3382;
wire n_13300;
wire n_16461;
wire n_7117;
wire n_11743;
wire n_3930;
wire n_3808;
wire n_12765;
wire n_9610;
wire n_5471;
wire n_2248;
wire n_13087;
wire n_813;
wire n_4660;
wire n_8503;
wire n_10082;
wire n_10870;
wire n_12796;
wire n_11914;
wire n_15364;
wire n_3081;
wire n_6446;
wire n_10756;
wire n_5497;
wire n_9139;
wire n_13287;
wire n_5519;
wire n_6071;
wire n_995;
wire n_2579;
wire n_12028;
wire n_8315;
wire n_16531;
wire n_11175;
wire n_15563;
wire n_1961;
wire n_10411;
wire n_1535;
wire n_6849;
wire n_2960;
wire n_3270;
wire n_871;
wire n_6807;
wire n_15236;
wire n_2844;
wire n_11753;
wire n_8197;
wire n_13726;
wire n_17153;
wire n_11790;
wire n_402;
wire n_1979;
wire n_12294;
wire n_6616;
wire n_6719;
wire n_9407;
wire n_14621;
wire n_15883;
wire n_10423;
wire n_829;
wire n_4814;
wire n_8801;
wire n_8019;
wire n_12190;
wire n_14396;
wire n_339;
wire n_15134;
wire n_6178;
wire n_11249;
wire n_8707;
wire n_6677;
wire n_11791;
wire n_2221;
wire n_12786;
wire n_7875;
wire n_15983;
wire n_5502;
wire n_8962;
wire n_13665;
wire n_8931;
wire n_14177;
wire n_8248;
wire n_1283;
wire n_14533;
wire n_7550;
wire n_8554;
wire n_2317;
wire n_2838;
wire n_13242;
wire n_1736;
wire n_11879;
wire n_13900;
wire n_15269;
wire n_10782;
wire n_13837;
wire n_2200;
wire n_7302;
wire n_2781;
wire n_6191;
wire n_12386;
wire n_13121;
wire n_13679;
wire n_13680;
wire n_9357;
wire n_2442;
wire n_9477;
wire n_11911;
wire n_16274;
wire n_13734;
wire n_14591;
wire n_15756;
wire n_7238;
wire n_6862;
wire n_8501;
wire n_3657;
wire n_5706;
wire n_11842;
wire n_12746;
wire n_14023;
wire n_2634;
wire n_13047;
wire n_11304;
wire n_11320;
wire n_2746;
wire n_15728;
wire n_7292;
wire n_242;
wire n_645;
wire n_13146;
wire n_7804;
wire n_10251;
wire n_15780;
wire n_12128;
wire n_11776;
wire n_14544;
wire n_11471;
wire n_14904;
wire n_5098;
wire n_16658;
wire n_15253;
wire n_13475;
wire n_721;
wire n_1084;
wire n_6000;
wire n_6774;
wire n_9289;
wire n_11794;
wire n_6443;
wire n_16478;
wire n_9828;
wire n_1276;
wire n_8263;
wire n_5145;
wire n_6072;
wire n_13236;
wire n_2878;
wire n_15656;
wire n_7248;
wire n_10737;
wire n_3830;
wire n_10475;
wire n_3252;
wire n_6647;
wire n_11198;
wire n_8040;
wire n_13336;
wire n_5466;
wire n_14465;
wire n_1528;
wire n_6941;
wire n_9797;
wire n_7239;
wire n_15015;
wire n_16523;
wire n_6552;
wire n_7826;
wire n_10665;
wire n_9981;
wire n_3315;
wire n_6094;
wire n_12761;
wire n_14482;
wire n_3523;
wire n_12113;
wire n_8102;
wire n_3999;
wire n_14440;
wire n_10541;
wire n_13393;
wire n_14765;
wire n_9793;
wire n_16380;
wire n_518;
wire n_11419;
wire n_14214;
wire n_13202;
wire n_8196;
wire n_11171;
wire n_7112;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_8822;
wire n_12017;
wire n_3474;
wire n_5738;
wire n_14483;
wire n_9514;
wire n_2458;
wire n_7971;
wire n_12139;
wire n_8885;
wire n_11564;
wire n_5592;
wire n_11078;
wire n_5620;
wire n_12802;
wire n_3150;
wire n_5491;
wire n_1542;
wire n_4831;
wire n_10633;
wire n_12592;
wire n_4782;
wire n_9825;
wire n_1539;
wire n_2859;
wire n_10573;
wire n_5216;
wire n_3412;
wire n_11218;
wire n_16983;
wire n_1851;
wire n_2162;
wire n_5953;
wire n_15799;
wire n_1415;
wire n_8474;
wire n_15315;
wire n_16623;
wire n_1034;
wire n_1652;
wire n_5703;
wire n_10258;
wire n_6886;
wire n_17029;
wire n_7078;
wire n_16439;
wire n_16765;
wire n_1636;
wire n_4597;
wire n_12791;
wire n_9501;
wire n_12352;
wire n_13811;
wire n_12296;
wire n_11459;
wire n_9043;
wire n_8152;
wire n_12491;
wire n_17166;
wire n_11998;
wire n_16279;
wire n_8269;
wire n_4546;
wire n_11775;
wire n_5187;
wire n_7006;
wire n_4031;
wire n_5119;
wire n_11288;
wire n_1254;
wire n_4147;
wire n_16066;
wire n_1703;
wire n_12454;
wire n_10042;
wire n_12162;
wire n_10570;
wire n_13151;
wire n_3073;
wire n_6531;
wire n_9481;
wire n_3571;
wire n_11768;
wire n_238;
wire n_4576;
wire n_7577;
wire n_12992;
wire n_7354;
wire n_6098;
wire n_5995;
wire n_17121;
wire n_3297;
wire n_11456;
wire n_14706;
wire n_11708;
wire n_15407;
wire n_14330;
wire n_12960;
wire n_8144;
wire n_5148;
wire n_3003;
wire n_11662;
wire n_13617;
wire n_6726;
wire n_16013;
wire n_6983;
wire n_7513;
wire n_10098;
wire n_4340;
wire n_3136;
wire n_15320;
wire n_2867;
wire n_9766;
wire n_5330;
wire n_9351;
wire n_13935;
wire n_7812;
wire n_13930;
wire n_6935;
wire n_1560;
wire n_2899;
wire n_6984;
wire n_6778;
wire n_10106;
wire n_8058;
wire n_12046;
wire n_11877;
wire n_16338;
wire n_8909;
wire n_16811;
wire n_6897;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_16747;
wire n_5202;
wire n_12074;
wire n_15819;
wire n_14380;
wire n_3817;
wire n_6345;
wire n_9242;
wire n_10754;
wire n_6386;
wire n_2722;
wire n_3728;
wire n_12749;
wire n_14630;
wire n_612;
wire n_333;
wire n_15303;
wire n_6596;
wire n_5107;
wire n_7165;
wire n_512;
wire n_15598;
wire n_9777;
wire n_15302;
wire n_4680;
wire n_5067;
wire n_11932;
wire n_11821;
wire n_12485;
wire n_14464;
wire n_15188;
wire n_15183;
wire n_9522;
wire n_15904;
wire n_15113;
wire n_14560;
wire n_6830;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_9748;
wire n_16737;
wire n_5987;
wire n_2512;
wire n_1790;
wire n_12488;
wire n_14028;
wire n_12252;
wire n_10851;
wire n_9005;
wire n_12090;
wire n_11395;
wire n_2788;
wire n_10387;
wire n_9666;
wire n_6291;
wire n_6642;
wire n_10615;
wire n_1443;
wire n_6510;
wire n_5264;
wire n_14081;
wire n_14281;
wire n_2595;
wire n_10790;
wire n_1465;
wire n_3084;
wire n_10028;
wire n_15842;
wire n_705;
wire n_10555;
wire n_12896;
wire n_7667;
wire n_6781;
wire n_4593;
wire n_11532;
wire n_8024;
wire n_7123;
wire n_14670;
wire n_4562;
wire n_17145;
wire n_3860;
wire n_10222;
wire n_16299;
wire n_2909;
wire n_461;
wire n_3554;
wire n_12868;
wire n_15233;
wire n_6509;
wire n_10671;
wire n_2717;
wire n_6376;
wire n_1391;
wire n_8107;
wire n_16610;
wire n_9605;
wire n_2981;
wire n_10498;
wire n_225;
wire n_13959;
wire n_15747;
wire n_9947;
wire n_1006;
wire n_16033;
wire n_546;
wire n_9930;
wire n_14921;
wire n_14755;
wire n_13292;
wire n_4995;
wire n_15250;
wire n_1159;
wire n_5873;
wire n_6514;
wire n_4498;
wire n_10420;
wire n_772;
wire n_6741;
wire n_10083;
wire n_1245;
wire n_10520;
wire n_14839;
wire n_6434;
wire n_9662;
wire n_5741;
wire n_16592;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_9768;
wire n_1675;
wire n_2466;
wire n_12583;
wire n_676;
wire n_15934;
wire n_3758;
wire n_7631;
wire n_6593;
wire n_7827;
wire n_8748;
wire n_14420;
wire n_8452;
wire n_6690;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_10255;
wire n_8742;
wire n_3777;
wire n_8393;
wire n_9835;
wire n_11117;
wire n_11494;
wire n_1872;
wire n_9656;
wire n_1585;
wire n_11643;
wire n_14613;
wire n_3767;
wire n_12462;
wire n_12618;
wire n_14090;
wire n_14604;
wire n_6056;
wire n_5926;
wire n_5866;
wire n_9475;
wire n_212;
wire n_3692;
wire n_16226;
wire n_1351;
wire n_3234;
wire n_14347;
wire n_2216;
wire n_11475;
wire n_8122;
wire n_11004;
wire n_9724;
wire n_2426;
wire n_652;
wire n_6947;
wire n_8403;
wire n_8912;
wire n_16329;
wire n_10612;
wire n_4850;
wire n_15613;
wire n_15676;
wire n_10007;
wire n_9154;
wire n_12127;
wire n_13651;
wire n_16614;
wire n_1260;
wire n_3716;
wire n_15773;
wire n_11223;
wire n_11570;
wire n_7157;
wire n_15945;
wire n_16667;
wire n_2926;
wire n_10937;
wire n_4937;
wire n_798;
wire n_8740;
wire n_10493;
wire n_13631;
wire n_5574;
wire n_13264;
wire n_15012;
wire n_13678;
wire n_8310;
wire n_3391;
wire n_5877;
wire n_14406;
wire n_912;
wire n_10104;
wire n_6375;
wire n_460;
wire n_11212;
wire n_10552;
wire n_7781;
wire n_13294;
wire n_16820;
wire n_4786;
wire n_6042;
wire n_14746;
wire n_8238;
wire n_5203;
wire n_16443;
wire n_7908;
wire n_10295;
wire n_8296;
wire n_16408;
wire n_16359;
wire n_10954;
wire n_7091;
wire n_9833;
wire n_9788;
wire n_4354;
wire n_9589;
wire n_4235;
wire n_6429;
wire n_3159;
wire n_6315;
wire n_16133;
wire n_17072;
wire n_7855;
wire n_15314;
wire n_15560;
wire n_14590;
wire n_8850;
wire n_9861;
wire n_15526;
wire n_2855;
wire n_794;
wire n_2848;
wire n_16534;
wire n_7886;
wire n_14740;
wire n_7675;
wire n_16328;
wire n_11122;
wire n_6775;
wire n_8943;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_8993;
wire n_11159;
wire n_12329;
wire n_9205;
wire n_15450;
wire n_11631;
wire n_9946;
wire n_9418;
wire n_288;
wire n_10376;
wire n_1292;
wire n_7774;
wire n_8634;
wire n_12611;
wire n_11715;
wire n_13625;
wire n_8831;
wire n_6970;
wire n_13034;
wire n_1026;
wire n_9979;
wire n_12205;
wire n_13122;
wire n_6948;
wire n_3460;
wire n_14324;
wire n_16476;
wire n_14956;
wire n_13210;
wire n_1610;
wire n_5155;
wire n_8676;
wire n_14337;
wire n_15119;
wire n_2202;
wire n_11889;
wire n_16746;
wire n_14509;
wire n_306;
wire n_2952;
wire n_3530;
wire n_6133;
wire n_6920;
wire n_2693;
wire n_7409;
wire n_10087;
wire n_5408;
wire n_10341;
wire n_11278;
wire n_12606;
wire n_14692;
wire n_8758;
wire n_11671;
wire n_5812;
wire n_15008;
wire n_9973;
wire n_5540;
wire n_11782;
wire n_7381;
wire n_5804;
wire n_9007;
wire n_8544;
wire n_3240;
wire n_7999;
wire n_16882;
wire n_5066;
wire n_14253;
wire n_931;
wire n_16520;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_7087;
wire n_967;
wire n_9020;
wire n_10027;
wire n_14212;
wire n_5130;
wire n_9260;
wire n_4175;
wire n_10154;
wire n_6241;
wire n_13597;
wire n_9619;
wire n_14392;
wire n_13510;
wire n_1079;
wire n_5200;
wire n_9235;
wire n_14973;
wire n_15822;
wire n_3393;
wire n_10161;
wire n_13003;
wire n_8652;
wire n_16708;
wire n_15203;
wire n_9112;
wire n_12365;
wire n_2836;
wire n_12423;
wire n_7873;
wire n_12843;
wire n_2864;
wire n_4456;
wire n_11372;
wire n_16401;
wire n_15219;
wire n_1717;
wire n_9691;
wire n_5992;
wire n_8646;
wire n_15782;
wire n_13573;
wire n_2172;
wire n_2601;
wire n_12518;
wire n_12861;
wire n_7754;
wire n_17083;
wire n_1880;
wire n_2365;
wire n_9133;
wire n_5684;
wire n_1399;
wire n_13708;
wire n_7228;
wire n_5981;
wire n_14987;
wire n_7784;
wire n_9752;
wire n_1855;
wire n_16965;
wire n_6632;
wire n_2333;
wire n_8999;
wire n_3629;
wire n_4948;
wire n_15041;
wire n_10902;
wire n_5413;
wire n_15477;
wire n_1903;
wire n_2147;
wire n_7713;
wire n_6623;
wire n_9395;
wire n_4020;
wire n_5111;
wire n_5150;
wire n_1226;
wire n_2224;
wire n_6933;
wire n_1970;
wire n_15770;
wire n_10294;
wire n_3724;
wire n_16578;
wire n_9353;
wire n_11155;
wire n_3287;
wire n_11714;
wire n_12293;
wire n_2167;
wire n_13947;
wire n_16433;
wire n_2293;
wire n_3046;
wire n_15908;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_11590;
wire n_3257;
wire n_8031;
wire n_9804;
wire n_12450;
wire n_5737;
wire n_9125;
wire n_8015;
wire n_8412;
wire n_425;
wire n_3730;
wire n_16640;
wire n_8439;
wire n_8575;
wire n_5615;
wire n_3979;
wire n_6908;
wire n_13648;
wire n_17157;
wire n_5097;
wire n_10323;
wire n_2695;
wire n_7084;
wire n_11976;
wire n_13274;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_6537;
wire n_976;
wire n_17025;
wire n_4003;
wire n_1832;
wire n_767;
wire n_8499;
wire n_10969;
wire n_9397;
wire n_13015;
wire n_13472;
wire n_13322;
wire n_13870;
wire n_6390;
wire n_7640;
wire n_12000;
wire n_16278;
wire n_2302;
wire n_6799;
wire n_8772;
wire n_10806;
wire n_9767;
wire n_12903;
wire n_3014;
wire n_7912;
wire n_2294;
wire n_6278;
wire n_11430;
wire n_2274;
wire n_7195;
wire n_12309;
wire n_15072;
wire n_5640;
wire n_3342;
wire n_13401;
wire n_2895;
wire n_6101;
wire n_7298;
wire n_8557;
wire n_13891;
wire n_16007;
wire n_3796;
wire n_9384;
wire n_16488;
wire n_3884;
wire n_4492;
wire n_15284;
wire n_13850;
wire n_15894;
wire n_16411;
wire n_3625;
wire n_13835;
wire n_5550;
wire n_397;
wire n_3375;
wire n_15224;
wire n_2768;
wire n_351;
wire n_10666;
wire n_12895;
wire n_155;
wire n_3760;
wire n_5661;
wire n_16420;
wire n_7641;
wire n_15029;
wire n_4975;
wire n_11638;
wire n_3515;
wire n_16654;
wire n_2363;
wire n_12687;
wire n_12023;
wire n_14460;
wire n_5306;
wire n_5905;
wire n_13908;
wire n_8815;
wire n_7949;
wire n_6112;
wire n_11659;
wire n_16287;
wire n_2728;
wire n_9906;
wire n_15942;
wire n_2025;
wire n_8679;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_11948;
wire n_15640;
wire n_4022;
wire n_7115;
wire n_17123;
wire n_1020;
wire n_16216;
wire n_11843;
wire n_9310;
wire n_15382;
wire n_16196;
wire n_10659;
wire n_16976;
wire n_11689;
wire n_7764;
wire n_16853;
wire n_8446;
wire n_9163;
wire n_172;
wire n_11535;
wire n_2495;
wire n_12022;
wire n_17021;
wire n_1058;
wire n_12624;
wire n_4336;
wire n_11808;
wire n_8789;
wire n_8128;
wire n_7520;
wire n_5314;
wire n_9322;
wire n_12719;
wire n_7616;
wire n_14493;
wire n_10793;
wire n_14868;
wire n_14491;
wire n_8359;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_6412;
wire n_1279;
wire n_15495;
wire n_6271;
wire n_11108;
wire n_9377;
wire n_7235;
wire n_2511;
wire n_564;
wire n_6572;
wire n_9224;
wire n_10837;
wire n_10211;
wire n_3981;
wire n_16958;
wire n_14381;
wire n_17065;
wire n_12664;
wire n_13020;
wire n_11577;
wire n_15045;
wire n_16577;
wire n_7271;
wire n_16802;
wire n_9055;
wire n_15686;
wire n_13749;
wire n_13311;
wire n_2681;
wire n_7222;
wire n_8678;
wire n_9971;
wire n_1689;
wire n_8605;
wire n_2535;
wire n_12981;
wire n_13945;
wire n_1255;
wire n_3031;
wire n_345;
wire n_10976;
wire n_9624;
wire n_14766;
wire n_6930;
wire n_10045;
wire n_15026;
wire n_14172;
wire n_16501;
wire n_2335;
wire n_10289;
wire n_16761;
wire n_5482;
wire n_9145;
wire n_12716;
wire n_10232;
wire n_13079;
wire n_11098;
wire n_15177;
wire n_3215;
wire n_15130;
wire n_8443;
wire n_8525;
wire n_12166;
wire n_12507;
wire n_1401;
wire n_3138;
wire n_8312;
wire n_10819;
wire n_16035;
wire n_776;
wire n_15968;
wire n_2860;
wire n_8901;
wire n_2041;
wire n_13786;
wire n_1933;
wire n_13645;
wire n_6584;
wire n_4494;
wire n_9887;
wire n_12044;
wire n_6387;
wire n_466;
wire n_9373;
wire n_4201;
wire n_346;
wire n_16384;
wire n_15359;
wire n_14374;
wire n_6470;
wire n_7206;
wire n_16019;
wire n_8869;
wire n_552;
wire n_11279;
wire n_11729;
wire n_14012;
wire n_9770;
wire n_11514;
wire n_5287;
wire n_8272;
wire n_4719;
wire n_15440;
wire n_5651;
wire n_15587;
wire n_264;
wire n_15401;
wire n_3577;
wire n_6625;
wire n_14569;
wire n_4074;
wire n_7383;
wire n_12430;
wire n_3994;
wire n_4636;
wire n_11606;
wire n_4983;
wire n_3185;
wire n_10306;
wire n_12902;
wire n_14664;
wire n_12257;
wire n_1217;
wire n_11727;
wire n_13299;
wire n_10103;
wire n_17014;
wire n_11337;
wire n_327;
wire n_2662;
wire n_4386;
wire n_6341;
wire n_6374;
wire n_3917;
wire n_12839;
wire n_1231;
wire n_10183;
wire n_13693;
wire n_5623;
wire n_16255;
wire n_16963;
wire n_11778;
wire n_12925;
wire n_11658;
wire n_10710;
wire n_8870;
wire n_9753;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_10931;
wire n_9468;
wire n_11433;
wire n_8178;
wire n_5524;
wire n_7854;
wire n_9517;
wire n_15821;
wire n_16179;
wire n_926;
wire n_9544;
wire n_2296;
wire n_5735;
wire n_7959;
wire n_14338;
wire n_14728;
wire n_16502;
wire n_15009;
wire n_13434;
wire n_6363;
wire n_8234;
wire n_6588;
wire n_11369;
wire n_2178;
wire n_14865;
wire n_15642;
wire n_4243;
wire n_2765;
wire n_7897;
wire n_12759;
wire n_11720;
wire n_14418;
wire n_186;
wire n_15197;
wire n_4225;
wire n_6811;
wire n_6687;
wire n_4658;
wire n_13500;
wire n_14815;
wire n_7135;
wire n_6037;
wire n_4186;
wire n_1501;
wire n_8488;
wire n_11840;
wire n_2241;
wire n_6865;
wire n_11284;
wire n_12553;
wire n_7211;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_9774;
wire n_2531;
wire n_16194;
wire n_12016;
wire n_11987;
wire n_12496;
wire n_7132;
wire n_1570;
wire n_11052;
wire n_9586;
wire n_13655;
wire n_10670;
wire n_7533;
wire n_10150;
wire n_16042;
wire n_3377;
wire n_6722;
wire n_9780;
wire n_1518;
wire n_13476;
wire n_11177;
wire n_6420;
wire n_14900;
wire n_14803;
wire n_16638;
wire n_10004;
wire n_4907;
wire n_11169;
wire n_3961;
wire n_5153;
wire n_7766;
wire n_855;
wire n_8862;
wire n_13229;
wire n_17037;
wire n_2059;
wire n_14092;
wire n_8184;
wire n_13950;
wire n_5787;
wire n_4713;
wire n_6911;
wire n_11221;
wire n_14219;
wire n_13344;
wire n_16573;
wire n_10353;
wire n_10151;
wire n_16111;
wire n_1287;
wire n_11095;
wire n_10187;
wire n_1611;
wire n_10171;
wire n_16353;
wire n_11211;
wire n_7129;
wire n_12138;
wire n_7080;
wire n_3374;
wire n_4870;
wire n_6981;
wire n_7776;
wire n_4818;
wire n_8001;
wire n_10406;
wire n_8695;
wire n_12230;
wire n_12521;
wire n_11236;
wire n_11931;
wire n_7436;
wire n_8767;
wire n_11036;
wire n_12562;
wire n_8571;
wire n_7020;
wire n_11600;
wire n_15517;
wire n_5935;
wire n_14117;
wire n_8064;
wire n_15925;
wire n_14588;
wire n_6696;
wire n_13721;
wire n_4916;
wire n_8472;
wire n_13302;
wire n_5967;
wire n_15334;
wire n_15295;
wire n_6095;
wire n_4323;
wire n_5934;
wire n_529;
wire n_1899;
wire n_6045;
wire n_5376;
wire n_12217;
wire n_13535;
wire n_16605;
wire n_17142;
wire n_14261;
wire n_17136;
wire n_15581;
wire n_3508;
wire n_17171;
wire n_6300;
wire n_17026;
wire n_13704;
wire n_6653;
wire n_6372;
wire n_13969;
wire n_4129;
wire n_7120;
wire n_11114;
wire n_16745;
wire n_16648;
wire n_10479;
wire n_7978;
wire n_10033;
wire n_5488;
wire n_11336;
wire n_1105;
wire n_6900;
wire n_10034;
wire n_5727;
wire n_9099;
wire n_15344;
wire n_15137;
wire n_3599;
wire n_6660;
wire n_8787;
wire n_11009;
wire n_9543;
wire n_8131;
wire n_5988;
wire n_16248;
wire n_6424;
wire n_10696;
wire n_14633;
wire n_16264;
wire n_11480;
wire n_5646;
wire n_14538;
wire n_16209;
wire n_7448;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_7694;
wire n_8771;
wire n_9245;
wire n_6787;
wire n_15142;
wire n_5832;
wire n_15418;
wire n_13269;
wire n_6254;
wire n_7460;
wire n_3401;
wire n_983;
wire n_7142;
wire n_10360;
wire n_6423;
wire n_16230;
wire n_16866;
wire n_6526;
wire n_699;
wire n_3542;
wire n_16794;
wire n_301;
wire n_3263;
wire n_5891;
wire n_8150;
wire n_14891;
wire n_2523;
wire n_1945;
wire n_11423;
wire n_9168;
wire n_16136;
wire n_12691;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_5328;
wire n_3819;
wire n_9074;
wire n_12159;
wire n_16378;
wire n_3222;
wire n_325;
wire n_1740;
wire n_5016;
wire n_4616;
wire n_6011;
wire n_11665;
wire n_12259;
wire n_12975;
wire n_9367;
wire n_9330;
wire n_11556;
wire n_7465;
wire n_11685;
wire n_13402;
wire n_14231;
wire n_15662;
wire n_5470;
wire n_11801;
wire n_12117;
wire n_10230;
wire n_16923;
wire n_8917;
wire n_12587;
wire n_15995;
wire n_1092;
wire n_11573;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_6176;
wire n_16330;
wire n_1963;
wire n_9300;
wire n_16011;
wire n_14489;
wire n_13619;
wire n_14663;
wire n_3868;
wire n_11589;
wire n_11667;
wire n_14395;
wire n_729;
wire n_8230;
wire n_10414;
wire n_6222;
wire n_13110;
wire n_2218;
wire n_12422;
wire n_8352;
wire n_1122;
wire n_7760;
wire n_1408;
wire n_2593;
wire n_15042;
wire n_1693;
wire n_9918;
wire n_12977;
wire n_13060;
wire n_390;
wire n_6969;
wire n_2741;
wire n_15651;
wire n_2184;
wire n_2714;
wire n_9496;
wire n_13177;
wire n_15214;
wire n_8914;
wire n_10953;
wire n_14082;
wire n_8821;
wire n_16430;
wire n_11446;
wire n_13853;
wire n_8465;
wire n_15285;
wire n_6587;
wire n_6688;
wire n_17064;
wire n_8360;
wire n_6505;
wire n_13586;
wire n_15163;
wire n_9837;
wire n_12772;
wire n_15979;
wire n_5362;
wire n_8209;
wire n_15421;
wire n_388;
wire n_8986;
wire n_14701;
wire n_2754;
wire n_4580;
wire n_15867;
wire n_6762;
wire n_16795;
wire n_16632;
wire n_1218;
wire n_15191;
wire n_3611;
wire n_11633;
wire n_5147;
wire n_15697;
wire n_4826;
wire n_3959;
wire n_11011;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_7629;
wire n_12145;
wire n_10787;
wire n_6987;
wire n_877;
wire n_3995;
wire n_7567;
wire n_8743;
wire n_11342;
wire n_8963;
wire n_9191;
wire n_3908;
wire n_11812;
wire n_6453;
wire n_9114;
wire n_6308;
wire n_11142;
wire n_13074;
wire n_1055;
wire n_10896;
wire n_8396;
wire n_1395;
wire n_3892;
wire n_13773;
wire n_15582;
wire n_1346;
wire n_8514;
wire n_12196;
wire n_16177;
wire n_16617;
wire n_13482;
wire n_8550;
wire n_1089;
wire n_7449;
wire n_11959;
wire n_8151;
wire n_16774;
wire n_13927;
wire n_17009;
wire n_14688;
wire n_1502;
wire n_16242;
wire n_16862;
wire n_3501;
wire n_15579;
wire n_12889;
wire n_1478;
wire n_15793;
wire n_13096;
wire n_16857;
wire n_2555;
wire n_3216;
wire n_3568;
wire n_12493;
wire n_9913;
wire n_2708;
wire n_6187;
wire n_735;
wire n_15436;
wire n_11626;
wire n_6597;
wire n_13810;
wire n_11178;
wire n_12440;
wire n_4844;
wire n_9329;
wire n_6220;
wire n_13684;
wire n_14452;
wire n_12608;
wire n_15439;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_10598;
wire n_845;
wire n_13008;
wire n_13800;
wire n_7479;
wire n_7882;
wire n_16818;
wire n_13607;
wire n_1649;
wire n_2470;
wire n_11750;
wire n_13742;
wire n_7517;
wire n_1297;
wire n_16002;
wire n_9627;
wire n_3551;
wire n_417;
wire n_13412;
wire n_1708;
wire n_11283;
wire n_10271;
wire n_11338;
wire n_5037;
wire n_11295;
wire n_15668;
wire n_7305;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_8070;
wire n_15342;
wire n_14896;
wire n_4525;
wire n_8866;
wire n_10402;
wire n_6149;
wire n_11191;
wire n_15595;
wire n_10064;
wire n_3364;
wire n_11661;
wire n_13329;
wire n_10137;
wire n_2643;
wire n_755;
wire n_9585;
wire n_14863;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_7878;
wire n_9376;
wire n_4369;
wire n_12515;
wire n_15232;
wire n_16135;
wire n_17151;
wire n_3826;
wire n_5648;
wire n_278;
wire n_2266;
wire n_11644;
wire n_12249;
wire n_15742;
wire n_6439;
wire n_11354;
wire n_4324;
wire n_842;
wire n_15298;
wire n_148;
wire n_13537;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_8797;
wire n_14247;
wire n_14462;
wire n_6547;
wire n_13075;
wire n_11126;
wire n_9524;
wire n_7177;
wire n_7902;
wire n_11408;
wire n_16574;
wire n_12623;
wire n_742;
wire n_5160;
wire n_12971;
wire n_1719;
wire n_2742;
wire n_13051;
wire n_769;
wire n_3671;
wire n_12674;
wire n_15193;
wire n_15206;
wire n_2366;
wire n_9606;
wire n_5762;
wire n_1753;
wire n_15768;
wire n_14419;
wire n_10800;
wire n_5484;
wire n_1372;
wire n_476;
wire n_12026;
wire n_13038;
wire n_14514;
wire n_13812;
wire n_14733;
wire n_10019;
wire n_16391;
wire n_10762;
wire n_14135;
wire n_1895;
wire n_7353;
wire n_4104;
wire n_11935;
wire n_8054;
wire n_982;
wire n_3791;
wire n_915;
wire n_10047;
wire n_6478;
wire n_16221;
wire n_16457;
wire n_11037;
wire n_2008;
wire n_454;
wire n_298;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_13977;
wire n_16980;
wire n_3199;
wire n_8841;
wire n_11396;
wire n_9084;
wire n_2127;
wire n_14681;
wire n_7050;
wire n_3151;
wire n_7590;
wire n_14453;
wire n_6906;
wire n_403;
wire n_3016;
wire n_2460;
wire n_6739;
wire n_15657;
wire n_15720;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_10995;
wire n_3956;
wire n_4898;
wire n_17104;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_14869;
wire n_606;
wire n_4528;
wire n_2772;
wire n_14036;
wire n_17101;
wire n_1700;
wire n_15490;
wire n_10597;
wire n_659;
wire n_1332;
wire n_10561;
wire n_14994;
wire n_7818;
wire n_509;
wire n_12345;
wire n_16789;
wire n_7645;
wire n_15655;
wire n_5385;
wire n_7482;
wire n_1747;
wire n_3990;
wire n_13841;
wire n_14312;
wire n_16555;
wire n_11726;
wire n_12346;
wire n_5622;
wire n_14522;
wire n_14110;
wire n_15647;
wire n_10523;
wire n_10377;
wire n_8618;
wire n_1171;
wire n_10243;
wire n_5635;
wire n_16568;
wire n_4069;
wire n_8538;
wire n_3582;
wire n_8590;
wire n_13883;
wire n_14945;
wire n_7907;
wire n_9204;
wire n_16492;
wire n_8970;
wire n_17117;
wire n_4280;
wire n_1867;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_15558;
wire n_2576;
wire n_3459;
wire n_8791;
wire n_15013;
wire n_14739;
wire n_13724;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_521;
wire n_5910;
wire n_17030;
wire n_2140;
wire n_10165;
wire n_14776;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_9616;
wire n_9708;
wire n_1400;
wire n_10153;
wire n_7862;
wire n_9130;
wire n_9988;
wire n_3735;
wire n_8703;
wire n_12265;
wire n_7565;
wire n_7410;
wire n_6422;
wire n_1527;
wire n_1513;
wire n_3656;
wire n_12147;
wire n_7721;
wire n_4524;
wire n_9209;
wire n_16987;
wire n_15374;
wire n_8061;
wire n_2831;
wire n_10775;
wire n_10173;
wire n_10585;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_12075;
wire n_8754;
wire n_15755;
wire n_14996;
wire n_8864;
wire n_5941;
wire n_15478;
wire n_10985;
wire n_4891;
wire n_11300;
wire n_14294;
wire n_8837;
wire n_12108;
wire n_10999;
wire n_13425;
wire n_2629;
wire n_3369;
wire n_13791;
wire n_8915;
wire n_15251;
wire n_1257;
wire n_10587;
wire n_1954;
wire n_8784;
wire n_11219;
wire n_6604;
wire n_3964;
wire n_6611;
wire n_5364;
wire n_3302;
wire n_15833;
wire n_15415;
wire n_8036;
wire n_11857;
wire n_5597;
wire n_11735;
wire n_2486;
wire n_11986;
wire n_12102;
wire n_1897;
wire n_8768;
wire n_8086;
wire n_9014;
wire n_9086;
wire n_8072;
wire n_15205;
wire n_6999;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_6019;
wire n_7539;
wire n_16447;
wire n_16485;
wire n_14611;
wire n_9010;
wire n_11637;
wire n_13925;
wire n_16100;
wire n_16760;
wire n_6440;
wire n_4977;
wire n_8774;
wire n_14417;
wire n_16878;
wire n_16508;
wire n_2492;
wire n_6976;
wire n_11072;
wire n_7234;
wire n_12183;
wire n_7608;
wire n_2939;
wire n_3425;
wire n_13432;
wire n_15860;
wire n_4876;
wire n_16022;
wire n_15084;
wire n_16193;
wire n_15217;
wire n_241;
wire n_5021;
wire n_1449;
wire n_12519;
wire n_16344;
wire n_2900;
wire n_12955;
wire n_797;
wire n_9044;
wire n_2912;
wire n_13538;
wire n_14176;
wire n_5936;
wire n_14650;
wire n_8307;
wire n_595;
wire n_14939;
wire n_1405;
wire n_3813;
wire n_13774;
wire n_14789;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_15290;
wire n_6784;
wire n_9694;
wire n_1757;
wire n_16237;
wire n_11421;
wire n_13323;
wire n_10718;
wire n_13214;
wire n_10951;
wire n_10412;
wire n_8470;
wire n_1950;
wire n_2264;
wire n_15216;
wire n_805;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_7830;
wire n_8050;
wire n_3124;
wire n_16427;
wire n_3811;
wire n_16642;
wire n_14980;
wire n_295;
wire n_10310;
wire n_4200;
wire n_190;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_10655;
wire n_9633;
wire n_6165;
wire n_10133;
wire n_12793;
wire n_3463;
wire n_11989;
wire n_15399;
wire n_10942;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_6114;
wire n_1856;
wire n_463;
wire n_1524;
wire n_13192;
wire n_15189;
wire n_2928;
wire n_13433;
wire n_5505;
wire n_13392;
wire n_12865;
wire n_1118;
wire n_14662;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_469;
wire n_9261;
wire n_11331;
wire n_12285;
wire n_726;
wire n_5504;
wire n_878;
wire n_7348;
wire n_9345;
wire n_14894;
wire n_11953;
wire n_4118;
wire n_6829;
wire n_11820;
wire n_12478;
wire n_3857;
wire n_3110;
wire n_9375;
wire n_4239;
wire n_9472;
wire n_9764;
wire n_10509;
wire n_16294;
wire n_8010;
wire n_3157;
wire n_13059;
wire n_12522;
wire n_13451;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_9448;
wire n_6464;
wire n_8802;
wire n_8950;
wire n_5129;
wire n_13199;
wire n_806;
wire n_1350;
wire n_7320;
wire n_4704;
wire n_2720;
wire n_649;
wire n_1561;
wire n_8603;
wire n_9487;
wire n_15654;
wire n_15691;
wire n_10639;
wire n_13588;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_15531;
wire n_11358;
wire n_12413;
wire n_6838;
wire n_13191;
wire n_16102;
wire n_2700;
wire n_6368;
wire n_14133;
wire n_10690;
wire n_16699;
wire n_12369;
wire n_12681;
wire n_1616;
wire n_11118;
wire n_2416;
wire n_7935;
wire n_8143;
wire n_11844;
wire n_2064;
wire n_3640;
wire n_9271;
wire n_17086;
wire n_5663;
wire n_15332;
wire n_12084;
wire n_5161;
wire n_14132;
wire n_7933;
wire n_12152;
wire n_12726;
wire n_12784;
wire n_16704;
wire n_1557;
wire n_7155;
wire n_6640;
wire n_9851;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_15281;
wire n_5626;
wire n_349;
wire n_4706;
wire n_3879;
wire n_2022;
wire n_4343;
wire n_6850;
wire n_12520;
wire n_12705;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_7743;
wire n_11861;
wire n_13899;
wire n_14443;
wire n_4990;
wire n_2986;
wire n_8584;
wire n_14934;
wire n_11370;
wire n_13017;
wire n_949;
wire n_2454;
wire n_9101;
wire n_15186;
wire n_16266;
wire n_6550;
wire n_6656;
wire n_8153;
wire n_6972;
wire n_3591;
wire n_8574;
wire n_198;
wire n_12832;
wire n_15461;
wire n_2760;
wire n_4919;
wire n_15145;
wire n_13422;
wire n_15448;
wire n_15834;
wire n_1208;
wire n_7043;
wire n_7986;
wire n_3317;
wire n_8049;
wire n_9927;
wire n_12207;
wire n_13666;
wire n_12782;
wire n_7266;
wire n_13042;
wire n_15875;
wire n_10621;
wire n_11884;
wire n_15664;
wire n_5653;
wire n_14860;
wire n_4835;
wire n_1151;
wire n_554;
wire n_4420;
wire n_15299;
wire n_7996;
wire n_14513;
wire n_12970;
wire n_15507;
wire n_10789;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_354;
wire n_5266;
wire n_10496;
wire n_4559;
wire n_4742;
wire n_12384;
wire n_12605;
wire n_5038;
wire n_14724;
wire n_15011;
wire n_15683;
wire n_3566;
wire n_10319;
wire n_15679;
wire n_15871;
wire n_5800;
wire n_16936;
wire n_14021;
wire n_8509;
wire n_14830;
wire n_12408;
wire n_1133;
wire n_883;
wire n_16223;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_9850;
wire n_4162;
wire n_5766;
wire n_10499;
wire n_14223;
wire n_17024;
wire n_11717;
wire n_5293;
wire n_10224;
wire n_13234;
wire n_15155;
wire n_779;
wire n_4790;
wire n_594;
wire n_7035;
wire n_10970;
wire n_4173;
wire n_8354;
wire n_12651;
wire n_5309;
wire n_15501;
wire n_15059;
wire n_6047;
wire n_9432;
wire n_16856;
wire n_3573;
wire n_2943;
wire n_12160;
wire n_13829;
wire n_16943;
wire n_11464;
wire n_3319;
wire n_16263;
wire n_11243;
wire n_2247;
wire n_2230;
wire n_9824;
wire n_422;
wire n_14582;
wire n_1269;
wire n_8277;
wire n_7442;
wire n_4727;
wire n_10827;
wire n_14880;
wire n_16448;
wire n_1547;
wire n_1438;
wire n_6568;
wire n_16472;
wire n_3654;
wire n_11473;
wire n_14508;
wire n_5627;
wire n_1047;
wire n_3783;
wire n_10055;
wire n_12638;
wire n_12698;
wire n_17071;
wire n_4008;
wire n_11654;
wire n_13878;
wire n_10783;
wire n_15208;
wire n_2158;
wire n_14562;
wire n_8583;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_7153;
wire n_8681;
wire n_6258;
wire n_1288;
wire n_8644;
wire n_10148;
wire n_7939;
wire n_9884;
wire n_7715;
wire n_11534;
wire n_2173;
wire n_3982;
wire n_10465;
wire n_14040;
wire n_14361;
wire n_11749;
wire n_7350;
wire n_3647;
wire n_16383;
wire n_15972;
wire n_7314;
wire n_6026;
wire n_10610;
wire n_8609;
wire n_13955;
wire n_1143;
wire n_9144;
wire n_3973;
wire n_15453;
wire n_16484;
wire n_8052;
wire n_12481;
wire n_4799;
wire n_8733;
wire n_9758;
wire n_12078;
wire n_8082;
wire n_5882;
wire n_6700;
wire n_12815;
wire n_16395;
wire n_7136;
wire n_4534;
wire n_12129;
wire n_5636;
wire n_4960;
wire n_9931;
wire n_7699;
wire n_9693;
wire n_12502;
wire n_11546;
wire n_10830;
wire n_1153;
wire n_9273;
wire n_271;
wire n_15530;
wire n_16126;
wire n_465;
wire n_9196;
wire n_1103;
wire n_5707;
wire n_15474;
wire n_5594;
wire n_16530;
wire n_9029;
wire n_10086;
wire n_15614;
wire n_3738;
wire n_894;
wire n_5697;
wire n_1380;
wire n_13763;
wire n_6255;
wire n_562;
wire n_2020;
wire n_7580;
wire n_5606;
wire n_15737;
wire n_11785;
wire n_6727;
wire n_2310;
wire n_510;
wire n_5911;
wire n_12697;
wire n_7340;
wire n_8080;
wire n_256;
wire n_13437;
wire n_16766;
wire n_3600;
wire n_10279;
wire n_7303;
wire n_1023;
wire n_10932;
wire n_11440;
wire n_9967;
wire n_15849;
wire n_12908;
wire n_16078;
wire n_8819;
wire n_914;
wire n_7870;
wire n_689;
wire n_6139;
wire n_7568;
wire n_7399;
wire n_5382;
wire n_4327;
wire n_14799;
wire n_7387;
wire n_3190;
wire n_8487;
wire n_13293;
wire n_3027;
wire n_6454;
wire n_11545;
wire n_4011;
wire n_11697;
wire n_16183;
wire n_3695;
wire n_13555;
wire n_3800;
wire n_13487;
wire n_15591;
wire n_13239;
wire n_3462;
wire n_17018;
wire n_10487;
wire n_14579;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_14853;
wire n_9881;
wire n_16390;
wire n_2820;
wire n_497;
wire n_3733;
wire n_1165;
wire n_11645;
wire n_3967;
wire n_12512;
wire n_11263;
wire n_12199;
wire n_15043;
wire n_6333;
wire n_11937;
wire n_7004;
wire n_15538;
wire n_16900;
wire n_12584;
wire n_455;
wire n_16596;
wire n_13854;
wire n_588;
wire n_13361;
wire n_638;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_10910;
wire n_16881;
wire n_5058;
wire n_8382;
wire n_1417;
wire n_9733;
wire n_3096;
wire n_16139;
wire n_8517;
wire n_7207;
wire n_8827;
wire n_13558;
wire n_9075;
wire n_11324;
wire n_13954;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_11763;
wire n_13803;
wire n_7167;
wire n_2234;
wire n_1341;
wire n_5849;
wire n_16754;
wire n_3233;
wire n_11853;
wire n_2431;
wire n_3322;
wire n_12988;
wire n_14537;
wire n_8906;
wire n_1603;
wire n_5841;
wire n_10109;
wire n_7146;
wire n_14542;
wire n_7030;
wire n_10857;
wire n_17089;
wire n_4478;
wire n_8203;
wire n_413;
wire n_2935;
wire n_9442;
wire n_15096;
wire n_4246;
wire n_715;
wire n_7618;
wire n_14625;
wire n_1066;
wire n_2863;
wire n_13244;
wire n_2331;
wire n_4632;
wire n_13305;
wire n_15741;
wire n_12284;
wire n_11364;
wire n_16372;
wire n_11941;
wire n_16513;
wire n_685;
wire n_9630;
wire n_4061;
wire n_11359;
wire n_16864;
wire n_12031;
wire n_14203;
wire n_9898;
wire n_15926;
wire n_11323;
wire n_11504;
wire n_15146;
wire n_11704;
wire n_2920;
wire n_11587;
wire n_1712;
wire n_11620;
wire n_13697;
wire n_3344;
wire n_8340;
wire n_4754;
wire n_12652;
wire n_16543;
wire n_9582;
wire n_1534;
wire n_10865;
wire n_8268;
wire n_17067;
wire n_15291;
wire n_16029;
wire n_8171;
wire n_16812;
wire n_1290;
wire n_16932;
wire n_4375;
wire n_12850;
wire n_15244;
wire n_617;
wire n_9877;
wire n_14578;
wire n_10179;
wire n_12969;
wire n_2396;
wire n_10925;
wire n_12607;
wire n_12379;
wire n_3368;
wire n_13743;
wire n_9986;
wire n_1559;
wire n_13951;
wire n_14222;
wire n_16528;
wire n_13695;
wire n_8008;
wire n_7633;
wire n_10246;
wire n_9636;
wire n_3117;
wire n_4684;
wire n_10439;
wire n_743;
wire n_13376;
wire n_16888;
wire n_14377;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_7159;
wire n_8553;
wire n_2592;
wire n_8824;
wire n_11902;
wire n_3490;
wire n_7280;
wire n_8369;
wire n_962;
wire n_5043;
wire n_12701;
wire n_14008;
wire n_7339;
wire n_7597;
wire n_16581;
wire n_8884;
wire n_12898;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_9225;
wire n_4183;
wire n_7768;
wire n_918;
wire n_1968;
wire n_11282;
wire n_5645;
wire n_639;
wire n_5020;
wire n_673;
wire n_6455;
wire n_13639;
wire n_16947;
wire n_2842;
wire n_7615;
wire n_2196;
wire n_16015;
wire n_12475;
wire n_16208;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_10182;
wire n_14795;
wire n_8271;
wire n_9091;
wire n_3720;
wire n_6183;
wire n_13772;
wire n_14643;
wire n_12027;
wire n_8392;
wire n_15835;
wire n_8309;
wire n_14986;
wire n_6107;
wire n_15685;
wire n_12218;
wire n_10795;
wire n_13602;
wire n_6476;
wire n_5232;
wire n_16197;
wire n_10046;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_9412;
wire n_11834;
wire n_8874;
wire n_8228;
wire n_16750;
wire n_12174;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_11405;
wire n_11028;
wire n_3037;
wire n_11663;
wire n_16989;
wire n_1336;
wire n_16692;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_15645;
wire n_5339;
wire n_8483;
wire n_6003;
wire n_5443;
wire n_8133;
wire n_7612;
wire n_15646;
wire n_12385;
wire n_17003;
wire n_1166;
wire n_2007;
wire n_14407;
wire n_3363;
wire n_15321;
wire n_15882;
wire n_17080;
wire n_6636;
wire n_9525;
wire n_1158;
wire n_11071;
wire n_12289;
wire n_11625;
wire n_1803;
wire n_15626;
wire n_872;
wire n_11187;
wire n_12041;
wire n_12565;
wire n_3522;
wire n_12882;
wire n_13736;
wire n_15075;
wire n_13254;
wire n_12819;
wire n_8172;
wire n_17098;
wire n_14810;
wire n_4455;
wire n_13341;
wire n_3241;
wire n_3899;
wire n_6554;
wire n_16322;
wire n_9575;
wire n_5631;
wire n_3481;
wire n_280;
wire n_7401;
wire n_10456;
wire n_10413;
wire n_11566;
wire n_12164;
wire n_11271;
wire n_12433;
wire n_6994;
wire n_15383;
wire n_11649;
wire n_12224;
wire n_13061;
wire n_5101;
wire n_9738;
wire n_10735;
wire n_6020;
wire n_2236;
wire n_13328;
wire n_14908;
wire n_9252;
wire n_16259;
wire n_12550;
wire n_6185;
wire n_8344;
wire n_12800;
wire n_14568;
wire n_15452;
wire n_16012;
wire n_692;
wire n_14259;
wire n_7594;
wire n_7711;
wire n_7321;
wire n_4457;
wire n_17173;
wire n_12561;
wire n_223;
wire n_2150;
wire n_8738;
wire n_8936;
wire n_10822;
wire n_9739;
wire n_6785;
wire n_14871;
wire n_1816;
wire n_2803;
wire n_9727;
wire n_2887;
wire n_10508;
wire n_2648;
wire n_4735;
wire n_6870;
wire n_17051;
wire n_3305;
wire n_6643;
wire n_13281;
wire n_15323;
wire n_7574;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_8226;
wire n_15272;
wire n_14874;
wire n_6695;
wire n_7529;
wire n_3354;
wire n_6501;
wire n_5608;
wire n_17022;
wire n_2204;
wire n_11308;
wire n_11739;
wire n_11593;
wire n_9148;
wire n_10858;
wire n_1481;
wire n_2040;
wire n_6466;
wire n_10736;
wire n_11828;
wire n_9958;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_6467;
wire n_9323;
wire n_2231;
wire n_14138;
wire n_4212;
wire n_622;
wire n_4584;
wire n_7522;
wire n_7188;
wire n_9779;
wire n_15074;
wire n_8088;
wire n_5702;
wire n_14244;
wire n_9545;
wire n_16706;
wire n_8930;
wire n_9155;
wire n_12563;
wire n_8662;
wire n_13114;
wire n_11291;
wire n_16286;
wire n_3574;
wire n_11425;
wire n_13566;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_9046;
wire n_9430;
wire n_16470;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_11890;
wire n_4110;
wire n_9625;
wire n_13621;
wire n_5806;
wire n_8783;
wire n_12398;
wire n_16639;
wire n_13624;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_8663;
wire n_14015;
wire n_10928;
wire n_16956;
wire n_5277;
wire n_792;
wire n_1262;
wire n_6507;
wire n_10842;
wire n_1942;
wire n_12941;
wire n_9447;
wire n_13407;
wire n_15865;
wire n_6618;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_13404;
wire n_16195;
wire n_8364;
wire n_1579;
wire n_9485;
wire n_6213;
wire n_4949;
wire n_2181;
wire n_17023;
wire n_15857;
wire n_2014;
wire n_16306;
wire n_14818;
wire n_2974;
wire n_9129;
wire n_8490;
wire n_229;
wire n_8981;
wire n_923;
wire n_12461;
wire n_1124;
wire n_11832;
wire n_7872;
wire n_1326;
wire n_3969;
wire n_6873;
wire n_7958;
wire n_2282;
wire n_4605;
wire n_8118;
wire n_981;
wire n_3873;
wire n_4649;
wire n_5747;
wire n_8671;
wire n_7101;
wire n_12095;
wire n_15714;
wire n_14191;
wire n_8785;
wire n_11294;
wire n_11470;
wire n_11744;
wire n_1204;
wire n_10210;
wire n_13994;
wire n_14841;
wire n_15817;
wire n_7843;
wire n_12998;
wire n_994;
wire n_2428;
wire n_9047;
wire n_13219;
wire n_15952;
wire n_10057;
wire n_1360;
wire n_6063;
wire n_13737;
wire n_2858;
wire n_16245;
wire n_12630;
wire n_11641;
wire n_15141;
wire n_15464;
wire n_15181;
wire n_3076;
wire n_7578;
wire n_12789;
wire n_12679;
wire n_14146;
wire n_3410;
wire n_13372;
wire n_5415;
wire n_14084;
wire n_856;
wire n_7261;
wire n_8982;
wire n_10739;
wire n_4999;
wire n_4592;
wire n_16656;
wire n_1564;
wire n_12327;
wire n_6993;
wire n_9745;
wire n_14288;
wire n_12038;
wire n_508;
wire n_13932;
wire n_10533;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_16585;
wire n_13978;
wire n_11875;
wire n_8100;
wire n_1858;
wire n_10878;
wire n_353;
wire n_1678;
wire n_16351;
wire n_2589;
wire n_15600;
wire n_4086;
wire n_10988;
wire n_1482;
wire n_8522;
wire n_13563;
wire n_1361;
wire n_15733;
wire n_13141;
wire n_12338;
wire n_10993;
wire n_13249;
wire n_8381;
wire n_9320;
wire n_16777;
wire n_8835;
wire n_6767;
wire n_11014;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_12030;
wire n_14553;
wire n_15258;
wire n_5687;
wire n_1411;
wire n_1359;
wire n_6558;
wire n_13517;
wire n_6755;
wire n_9108;
wire n_9457;
wire n_15001;
wire n_17169;
wire n_16602;
wire n_9907;
wire n_10959;
wire n_6153;
wire n_15545;
wire n_11310;
wire n_3536;
wire n_1721;
wire n_16670;
wire n_11062;
wire n_7263;
wire n_3782;
wire n_10940;
wire n_12067;
wire n_16786;
wire n_13783;
wire n_16354;
wire n_1317;
wire n_12675;
wire n_16821;
wire n_6608;
wire n_11400;
wire n_11040;
wire n_15797;
wire n_6202;
wire n_15353;
wire n_6780;
wire n_7688;
wire n_13968;
wire n_16073;
wire n_12870;
wire n_14038;
wire n_3594;
wire n_12291;
wire n_5383;
wire n_2385;
wire n_6635;
wire n_7245;
wire n_7925;
wire n_16899;
wire n_7310;
wire n_9567;
wire n_294;
wire n_6359;
wire n_11773;
wire n_14385;
wire n_5690;
wire n_10583;
wire n_14027;
wire n_11332;
wire n_1980;
wire n_5740;
wire n_7093;
wire n_4177;
wire n_2501;
wire n_7585;
wire n_8356;
wire n_1385;
wire n_16146;
wire n_1998;
wire n_5029;
wire n_13279;
wire n_13731;
wire n_12013;
wire n_13007;
wire n_16781;
wire n_2675;
wire n_16317;
wire n_2604;
wire n_15818;
wire n_3521;
wire n_9852;
wire n_10881;
wire n_16037;
wire n_12395;
wire n_3855;
wire n_16268;
wire n_7418;
wire n_16192;
wire n_6353;
wire n_14049;
wire n_13160;
wire n_2985;
wire n_11943;
wire n_5218;
wire n_10544;
wire n_12933;
wire n_16271;
wire n_2630;
wire n_6577;
wire n_7772;
wire n_13895;
wire n_14403;
wire n_13213;
wire n_8736;
wire n_15899;
wire n_2028;
wire n_919;
wire n_3114;
wire n_10491;
wire n_12131;
wire n_17069;
wire n_2092;
wire n_13507;
wire n_6082;
wire n_15625;
wire n_11144;
wire n_13385;
wire n_10926;
wire n_3622;
wire n_2817;
wire n_2773;
wire n_11841;
wire n_8918;
wire n_11766;
wire n_2402;
wire n_1458;
wire n_12766;
wire n_16465;
wire n_679;
wire n_10839;
wire n_16342;
wire n_220;
wire n_3047;
wire n_10603;
wire n_3163;
wire n_5361;
wire n_7312;
wire n_9022;
wire n_13790;
wire n_16854;
wire n_7514;
wire n_15985;
wire n_1550;
wire n_16634;
wire n_12399;
wire n_1358;
wire n_8616;
wire n_1200;
wire n_6105;
wire n_387;
wire n_12762;
wire n_10400;
wire n_11518;
wire n_826;
wire n_5512;
wire n_13567;
wire n_14346;
wire n_7738;
wire n_2808;
wire n_14787;
wire n_2344;
wire n_16928;
wire n_8838;
wire n_8908;
wire n_13687;
wire n_3520;
wire n_11960;
wire n_2392;
wire n_7609;
wire n_13580;
wire n_9161;
wire n_3272;
wire n_12241;
wire n_10792;
wire n_3122;
wire n_5898;
wire n_15336;
wire n_7113;
wire n_11274;
wire n_8607;
wire n_6548;
wire n_13779;
wire n_15473;
wire n_16124;
wire n_607;
wire n_8213;
wire n_14487;
wire n_13722;
wire n_13225;
wire n_14615;
wire n_15699;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_6657;
wire n_10994;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_13514;
wire n_1268;
wire n_13806;
wire n_2676;
wire n_9903;
wire n_9831;
wire n_14595;
wire n_15460;
wire n_10032;
wire n_8436;
wire n_7282;
wire n_17168;
wire n_372;
wire n_13261;
wire n_8551;
wire n_14638;
wire n_16552;
wire n_13039;
wire n_15524;
wire n_2770;
wire n_4550;
wire n_14717;
wire n_9238;
wire n_12137;
wire n_14167;
wire n_4347;
wire n_11624;
wire n_10580;
wire n_7921;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_10512;
wire n_9248;
wire n_12495;
wire n_5514;
wire n_11917;
wire n_5611;
wire n_2375;
wire n_3278;
wire n_12790;
wire n_6380;
wire n_4167;
wire n_5579;
wire n_3608;
wire n_4895;
wire n_14924;
wire n_15288;
wire n_9867;
wire n_12106;
wire n_1282;
wire n_11130;
wire n_6163;
wire n_7170;
wire n_4726;
wire n_11053;
wire n_10005;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_1755;
wire n_11872;
wire n_12434;
wire n_15881;
wire n_6674;
wire n_5188;
wire n_13669;
wire n_5049;
wire n_12710;
wire n_2212;
wire n_16403;
wire n_7489;
wire n_9056;
wire n_6331;
wire n_5308;
wire n_9106;
wire n_311;
wire n_4434;
wire n_13303;
wire n_5068;
wire n_12881;
wire n_7863;
wire n_15906;
wire n_6493;
wire n_7363;
wire n_14496;
wire n_7281;
wire n_5739;
wire n_2569;
wire n_10596;
wire n_12920;
wire n_4019;
wire n_4199;
wire n_14260;
wire n_7968;
wire n_16451;
wire n_11220;
wire n_16398;
wire n_10061;
wire n_16790;
wire n_10507;
wire n_6023;
wire n_7820;
wire n_8437;
wire n_269;
wire n_816;
wire n_12086;
wire n_7833;
wire n_1322;
wire n_11887;
wire n_3829;
wire n_14189;
wire n_12281;
wire n_15437;
wire n_12991;
wire n_4510;
wire n_14552;
wire n_7750;
wire n_5057;
wire n_446;
wire n_9071;
wire n_6196;
wire n_12995;
wire n_16247;
wire n_5425;
wire n_5273;
wire n_10136;
wire n_5839;
wire n_2469;
wire n_7588;
wire n_1125;
wire n_10967;
wire n_11551;
wire n_2358;
wire n_1710;
wire n_14339;
wire n_13368;
wire n_10369;
wire n_3546;
wire n_14971;
wire n_2355;
wire n_1390;
wire n_10708;
wire n_11703;
wire n_10025;
wire n_7697;
wire n_5887;
wire n_16996;
wire n_16053;
wire n_13948;
wire n_7808;
wire n_3068;
wire n_9519;
wire n_1629;
wire n_15960;
wire n_9027;
wire n_7603;
wire n_13598;
wire n_1094;
wire n_6321;
wire n_14180;
wire n_5683;
wire n_1510;
wire n_8704;
wire n_14341;
wire n_3002;
wire n_8984;
wire n_9786;
wire n_10194;
wire n_7192;
wire n_1099;
wire n_12807;
wire n_5248;
wire n_4899;
wire n_11153;
wire n_10833;
wire n_3146;
wire n_10685;
wire n_3038;
wire n_759;
wire n_10513;
wire n_16516;
wire n_567;
wire n_4156;
wire n_8613;
wire n_13611;
wire n_1727;
wire n_11030;
wire n_14704;
wire n_3693;
wire n_13178;
wire n_14293;
wire n_10223;
wire n_5880;
wire n_13495;
wire n_15417;
wire n_8012;
wire n_12012;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_8881;
wire n_5531;
wire n_16016;
wire n_16459;
wire n_9404;
wire n_831;
wire n_13777;
wire n_3681;
wire n_5666;
wire n_13301;
wire n_3970;
wire n_11368;
wire n_778;
wire n_2351;
wire n_1619;
wire n_12098;
wire n_7988;
wire n_12025;
wire n_550;
wire n_12669;
wire n_15468;
wire n_13205;
wire n_15617;
wire n_3188;
wire n_4448;
wire n_10410;
wire n_13049;
wire n_3218;
wire n_6824;
wire n_6954;
wire n_8763;
wire n_6450;
wire n_9370;
wire n_16917;
wire n_1152;
wire n_15553;
wire n_6995;
wire n_2447;
wire n_13009;
wire n_16175;
wire n_2101;
wire n_4193;
wire n_17114;
wire n_1236;
wire n_4579;
wire n_14885;
wire n_6347;
wire n_13748;
wire n_14878;
wire n_16438;
wire n_13338;
wire n_6496;
wire n_13747;
wire n_4776;
wire n_671;
wire n_8387;
wire n_9352;
wire n_14972;
wire n_17179;
wire n_11716;
wire n_14083;
wire n_8105;
wire n_10984;
wire n_13485;
wire n_10144;
wire n_16167;
wire n_12019;
wire n_2704;
wire n_1334;
wire n_6745;
wire n_7943;
wire n_3729;
wire n_6698;
wire n_16848;
wire n_4471;
wire n_6968;
wire n_13416;
wire n_11967;
wire n_7377;
wire n_12255;
wire n_8900;
wire n_4392;
wire n_3103;
wire n_488;
wire n_6064;
wire n_9681;
wire n_14439;
wire n_8353;
wire n_12503;
wire n_505;
wire n_17077;
wire n_9051;
wire n_2048;
wire n_16352;
wire n_7723;
wire n_498;
wire n_3028;
wire n_4691;
wire n_7904;
wire n_3148;
wire n_3775;
wire n_5682;
wire n_16687;
wire n_684;
wire n_5461;
wire n_9098;
wire n_12415;
wire n_8323;
wire n_3966;
wire n_4397;
wire n_13053;
wire n_13752;
wire n_7296;
wire n_10459;
wire n_12951;
wire n_14125;
wire n_6164;
wire n_11426;
wire n_8711;
wire n_13273;
wire n_15787;
wire n_3616;
wire n_11628;
wire n_4753;
wire n_12704;
wire n_9484;
wire n_4803;
wire n_8731;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_10155;
wire n_11367;
wire n_6292;
wire n_7759;
wire n_6743;
wire n_4165;
wire n_16020;
wire n_2056;
wire n_5754;
wire n_11418;
wire n_2852;
wire n_8597;
wire n_2515;
wire n_6330;
wire n_15289;
wire n_1600;
wire n_1144;
wire n_7178;
wire n_838;
wire n_11026;
wire n_15672;
wire n_1941;
wire n_7045;
wire n_11576;
wire n_175;
wire n_3637;
wire n_9853;
wire n_8534;
wire n_1017;
wire n_15046;
wire n_9210;
wire n_8655;
wire n_12884;
wire n_16165;
wire n_734;
wire n_16056;
wire n_13324;
wire n_4893;
wire n_10915;
wire n_13414;
wire n_13894;
wire n_2240;
wire n_16967;
wire n_10949;
wire n_12339;
wire n_7777;
wire n_16482;
wire n_8302;
wire n_14616;
wire n_4258;
wire n_5756;
wire n_14784;
wire n_14695;
wire n_14455;
wire n_310;
wire n_12911;
wire n_15301;
wire n_8496;
wire n_7693;
wire n_11150;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2432;
wire n_2085;
wire n_10156;
wire n_5033;
wire n_11123;
wire n_14414;
wire n_16527;
wire n_10248;
wire n_14941;
wire n_6015;
wire n_1686;
wire n_6408;
wire n_4232;
wire n_5075;
wire n_8078;
wire n_14449;
wire n_16273;
wire n_2097;
wire n_662;
wire n_11733;
wire n_3461;
wire n_15903;
wire n_10215;
wire n_17125;
wire n_10624;
wire n_12915;
wire n_7682;
wire n_7300;
wire n_939;
wire n_1410;
wire n_2297;
wire n_10152;
wire n_12888;
wire n_15811;
wire n_6861;
wire n_16844;
wire n_4203;
wire n_12105;
wire n_9756;
wire n_16132;
wire n_5789;
wire n_12034;
wire n_5400;
wire n_1325;
wire n_7558;
wire n_1223;
wire n_5347;
wire n_14744;
wire n_2957;
wire n_572;
wire n_11188;
wire n_9166;
wire n_8103;
wire n_8719;
wire n_1983;
wire n_10877;
wire n_15954;
wire n_7798;
wire n_9778;
wire n_8879;
wire n_13906;
wire n_4767;
wire n_16615;
wire n_15218;
wire n_8969;
wire n_9141;
wire n_4569;
wire n_11209;
wire n_948;
wire n_448;
wire n_6528;
wire n_14441;
wire n_13159;
wire n_9700;
wire n_10316;
wire n_8896;
wire n_3820;
wire n_5144;
wire n_11503;
wire n_6895;
wire n_3072;
wire n_10385;
wire n_14769;
wire n_15192;
wire n_15775;
wire n_14732;
wire n_8335;
wire n_2961;
wire n_16607;
wire n_13337;
wire n_5509;
wire n_4468;
wire n_15917;
wire n_1923;
wire n_3848;
wire n_15433;
wire n_7400;
wire n_14230;
wire n_11699;
wire n_13145;
wire n_16014;
wire n_3631;
wire n_7393;
wire n_6590;
wire n_8116;
wire n_12549;
wire n_6523;
wire n_11817;
wire n_5169;
wire n_4885;
wire n_14618;
wire n_7475;
wire n_1479;
wire n_11469;
wire n_9363;
wire n_11971;
wire n_4698;
wire n_14199;
wire n_1031;
wire n_16003;
wire n_3674;
wire n_1638;
wire n_853;
wire n_16842;
wire n_15497;
wire n_716;
wire n_1571;
wire n_14722;
wire n_5349;
wire n_14101;
wire n_16519;
wire n_6472;
wire n_3763;
wire n_9532;
wire n_10823;
wire n_12237;
wire n_933;
wire n_14001;
wire n_6389;
wire n_14586;
wire n_3499;
wire n_14623;
wire n_14635;
wire n_15586;
wire n_10680;
wire n_5534;
wire n_1821;
wire n_9307;
wire n_16462;
wire n_13922;
wire n_16711;
wire n_9876;
wire n_12220;
wire n_3947;
wire n_3910;
wire n_12564;
wire n_492;
wire n_10814;
wire n_12375;
wire n_13333;
wire n_252;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_8462;
wire n_9959;
wire n_3228;
wire n_8834;
wire n_9989;
wire n_10651;
wire n_14495;
wire n_8286;
wire n_8417;
wire n_2164;
wire n_1732;
wire n_13872;
wire n_12809;
wire n_2678;
wire n_8964;
wire n_10611;
wire n_1186;
wire n_6869;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_10549;
wire n_10370;
wire n_11621;
wire n_16590;
wire n_7672;
wire n_10770;
wire n_14171;
wire n_4556;
wire n_6137;
wire n_9467;
wire n_2205;
wire n_2183;
wire n_15635;
wire n_11558;
wire n_389;
wire n_12043;
wire n_1724;
wire n_3088;
wire n_12513;
wire n_14988;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_12337;
wire n_1126;
wire n_10393;
wire n_5079;
wire n_14975;
wire n_9406;
wire n_2761;
wire n_2357;
wire n_10089;
wire n_8247;
wire n_11417;
wire n_11113;
wire n_14182;
wire n_4520;
wire n_10543;
wire n_895;
wire n_13355;
wire n_15639;
wire n_8639;
wire n_12504;
wire n_15246;
wire n_1639;
wire n_11301;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_9160;
wire n_5751;
wire n_11051;
wire n_12489;
wire n_626;
wire n_10321;
wire n_12886;
wire n_13308;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_7712;
wire n_7681;
wire n_6885;
wire n_15173;
wire n_5039;
wire n_1818;
wire n_6580;
wire n_6613;
wire n_8566;
wire n_8727;
wire n_15492;
wire n_14791;
wire n_4265;
wire n_8482;
wire n_6404;
wire n_6120;
wire n_3557;
wire n_13923;
wire n_1598;
wire n_11018;
wire n_13905;
wire n_14884;
wire n_15956;
wire n_2269;
wire n_10259;
wire n_14927;
wire n_7491;
wire n_15194;
wire n_12836;
wire n_265;
wire n_1583;
wire n_14243;
wire n_13936;
wire n_15419;
wire n_10909;
wire n_10094;
wire n_8599;
wire n_4612;
wire n_14386;
wire n_5997;
wire n_10302;
wire n_11328;
wire n_15243;
wire n_8781;
wire n_5375;
wire n_5438;
wire n_9167;
wire n_11276;
wire n_15796;
wire n_7150;
wire n_7954;
wire n_7974;
wire n_1264;
wire n_6530;
wire n_6602;
wire n_15845;
wire n_7915;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_6135;
wire n_246;
wire n_12655;
wire n_10623;
wire n_8839;
wire n_11326;
wire n_13627;
wire n_14359;
wire n_14786;
wire n_1752;
wire n_2361;
wire n_3030;
wire n_4538;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_13882;
wire n_12779;
wire n_8365;
wire n_1102;
wire n_15973;
wire n_13144;
wire n_14085;
wire n_2239;
wire n_6942;
wire n_16466;
wire n_7860;
wire n_14108;
wire n_6892;
wire n_1296;
wire n_4730;
wire n_7357;
wire n_8489;
wire n_8112;
wire n_13364;
wire n_8859;
wire n_8060;
wire n_9290;
wire n_6782;
wire n_4421;
wire n_6230;
wire n_2464;
wire n_3697;
wire n_15319;
wire n_15427;
wire n_882;
wire n_13134;
wire n_2304;
wire n_8244;
wire n_13340;
wire n_2514;
wire n_6977;
wire n_7229;
wire n_16832;
wire n_12688;
wire n_11732;
wire n_7663;
wire n_10485;
wire n_8096;
wire n_11946;
wire n_7336;
wire n_5932;
wire n_11334;
wire n_289;
wire n_6598;
wire n_16850;
wire n_10105;
wire n_6795;
wire n_6121;
wire n_12321;
wire n_11855;
wire n_457;
wire n_1299;
wire n_3430;
wire n_5919;
wire n_2063;
wire n_8346;
wire n_3489;
wire n_5012;
wire n_6614;
wire n_6506;
wire n_11781;
wire n_13310;
wire n_14548;
wire n_14427;
wire n_14306;
wire n_15765;
wire n_11080;
wire n_2079;
wire n_9705;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_8367;
wire n_9113;
wire n_10761;
wire n_12104;
wire n_3484;
wire n_6001;
wire n_13445;
wire n_411;
wire n_14074;
wire n_4971;
wire n_9521;
wire n_9682;
wire n_2095;
wire n_14043;
wire n_14676;
wire n_7493;
wire n_9278;
wire n_5664;
wire n_2738;
wire n_15967;
wire n_16719;
wire n_6406;
wire n_5890;
wire n_14355;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_357;
wire n_3041;
wire n_412;
wire n_5823;
wire n_8898;
wire n_8658;
wire n_1421;
wire n_2423;
wire n_2208;
wire n_5944;
wire n_5422;
wire n_8905;
wire n_9222;
wire n_15174;
wire n_15939;
wire n_12643;
wire n_8237;
wire n_11445;
wire n_6299;
wire n_6989;
wire n_8145;
wire n_16836;
wire n_10592;
wire n_9813;
wire n_7424;
wire n_10216;
wire n_5246;
wire n_8562;
wire n_4376;
wire n_9863;
wire n_3832;
wire n_15348;
wire n_10616;
wire n_11350;
wire n_14527;
wire n_12799;
wire n_3525;
wire n_13833;
wire n_3712;
wire n_15022;
wire n_12202;
wire n_12694;
wire n_11057;
wire n_9394;
wire n_10170;
wire n_11182;
wire n_1069;
wire n_4305;
wire n_11140;
wire n_2037;
wire n_16213;
wire n_2953;
wire n_573;
wire n_2823;
wire n_11082;
wire n_15754;
wire n_7273;
wire n_9663;
wire n_7901;
wire n_3684;
wire n_14371;
wire n_15759;
wire n_5725;
wire n_10146;
wire n_5404;
wire n_15378;
wire n_16060;
wire n_913;
wire n_15287;
wire n_10175;
wire n_1681;
wire n_11949;
wire n_13576;
wire n_12055;
wire n_4834;
wire n_9994;
wire n_1507;
wire n_5332;
wire n_7149;
wire n_9723;
wire n_15095;
wire n_16791;
wire n_589;
wire n_2866;
wire n_7116;
wire n_3153;
wire n_1174;
wire n_16270;
wire n_2346;
wire n_4692;
wire n_15153;
wire n_1353;
wire n_11693;
wire n_12506;
wire n_8211;
wire n_3268;
wire n_2559;
wire n_8537;
wire n_15670;
wire n_15717;
wire n_8946;
wire n_16515;
wire n_5616;
wire n_16621;
wire n_1383;
wire n_17116;
wire n_603;
wire n_8055;
wire n_16763;
wire n_10848;
wire n_373;
wire n_4259;
wire n_5870;
wire n_7909;
wire n_12788;
wire n_12894;
wire n_2030;
wire n_6053;
wire n_11024;
wire n_850;
wire n_6233;
wire n_10918;
wire n_10450;
wire n_12333;
wire n_13502;
wire n_4299;
wire n_15254;
wire n_14879;
wire n_13131;
wire n_5625;
wire n_245;
wire n_13238;
wire n_14597;
wire n_319;
wire n_6758;
wire n_14801;
wire n_2407;
wire n_690;
wire n_5367;
wire n_9069;
wire n_525;
wire n_2243;
wire n_12866;
wire n_6629;
wire n_5288;
wire n_16122;
wire n_13247;
wire n_11158;
wire n_16720;
wire n_2694;
wire n_6356;
wire n_8332;
wire n_5601;
wire n_3742;
wire n_4965;
wire n_7601;
wire n_8998;
wire n_13391;
wire n_15561;
wire n_14190;
wire n_11046;
wire n_1837;
wire n_15529;
wire n_7033;
wire n_16092;
wire n_16009;
wire n_4178;
wire n_6010;
wire n_11390;
wire n_15296;
wire n_12551;
wire n_11224;
wire n_13970;
wire n_10536;
wire n_15604;
wire n_14696;
wire n_189;
wire n_8157;
wire n_2006;
wire n_9284;
wire n_4953;
wire n_10990;
wire n_8484;
wire n_4813;
wire n_3352;
wire n_12223;
wire n_12627;
wire n_12390;
wire n_16469;
wire n_15794;
wire n_2367;
wire n_7147;
wire n_7596;
wire n_9556;
wire n_12226;
wire n_14546;
wire n_5294;
wire n_11380;
wire n_8161;
wire n_5570;
wire n_11101;
wire n_6411;
wire n_11578;
wire n_9337;
wire n_2731;
wire n_3703;
wire n_5670;
wire n_5411;
wire n_16041;
wire n_1246;
wire n_13256;
wire n_11015;
wire n_11214;
wire n_9211;
wire n_12378;
wire n_5265;
wire n_5955;
wire n_7549;
wire n_10278;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_10482;
wire n_14174;
wire n_6032;
wire n_1196;
wire n_10996;
wire n_5733;
wire n_8692;
wire n_3435;
wire n_12794;
wire n_410;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_9243;
wire n_14046;
wire n_12436;
wire n_16341;
wire n_6918;
wire n_1298;
wire n_10733;
wire n_16244;
wire n_1745;
wire n_9773;
wire n_14158;
wire n_4674;
wire n_15127;
wire n_15724;
wire n_8812;
wire n_14218;
wire n_568;
wire n_11033;
wire n_8682;
wire n_13170;
wire n_4796;
wire n_8290;
wire n_1088;
wire n_13664;
wire n_7138;
wire n_766;
wire n_6401;
wire n_7279;
wire n_5184;
wire n_9928;
wire n_377;
wire n_7976;
wire n_10975;
wire n_2750;
wire n_11950;
wire n_16437;
wire n_16647;
wire n_8890;
wire n_17039;
wire n_10484;
wire n_2547;
wire n_12962;
wire n_8747;
wire n_7617;
wire n_12094;
wire n_279;
wire n_945;
wire n_4575;
wire n_9784;
wire n_10641;
wire n_11115;
wire n_12964;
wire n_3665;
wire n_3063;
wire n_8062;
wire n_14120;
wire n_3281;
wire n_16690;
wire n_7137;
wire n_3535;
wire n_5061;
wire n_14652;
wire n_16566;
wire n_2288;
wire n_14412;
wire n_3858;
wire n_14499;
wire n_4653;
wire n_7700;
wire n_11709;
wire n_15431;
wire n_15491;
wire n_8275;
wire n_7474;
wire n_4589;
wire n_7124;
wire n_5978;
wire n_14938;
wire n_6853;
wire n_10584;
wire n_16911;
wire n_16222;
wire n_14609;
wire n_8667;
wire n_3220;
wire n_4581;
wire n_9192;
wire n_10365;
wire n_14466;
wire n_6008;
wire n_500;
wire n_665;
wire n_10778;
wire n_4625;
wire n_11607;
wire n_11542;
wire n_7098;
wire n_6181;
wire n_14668;
wire n_2107;
wire n_16334;
wire n_5070;
wire n_4845;
wire n_13105;
wire n_4148;
wire n_9134;
wire n_12838;
wire n_13964;
wire n_16785;
wire n_3679;
wire n_738;
wire n_5575;
wire n_6654;
wire n_11491;
wire n_7661;
wire n_672;
wire n_16631;
wire n_4968;
wire n_8807;
wire n_7801;
wire n_17054;
wire n_9975;
wire n_13766;
wire n_9765;
wire n_11896;
wire n_13525;
wire n_6907;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_11371;
wire n_11939;
wire n_5316;
wire n_7876;
wire n_2735;
wire n_953;
wire n_14332;
wire n_4214;
wire n_13081;
wire n_10378;
wire n_143;
wire n_1888;
wire n_5290;
wire n_13057;
wire n_1224;
wire n_15067;
wire n_10324;
wire n_11563;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_557;
wire n_3419;
wire n_7323;
wire n_13861;
wire n_15223;
wire n_989;
wire n_10850;
wire n_5048;
wire n_11565;
wire n_2233;
wire n_13129;
wire n_13257;
wire n_15395;
wire n_5363;
wire n_14583;
wire n_11164;
wire n_12633;
wire n_5665;
wire n_6517;
wire n_11401;
wire n_16806;
wire n_11414;
wire n_795;
wire n_4892;
wire n_6339;
wire n_12514;
wire n_10330;
wire n_15136;
wire n_14659;
wire n_14408;
wire n_16034;
wire n_16389;
wire n_16892;
wire n_1936;
wire n_9564;
wire n_14267;
wire n_9127;
wire n_11199;
wire n_15540;
wire n_3890;
wire n_6170;
wire n_7247;
wire n_6394;
wire n_8048;
wire n_821;
wire n_770;
wire n_14370;
wire n_5607;
wire n_1514;
wire n_7929;
wire n_14516;
wire n_16456;
wire n_486;
wire n_2782;
wire n_14840;
wire n_569;
wire n_15692;
wire n_3929;
wire n_11319;
wire n_9306;
wire n_971;
wire n_4353;
wire n_2201;
wire n_8212;
wire n_4950;
wire n_10442;
wire n_1650;
wire n_7755;
wire n_14970;
wire n_13865;
wire n_9891;
wire n_6504;
wire n_13135;
wire n_10962;
wire n_10022;
wire n_13973;
wire n_4176;
wire n_9078;
wire n_7556;
wire n_222;
wire n_11415;
wire n_13553;
wire n_4124;
wire n_4431;
wire n_15005;
wire n_17156;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_10972;
wire n_7216;
wire n_6814;
wire n_13248;
wire n_16326;
wire n_4488;
wire n_10127;
wire n_17050;
wire n_5278;
wire n_15123;
wire n_14278;
wire n_2779;
wire n_3627;
wire n_10824;
wire n_3596;
wire n_5214;
wire n_11128;
wire n_9332;
wire n_12262;
wire n_3756;
wire n_12391;
wire n_8223;
wire n_8043;
wire n_16941;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_8159;
wire n_5845;
wire n_8868;
wire n_9889;
wire n_4608;
wire n_9294;
wire n_12731;
wire n_6691;
wire n_13623;
wire n_432;
wire n_293;
wire n_13775;
wire n_12235;
wire n_3948;
wire n_4839;
wire n_9174;
wire n_1074;
wire n_5969;
wire n_10375;
wire n_1765;
wire n_13464;
wire n_9132;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_11669;
wire n_4184;
wire n_15609;
wire n_206;
wire n_2332;
wire n_9547;
wire n_2391;
wire n_6343;
wire n_12406;
wire n_15213;
wire n_6005;
wire n_611;
wire n_1295;
wire n_2060;
wire n_4988;
wire n_3883;
wire n_1013;
wire n_6686;
wire n_4032;
wire n_12929;
wire n_16217;
wire n_2571;
wire n_136;
wire n_6437;
wire n_5736;
wire n_4929;
wire n_14067;
wire n_2874;
wire n_6029;
wire n_6536;
wire n_6684;
wire n_4117;
wire n_300;
wire n_6025;
wire n_12229;
wire n_15252;
wire n_3049;
wire n_8434;
wire n_16740;
wire n_14264;
wire n_3634;
wire n_15969;
wire n_12508;
wire n_5436;
wire n_7962;
wire n_2341;
wire n_1654;
wire n_6697;
wire n_11262;
wire n_16121;
wire n_12271;
wire n_3066;
wire n_11110;
wire n_13084;
wire n_2045;
wire n_12803;
wire n_14451;
wire n_14614;
wire n_10122;
wire n_6085;
wire n_10898;
wire n_3913;
wire n_14785;
wire n_9762;
wire n_11849;
wire n_5341;
wire n_8608;
wire n_2575;
wire n_13583;
wire n_3739;
wire n_1230;
wire n_16874;
wire n_5140;
wire n_376;
wire n_13470;
wire n_16481;
wire n_1597;
wire n_12245;
wire n_16218;
wire n_2942;
wire n_15430;
wire n_1771;
wire n_4541;
wire n_14394;
wire n_6062;
wire n_6715;
wire n_3271;
wire n_15872;
wire n_16110;
wire n_16902;
wire n_3164;
wire n_8656;
wire n_3861;
wire n_15414;
wire n_5096;
wire n_9183;
wire n_2043;
wire n_11287;
wire n_7905;
wire n_6771;
wire n_4171;
wire n_11247;
wire n_5847;
wire n_7204;
wire n_12376;
wire n_9461;
wire n_9117;
wire n_7022;
wire n_6383;
wire n_4815;
wire n_12773;
wire n_4665;
wire n_5639;
wire n_6877;
wire n_7308;
wire n_7476;
wire n_10116;
wire n_10590;
wire n_10991;
wire n_11945;
wire n_14743;
wire n_16985;
wire n_11769;
wire n_4884;
wire n_16185;
wire n_3580;
wire n_12720;
wire n_1437;
wire n_12736;
wire n_8249;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_9062;
wire n_209;
wire n_5240;
wire n_5718;
wire n_1461;
wire n_5503;
wire n_7208;
wire n_10265;
wire n_7718;
wire n_9915;
wire n_13006;
wire n_17163;
wire n_11277;
wire n_1876;
wire n_1830;
wire n_12459;
wire n_11075;
wire n_5001;
wire n_12708;
wire n_6567;
wire n_11919;
wire n_16063;
wire n_503;
wire n_12387;
wire n_13705;
wire n_5658;
wire n_1112;
wire n_700;
wire n_16934;
wire n_4174;
wire n_9001;
wire n_13599;
wire n_15211;
wire n_16910;
wire n_6868;
wire n_7290;
wire n_5131;
wire n_13077;
wire n_9081;
wire n_6813;
wire n_7756;
wire n_5546;
wire n_9156;
wire n_6294;
wire n_7795;
wire n_7822;
wire n_8717;
wire n_10159;
wire n_15643;
wire n_5174;
wire n_9024;
wire n_9198;
wire n_10178;
wire n_2145;
wire n_4801;
wire n_10571;
wire n_15516;
wire n_6079;
wire n_6260;
wire n_680;
wire n_4582;
wire n_14268;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_6520;
wire n_13892;
wire n_7623;
wire n_380;
wire n_14251;
wire n_17106;
wire n_15911;
wire n_12239;
wire n_15567;
wire n_14136;
wire n_12636;
wire n_14002;
wire n_16628;
wire n_3119;
wire n_6671;
wire n_11085;
wire n_9335;
wire n_4740;
wire n_16047;
wire n_1108;
wire n_10550;
wire n_16297;
wire n_9488;
wire n_16090;
wire n_1274;
wire n_7632;
wire n_4394;
wire n_257;
wire n_15850;
wire n_5544;
wire n_6444;
wire n_6637;
wire n_16112;
wire n_11510;
wire n_16843;
wire n_9725;
wire n_8842;
wire n_475;
wire n_16473;
wire n_17075;
wire n_6729;
wire n_5660;
wire n_6958;
wire n_8073;
wire n_10185;
wire n_12648;
wire n_17177;
wire n_9526;
wire n_4920;
wire n_3909;
wire n_10809;
wire n_13316;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_13140;
wire n_5541;
wire n_6314;
wire n_10660;
wire n_13162;
wire n_15308;
wire n_12501;
wire n_577;
wire n_5610;
wire n_407;
wire n_9962;
wire n_15848;
wire n_8576;
wire n_916;
wire n_2810;
wire n_12755;
wire n_15869;
wire n_6703;
wire n_1884;
wire n_14262;
wire n_1555;
wire n_10657;
wire n_10627;
wire n_8799;
wire n_762;
wire n_1253;
wire n_1468;
wire n_4378;
wire n_9667;
wire n_5166;
wire n_2683;
wire n_11256;
wire n_6065;
wire n_7265;
wire n_12441;
wire n_14018;
wire n_14805;
wire n_14935;
wire n_4180;
wire n_11516;
wire n_11520;
wire n_15376;
wire n_4459;
wire n_11461;
wire n_6878;
wire n_11137;
wire n_3624;
wire n_6725;
wire n_8181;
wire n_5808;
wire n_1182;
wire n_15309;
wire n_6527;
wire n_16733;
wire n_4594;
wire n_13604;
wire n_14877;
wire n_8447;
wire n_8045;
wire n_7289;
wire n_7538;
wire n_14029;
wire n_13157;
wire n_2748;
wire n_11536;
wire n_15790;
wire n_16521;
wire n_11544;
wire n_14488;
wire n_10897;
wire n_4642;
wire n_13952;
wire n_14234;
wire n_9716;
wire n_6913;
wire n_15502;
wire n_1376;
wire n_7473;
wire n_7242;
wire n_9253;
wire n_6533;
wire n_513;
wire n_11305;
wire n_14126;
wire n_15352;
wire n_179;
wire n_7164;
wire n_15890;
wire n_2925;
wire n_1435;
wire n_15164;
wire n_15804;
wire n_1750;
wire n_1506;
wire n_15959;
wire n_16468;
wire n_8022;
wire n_10617;
wire n_12011;
wire n_3544;
wire n_6845;
wire n_10451;
wire n_5300;
wire n_8227;
wire n_14438;
wire n_10768;
wire n_7853;
wire n_2072;
wire n_3852;
wire n_11268;
wire n_16429;
wire n_13707;
wire n_5233;
wire n_16611;
wire n_12742;
wire n_10309;
wire n_5381;
wire n_15569;
wire n_436;
wire n_9796;
wire n_5770;
wire n_7483;
wire n_13868;
wire n_8756;
wire n_5710;
wire n_10021;
wire n_324;
wire n_9953;
wire n_1491;
wire n_2628;
wire n_7389;
wire n_3219;
wire n_10053;
wire n_10315;
wire n_16125;
wire n_274;
wire n_1083;
wire n_5799;
wire n_5333;
wire n_10765;
wire n_6265;
wire n_4914;
wire n_12317;
wire n_8604;
wire n_12831;
wire n_8809;
wire n_16824;
wire n_13092;
wire n_8976;
wire n_11815;
wire n_13694;
wire n_3510;
wire n_10907;
wire n_7046;
wire n_13928;
wire n_15135;
wire n_7834;
wire n_10312;
wire n_11299;
wire n_16116;
wire n_4587;
wire n_16085;
wire n_1139;
wire n_3688;
wire n_11273;
wire n_8940;
wire n_15416;
wire n_16512;
wire n_5008;
wire n_1312;
wire n_9077;
wire n_12872;
wire n_16682;
wire n_15541;
wire n_13147;
wire n_15879;
wire n_12871;
wire n_3871;
wire n_13212;
wire n_16727;
wire n_12590;
wire n_14503;
wire n_892;
wire n_14325;
wire n_3757;
wire n_15644;
wire n_1567;
wire n_16453;
wire n_563;
wire n_11213;
wire n_13519;
wire n_2219;
wire n_8844;
wire n_14998;
wire n_6148;
wire n_8995;
wire n_2100;
wire n_8255;
wire n_3666;
wire n_5538;
wire n_16370;
wire n_990;
wire n_17011;
wire n_6357;
wire n_867;
wire n_12785;
wire n_8693;
wire n_8216;
wire n_3479;
wire n_14808;
wire n_16314;
wire n_944;
wire n_5499;
wire n_749;
wire n_13661;
wire n_9123;
wire n_2888;
wire n_3998;
wire n_16509;
wire n_16960;
wire n_4150;
wire n_1920;
wire n_7811;
wire n_12545;
wire n_6522;
wire n_8669;
wire n_4285;
wire n_7097;
wire n_12531;
wire n_7000;
wire n_2668;
wire n_10486;
wire n_11290;
wire n_16570;
wire n_2701;
wire n_2400;
wire n_15228;
wire n_10357;
wire n_650;
wire n_3741;
wire n_9922;
wire n_5582;
wire n_2567;
wire n_9177;
wire n_14348;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_7880;
wire n_14130;
wire n_712;
wire n_8769;
wire n_9463;
wire n_909;
wire n_12916;
wire n_6713;
wire n_8149;
wire n_1392;
wire n_13163;
wire n_10067;
wire n_12953;
wire n_15198;
wire n_17044;
wire n_10698;
wire n_2066;
wire n_16860;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_964;
wire n_13874;
wire n_13106;
wire n_7851;
wire n_2220;
wire n_13246;
wire n_7342;
wire n_7044;
wire n_16490;
wire n_7810;
wire n_10135;
wire n_13776;
wire n_6108;
wire n_12222;
wire n_10260;
wire n_7664;
wire n_12370;
wire n_6100;
wire n_14329;
wire n_6800;
wire n_7364;
wire n_6866;
wire n_7114;
wire n_6373;
wire n_16782;
wire n_4433;
wire n_11412;
wire n_2829;
wire n_16432;
wire n_7332;
wire n_14428;
wire n_14813;
wire n_8990;
wire n_5862;
wire n_471;
wire n_7477;
wire n_1914;
wire n_14617;
wire n_10268;
wire n_8208;
wire n_2253;
wire n_7468;
wire n_11550;
wire n_12692;
wire n_13640;
wire n_15965;
wire n_5886;
wire n_9451;
wire n_7714;
wire n_7899;
wire n_8710;
wire n_12976;
wire n_6415;
wire n_8479;
wire n_14660;
wire n_6783;
wire n_2130;
wire n_4861;
wire n_13984;
wire n_12397;
wire n_16787;
wire n_2021;
wire n_8512;
wire n_14524;
wire n_13093;
wire n_9843;
wire n_16990;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_9710;
wire n_2507;
wire n_12634;
wire n_16535;
wire n_13288;
wire n_16104;
wire n_1633;
wire n_9087;
wire n_4621;
wire n_15896;
wire n_14287;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_7845;
wire n_11619;
wire n_13086;
wire n_347;
wire n_2434;
wire n_14052;
wire n_183;
wire n_14216;
wire n_1234;
wire n_3936;
wire n_479;
wire n_5564;
wire n_15044;
wire n_16913;
wire n_2261;
wire n_12613;
wire n_16779;
wire n_9956;
wire n_3082;
wire n_9079;
wire n_5162;
wire n_14925;
wire n_15641;
wire n_5442;
wire n_2473;
wire n_12946;
wire n_5802;
wire n_16298;
wire n_9782;
wire n_10049;
wire n_4784;
wire n_14206;
wire n_13012;
wire n_16830;
wire n_13606;
wire n_2438;
wire n_12901;
wire n_13449;
wire n_10589;
wire n_3210;
wire n_6340;
wire n_13099;
wire n_14475;
wire n_9950;
wire n_11019;
wire n_14620;
wire n_7858;
wire n_11580;
wire n_17109;
wire n_3867;
wire n_3397;
wire n_13699;
wire n_12683;
wire n_6103;
wire n_15829;
wire n_14837;
wire n_1646;
wire n_6513;
wire n_6392;
wire n_11642;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_13389;
wire n_14978;
wire n_9197;
wire n_1237;
wire n_6720;
wire n_12286;
wire n_11076;
wire n_11752;
wire n_5883;
wire n_9140;
wire n_14134;
wire n_13995;
wire n_10785;
wire n_14726;
wire n_13439;
wire n_8401;
wire n_1095;
wire n_3078;
wire n_6078;
wire n_14122;
wire n_3971;
wire n_12146;
wire n_370;
wire n_7680;
wire n_14415;
wire n_5630;
wire n_6666;
wire n_286;
wire n_9364;
wire n_9452;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_9362;
wire n_9398;
wire n_13675;
wire n_13483;
wire n_1531;
wire n_2113;
wire n_14977;
wire n_6815;
wire n_14321;
wire n_15275;
wire n_9203;
wire n_1387;
wire n_6207;
wire n_6381;
wire n_3711;
wire n_9712;
wire n_14903;
wire n_15201;
wire n_9536;
wire n_12054;
wire n_8450;
wire n_16981;
wire n_9848;
wire n_12081;
wire n_13614;
wire n_14095;
wire n_11202;
wire n_5054;
wire n_9460;
wire n_3171;
wire n_5929;
wire n_6571;
wire n_7710;
wire n_8788;
wire n_5394;
wire n_14080;
wire n_8324;
wire n_16159;
wire n_11227;
wire n_4751;
wire n_4242;
wire n_5975;
wire n_13814;
wire n_10381;
wire n_9841;
wire n_14502;
wire n_15367;
wire n_16324;
wire n_1951;
wire n_12557;
wire n_2490;
wire n_2558;
wire n_10147;
wire n_1496;
wire n_9772;
wire n_2812;
wire n_10554;
wire n_9057;
wire n_14847;
wire n_3300;
wire n_7061;
wire n_8104;
wire n_11860;
wire n_9068;
wire n_7066;
wire n_5496;
wire n_7485;
wire n_3104;
wire n_7174;
wire n_8014;
wire n_12213;
wire n_4122;
wire n_6661;
wire n_16265;
wire n_10919;
wire n_12646;
wire n_2132;
wire n_14750;
wire n_4522;
wire n_15350;
wire n_10228;
wire n_14159;
wire n_5991;
wire n_8623;
wire n_14077;
wire n_14518;
wire n_4952;
wire n_9634;
wire n_6967;
wire n_4426;
wire n_15704;
wire n_5956;
wire n_5699;
wire n_15766;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_11125;
wire n_9348;
wire n_15209;
wire n_15554;
wire n_3946;
wire n_5920;
wire n_13011;
wire n_12737;
wire n_2112;
wire n_2640;
wire n_6125;
wire n_8651;
wire n_5000;
wire n_10699;
wire n_4634;
wire n_9632;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_14358;
wire n_12092;
wire n_2237;
wire n_11951;
wire n_2983;
wire n_5211;
wire n_9257;
wire n_4089;
wire n_15017;
wire n_11451;
wire n_11816;
wire n_9500;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_9747;
wire n_2350;
wire n_9470;
wire n_11508;
wire n_6414;
wire n_5535;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_6097;
wire n_14467;
wire n_7783;
wire n_11232;
wire n_7662;
wire n_6057;
wire n_6936;
wire n_13531;
wire n_10188;
wire n_14898;
wire n_9591;
wire n_11138;
wire n_14373;
wire n_9049;
wire n_487;
wire n_14912;
wire n_4728;
wire n_7171;
wire n_7990;
wire n_1886;
wire n_4346;
wire n_13585;
wire n_1648;
wire n_7003;
wire n_10433;
wire n_8137;
wire n_2187;
wire n_10231;
wire n_1413;
wire n_8413;
wire n_10841;
wire n_2481;
wire n_3863;
wire n_6302;
wire n_10929;
wire n_12642;
wire n_13142;
wire n_15300;
wire n_2327;
wire n_158;
wire n_16912;
wire n_3882;
wire n_13974;
wire n_9471;
wire n_3916;
wire n_6922;
wire n_14656;
wire n_15185;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_14070;
wire n_14909;
wire n_15772;
wire n_16004;
wire n_15294;
wire n_10582;
wire n_16660;
wire n_13494;
wire n_12601;
wire n_16361;
wire n_2841;
wire n_405;
wire n_15210;
wire n_10719;
wire n_3332;
wire n_8300;
wire n_8069;
wire n_10934;
wire n_10747;
wire n_11383;
wire n_7501;
wire n_320;
wire n_9409;
wire n_10711;
wire n_10743;
wire n_11088;
wire n_6432;
wire n_12959;
wire n_7984;
wire n_12899;
wire n_2055;
wire n_15447;
wire n_12616;
wire n_17040;
wire n_2998;
wire n_7366;
wire n_1423;
wire n_8173;
wire n_4359;
wire n_10481;
wire n_13562;
wire n_481;
wire n_1609;
wire n_13540;
wire n_12919;
wire n_15895;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_14953;
wire n_7589;
wire n_13568;
wire n_13642;
wire n_15379;
wire n_16775;
wire n_4447;
wire n_14764;
wire n_2937;
wire n_4293;
wire n_218;
wire n_12511;
wire n_16290;
wire n_6880;
wire n_5176;
wire n_6223;
wire n_9832;
wire n_4039;
wire n_12010;
wire n_12314;
wire n_5793;
wire n_14632;
wire n_6926;
wire n_1798;
wire n_13751;
wire n_8091;
wire n_3057;
wire n_1608;
wire n_12394;
wire n_12856;
wire n_5761;
wire n_13465;
wire n_6699;
wire n_12797;
wire n_547;
wire n_13683;
wire n_16231;
wire n_13630;
wire n_439;
wire n_677;
wire n_3983;
wire n_9067;
wire n_8254;
wire n_703;
wire n_8400;
wire n_10141;
wire n_11090;
wire n_14661;
wire n_10305;
wire n_3318;
wire n_7232;
wire n_3385;
wire n_16728;
wire n_16801;
wire n_15372;
wire n_9858;
wire n_7511;
wire n_326;
wire n_10936;
wire n_12134;
wire n_227;
wire n_13824;
wire n_12730;
wire n_3773;
wire n_17103;
wire n_3494;
wire n_9482;
wire n_1278;
wire n_11429;
wire n_6957;
wire n_9033;
wire n_15570;
wire n_5074;
wire n_14624;
wire n_17147;
wire n_12735;
wire n_14510;
wire n_7917;
wire n_11908;
wire n_3788;
wire n_3939;
wire n_727;
wire n_590;
wire n_16494;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_8368;
wire n_15388;
wire n_6694;
wire n_545;
wire n_9247;
wire n_2496;
wire n_3260;
wire n_8463;
wire n_536;
wire n_10425;
wire n_9965;
wire n_15226;
wire n_15927;
wire n_3349;
wire n_6449;
wire n_16944;
wire n_10862;
wire n_12254;
wire n_14333;
wire n_4348;
wire n_1602;
wire n_16739;
wire n_7422;
wire n_9299;
wire n_13357;
wire n_3139;
wire n_8889;
wire n_427;
wire n_3801;
wire n_5681;
wire n_9785;
wire n_11298;
wire n_9244;
wire n_14667;
wire n_16232;
wire n_2338;
wire n_5261;
wire n_16871;
wire n_12427;
wire n_1080;
wire n_12124;
wire n_9195;
wire n_8322;
wire n_11353;
wire n_12494;
wire n_15623;
wire n_3636;
wire n_6591;
wire n_7466;
wire n_8987;
wire n_13454;
wire n_3653;
wire n_16529;
wire n_3823;
wire n_9280;
wire n_3403;
wire n_7621;
wire n_9911;
wire n_12051;
wire n_13958;
wire n_8274;
wire n_2057;
wire n_6594;
wire n_6342;
wire n_1205;
wire n_6195;
wire n_14802;
wire n_163;
wire n_6826;
wire n_2716;
wire n_10373;
wire n_6441;
wire n_11116;
wire n_7158;
wire n_13637;
wire n_7572;
wire n_11173;
wire n_16603;
wire n_314;
wire n_2944;
wire n_11660;
wire n_15675;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_7500;
wire n_1202;
wire n_4084;
wire n_627;
wire n_12355;
wire n_17052;
wire n_7985;
wire n_9687;
wire n_1371;
wire n_4240;
wire n_8657;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_11567;
wire n_233;
wire n_8954;
wire n_16838;
wire n_2774;
wire n_6354;
wire n_11881;
wire n_10563;
wire n_12458;
wire n_2799;
wire n_8311;
wire n_15786;
wire n_5748;
wire n_4393;
wire n_11363;
wire n_321;
wire n_17152;
wire n_6662;
wire n_7494;
wire n_9088;
wire n_3984;
wire n_1586;
wire n_16250;
wire n_14050;
wire n_8728;
wire n_17094;
wire n_9580;
wire n_11280;
wire n_9569;
wire n_16435;
wire n_1431;
wire n_8994;
wire n_4389;
wire n_6433;
wire n_16589;
wire n_9680;
wire n_1763;
wire n_8398;
wire n_6200;
wire n_5641;
wire n_12463;
wire n_12612;
wire n_8407;
wire n_8071;
wire n_13423;
wire n_13046;
wire n_16292;
wire n_4461;
wire n_2763;
wire n_11636;
wire n_3156;
wire n_14926;
wire n_16355;
wire n_17048;
wire n_10530;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_6902;
wire n_4615;
wire n_3492;
wire n_3044;
wire n_12798;
wire n_7197;
wire n_3737;
wire n_6369;
wire n_8528;
wire n_14088;
wire n_16993;
wire n_9227;
wire n_13644;
wire n_5657;
wire n_16685;
wire n_12510;
wire n_11313;
wire n_14364;
wire n_8475;
wire n_297;
wire n_9951;
wire n_15182;
wire n_9855;
wire n_2379;
wire n_3579;
wire n_9072;
wire n_12635;
wire n_10102;
wire n_13545;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_12537;
wire n_14913;
wire n_4067;
wire n_13197;
wire n_1677;
wire n_5244;
wire n_5765;
wire n_12076;
wire n_5114;
wire n_9054;
wire n_4551;
wire n_15836;
wire n_178;
wire n_10117;
wire n_551;
wire n_4521;
wire n_13252;
wire n_13139;
wire n_6956;
wire n_10126;
wire n_7587;
wire n_2284;
wire n_6451;
wire n_12874;
wire n_11920;
wire n_3005;
wire n_7704;
wire n_10604;
wire n_6497;
wire n_5420;
wire n_8511;
wire n_16915;
wire n_16289;
wire n_7865;
wire n_2283;
wire n_5206;
wire n_582;
wire n_2526;
wire n_13356;
wire n_1097;
wire n_14447;
wire n_16039;
wire n_1711;
wire n_4387;
wire n_14237;
wire n_14745;
wire n_9584;
wire n_9287;
wire n_534;
wire n_2508;
wire n_3186;
wire n_10344;
wire n_10568;
wire n_9459;
wire n_6701;
wire n_2594;
wire n_1239;
wire n_5298;
wire n_9490;
wire n_10209;
wire n_16770;
wire n_8867;
wire n_3417;
wire n_8246;
wire n_560;
wire n_8558;
wire n_890;
wire n_9655;
wire n_13769;
wire n_9846;
wire n_3626;
wire n_12048;
wire n_451;
wire n_9593;
wire n_4598;
wire n_4464;
wire n_12072;
wire n_8925;
wire n_5106;
wire n_7881;
wire n_11317;
wire n_9147;
wire n_13339;
wire n_15854;
wire n_4789;
wire n_16394;
wire n_3180;
wire n_14433;
wire n_12829;
wire n_3423;
wire n_14672;
wire n_1081;
wire n_9678;
wire n_16988;
wire n_10803;
wire n_2119;
wire n_12132;
wire n_13626;
wire n_11903;
wire n_8641;
wire n_9658;
wire n_10299;
wire n_2493;
wire n_9560;
wire n_15036;
wire n_12528;
wire n_9578;
wire n_16732;
wire n_11813;
wire n_14195;
wire n_5080;
wire n_535;
wire n_9396;
wire n_4565;
wire n_7032;
wire n_12745;
wire n_16061;
wire n_9303;
wire n_3392;
wire n_12371;
wire n_1800;
wire n_11811;
wire n_12841;
wire n_7198;
wire n_12417;
wire n_14866;
wire n_6884;
wire n_7752;
wire n_10618;
wire n_11378;
wire n_10836;
wire n_5081;
wire n_8201;
wire n_6921;
wire n_2904;
wire n_12180;
wire n_16743;
wire n_12049;
wire n_3353;
wire n_2946;
wire n_16691;
wire n_7953;
wire n_6106;
wire n_14434;
wire n_16086;
wire n_6876;
wire n_15746;
wire n_16446;
wire n_3512;
wire n_9553;
wire n_12603;
wire n_1734;
wire n_1860;
wire n_4552;
wire n_8046;
wire n_14964;
wire n_12978;
wire n_7193;
wire n_6287;
wire n_2840;
wire n_14575;
wire n_10930;
wire n_6172;
wire n_14005;
wire n_9942;
wire n_9805;
wire n_13686;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_5957;
wire n_12466;
wire n_13842;
wire n_4040;
wire n_16220;
wire n_8414;
wire n_3024;
wire n_5567;
wire n_8292;
wire n_9138;
wire n_9879;
wire n_5406;
wire n_8647;
wire n_11936;
wire n_6362;
wire n_9213;
wire n_12071;
wire n_17119;
wire n_4328;
wire n_12982;
wire n_8543;
wire n_14680;
wire n_13459;
wire n_1854;
wire n_666;
wire n_11543;
wire n_15637;
wire n_11184;
wire n_11795;
wire n_5191;
wire n_11391;
wire n_1206;
wire n_1729;
wire n_17149;
wire n_1508;
wire n_6067;
wire n_2893;
wire n_11646;
wire n_6833;
wire n_4940;
wire n_15156;
wire n_9374;
wire n_785;
wire n_3161;
wire n_13649;
wire n_2389;
wire n_14720;
wire n_14497;
wire n_1309;
wire n_8331;
wire n_999;
wire n_2280;
wire n_8317;
wire n_7126;
wire n_12578;
wire n_12311;
wire n_11963;
wire n_5867;
wire n_14109;
wire n_13253;
wire n_456;
wire n_12985;
wire n_12232;
wire n_1394;
wire n_15316;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_12640;
wire n_13729;
wire n_7496;
wire n_15027;
wire n_6430;
wire n_11435;
wire n_13647;
wire n_9179;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_6296;
wire n_11056;
wire n_4112;
wire n_342;
wire n_10014;
wire n_10714;
wire n_5602;
wire n_2035;
wire n_4928;
wire n_7196;
wire n_14241;
wire n_2614;
wire n_12101;
wire n_14855;
wire n_16275;
wire n_16514;
wire n_11120;
wire n_11185;
wire n_7360;
wire n_5428;
wire n_10895;
wire n_6325;
wire n_10916;
wire n_14693;
wire n_12497;
wire n_2494;
wire n_12197;
wire n_1538;
wire n_4865;
wire n_15611;
wire n_6678;
wire n_7982;
wire n_10838;
wire n_13002;
wire n_2128;
wire n_4071;
wire n_7268;
wire n_8929;
wire n_8174;
wire n_8187;
wire n_10108;
wire n_14069;
wire n_6564;
wire n_4436;
wire n_15196;
wire n_5786;
wire n_5822;
wire n_15964;
wire n_17095;
wire n_3586;
wire n_10661;
wire n_8846;
wire n_5817;
wire n_16587;
wire n_9277;
wire n_4160;
wire n_14754;
wire n_15111;
wire n_15151;
wire n_6109;
wire n_9611;
wire n_6385;
wire n_1668;
wire n_16400;
wire n_12571;
wire n_9744;
wire n_5798;
wire n_10123;
wire n_4137;
wire n_1078;
wire n_13022;
wire n_15949;
wire n_9504;
wire n_8032;
wire n_16865;
wire n_5417;
wire n_14118;
wire n_14445;
wire n_11147;
wire n_10048;
wire n_4545;
wire n_11194;
wire n_8200;
wire n_9285;
wire n_1161;
wire n_15068;
wire n_15590;
wire n_15771;
wire n_4758;
wire n_4840;
wire n_5713;
wire n_9905;
wire n_10963;
wire n_11016;
wire n_12228;
wire n_11146;
wire n_3097;
wire n_13088;
wire n_16971;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_10788;
wire n_16161;
wire n_14142;
wire n_9190;
wire n_8586;
wire n_15937;
wire n_8524;
wire n_618;
wire n_1191;
wire n_11924;
wire n_12540;
wire n_4535;
wire n_8828;
wire n_9639;
wire n_10422;
wire n_7518;
wire n_4385;
wire n_12001;
wire n_15916;
wire n_7779;
wire n_12059;
wire n_9664;
wire n_1215;
wire n_13275;
wire n_16434;
wire n_11830;
wire n_14577;
wire n_3748;
wire n_4731;
wire n_11489;
wire n_7575;
wire n_2337;
wire n_7073;
wire n_13026;
wire n_15753;
wire n_8092;
wire n_10471;
wire n_16582;
wire n_13760;
wire n_12479;
wire n_16087;
wire n_10979;
wire n_1786;
wire n_6309;
wire n_8370;
wire n_16894;
wire n_3732;
wire n_9109;
wire n_211;
wire n_1804;
wire n_10189;
wire n_408;
wire n_13820;
wire n_8135;
wire n_12702;
wire n_6519;
wire n_4671;
wire n_14366;
wire n_9741;
wire n_2272;
wire n_5571;
wire n_4766;
wire n_5989;
wire n_592;
wire n_4558;
wire n_10569;
wire n_13116;
wire n_13663;
wire n_10686;
wire n_1318;
wire n_14055;
wire n_14197;
wire n_16153;
wire n_8764;
wire n_14454;
wire n_1769;
wire n_1632;
wire n_7349;
wire n_1929;
wire n_9875;
wire n_8502;
wire n_10713;
wire n_11411;
wire n_4319;
wire n_12211;
wire n_6585;
wire n_9360;
wire n_14323;
wire n_7786;
wire n_10913;
wire n_9021;
wire n_8454;
wire n_2929;
wire n_16325;
wire n_12306;
wire n_4358;
wire n_11145;
wire n_9122;
wire n_1526;
wire n_7579;
wire n_10099;
wire n_7122;
wire n_12637;
wire n_12335;
wire n_10193;
wire n_14096;
wire n_4874;
wire n_180;
wire n_2656;
wire n_4904;
wire n_516;
wire n_1997;
wire n_10203;
wire n_10140;
wire n_13982;
wire n_1137;
wire n_16979;
wire n_1258;
wire n_640;
wire n_1733;
wire n_6490;
wire n_7867;
wire n_4651;
wire n_10920;
wire n_11000;
wire n_943;
wire n_11712;
wire n_10149;
wire n_14068;
wire n_3167;
wire n_4748;
wire n_14019;
wire n_7624;
wire n_13405;
wire n_9803;
wire n_13828;
wire n_14397;
wire n_16895;
wire n_16441;
wire n_1807;
wire n_1123;
wire n_15738;
wire n_8776;
wire n_10576;
wire n_2857;
wire n_8564;
wire n_16744;
wire n_12114;
wire n_8343;
wire n_7828;
wire n_14319;
wire n_1784;
wire n_4618;
wire n_6721;
wire n_3787;
wire n_4025;
wire n_15106;
wire n_1321;
wire n_16984;
wire n_3050;
wire n_3919;
wire n_8718;
wire n_13102;
wire n_13550;
wire n_14301;
wire n_10682;
wire n_752;
wire n_14910;
wire n_16198;
wire n_985;
wire n_5506;
wire n_7543;
wire n_9659;
wire n_12204;
wire n_13643;
wire n_15997;
wire n_15812;
wire n_16252;
wire n_5475;
wire n_8042;
wire n_7727;
wire n_2412;
wire n_16382;
wire n_14774;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_1352;
wire n_9013;
wire n_5431;
wire n_9427;
wire n_12325;
wire n_8379;
wire n_643;
wire n_8034;
wire n_12143;
wire n_226;
wire n_7778;
wire n_5100;
wire n_2383;
wire n_10225;
wire n_2764;
wire n_1822;
wire n_1441;
wire n_7019;
wire n_682;
wire n_9126;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_5752;
wire n_2907;
wire n_8441;
wire n_9474;
wire n_14026;
wire n_14362;
wire n_1429;
wire n_2353;
wire n_7702;
wire n_14114;
wire n_2528;
wire n_1778;
wire n_5746;
wire n_686;
wire n_10368;
wire n_1154;
wire n_584;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_10237;
wire n_14504;
wire n_9538;
wire n_3718;
wire n_6685;
wire n_14930;
wire n_756;
wire n_3390;
wire n_16374;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_8569;
wire n_9574;
wire n_10531;
wire n_12032;
wire n_4666;
wire n_3140;
wire n_2320;
wire n_4082;
wire n_979;
wire n_12066;
wire n_14471;
wire n_8865;
wire n_8592;
wire n_3976;
wire n_2813;
wire n_897;
wire n_2546;
wire n_3381;
wire n_7952;
wire n_11170;
wire n_7347;
wire n_9450;
wire n_3736;
wire n_10031;
wire n_4466;
wire n_6016;
wire n_9998;
wire n_891;
wire n_13963;
wire n_885;
wire n_1659;
wire n_3955;
wire n_15568;
wire n_15948;
wire n_5366;
wire n_11523;
wire n_5322;
wire n_1864;
wire n_11121;
wire n_12176;
wire n_5414;
wire n_11805;
wire n_3086;
wire n_13266;
wire n_1887;
wire n_3165;
wire n_7791;
wire n_8362;
wire n_6971;
wire n_10847;
wire n_3336;
wire n_8632;
wire n_10035;
wire n_14242;
wire n_14523;
wire n_16295;
wire n_15660;
wire n_7739;
wire n_396;
wire n_12740;
wire n_9372;
wire n_15040;
wire n_9045;
wire n_7945;
wire n_16233;
wire n_8361;
wire n_9657;
wire n_14883;
wire n_11457;
wire n_7656;
wire n_5903;
wire n_7199;
wire n_10107;
wire n_3635;
wire n_11725;
wire n_3541;
wire n_2502;
wire n_10283;
wire n_5151;
wire n_15731;
wire n_714;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_9904;
wire n_12344;
wire n_14937;
wire n_9924;
wire n_17154;
wire n_9159;
wire n_8561;
wire n_6549;
wire n_725;
wire n_8611;
wire n_9326;
wire n_8410;
wire n_1577;
wire n_15486;
wire n_16225;
wire n_16662;
wire n_5003;
wire n_3840;
wire n_6540;
wire n_7166;
wire n_2198;
wire n_11694;
wire n_6658;
wire n_5369;
wire n_9476;
wire n_16360;
wire n_6683;
wire n_15634;
wire n_3067;
wire n_154;
wire n_16496;
wire n_3809;
wire n_4921;
wire n_473;
wire n_1852;
wire n_801;
wire n_5912;
wire n_11540;
wire n_5745;
wire n_7923;
wire n_6086;
wire n_4377;
wire n_818;
wire n_10050;
wire n_14800;
wire n_11058;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_15743;
wire n_5803;
wire n_8878;
wire n_6327;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_3468;
wire n_5779;
wire n_12203;
wire n_15606;
wire n_16156;
wire n_1877;
wire n_11403;
wire n_272;
wire n_9301;
wire n_8492;
wire n_14099;
wire n_7213;
wire n_16964;
wire n_4301;
wire n_5313;
wire n_10392;
wire n_2133;
wire n_14041;
wire n_12769;
wire n_15076;
wire n_8888;
wire n_6820;
wire n_2497;
wire n_879;
wire n_5446;
wire n_11741;
wire n_11245;
wire n_7107;
wire n_7610;
wire n_4561;
wire n_14225;
wire n_1541;
wire n_597;
wire n_3291;
wire n_9382;
wire n_15426;
wire n_11784;
wire n_7456;
wire n_8095;
wire n_11365;
wire n_13291;
wire n_14756;
wire n_9921;
wire n_7369;
wire n_15559;
wire n_1472;
wire n_14888;
wire n_9325;
wire n_1050;
wire n_11005;
wire n_9643;
wire n_13016;
wire n_9945;
wire n_7548;
wire n_2578;
wire n_12820;
wire n_152;
wire n_1201;
wire n_8735;
wire n_15073;
wire n_7598;
wire n_1185;
wire n_2475;
wire n_7250;
wire n_8808;
wire n_9201;
wire n_8902;
wire n_7823;
wire n_9771;
wire n_8833;
wire n_14605;
wire n_12869;
wire n_4715;
wire n_6157;
wire n_8796;
wire n_2715;
wire n_335;
wire n_14413;
wire n_16154;
wire n_2665;
wire n_4879;
wire n_344;
wire n_13435;
wire n_16031;
wire n_8794;
wire n_12689;
wire n_11074;
wire n_5044;
wire n_210;
wire n_1090;
wire n_3755;
wire n_4536;
wire n_9894;
wire n_11141;
wire n_12750;
wire n_9274;
wire n_14753;
wire n_8549;
wire n_15936;
wire n_14161;
wire n_16827;
wire n_6676;
wire n_4304;
wire n_10095;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_14285;
wire n_10716;
wire n_11102;
wire n_12171;
wire n_14812;
wire n_14000;
wire n_224;
wire n_10088;
wire n_11238;
wire n_11406;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_16000;
wire n_10443;
wire n_10488;
wire n_7525;
wire n_16251;
wire n_4418;
wire n_7924;
wire n_3341;
wire n_11103;
wire n_12420;
wire n_9232;
wire n_8690;
wire n_16826;
wire n_4125;
wire n_5390;
wire n_16924;
wire n_16557;
wire n_12954;
wire n_17032;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_11852;
wire n_5024;
wire n_7012;
wire n_3043;
wire n_2747;
wire n_12500;
wire n_1511;
wire n_15393;
wire n_16599;
wire n_8593;
wire n_11837;
wire n_10912;
wire n_13501;
wire n_10469;
wire n_276;
wire n_15958;
wire n_13533;
wire n_9649;
wire n_11684;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_12112;
wire n_15377;
wire n_1641;
wire n_15864;
wire n_3731;
wire n_4527;
wire n_16562;
wire n_4291;
wire n_538;
wire n_2845;
wire n_4151;
wire n_4412;
wire n_2036;
wire n_6923;
wire n_7649;
wire n_843;
wire n_8588;
wire n_8009;
wire n_8195;
wire n_16027;
wire n_15628;
wire n_9839;
wire n_10887;
wire n_16788;
wire n_3358;
wire n_12004;
wire n_7634;
wire n_9090;
wire n_6704;
wire n_2533;
wire n_2003;
wire n_1307;
wire n_7406;
wire n_13520;
wire n_4682;
wire n_1128;
wire n_9346;
wire n_11012;
wire n_6673;
wire n_14480;
wire n_9696;
wire n_2419;
wire n_11041;
wire n_14181;
wire n_10742;
wire n_2330;
wire n_14024;
wire n_11798;
wire n_12614;
wire n_13165;
wire n_15312;
wire n_9996;
wire n_6534;
wire n_9968;
wire n_8805;
wire n_5078;
wire n_4810;
wire n_7659;
wire n_6162;
wire n_3189;
wire n_2309;
wire n_16575;
wire n_4957;
wire n_15576;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_6127;
wire n_9383;
wire n_9498;
wire n_10405;
wire n_1440;
wire n_6246;
wire n_10390;
wire n_11978;
wire n_1370;
wire n_10989;
wire n_305;
wire n_9836;
wire n_5005;
wire n_14570;
wire n_14702;
wire n_11827;
wire n_10328;
wire n_16191;
wire n_13315;
wire n_10692;
wire n_15118;
wire n_6126;
wire n_8596;
wire n_12912;
wire n_9938;
wire n_7372;
wire n_1549;
wire n_7427;
wire n_16467;
wire n_6151;
wire n_6828;
wire n_15592;
wire n_10867;
wire n_6841;
wire n_11847;
wire n_10206;
wire n_16697;
wire n_7844;
wire n_5207;
wire n_7934;
wire n_11281;
wire n_16837;
wire n_361;
wire n_2658;
wire n_12957;
wire n_5624;
wire n_10092;
wire n_3620;
wire n_4601;
wire n_16377;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_5474;
wire n_7009;
wire n_3376;
wire n_11772;
wire n_16371;
wire n_181;
wire n_15837;
wire n_9743;
wire n_9121;
wire n_7371;
wire n_13448;
wire n_1362;
wire n_16661;
wire n_11237;
wire n_14752;
wire n_9509;
wire n_3123;
wire n_5447;
wire n_12153;
wire n_2692;
wire n_12005;
wire n_683;
wire n_16493;
wire n_7463;
wire n_9621;
wire n_1300;
wire n_1960;
wire n_15966;
wire n_4102;
wire n_10738;
wire n_5700;
wire n_5755;
wire n_11851;
wire n_4308;
wire n_16961;
wire n_9158;
wire n_2862;
wire n_4325;
wire n_14239;
wire n_14501;
wire n_1420;
wire n_2645;
wire n_2553;
wire n_4711;
wire n_16068;
wire n_6889;
wire n_2749;
wire n_12586;
wire n_11993;
wire n_5962;
wire n_660;
wire n_464;
wire n_15710;
wire n_4413;
wire n_16780;
wire n_11131;
wire n_12221;
wire n_17074;
wire n_8627;
wire n_1210;
wire n_14318;
wire n_11432;
wire n_12302;
wire n_3307;
wire n_8945;
wire n_9142;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_13628;
wire n_2833;
wire n_9216;
wire n_9189;
wire n_6723;
wire n_7398;
wire n_1038;
wire n_3723;
wire n_9563;
wire n_4135;
wire n_7941;
wire n_12757;
wire n_13010;
wire n_6154;
wire n_15229;
wire n_5223;
wire n_5662;
wire n_13251;
wire n_14738;
wire n_8858;
wire n_12107;
wire n_414;
wire n_571;
wire n_11738;
wire n_11595;
wire n_3880;
wire n_13504;
wire n_13521;
wire n_14404;
wire n_16886;
wire n_12695;
wire n_11512;
wire n_5801;
wire n_14163;
wire n_16723;
wire n_3904;
wire n_15504;
wire n_12349;
wire n_6054;
wire n_13703;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_14758;
wire n_13161;
wire n_7011;
wire n_10813;
wire n_3405;
wire n_15403;
wire n_2313;
wire n_14076;
wire n_10986;
wire n_11603;
wire n_15573;
wire n_6393;
wire n_14291;
wire n_14761;
wire n_17167;
wire n_12380;
wire n_7074;
wire n_10853;
wire n_8916;
wire n_10899;
wire n_11707;
wire n_11728;
wire n_613;
wire n_13352;
wire n_11521;
wire n_1022;
wire n_13309;
wire n_5465;
wire n_16137;
wire n_12577;
wire n_10575;
wire n_171;
wire n_8745;
wire n_3532;
wire n_5154;
wire n_14388;
wire n_5721;
wire n_2609;
wire n_8169;
wire n_14932;
wire n_6184;
wire n_8018;
wire n_11802;
wire n_1767;
wire n_9984;
wire n_1040;
wire n_4138;
wire n_3131;
wire n_7083;
wire n_316;
wire n_1973;
wire n_1444;
wire n_15889;
wire n_820;
wire n_8260;
wire n_12723;
wire n_10334;
wire n_14153;
wire n_12135;
wire n_254;
wire n_2882;
wire n_14674;
wire n_7143;
wire n_2303;
wire n_7701;
wire n_11688;
wire n_16419;
wire n_13484;
wire n_16939;
wire n_9794;
wire n_8688;
wire n_15761;
wire n_7969;
wire n_16062;
wire n_10726;
wire n_16210;
wire n_8279;
wire n_4384;
wire n_16712;
wire n_8793;
wire n_4639;
wire n_1664;
wire n_12864;
wire n_13486;
wire n_10388;
wire n_4577;
wire n_6312;
wire n_13478;
wire n_7683;
wire n_9550;
wire n_13108;
wire n_532;
wire n_11042;
wire n_2154;
wire n_15701;
wire n_12570;
wire n_14124;
wire n_15932;
wire n_10510;
wire n_6955;
wire n_14344;
wire n_7669;
wire n_1986;
wire n_8298;
wire n_6711;
wire n_2624;
wire n_6818;
wire n_11696;
wire n_15802;
wire n_6438;
wire n_2054;
wire n_1857;
wire n_11761;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_10635;
wire n_17047;
wire n_11681;
wire n_1552;
wire n_2938;
wire n_7209;
wire n_2498;
wire n_13429;
wire n_6193;
wire n_3992;
wire n_13897;
wire n_8023;
wire n_9319;
wire n_7330;
wire n_6007;
wire n_13374;
wire n_16906;
wire n_621;
wire n_13182;
wire n_16969;
wire n_10852;
wire n_14867;
wire n_6535;
wire n_14893;
wire n_6734;
wire n_17174;
wire n_13789;
wire n_15893;
wire n_11407;
wire n_8053;
wire n_8059;
wire n_1772;
wire n_9871;
wire n_14354;
wire n_6879;
wire n_9562;
wire n_15442;
wire n_15632;
wire n_9896;
wire n_9612;
wire n_493;
wire n_1311;
wire n_3106;
wire n_6208;
wire n_7190;
wire n_9698;
wire n_2881;
wire n_6303;
wire n_3092;
wire n_6014;
wire n_15840;
wire n_4270;
wire n_7692;
wire n_697;
wire n_10241;
wire n_13690;
wire n_4620;
wire n_5397;
wire n_6457;
wire n_9528;
wire n_14016;
wire n_9272;
wire n_13055;
wire n_14379;
wire n_9955;
wire n_15451;
wire n_9645;
wire n_15953;
wire n_4924;
wire n_4044;
wire n_8372;
wire n_6270;
wire n_14283;
wire n_2305;
wire n_8737;
wire n_10026;
wire n_9731;
wire n_15999;
wire n_5996;
wire n_880;
wire n_13577;
wire n_5566;
wire n_16392;
wire n_9697;
wire n_3304;
wire n_7288;
wire n_15307;
wire n_10772;
wire n_4388;
wire n_13098;
wire n_10901;
wire n_7362;
wire n_15855;
wire n_14942;
wire n_7237;
wire n_7082;
wire n_8988;
wire n_3247;
wire n_10664;
wire n_7131;
wire n_6276;
wire n_739;
wire n_1028;
wire n_15661;
wire n_12328;
wire n_13839;
wire n_9642;
wire n_530;
wire n_8723;
wire n_11189;
wire n_12559;
wire n_9929;
wire n_9050;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_12056;
wire n_13898;
wire n_15030;
wire n_16204;
wire n_7042;
wire n_9859;
wire n_8419;
wire n_2809;
wire n_10767;
wire n_10320;
wire n_5652;
wire n_13380;
wire n_8893;
wire n_975;
wire n_1645;
wire n_5805;
wire n_16375;
wire n_7304;
wire n_932;
wire n_11910;
wire n_16235;
wire n_6266;
wire n_2276;
wire n_15386;
wire n_3301;
wire n_12109;
wire n_2910;
wire n_14457;
wire n_2503;
wire n_14905;
wire n_9531;
wire n_10521;
wire n_3785;
wire n_5492;
wire n_8077;
wire n_11242;
wire n_2465;
wire n_5501;
wire n_12917;
wire n_14711;
wire n_15445;
wire n_6934;
wire n_16586;
wire n_13188;
wire n_17158;
wire n_14179;
wire n_13362;
wire n_15259;
wire n_2972;
wire n_7386;
wire n_7391;
wire n_4401;
wire n_11361;
wire n_2586;
wire n_2989;
wire n_12058;
wire n_8826;
wire n_3178;
wire n_11894;
wire n_13819;
wire n_268;
wire n_15631;
wire n_13990;
wire n_10872;
wire n_7023;
wire n_15745;
wire n_2251;
wire n_9732;
wire n_5758;
wire n_12083;
wire n_5842;
wire n_9685;
wire n_12529;
wire n_3100;
wire n_15521;
wire n_3721;
wire n_10374;
wire n_11253;
wire n_13983;
wire n_12045;
wire n_13193;
wire n_14995;
wire n_15856;
wire n_7404;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_17113;
wire n_10345;
wire n_8959;
wire n_15648;
wire n_6147;
wire n_5692;
wire n_6765;
wire n_12471;
wire n_4973;
wire n_13802;
wire n_13781;
wire n_15887;
wire n_7981;
wire n_4792;
wire n_1601;
wire n_13037;
wire n_3537;
wire n_4402;
wire n_14252;
wire n_14736;
wire n_15058;
wire n_15351;
wire n_12188;
wire n_191;
wire n_14851;
wire n_2487;
wire n_5473;
wire n_12575;
wire n_1834;
wire n_10601;
wire n_14698;
wire n_16619;
wire n_16869;
wire n_11623;
wire n_8712;
wire n_12473;
wire n_10372;
wire n_1011;
wire n_15394;
wire n_2534;
wire n_11124;
wire n_14295;
wire n_6352;
wire n_2941;
wire n_4286;
wire n_9378;
wire n_3638;
wire n_6211;
wire n_17112;
wire n_10448;
wire n_15100;
wire n_8109;
wire n_10301;
wire n_11977;
wire n_15487;
wire n_3576;
wire n_10074;
wire n_12040;
wire n_14025;
wire n_13127;
wire n_9389;
wire n_12598;
wire n_5562;
wire n_4858;
wire n_1445;
wire n_6093;
wire n_5370;
wire n_16859;
wire n_10001;
wire n_13561;
wire n_7378;
wire n_15922;
wire n_9623;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_14944;
wire n_15987;
wire n_15562;
wire n_7877;
wire n_14336;
wire n_16938;
wire n_11351;
wire n_7787;
wire n_7836;
wire n_8515;
wire n_8725;
wire n_12626;
wire n_11094;
wire n_10960;
wire n_10712;
wire n_8007;
wire n_13911;
wire n_14313;
wire n_2387;
wire n_15578;
wire n_4318;
wire n_332;
wire n_13961;
wire n_16849;
wire n_13343;
wire n_12546;
wire n_8910;
wire n_16412;
wire n_16070;
wire n_5227;
wire n_14091;
wire n_830;
wire n_14842;
wire n_15981;
wire n_10100;
wire n_5902;
wire n_987;
wire n_2510;
wire n_9164;
wire n_6402;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_11366;
wire n_2793;
wire n_5282;
wire n_9387;
wire n_8301;
wire n_7871;
wire n_14512;
wire n_6764;
wire n_541;
wire n_499;
wire n_13539;
wire n_10162;
wire n_16679;
wire n_2639;
wire n_9840;
wire n_15982;
wire n_15471;
wire n_7016;
wire n_4738;
wire n_17019;
wire n_12100;
wire n_2603;
wire n_8892;
wire n_11399;
wire n_16835;
wire n_9637;
wire n_5386;
wire n_1167;
wire n_12676;
wire n_4554;
wire n_13584;
wire n_8252;
wire n_4526;
wire n_4105;
wire n_10535;
wire n_10674;
wire n_7571;
wire n_6215;
wire n_969;
wire n_3663;
wire n_9491;
wire n_1663;
wire n_7563;
wire n_10774;
wire n_13107;
wire n_10337;
wire n_5952;
wire n_7180;
wire n_14655;
wire n_10407;
wire n_14850;
wire n_16253;
wire n_10577;
wire n_2086;
wire n_14481;
wire n_13778;
wire n_16171;
wire n_1926;
wire n_8972;
wire n_14531;
wire n_8494;
wire n_12999;
wire n_14709;
wire n_10264;
wire n_15148;
wire n_6569;
wire n_1630;
wire n_16710;
wire n_7919;
wire n_13740;
wire n_15355;
wire n_9992;
wire n_14606;
wire n_14089;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_8278;
wire n_443;
wire n_3431;
wire n_8180;
wire n_11549;
wire n_14437;
wire n_12362;
wire n_3355;
wire n_7031;
wire n_13913;
wire n_1738;
wire n_13367;
wire n_5716;
wire n_10313;
wire n_10843;
wire n_12983;
wire n_14003;
wire n_8941;
wire n_10771;
wire n_8891;
wire n_406;
wire n_3897;
wire n_7103;
wire n_12360;
wire n_139;
wire n_13570;
wire n_6605;
wire n_10724;
wire n_1735;
wire n_391;
wire n_16356;
wire n_5888;
wire n_9266;
wire n_4005;
wire n_14409;
wire n_16182;
wire n_8270;
wire n_16103;
wire n_8231;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_11983;
wire n_12313;
wire n_12604;
wire n_15885;
wire n_5980;
wire n_8683;
wire n_956;
wire n_6832;
wire n_15114;
wire n_9391;
wire n_16594;
wire n_765;
wire n_4092;
wire n_12558;
wire n_15503;
wire n_15053;
wire n_10445;
wire n_4875;
wire n_7771;
wire n_8903;
wire n_4255;
wire n_13284;
wire n_16946;
wire n_2758;
wire n_385;
wire n_8810;
wire n_12596;
wire n_6544;
wire n_6469;
wire n_12840;
wire n_17155;
wire n_5036;
wire n_1271;
wire n_11119;
wire n_12696;
wire n_6332;
wire n_15241;
wire n_10863;
wire n_10958;
wire n_2186;
wire n_11215;
wire n_16335;
wire n_13730;
wire n_5790;
wire n_399;
wire n_10174;
wire n_7130;
wire n_15729;
wire n_6680;
wire n_4647;
wire n_3575;
wire n_13960;
wire n_6310;
wire n_8932;
wire n_8264;
wire n_12435;
wire n_2471;
wire n_9695;
wire n_7134;
wire n_3042;
wire n_8288;
wire n_13411;
wire n_1067;
wire n_11954;
wire n_14629;
wire n_14778;
wire n_15891;
wire n_16240;
wire n_1323;
wire n_11526;
wire n_13438;
wire n_14010;
wire n_11591;
wire n_10403;
wire n_1937;
wire n_16813;
wire n_11972;
wire n_4142;
wire n_5118;
wire n_9834;
wire n_900;
wire n_5485;
wire n_9901;
wire n_5525;
wire n_10076;
wire n_10015;
wire n_7102;
wire n_6259;
wire n_3004;
wire n_14432;
wire n_15371;
wire n_1551;
wire n_4849;
wire n_5271;
wire n_13410;
wire n_2039;
wire n_7133;
wire n_9800;
wire n_1285;
wire n_10745;
wire n_17140;
wire n_193;
wire n_761;
wire n_733;
wire n_3838;
wire n_6289;
wire n_6651;
wire n_9255;
wire n_8882;
wire n_14308;
wire n_12460;
wire n_4059;
wire n_6565;
wire n_5194;
wire n_12733;
wire n_15532;
wire n_8388;
wire n_5445;
wire n_2734;
wire n_13600;
wire n_8067;
wire n_8385;
wire n_5948;
wire n_7227;
wire n_4499;
wire n_15061;
wire n_8670;
wire n_4504;
wire n_16650;
wire n_10460;
wire n_14299;
wire n_14215;
wire n_3598;
wire n_4917;
wire n_7706;
wire n_7813;
wire n_8142;
wire n_13332;
wire n_14265;
wire n_15266;
wire n_13942;
wire n_16280;
wire n_2420;
wire n_7992;
wire n_9085;
wire n_7643;
wire n_15381;
wire n_15090;
wire n_11204;
wire n_153;
wire n_648;
wire n_12939;
wire n_6836;
wire n_3273;
wire n_9120;
wire n_2918;
wire n_6595;
wire n_10415;
wire n_11302;
wire n_835;
wire n_17105;
wire n_16089;
wire n_9899;
wire n_12374;
wire n_15054;
wire n_17150;
wire n_15398;
wire n_9136;
wire n_16898;
wire n_16081;
wire n_12261;
wire n_6186;
wire n_11561;
wire n_10227;
wire n_1865;
wire n_2641;
wire n_13490;
wire n_16767;
wire n_2463;
wire n_14198;
wire n_2580;
wire n_14836;
wire n_401;
wire n_7628;
wire n_1792;
wire n_13381;
wire n_5628;
wire n_504;
wire n_5245;
wire n_2062;
wire n_483;
wire n_4489;
wire n_9436;
wire n_14013;
wire n_15220;
wire n_16684;
wire n_11385;
wire n_822;
wire n_1459;
wire n_2153;
wire n_14989;
wire n_12065;
wire n_13204;
wire n_5329;
wire n_12275;
wire n_8224;
wire n_5472;
wire n_6035;
wire n_10884;
wire n_9042;
wire n_13375;
wire n_839;
wire n_15669;
wire n_1754;
wire n_7236;
wire n_9570;
wire n_4833;
wire n_3394;
wire n_9239;
wire n_6405;
wire n_8345;
wire n_11054;
wire n_11777;
wire n_16722;
wire n_9644;
wire n_2235;
wire n_5850;
wire n_1575;
wire n_9343;
wire n_8614;
wire n_16751;
wire n_8242;
wire n_6786;
wire n_4564;
wire n_8299;
wire n_1848;
wire n_9131;
wire n_1172;
wire n_13286;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_9060;
wire n_9792;
wire n_15826;
wire n_3581;
wire n_8110;
wire n_5072;
wire n_8529;
wire n_3778;
wire n_14204;
wire n_13384;
wire n_11325;
wire n_10801;
wire n_6769;
wire n_10325;
wire n_16301;
wire n_13013;
wire n_6844;
wire n_4322;
wire n_6361;
wire n_8951;
wire n_2260;
wire n_323;
wire n_1660;
wire n_1315;
wire n_11217;
wire n_15744;
wire n_4080;
wire n_2206;
wire n_997;
wire n_635;
wire n_13582;
wire n_12752;
wire n_10327;
wire n_8700;
wire n_6766;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_5940;
wire n_3001;
wire n_14157;
wire n_5260;
wire n_6751;
wire n_4981;
wire n_11651;
wire n_6232;
wire n_2347;
wire n_13255;
wire n_4676;
wire n_2657;
wire n_15144;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_7802;
wire n_10505;
wire n_7519;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_12979;
wire n_14140;
wire n_2362;
wire n_7457;
wire n_14723;
wire n_11196;
wire n_5372;
wire n_6736;
wire n_4507;
wire n_14933;
wire n_4756;
wire n_15851;
wire n_1576;
wire n_5860;
wire n_15262;
wire n_11672;
wire n_11557;
wire n_9982;
wire n_2422;
wire n_11552;
wire n_6416;
wire n_654;
wire n_13682;
wire n_2933;
wire n_8468;
wire n_9031;
wire n_12715;
wire n_12910;
wire n_7515;
wire n_3387;
wire n_7639;
wire n_11084;
wire n_12787;
wire n_8933;
wire n_6214;
wire n_3952;
wire n_9006;
wire n_8636;
wire n_10408;
wire n_16345;
wire n_11442;
wire n_9221;
wire n_13424;
wire n_4365;
wire n_3584;
wire n_14102;
wire n_4349;
wire n_3446;
wire n_10514;
wire n_1059;
wire n_7049;
wire n_7884;
wire n_6945;
wire n_8378;
wire n_6143;
wire n_14603;
wire n_2736;
wire n_6491;
wire n_7749;
wire n_10091;
wire n_7592;
wire n_11195;
wire n_3825;
wire n_4198;
wire n_7172;
wire n_10562;
wire n_539;
wire n_10586;
wire n_10893;
wire n_8283;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_6225;
wire n_2532;
wire n_4373;
wire n_7914;
wire n_17017;
wire n_1866;
wire n_8860;
wire n_2664;
wire n_16243;
wire n_15052;
wire n_12401;
wire n_4154;
wire n_7344;
wire n_5859;
wire n_6447;
wire n_14104;
wire n_4390;
wire n_459;
wire n_10593;
wire n_13304;
wire n_17088;
wire n_1782;
wire n_11517;
wire n_7892;
wire n_1558;
wire n_4107;
wire n_15078;
wire n_12722;
wire n_13716;
wire n_2519;
wire n_9523;
wire n_10821;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_16608;
wire n_7325;
wire n_11918;
wire n_14561;
wire n_13460;
wire n_2360;
wire n_4453;
wire n_15484;
wire n_6219;
wire n_723;
wire n_1393;
wire n_7674;
wire n_8686;
wire n_13590;
wire n_12712;
wire n_15494;
wire n_10961;
wire n_6175;
wire n_6445;
wire n_9829;
wire n_15778;
wire n_8563;
wire n_11077;
wire n_4571;
wire n_13914;
wire n_3137;
wire n_2544;
wire n_11579;
wire n_809;
wire n_14887;
wire n_10197;
wire n_3032;
wire n_16207;
wire n_5612;
wire n_4886;
wire n_8493;
wire n_6198;
wire n_5172;
wire n_14119;
wire n_13670;
wire n_13148;
wire n_14962;
wire n_15792;
wire n_10950;
wire n_881;
wire n_1019;
wire n_1477;
wire n_6499;
wire n_9411;
wire n_1982;
wire n_12209;
wire n_7983;
wire n_641;
wire n_5311;
wire n_8765;
wire n_14168;
wire n_14494;
wire n_15946;
wire n_910;
wire n_13452;
wire n_290;
wire n_16397;
wire n_14506;
wire n_5164;
wire n_11640;
wire n_13688;
wire n_4964;
wire n_10180;
wire n_9153;
wire n_4700;
wire n_6842;
wire n_4002;
wire n_217;
wire n_10079;
wire n_7361;
wire n_14825;
wire n_1114;
wire n_11656;
wire n_1742;
wire n_4679;
wire n_6397;
wire n_3815;
wire n_6827;
wire n_201;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_11845;
wire n_1199;
wire n_11679;
wire n_14007;
wire n_13671;
wire n_1273;
wire n_2982;
wire n_15839;
wire n_8653;
wire n_17058;
wire n_5495;
wire n_6281;
wire n_13005;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_13313;
wire n_15884;
wire n_5547;
wire n_4693;
wire n_10361;
wire n_15708;
wire n_14154;
wire n_16454;
wire n_11635;
wire n_8601;
wire n_1043;
wire n_9675;
wire n_6822;
wire n_5121;
wire n_4956;
wire n_255;
wire n_2869;
wire n_8333;
wire n_9571;
wire n_9097;
wire n_12323;
wire n_12835;
wire n_5379;
wire n_7079;
wire n_15703;
wire n_16503;
wire n_4487;
wire n_5878;
wire n_10075;
wire n_11572;
wire n_9789;
wire n_2674;
wire n_16694;
wire n_13387;
wire n_5820;
wire n_13068;
wire n_16893;
wire n_11529;
wire n_17045;
wire n_9925;
wire n_1737;
wire n_7309;
wire n_7119;
wire n_1613;
wire n_15139;
wire n_14426;
wire n_3026;
wire n_7184;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_7696;
wire n_4010;
wire n_4501;
wire n_16653;
wire n_4808;
wire n_13173;
wire n_10012;
wire n_3902;
wire n_14351;
wire n_196;
wire n_14957;
wire n_12873;
wire n_12830;
wire n_12015;
wire n_12348;
wire n_12767;
wire n_3244;
wire n_10939;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_11384;
wire n_10008;
wire n_14382;
wire n_9511;
wire n_15992;
wire n_9795;
wire n_16538;
wire n_3196;
wire n_231;
wire n_16834;
wire n_11134;
wire n_16386;
wire n_8708;
wire n_10503;
wire n_5964;
wire n_2673;
wire n_6076;
wire n_10982;
wire n_10798;
wire n_11630;
wire n_4678;
wire n_664;
wire n_1591;
wire n_12867;
wire n_13479;
wire n_13710;
wire n_5301;
wire n_13203;
wire n_13263;
wire n_14700;
wire n_5126;
wire n_13211;
wire n_8659;
wire n_15469;
wire n_8759;
wire n_6732;
wire n_16937;
wire n_2548;
wire n_3488;
wire n_9622;
wire n_2381;
wire n_12198;
wire n_9761;
wire n_14707;
wire n_2744;
wire n_6817;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_1280;
wire n_15408;
wire n_544;
wire n_7646;
wire n_14249;
wire n_9954;
wire n_14530;
wire n_3779;
wire n_599;
wire n_14870;
wire n_13848;
wire n_6982;
wire n_12617;
wire n_15184;
wire n_537;
wire n_1063;
wire n_7291;
wire n_10669;
wire n_8790;
wire n_991;
wire n_2275;
wire n_13052;
wire n_8832;
wire n_7435;
wire n_4606;
wire n_13282;
wire n_7668;
wire n_17090;
wire n_8305;
wire n_14999;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_938;
wire n_1891;
wire n_8453;
wire n_15800;
wire n_6560;
wire n_6634;
wire n_14275;
wire n_5348;
wire n_583;
wire n_12666;
wire n_9847;
wire n_16564;
wire n_13818;
wire n_1000;
wire n_313;
wire n_4868;
wire n_7017;
wire n_13846;
wire n_378;
wire n_12845;
wire n_16649;
wire n_15961;
wire n_11617;
wire n_4072;
wire n_7848;
wire n_2792;
wire n_13312;
wire n_4465;
wire n_14969;
wire n_9640;
wire n_13565;
wire n_8127;
wire n_2596;
wire n_5217;
wire n_15764;
wire n_8337;
wire n_9115;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_12047;
wire n_7861;
wire n_10190;
wire n_12411;
wire n_9534;
wire n_472;
wire n_15274;
wire n_4026;
wire n_13788;
wire n_4245;
wire n_11422;
wire n_5520;
wire n_2524;
wire n_7889;
wire n_13295;
wire n_208;
wire n_3894;
wire n_1702;
wire n_12594;
wire n_10542;
wire n_14349;
wire n_5909;
wire n_16127;
wire n_4852;
wire n_275;
wire n_7554;
wire n_3202;
wire n_11289;
wire n_16550;
wire n_8508;
wire n_4290;
wire n_4945;
wire n_11376;
wire n_5750;
wire n_7648;
wire n_8968;
wire n_147;
wire n_1232;
wire n_1211;
wire n_996;
wire n_10752;
wire n_1082;
wire n_1725;
wire n_5654;
wire n_11157;
wire n_2318;
wire n_16178;
wire n_14718;
wire n_14819;
wire n_866;
wire n_10868;
wire n_11013;
wire n_2819;
wire n_1722;
wire n_9594;
wire n_11017;
wire n_2229;
wire n_7653;
wire n_11765;
wire n_6400;
wire n_12885;
wire n_1644;
wire n_11307;
wire n_7846;
wire n_4014;
wire n_3547;
wire n_2551;
wire n_8347;
wire n_2255;
wire n_5554;
wire n_9503;
wire n_1252;
wire n_12811;
wire n_3045;
wire n_9919;
wire n_250;
wire n_15596;
wire n_13346;
wire n_773;
wire n_13331;
wire n_16845;
wire n_5135;
wire n_16071;
wire n_15605;
wire n_7551;
wire n_11793;
wire n_11574;
wire n_4599;
wire n_13307;
wire n_2706;
wire n_4222;
wire n_6655;
wire n_10017;
wire n_13574;
wire n_718;
wire n_12073;
wire n_1434;
wire n_8093;
wire n_8899;
wire n_9385;
wire n_13027;
wire n_1905;
wire n_12913;
wire n_1569;
wire n_14563;
wire n_5448;
wire n_14357;
wire n_2573;
wire n_15104;
wire n_7737;
wire n_6480;
wire n_5837;
wire n_11836;
wire n_2336;
wire n_5412;
wire n_523;
wire n_1662;
wire n_8481;
wire n_14169;
wire n_3249;
wire n_15456;
wire n_15971;
wire n_16880;
wire n_3483;
wire n_11747;
wire n_6621;
wire n_4046;
wire n_6851;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_7606;
wire n_9963;
wire n_7420;
wire n_10572;
wire n_11193;
wire n_9885;
wire n_8115;
wire n_4869;
wire n_15914;
wire n_13939;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_11670;
wire n_16954;
wire n_1244;
wire n_1796;
wire n_14042;
wire n_484;
wire n_10642;
wire n_2719;
wire n_10115;
wire n_10517;
wire n_14429;
wire n_14098;
wire n_13289;
wire n_10247;
wire n_2876;
wire n_13851;
wire n_16749;
wire n_13852;
wire n_4063;
wire n_17102;
wire n_5224;
wire n_2778;
wire n_12585;
wire n_12451;
wire n_12029;
wire n_12963;
wire n_13616;
wire n_6226;
wire n_14490;
wire n_16769;
wire n_16982;
wire n_9827;
wire n_1574;
wire n_12169;
wire n_14748;
wire n_3033;
wire n_12801;
wire n_893;
wire n_9182;
wire n_10620;
wire n_17175;
wire n_1582;
wire n_9426;
wire n_8182;
wire n_9293;
wire n_1981;
wire n_2824;
wire n_10065;
wire n_15318;
wire n_7973;
wire n_7545;
wire n_5327;
wire n_4417;
wire n_796;
wire n_11762;
wire n_14030;
wire n_14500;
wire n_531;
wire n_1374;
wire n_16636;
wire n_2089;
wire n_7896;
wire n_6283;
wire n_16955;
wire n_17146;
wire n_4688;
wire n_7156;
wire n_4939;
wire n_9581;
wire n_5900;
wire n_12657;
wire n_8629;
wire n_8186;
wire n_7319;
wire n_15721;
wire n_1486;
wire n_11758;
wire n_15082;
wire n_3619;
wire n_6158;
wire n_13366;
wire n_9400;
wire n_4013;
wire n_15028;
wire n_10744;
wire n_3434;
wire n_9246;
wire n_4342;
wire n_691;
wire n_6819;
wire n_4903;
wire n_6122;
wire n_16977;
wire n_2131;
wire n_3853;
wire n_17004;
wire n_8233;
wire n_4382;
wire n_2509;
wire n_423;
wire n_4085;
wire n_6898;
wire n_14734;
wire n_14814;
wire n_6570;
wire n_5486;
wire n_2135;
wire n_9445;
wire n_8282;
wire n_7260;
wire n_6894;
wire n_4475;
wire n_6843;
wire n_5432;
wire n_5851;
wire n_7516;
wire n_14838;
wire n_15620;
wire n_6317;
wire n_6928;
wire n_10609;
wire n_15449;
wire n_13860;
wire n_16905;
wire n_11958;
wire n_6707;
wire n_10009;
wire n_16717;
wire n_13847;
wire n_7244;
wire n_16569;
wire n_187;
wire n_11314;
wire n_16293;
wire n_1463;
wire n_4626;
wire n_12210;
wire n_10072;
wire n_12443;
wire n_12699;
wire n_7625;
wire n_8750;
wire n_10130;
wire n_4997;
wire n_8183;
wire n_13657;
wire n_5065;
wire n_13450;
wire n_9104;
wire n_6806;
wire n_15752;
wire n_924;
wire n_10956;
wire n_15389;
wire n_7991;
wire n_781;
wire n_9542;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_8637;
wire n_11515;
wire n_11490;
wire n_16486;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_8792;
wire n_6835;
wire n_7286;
wire n_2436;
wire n_3517;
wire n_13610;
wire n_15813;
wire n_6269;
wire n_7857;
wire n_13871;
wire n_7970;
wire n_16021;
wire n_9302;
wire n_1706;
wire n_2461;
wire n_10829;
wire n_8258;
wire n_3719;
wire n_16840;
wire n_11356;
wire n_7154;
wire n_524;
wire n_12781;
wire n_15991;
wire n_634;
wire n_1214;
wire n_16753;
wire n_10506;
wire n_3526;
wire n_3888;
wire n_12573;
wire n_9960;
wire n_14843;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_8416;
wire n_8390;
wire n_13881;
wire n_6248;
wire n_11678;
wire n_12744;
wire n_6088;
wire n_10236;
wire n_11374;
wire n_14519;
wire n_1181;
wire n_1999;
wire n_11176;
wire n_7194;
wire n_16072;
wire n_4841;
wire n_11402;
wire n_4683;
wire n_5173;
wire n_11162;
wire n_2873;
wire n_10002;
wire n_8696;
wire n_9185;
wire n_9601;
wire n_13137;
wire n_2084;
wire n_15698;
wire n_13226;
wire n_3330;
wire n_3514;
wire n_11771;
wire n_15951;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_5855;
wire n_13431;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_7163;
wire n_14402;
wire n_14845;
wire n_14507;
wire n_14020;
wire n_3797;
wire n_1836;
wire n_13552;
wire n_13164;
wire n_7027;
wire n_3416;
wire n_8552;
wire n_12006;
wire n_4600;
wire n_5861;
wire n_1453;
wire n_6964;
wire n_3943;
wire n_10855;
wire n_3145;
wire n_14389;
wire n_7964;
wire n_5749;
wire n_6320;
wire n_9403;
wire n_14558;
wire n_16716;
wire n_11322;
wire n_16680;
wire n_6316;
wire n_8619;
wire n_419;
wire n_7068;
wire n_11484;
wire n_9972;
wire n_11711;
wire n_13227;
wire n_2908;
wire n_8594;
wire n_9878;
wire n_14541;
wire n_10139;
wire n_14183;
wire n_270;
wire n_4106;
wire n_9541;
wire n_16055;
wire n_10941;
wire n_14689;
wire n_285;
wire n_2156;
wire n_15667;
wire n_12548;
wire n_1184;
wire n_17084;
wire n_16797;
wire n_202;
wire n_8162;
wire n_9735;
wire n_754;
wire n_9576;
wire n_14528;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_7327;
wire n_16190;
wire n_12727;
wire n_15588;
wire n_1277;
wire n_1746;
wire n_12240;
wire n_13045;
wire n_13620;
wire n_6610;
wire n_1062;
wire n_15919;
wire n_5998;
wire n_8318;
wire n_14742;
wire n_4702;
wire n_5102;
wire n_16376;
wire n_9974;
wire n_4954;
wire n_15707;
wire n_740;
wire n_10992;
wire n_167;
wire n_16889;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_8425;
wire n_6752;
wire n_16281;
wire n_13001;
wire n_6959;
wire n_9704;
wire n_6250;
wire n_13919;
wire n_11392;
wire n_12372;
wire n_3283;
wire n_11803;
wire n_15597;
wire n_17034;
wire n_259;
wire n_4331;
wire n_7317;
wire n_4159;
wire n_16458;
wire n_11912;
wire n_13862;
wire n_15066;
wire n_13784;
wire n_7864;
wire n_11139;
wire n_3451;
wire n_10650;
wire n_8051;
wire n_4734;
wire n_11021;
wire n_6675;
wire n_15204;
wire n_7955;
wire n_2832;
wire n_1688;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_9039;
wire n_12914;
wire n_16141;
wire n_16919;
wire n_7384;
wire n_12844;
wire n_267;
wire n_2914;
wire n_5656;
wire n_7218;
wire n_1988;
wire n_12952;
wire n_15996;
wire n_5678;
wire n_6561;
wire n_11379;
wire n_6858;
wire n_16381;
wire n_5865;
wire n_6050;
wire n_13271;
wire n_7512;
wire n_1718;
wire n_7814;
wire n_12276;
wire n_12096;
wire n_8389;
wire n_4515;
wire n_10417;
wire n_2149;
wire n_2277;
wire n_200;
wire n_10029;
wire n_12150;
wire n_16507;
wire n_16873;
wire n_14271;
wire n_16664;
wire n_13595;
wire n_2539;
wire n_8620;
wire n_10125;
wire n_5555;
wire n_13757;
wire n_15711;
wire n_2078;
wire n_8886;
wire n_1145;
wire n_4809;
wire n_7152;
wire n_14770;
wire n_787;
wire n_4012;
wire n_10253;
wire n_11899;
wire n_16051;
wire n_16829;
wire n_1195;
wire n_15533;
wire n_13761;
wire n_15705;
wire n_15574;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_13136;
wire n_13190;
wire n_6823;
wire n_10693;
wire n_3606;
wire n_14461;
wire n_7062;
wire n_7090;
wire n_12449;
wire n_15261;
wire n_8202;
wire n_13633;
wire n_2232;
wire n_11966;
wire n_1847;
wire n_14205;
wire n_5815;
wire n_4320;
wire n_12118;
wire n_10599;
wire n_5084;
wire n_7223;
wire n_14266;
wire n_12770;
wire n_5251;
wire n_15014;
wire n_1314;
wire n_8755;
wire n_13174;
wire n_16028;
wire n_1512;
wire n_8668;
wire n_5965;
wire n_16748;
wire n_884;
wire n_4980;
wire n_3324;
wire n_10977;
wire n_13528;
wire n_2192;
wire n_6796;
wire n_8979;
wire n_5407;
wire n_2988;
wire n_12814;
wire n_11553;
wire n_4560;
wire n_14064;
wire n_14322;
wire n_13220;
wire n_12009;
wire n_15550;
wire n_13456;
wire n_13916;
wire n_7761;
wire n_10947;
wire n_8141;
wire n_10386;
wire n_3793;
wire n_3230;
wire n_859;
wire n_5042;
wire n_8199;
wire n_16918;
wire n_12826;
wire n_7055;
wire n_6024;
wire n_4768;
wire n_1889;
wire n_10267;
wire n_16953;
wire n_6090;
wire n_693;
wire n_5368;
wire n_929;
wire n_10401;
wire n_3207;
wire n_3641;
wire n_16707;
wire n_16674;
wire n_3828;
wire n_16773;
wire n_15666;
wire n_15511;
wire n_16160;
wire n_15171;
wire n_15933;
wire n_16973;
wire n_1850;
wire n_3183;
wire n_11127;
wire n_9908;
wire n_11926;
wire n_8004;
wire n_8383;
wire n_14763;
wire n_3607;
wire n_1637;
wire n_9688;
wire n_9864;
wire n_2427;
wire n_12144;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_7388;
wire n_1751;
wire n_7056;
wire n_10428;
wire n_14585;
wire n_10212;
wire n_7437;
wire n_11460;
wire n_6489;
wire n_11486;
wire n_9023;
wire n_16491;
wire n_5310;
wire n_2769;
wire n_8895;
wire n_438;
wire n_8680;
wire n_1548;
wire n_14208;
wire n_4987;
wire n_6714;
wire n_8394;
wire n_440;
wire n_10539;
wire n_14152;
wire n_7849;
wire n_7726;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_7417;
wire n_2739;
wire n_12937;
wire n_3962;
wire n_11148;
wire n_7446;
wire n_12312;
wire n_6038;
wire n_10728;
wire n_15109;
wire n_2902;
wire n_6030;
wire n_6620;
wire n_4360;
wire n_1544;
wire n_6791;
wire n_6245;
wire n_4540;
wire n_9220;
wire n_13929;
wire n_16676;
wire n_6821;
wire n_9317;
wire n_12580;
wire n_13965;
wire n_2094;
wire n_13796;
wire n_5588;
wire n_3854;
wire n_8198;
wire n_17130;
wire n_9993;
wire n_1354;
wire n_10879;
wire n_13474;
wire n_8665;
wire n_12393;
wire n_16168;
wire n_6583;
wire n_10545;
wire n_2349;
wire n_3652;
wire n_12201;
wire n_7859;
wire n_16755;
wire n_3449;
wire n_13240;
wire n_1021;
wire n_13187;
wire n_13594;
wire n_3089;
wire n_4854;
wire n_9561;
wire n_491;
wire n_10516;
wire n_14640;
wire n_9444;
wire n_1595;
wire n_8017;
wire n_1142;
wire n_10497;
wire n_16131;
wire n_11675;
wire n_5477;
wire n_260;
wire n_17134;
wire n_2727;
wire n_942;
wire n_10705;
wire n_7523;
wire n_12082;
wire n_13966;
wire n_14936;
wire n_11032;
wire n_5234;
wire n_14035;
wire n_12322;
wire n_1416;
wire n_6890;
wire n_10432;
wire n_11454;
wire n_9184;
wire n_7559;
wire n_14345;
wire n_9037;
wire n_16974;
wire n_7576;
wire n_6988;
wire n_10779;
wire n_8303;
wire n_11554;
wire n_1599;
wire n_5871;
wire n_11988;
wire n_13981;
wire n_4747;
wire n_14647;
wire n_16162;
wire n_8000;
wire n_11197;
wire n_14286;
wire n_3472;
wire n_14686;
wire n_16542;
wire n_2527;
wire n_6052;
wire n_7769;
wire n_15172;
wire n_15305;
wire n_11416;
wire n_9505;
wire n_9193;
wire n_14360;
wire n_7257;
wire n_3126;
wire n_12986;
wire n_15179;
wire n_2759;
wire n_6973;
wire n_10869;
wire n_8852;
wire n_5007;
wire n_17062;
wire n_8709;
wire n_4881;
wire n_10314;
wire n_2038;
wire n_10504;
wire n_6488;
wire n_3958;
wire n_4495;
wire n_10687;
wire n_13691;
wire n_16945;
wire n_4737;
wire n_1838;
wire n_9218;
wire n_9755;
wire n_4357;
wire n_11341;
wire n_7729;
wire n_2806;
wire n_4502;
wire n_11045;
wire n_287;
wire n_3191;
wire n_1716;
wire n_12373;
wire n_302;
wire n_12741;
wire n_7005;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_15544;
wire n_8782;
wire n_7081;
wire n_10882;
wire n_7742;
wire n_5253;
wire n_10293;
wire n_3588;
wire n_355;
wire n_6280;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_16897;
wire n_16942;
wire n_5274;
wire n_6399;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_14828;
wire n_1819;
wire n_15152;
wire n_9506;
wire n_9162;
wire n_13629;
wire n_3095;
wire n_15264;
wire n_15584;
wire n_947;
wire n_7341;
wire n_5792;
wire n_13155;
wire n_14581;
wire n_3698;
wire n_15493;
wire n_4513;
wire n_1179;
wire n_11569;
wire n_468;
wire n_13152;
wire n_10256;
wire n_182;
wire n_696;
wire n_1442;
wire n_4775;
wire n_6256;
wire n_482;
wire n_2620;
wire n_1833;
wire n_8716;
wire n_12412;
wire n_1691;
wire n_12677;
wire n_7264;
wire n_8250;
wire n_7842;
wire n_15976;
wire n_16142;
wire n_14315;
wire n_12181;
wire n_12833;
wire n_2499;
wire n_2549;
wire n_10298;
wire n_9415;
wire n_12631;
wire n_12115;
wire n_14829;
wire n_6648;
wire n_16091;
wire n_7492;
wire n_13194;
wire n_15331;
wire n_13546;
wire n_804;
wire n_6649;
wire n_8714;
wire n_1656;
wire n_8357;
wire n_12567;
wire n_15424;
wire n_1382;
wire n_3093;
wire n_12175;
wire n_15791;
wire n_2970;
wire n_14920;
wire n_9990;
wire n_6910;
wire n_3885;
wire n_955;
wire n_15687;
wire n_8466;
wire n_4264;
wire n_5954;
wire n_10326;
wire n_9015;
wire n_14827;
wire n_2166;
wire n_13446;
wire n_15482;
wire n_10235;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_514;
wire n_6431;
wire n_418;
wire n_8589;
wire n_12754;
wire n_3250;
wire n_4223;
wire n_14141;
wire n_12455;
wire n_3538;
wire n_13363;
wire n_3915;
wire n_11990;
wire n_8266;
wire n_3839;
wire n_8587;
wire n_7285;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_6324;
wire n_5489;
wire n_3407;
wire n_10725;
wire n_15653;
wire n_10274;
wire n_13728;
wire n_13601;
wire n_3875;
wire n_4029;
wire n_8876;
wire n_11541;
wire n_9214;
wire n_14780;
wire n_4206;
wire n_12340;
wire n_2415;
wire n_4099;
wire n_10799;
wire n_8922;
wire n_11680;
wire n_10090;
wire n_3120;
wire n_6512;
wire n_12686;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_9070;
wire n_15993;
wire n_16709;
wire n_8498;
wire n_4794;
wire n_9933;
wire n_4843;
wire n_12734;
wire n_669;
wire n_5580;
wire n_15108;
wire n_5215;
wire n_15870;
wire n_337;
wire n_437;
wire n_12331;
wire n_3937;
wire n_4763;
wire n_10874;
wire n_9339;
wire n_11596;
wire n_1418;
wire n_9991;
wire n_12880;
wire n_9486;
wire n_8457;
wire n_6243;
wire n_14113;
wire n_5795;
wire n_10763;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_12425;
wire n_8267;
wire n_12184;
wire n_10266;
wire n_2462;
wire n_13918;
wire n_14997;
wire n_7051;
wire n_11180;
wire n_6773;
wire n_16814;
wire n_10290;
wire n_2155;
wire n_6231;
wire n_15758;
wire n_12472;
wire n_615;
wire n_13048;
wire n_12266;
wire n_7503;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_12432;
wire n_517;
wire n_8124;
wire n_3604;
wire n_8545;
wire n_5430;
wire n_16890;
wire n_6041;
wire n_8526;
wire n_824;
wire n_12300;
wire n_159;
wire n_13593;
wire n_8319;
wire n_7997;
wire n_12527;
wire n_5659;
wire n_11839;
wire n_16510;
wire n_9279;
wire n_6859;
wire n_7716;
wire n_4272;
wire n_10732;
wire n_5195;
wire n_12110;
wire n_15354;
wire n_16851;
wire n_15310;
wire n_13744;
wire n_3176;
wire n_9790;
wire n_144;
wire n_11404;
wire n_3792;
wire n_7950;
wire n_11548;
wire n_6323;
wire n_13515;
wire n_5720;
wire n_4267;
wire n_8581;
wire n_12122;
wire n_14889;
wire n_10873;
wire n_16026;
wire n_8214;
wire n_15583;
wire n_7793;
wire n_9053;
wire n_16337;
wire n_8516;
wire n_2083;
wire n_815;
wire n_12310;
wire n_5598;
wire n_2753;
wire n_1340;
wire n_470;
wire n_11343;
wire n_3021;
wire n_8989;
wire n_13028;
wire n_7746;
wire n_477;
wire n_11362;
wire n_15941;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_11007;
wire n_3950;
wire n_7570;
wire n_9650;
wire n_16119;
wire n_9880;
wire n_11497;
wire n_2898;
wire n_1825;
wire n_15859;
wire n_16504;
wire n_10720;
wire n_6912;
wire n_3567;
wire n_14574;
wire n_7425;
wire n_15050;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_16693;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_14014;
wire n_12827;
wire n_14078;
wire n_10220;
wire n_9217;
wire n_9499;
wire n_5783;
wire n_7829;
wire n_6837;
wire n_15696;
wire n_13467;
wire n_13245;
wire n_6747;
wire n_2903;
wire n_5303;
wire n_10081;
wire n_12804;
wire n_3812;
wire n_3127;
wire n_9282;
wire n_1731;
wire n_799;
wire n_10145;
wire n_11347;
wire n_1147;
wire n_12892;
wire n_6916;
wire n_7894;
wire n_8262;
wire n_2378;
wire n_10167;
wire n_5530;
wire n_7957;
wire n_16440;
wire n_12656;
wire n_6718;
wire n_8289;
wire n_965;
wire n_13804;
wire n_5809;
wire n_10447;
wire n_12418;
wire n_934;
wire n_2213;
wire n_7121;
wire n_7531;
wire n_6410;
wire n_12448;
wire n_15180;
wire n_12219;
wire n_12729;
wire n_356;
wire n_13549;
wire n_13921;
wire n_6473;
wire n_8087;
wire n_4056;
wire n_10238;
wire n_13345;
wire n_4806;
wire n_11029;
wire n_7961;
wire n_1674;
wire n_9920;
wire n_5993;
wire n_4015;
wire n_15129;
wire n_6574;
wire n_2924;
wire n_6492;
wire n_4445;
wire n_7687;
wire n_9948;
wire n_4462;
wire n_5299;
wire n_13216;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_11226;
wire n_2142;
wire n_8863;
wire n_9371;
wire n_15396;
wire n_4517;
wire n_2896;
wire n_8701;
wire n_1913;
wire n_2069;
wire n_15551;
wire n_4043;
wire n_13036;
wire n_15603;
wire n_1042;
wire n_3170;
wire n_9237;
wire n_15038;
wire n_2311;
wire n_13398;
wire n_6857;
wire n_8705;
wire n_14148;
wire n_1455;
wire n_2287;
wire n_9815;
wire n_836;
wire n_3415;
wire n_16309;
wire n_10292;
wire n_12644;
wire n_6975;
wire n_15413;
wire n_10820;
wire n_7763;
wire n_13258;
wire n_16681;
wire n_3464;
wire n_6290;
wire n_3414;
wire n_6646;
wire n_16423;
wire n_205;
wire n_7703;
wire n_11760;
wire n_15781;
wire n_13827;
wire n_7928;
wire n_4234;
wire n_10395;
wire n_760;
wire n_1483;
wire n_12576;
wire n_10168;
wire n_14350;
wire n_1363;
wire n_8722;
wire n_1111;
wire n_970;
wire n_3467;
wire n_5821;
wire n_11664;
wire n_713;
wire n_3179;
wire n_15306;
wire n_598;
wire n_12187;
wire n_6622;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_7665;
wire n_5262;
wire n_7677;
wire n_13169;
wire n_14782;
wire n_15978;
wire n_16887;
wire n_3262;
wire n_10366;
wire n_5319;
wire n_10287;
wire n_14017;
wire n_15358;
wire n_927;
wire n_13940;
wire n_7469;
wire n_261;
wire n_3699;
wire n_16584;
wire n_10163;
wire n_6118;
wire n_706;
wire n_2120;
wire n_7125;
wire n_7856;
wire n_6028;
wire n_6663;
wire n_14145;
wire n_11006;
wire n_6532;
wire n_1419;
wire n_13406;
wire n_10431;
wire n_8622;
wire n_3816;
wire n_8099;
wire n_8729;
wire n_9479;
wire n_10876;
wire n_11485;
wire n_3528;
wire n_15092;
wire n_6267;
wire n_15397;
wire n_6682;
wire n_9480;
wire n_12453;
wire n_12593;
wire n_4207;
wire n_11449;
wire n_8085;
wire n_15984;
wire n_2404;
wire n_2757;
wire n_2168;
wire n_4725;
wire n_9597;
wire n_10614;
wire n_10786;
wire n_13873;
wire n_13335;
wire n_14273;
wire n_348;
wire n_10352;
wire n_9173;
wire n_15458;
wire n_16067;
wire n_2312;
wire n_7203;
wire n_9641;
wire n_8947;
wire n_13714;
wire n_7797;
wire n_1826;
wire n_9983;
wire n_9267;
wire n_14565;
wire n_5943;
wire n_6556;
wire n_10039;
wire n_15079;
wire n_4880;
wire n_15784;
wire n_2834;
wire n_4051;
wire n_13070;
wire n_6216;
wire n_13866;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_637;
wire n_15231;
wire n_9849;
wire n_15454;
wire n_11831;
wire n_7128;
wire n_5335;
wire n_1259;
wire n_6365;
wire n_8459;
wire n_7111;
wire n_2801;
wire n_11096;
wire n_1177;
wire n_4334;
wire n_8478;
wire n_5284;
wire n_12288;
wire n_8786;
wire n_16553;
wire n_16665;
wire n_9414;
wire n_4978;
wire n_11677;
wire n_13025;
wire n_14256;
wire n_5771;
wire n_3246;
wire n_9419;
wire n_3299;
wire n_8887;
wire n_980;
wire n_1618;
wire n_1869;
wire n_12091;
wire n_3623;
wire n_905;
wire n_2718;
wire n_14922;
wire n_11898;
wire n_4707;
wire n_14749;
wire n_2687;
wire n_8851;
wire n_6950;
wire n_4923;
wire n_4911;
wire n_15168;
wire n_15716;
wire n_3876;
wire n_8540;
wire n_5516;
wire n_7284;
wire n_3615;
wire n_8276;
wire n_7057;
wire n_16546;
wire n_1802;
wire n_14862;
wire n_13457;
wire n_9823;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_9152;
wire n_15915;
wire n_8706;
wire n_3200;
wire n_6167;
wire n_12357;
wire n_3642;
wire n_145;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_7064;
wire n_11826;
wire n_12629;
wire n_8532;
wire n_9533;
wire n_10750;
wire n_5433;
wire n_3682;
wire n_11825;
wire n_5429;
wire n_7278;
wire n_12893;
wire n_9281;
wire n_9103;
wire n_9111;
wire n_6772;
wire n_15499;
wire n_7088;
wire n_7799;
wire n_9618;
wire n_10383;
wire n_16134;
wire n_5698;
wire n_10856;
wire n_5731;
wire n_14532;
wire n_14105;
wire n_10883;
wire n_12935;
wire n_8871;
wire n_4007;
wire n_1456;
wire n_8433;
wire n_9065;
wire n_10429;
wire n_14627;
wire n_15552;
wire n_14463;
wire n_1879;
wire n_15727;
wire n_14735;
wire n_17124;
wire n_15808;
wire n_15103;
wire n_6159;
wire n_2129;
wire n_5857;
wire n_12732;
wire n_7048;
wire n_7979;
wire n_12569;
wire n_9674;
wire n_16673;
wire n_6617;
wire n_16629;
wire n_16885;
wire n_553;
wire n_7725;
wire n_13547;
wire n_814;
wire n_578;
wire n_10859;
wire n_5120;
wire n_3572;
wire n_8371;
wire n_16756;
wire n_2975;
wire n_2399;
wire n_8547;
wire n_11538;
wire n_10815;
wire n_16558;
wire n_17059;
wire n_1134;
wire n_11008;
wire n_4075;
wire n_3471;
wire n_1484;
wire n_8467;
wire n_12980;
wire n_647;
wire n_11093;
wire n_11585;
wire n_2932;
wire n_2027;
wire n_16205;
wire n_8409;
wire n_6217;
wire n_600;
wire n_3118;
wire n_11616;
wire n_10303;
wire n_9157;
wire n_5560;
wire n_16093;
wire n_15071;
wire n_14831;
wire n_16396;
wire n_9170;
wire n_4441;
wire n_10424;
wire n_16445;
wire n_3922;
wire n_3039;
wire n_2195;
wire n_5455;
wire n_502;
wire n_8640;
wire n_11001;
wire n_15500;
wire n_16303;
wire n_6777;
wire n_10196;
wire n_16522;
wire n_16951;
wire n_15543;
wire n_6742;
wire n_16444;
wire n_14823;
wire n_1467;
wire n_7447;
wire n_5209;
wire n_15807;
wire n_10684;
wire n_247;
wire n_13154;
wire n_6307;
wire n_5704;
wire n_14129;
wire n_16074;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_8431;
wire n_16049;
wire n_14547;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_13280;
wire n_3618;
wire n_5916;
wire n_8415;
wire n_10184;
wire n_3705;
wire n_3022;
wire n_13904;
wire n_10421;
wire n_13944;
wire n_15935;
wire n_13359;
wire n_1709;
wire n_6479;
wire n_11472;
wire n_14376;
wire n_13855;
wire n_13073;
wire n_5099;
wire n_11063;
wire n_681;
wire n_3286;
wire n_5781;
wire n_11179;
wire n_5619;
wire n_2023;
wire n_14777;
wire n_9416;
wire n_11885;
wire n_3974;
wire n_9368;
wire n_7365;
wire n_3443;
wire n_16644;
wire n_8329;
wire n_13083;
wire n_14201;
wire n_2599;
wire n_3988;
wire n_7792;
wire n_5022;
wire n_8089;
wire n_9208;
wire n_11657;
wire n_6370;
wire n_13124;
wire n_9223;
wire n_16327;
wire n_2075;
wire n_13771;
wire n_1726;
wire n_10329;
wire n_10924;
wire n_13845;
wire n_11921;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_15443;
wire n_14224;
wire n_10285;
wire n_16349;
wire n_7275;
wire n_15039;
wire n_5353;
wire n_4771;
wire n_12099;
wire n_2853;
wire n_14991;
wire n_3350;
wire n_6856;
wire n_1098;
wire n_9781;
wire n_3009;
wire n_13609;
wire n_13572;
wire n_13817;
wire n_8633;
wire n_12897;
wire n_777;
wire n_7095;
wire n_9392;
wire n_7390;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_9422;
wire n_920;
wire n_15338;
wire n_8541;
wire n_10084;
wire n_12924;
wire n_17148;
wire n_8762;
wire n_15866;
wire n_14162;
wire n_12619;
wire n_16930;
wire n_12541;
wire n_3951;
wire n_5518;
wire n_9970;
wire n_3035;
wire n_14882;
wire n_13428;
wire n_15880;
wire n_4261;
wire n_15488;
wire n_15508;
wire n_7037;
wire n_13104;
wire n_17133;
wire n_15292;
wire n_1132;
wire n_9338;
wire n_15176;
wire n_11647;
wire n_8125;
wire n_501;
wire n_1823;
wire n_6240;
wire n_15222;
wire n_5236;
wire n_4236;
wire n_10077;
wire n_3942;
wire n_3023;
wire n_10964;
wire n_14566;
wire n_9492;
wire n_2254;
wire n_3290;
wire n_14367;
wire n_6693;
wire n_15694;
wire n_10759;
wire n_9226;
wire n_6712;
wire n_10129;
wire n_16475;
wire n_10101;
wire n_1402;
wire n_7530;
wire n_3957;
wire n_13844;
wire n_11757;
wire n_3418;
wire n_10566;
wire n_1607;
wire n_7471;
wire n_9328;
wire n_17028;
wire n_6465;
wire n_221;
wire n_10192;
wire n_8188;
wire n_17137;
wire n_5673;
wire n_14363;
wire n_861;
wire n_16606;
wire n_11846;
wire n_11519;
wire n_16450;
wire n_14571;
wire n_8615;
wire n_16940;
wire n_5814;
wire n_16560;
wire n_1666;
wire n_6586;
wire n_7058;
wire n_14857;
wire n_5103;
wire n_17164;
wire n_4648;
wire n_8011;
wire n_12191;
wire n_10207;
wire n_2214;
wire n_11530;
wire n_6730;
wire n_17138;
wire n_13526;
wire n_13998;
wire n_6367;
wire n_2256;
wire n_8923;
wire n_11488;
wire n_281;
wire n_3326;
wire n_11389;
wire n_8624;
wire n_262;
wire n_8222;
wire n_11928;
wire n_15150;
wire n_12429;
wire n_12825;
wire n_6069;
wire n_2732;
wire n_1883;
wire n_8206;
wire n_15547;
wire n_15907;
wire n_6515;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_9513;
wire n_11315;
wire n_3224;
wire n_13267;
wire n_9393;
wire n_1969;
wire n_15249;
wire n_5671;
wire n_7429;
wire n_13506;
wire n_6940;
wire n_8065;
wire n_9914;
wire n_14833;
wire n_14398;
wire n_527;
wire n_2949;
wire n_16861;
wire n_7008;
wire n_12318;
wire n_12918;
wire n_14731;
wire n_6468;
wire n_7709;
wire n_4269;
wire n_1927;
wire n_7540;
wire n_16533;
wire n_10886;
wire n_12923;
wire n_15112;
wire n_13632;
wire n_14600;
wire n_10804;
wire n_16931;
wire n_7581;
wire n_12077;
wire n_343;
wire n_15132;
wire n_10362;
wire n_1222;
wire n_16875;
wire n_16313;
wire n_7139;
wire n_10384;
wire n_10437;
wire n_13834;
wire n_8935;
wire n_14213;
wire n_15081;
wire n_16158;
wire n_16044;
wire n_13444;
wire n_10885;
wire n_11962;
wire n_11002;
wire n_3803;
wire n_14331;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_13885;
wire n_12805;
wire n_1791;
wire n_14928;
wire n_7782;
wire n_7432;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_16620;
wire n_13067;
wire n_8155;
wire n_9334;
wire n_2449;
wire n_14059;
wire n_16565;
wire n_11648;
wire n_10093;
wire n_13924;
wire n_14289;
wire n_4428;
wire n_12808;
wire n_745;
wire n_6483;
wire n_1572;
wire n_7770;
wire n_12853;
wire n_9684;
wire n_12591;
wire n_16536;
wire n_8397;
wire n_8568;
wire n_4463;
wire n_10600;
wire n_17118;
wire n_10480;
wire n_11994;
wire n_5357;
wire n_8175;
wire n_10796;
wire n_3648;
wire n_10892;
wire n_9254;
wire n_6576;
wire n_6810;
wire n_11050;
wire n_1975;
wire n_5421;
wire n_9083;
wire n_11250;
wire n_10003;
wire n_16106;
wire n_16425;
wire n_1388;
wire n_1266;
wire n_11316;
wire n_14727;
wire n_14485;
wire n_15277;
wire n_12987;
wire n_4396;
wire n_15938;
wire n_13717;
wire n_1990;
wire n_6708;
wire n_12251;
wire n_10252;
wire n_16229;
wire n_17165;
wire n_12948;
wire n_16379;
wire n_8026;
wire n_16517;
wire n_6667;
wire n_9175;
wire n_9838;
wire n_3491;
wire n_15636;
wire n_2690;
wire n_3090;
wire n_11428;
wire n_2474;
wire n_12467;
wire n_12756;
wire n_2623;
wire n_11463;
wire n_15280;
wire n_1075;
wire n_6040;
wire n_10495;
wire n_1890;
wire n_8974;
wire n_6847;
wire n_6305;
wire n_8836;
wire n_10812;
wire n_4034;
wire n_12678;
wire n_14211;
wire n_4228;
wire n_14641;
wire n_12700;
wire n_1227;
wire n_11674;
wire n_11097;
wire n_11069;
wire n_7251;
wire n_10894;
wire n_3166;
wire n_12602;
wire n_14155;
wire n_12194;
wire n_15751;
wire n_7356;
wire n_16406;
wire n_3649;
wire n_7412;
wire n_16724;
wire n_3065;
wire n_16952;
wire n_8168;
wire n_7212;
wire n_5045;
wire n_16799;
wire n_5237;
wire n_15465;
wire n_11318;
wire n_7751;
wire n_12351;
wire n_7951;
wire n_12965;
wire n_657;
wire n_14184;
wire n_7060;
wire n_3924;
wire n_9336;
wire n_3997;
wire n_12367;
wire n_13603;
wire n_8873;
wire n_14111;
wire n_10311;
wire n_7591;
wire n_10490;
wire n_3564;
wire n_862;
wire n_5769;
wire n_2637;
wire n_7444;
wire n_10702;
wire n_6750;
wire n_15207;
wire n_7911;
wire n_3795;
wire n_7595;
wire n_4931;
wire n_2306;
wire n_7790;
wire n_11586;
wire n_2071;
wire n_7426;
wire n_11786;
wire n_430;
wire n_13571;
wire n_3953;
wire n_4400;
wire n_7502;
wire n_2414;
wire n_17066;
wire n_13492;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_10906;
wire n_1532;
wire n_6855;
wire n_10840;
wire n_10891;
wire n_14257;
wire n_15019;
wire n_8170;
wire n_1030;
wire n_5181;
wire n_6239;
wire n_10181;
wire n_3208;
wire n_13673;
wire n_12036;
wire n_9554;
wire n_14589;
wire n_15950;
wire n_16417;
wire n_5768;
wire n_1342;
wire n_11330;
wire n_6199;
wire n_16796;
wire n_2737;
wire n_3282;
wire n_8120;
wire n_12263;
wire n_9830;
wire n_9315;
wire n_9116;
wire n_8825;
wire n_14416;
wire n_852;
wire n_9169;
wire n_16776;
wire n_2916;
wire n_7252;
wire n_11201;
wire n_1060;
wire n_5963;
wire n_9999;
wire n_4424;
wire n_4351;
wire n_6543;
wire n_7532;
wire n_14899;
wire n_12703;
wire n_4192;
wire n_8003;
wire n_11979;
wire n_12253;
wire n_9215;
wire n_15380;
wire n_1748;
wire n_1301;
wire n_6789;
wire n_5972;
wire n_3400;
wire n_8395;
wire n_13986;
wire n_7065;
wire n_1466;
wire n_8083;
wire n_14963;
wire n_11888;
wire n_14596;
wire n_6177;
wire n_8057;
wire n_2581;
wire n_5937;
wire n_1783;
wire n_15902;
wire n_9259;
wire n_5146;
wire n_16366;
wire n_7367;
wire n_10755;
wire n_14274;
wire n_11835;
wire n_11537;
wire n_8164;
wire n_10525;
wire n_11583;
wire n_12776;
wire n_14714;
wire n_15897;
wire n_7405;
wire n_7267;
wire n_4646;
wire n_15069;
wire n_4221;
wire n_12445;
wire n_1037;
wire n_3650;
wire n_8877;
wire n_1329;
wire n_16477;
wire n_6825;
wire n_15282;
wire n_7614;
wire n_1993;
wire n_1545;
wire n_6460;
wire n_4035;
wire n_9150;
wire n_6952;
wire n_9595;
wire n_16385;
wire n_1480;
wire n_3670;
wire n_11420;
wire n_8366;
wire n_14907;
wire n_6173;
wire n_16588;
wire n_2540;
wire n_4190;
wire n_8476;
wire n_1605;
wire n_11527;
wire n_3060;
wire n_6218;
wire n_10435;
wire n_11048;
wire n_10342;
wire n_15133;
wire n_14584;
wire n_11933;
wire n_6486;
wire n_7685;
wire n_13826;
wire n_4009;
wire n_2984;
wire n_11900;
wire n_157;
wire n_12620;
wire n_7619;
wire n_11106;
wire n_2489;
wire n_15237;
wire n_15832;
wire n_12299;
wire n_13078;
wire n_5013;
wire n_4145;
wire n_10983;
wire n_11266;
wire n_6852;
wire n_11340;
wire n_11929;
wire n_15659;
wire n_624;
wire n_15709;
wire n_5577;
wire n_876;
wire n_12673;
wire n_13516;
wire n_9100;
wire n_5872;
wire n_7883;
wire n_13557;
wire n_10397;
wire n_15007;
wire n_15337;
wire n_6692;
wire n_13208;
wire n_9707;
wire n_5017;
wire n_16010;
wire n_8854;
wire n_736;
wire n_13523;
wire n_12834;
wire n_10202;
wire n_14549;
wire n_12821;
wire n_10677;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_7220;
wire n_7560;
wire n_1327;
wire n_10648;
wire n_1475;
wire n_2106;
wire n_9262;
wire n_5976;
wire n_4717;
wire n_9249;
wire n_6888;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_602;
wire n_14798;
wire n_11964;
wire n_12247;
wire n_15023;
wire n_17033;
wire n_13030;
wire n_854;
wire n_8256;
wire n_16643;
wire n_2091;
wire n_393;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_13065;
wire n_7270;
wire n_14751;
wire n_14217;
wire n_10273;
wire n_12927;
wire n_1658;
wire n_12324;
wire n_12817;
wire n_15627;
wire n_1072;
wire n_11255;
wire n_8621;
wire n_13753;
wire n_16511;
wire n_1305;
wire n_11751;
wire n_4750;
wire n_2348;
wire n_10978;
wire n_9806;
wire n_10834;
wire n_1873;
wire n_13430;
wire n_8577;
wire n_9019;
wire n_10097;
wire n_13880;
wire n_14796;
wire n_2667;
wire n_2725;
wire n_9361;
wire n_3746;
wire n_16828;
wire n_7731;
wire n_13050;
wire n_13175;
wire n_4537;
wire n_6626;
wire n_1046;
wire n_10890;
wire n_5838;
wire n_13732;
wire n_7034;
wire n_10816;
wire n_8654;
wire n_3694;
wire n_12887;
wire n_13133;
wire n_17087;
wire n_6854;
wire n_7940;
wire n_15496;
wire n_771;
wire n_16256;
wire n_14188;
wire n_6793;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_9814;
wire n_2307;
wire n_11930;
wire n_15361;
wire n_421;
wire n_3702;
wire n_5930;
wire n_11269;
wire n_10462;
wire n_12316;
wire n_12539;
wire n_13358;
wire n_8952;
wire n_13823;
wire n_12758;
wire n_1984;
wire n_12414;
wire n_3453;
wire n_9438;
wire n_1556;
wire n_7537;
wire n_12600;
wire n_6980;
wire n_7040;
wire n_5345;
wire n_2815;
wire n_14875;
wire n_15920;
wire n_15506;
wire n_11985;
wire n_4427;
wire n_7458;
wire n_1824;
wire n_7740;
wire n_17061;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_15572;
wire n_16689;
wire n_15149;
wire n_6794;
wire n_819;
wire n_12949;
wire n_1971;
wire n_2945;
wire n_586;
wire n_1324;
wire n_3543;
wire n_8421;
wire n_9856;
wire n_11205;
wire n_7179;
wire n_10832;
wire n_1776;
wire n_3448;
wire n_7433;
wire n_13499;
wire n_4279;
wire n_14057;
wire n_16925;
wire n_16500;
wire n_9327;
wire n_9313;
wire n_4330;
wire n_605;
wire n_2936;
wire n_3609;
wire n_6334;
wire n_13560;
wire n_6257;
wire n_16219;
wire n_10142;
wire n_4152;
wire n_6874;
wire n_14079;
wire n_14073;
wire n_10300;
wire n_15489;
wire n_8911;
wire n_15340;
wire n_16410;
wire n_5537;
wire n_9518;
wire n_2698;
wire n_5572;
wire n_15693;
wire n_4783;
wire n_7658;
wire n_3017;
wire n_10335;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_10753;
wire n_14220;
wire n_2525;
wire n_15783;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_12783;
wire n_13658;
wire n_807;
wire n_5142;
wire n_12431;
wire n_10921;
wire n_10177;
wire n_8971;
wire n_6355;
wire n_7015;
wire n_6039;
wire n_10567;
wire n_6286;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_15677;
wire n_4332;
wire n_17070;
wire n_7226;
wire n_11915;
wire n_9291;
wire n_7987;
wire n_1987;
wire n_7217;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_9009;
wire n_2368;
wire n_9882;
wire n_6377;
wire n_802;
wire n_10492;
wire n_14137;
wire n_15385;
wire n_12061;
wire n_5401;
wire n_16176;
wire n_4595;
wire n_960;
wire n_11873;
wire n_15505;
wire n_7272;
wire n_16048;
wire n_2352;
wire n_8215;
wire n_5201;
wire n_16959;
wire n_5816;
wire n_12628;
wire n_790;
wire n_5551;
wire n_9722;
wire n_16762;
wire n_5416;
wire n_14175;
wire n_4404;
wire n_15373;
wire n_2377;
wire n_14644;
wire n_151;
wire n_16302;
wire n_7906;
wire n_2652;
wire n_11260;
wire n_5498;
wire n_16172;
wire n_5543;
wire n_12359;
wire n_15328;
wire n_16305;
wire n_4054;
wire n_9760;
wire n_6018;
wire n_7765;
wire n_14320;
wire n_1286;
wire n_6021;
wire n_11880;
wire n_11605;
wire n_13615;
wire n_4617;
wire n_14022;
wire n_12974;
wire n_13156;
wire n_1685;
wire n_10741;
wire n_2477;
wire n_4611;
wire n_10037;
wire n_8949;
wire n_2279;
wire n_3169;
wire n_12136;
wire n_2222;
wire n_5797;
wire n_9454;
wire n_10760;
wire n_6511;
wire n_17010;
wire n_13849;
wire n_12121;
wire n_7815;
wire n_1052;
wire n_12658;
wire n_11838;
wire n_13956;
wire n_4732;
wire n_14768;
wire n_10607;
wire n_2076;
wire n_2203;
wire n_5942;
wire n_5764;
wire n_1426;
wire n_13702;
wire n_8983;
wire n_4969;
wire n_11089;
wire n_14314;
wire n_15088;
wire n_8121;
wire n_5252;
wire n_11629;
wire n_11259;
wire n_5777;
wire n_11100;
wire n_15283;
wire n_13119;
wire n_8942;
wire n_7785;
wire n_11608;
wire n_16883;
wire n_13756;
wire n_5063;
wire n_4641;
wire n_15564;
wire n_4399;
wire n_6867;
wire n_4140;
wire n_5171;
wire n_12364;
wire n_14628;
wire n_13867;
wire n_566;
wire n_7728;
wire n_8280;
wire n_2607;
wire n_11632;
wire n_16094;
wire n_3343;
wire n_4712;
wire n_7255;
wire n_3309;
wire n_169;
wire n_7181;
wire n_12156;
wire n_11443;
wire n_173;
wire n_2796;
wire n_858;
wire n_13409;
wire n_13832;
wire n_5393;
wire n_10658;
wire n_8328;
wire n_4817;
wire n_8861;
wire n_6863;
wire n_7352;
wire n_7355;
wire n_11161;
wire n_11770;
wire n_2136;
wire n_13509;
wire n_433;
wire n_8427;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_7328;
wire n_14399;
wire n_2771;
wire n_6322;
wire n_7359;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_11466;
wire n_15931;
wire n_10489;
wire n_15270;
wire n_9826;
wire n_253;
wire n_928;
wire n_9937;
wire n_10347;
wire n_12632;
wire n_3769;
wire n_11810;
wire n_7825;
wire n_13168;
wire n_1565;
wire n_4437;
wire n_6419;
wire n_7916;
wire n_16170;
wire n_13581;
wire n_10952;
wire n_3055;
wire n_8194;
wire n_15862;
wire n_420;
wire n_10758;
wire n_4070;
wire n_15798;
wire n_5346;
wire n_7283;
wire n_9453;
wire n_17126;
wire n_748;
wire n_7903;
wire n_9900;
wire n_12033;
wire n_16282;
wire n_7089;
wire n_1045;
wire n_16128;
wire n_14954;
wire n_8217;
wire n_14534;
wire n_14890;
wire n_16489;
wire n_16808;
wire n_10518;
wire n_9331;
wire n_1881;
wire n_2635;
wire n_7604;
wire n_11789;
wire n_2999;
wire n_988;
wire n_13447;
wire n_12465;
wire n_7647;
wire n_4139;
wire n_4769;
wire n_6130;
wire n_330;
wire n_15649;
wire n_14164;
wire n_14771;
wire n_5868;
wire n_16613;
wire n_6417;
wire n_328;
wire n_368;
wire n_8521;
wire n_7145;
wire n_10808;
wire n_1958;
wire n_12358;
wire n_8285;
wire n_4867;
wire n_3667;
wire n_12446;
wire n_9178;
wire n_9689;
wire n_7803;
wire n_13999;
wire n_2713;
wire n_1422;
wire n_8448;
wire n_14526;
wire n_1965;
wire n_644;
wire n_5167;
wire n_5257;
wire n_16497;
wire n_4450;
wire n_6979;
wire n_11690;
wire n_5986;
wire n_12684;
wire n_9355;
wire n_12851;
wire n_13725;
wire n_16206;
wire n_9489;
wire n_13319;
wire n_16876;
wire n_12307;
wire n_6932;
wire n_10971;
wire n_15757;
wire n_2934;
wire n_7258;
wire n_13019;
wire n_5104;
wire n_16236;
wire n_12341;
wire n_13807;
wire n_16730;
wire n_6961;
wire n_576;
wire n_8732;
wire n_511;
wire n_13297;
wire n_7622;
wire n_14610;
wire n_11968;
wire n_9359;
wire n_429;
wire n_13395;
wire n_7839;
wire n_11854;
wire n_6792;
wire n_7720;
wire n_2210;
wire n_4368;
wire n_16152;
wire n_5794;
wire n_8136;
wire n_10404;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_16816;
wire n_3476;
wire n_6919;
wire n_1049;
wire n_16455;
wire n_11797;
wire n_8420;
wire n_13672;
wire n_141;
wire n_4430;
wire n_8386;
wire n_16593;
wire n_16097;
wire n_6123;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_7440;
wire n_10802;
wire n_15317;
wire n_1356;
wire n_9568;
wire n_6831;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_14302;
wire n_2666;
wire n_5578;
wire n_12654;
wire n_312;
wire n_728;
wire n_4191;
wire n_4409;
wire n_12921;
wire n_11991;
wire n_2401;
wire n_7809;
wire n_16140;
wire n_3255;
wire n_10340;
wire n_16804;
wire n_2588;
wire n_5722;
wire n_16043;
wire n_5811;
wire n_14170;
wire n_935;
wire n_7072;
wire n_10681;
wire n_14303;
wire n_15077;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_11618;
wire n_911;
wire n_15202;
wire n_16498;
wire n_623;
wire n_3509;
wire n_11502;
wire n_10452;
wire n_10221;
wire n_8746;
wire n_10051;
wire n_1403;
wire n_5395;
wire n_453;
wire n_3006;
wire n_4531;
wire n_12498;
wire n_17120;
wire n_3770;
wire n_6458;
wire n_11465;
wire n_12768;
wire n_16935;
wire n_9401;
wire n_8857;
wire n_543;
wire n_11335;
wire n_6986;
wire n_9495;
wire n_3456;
wire n_12625;
wire n_13221;
wire n_10987;
wire n_4532;
wire n_15409;
wire n_236;
wire n_601;
wire n_10551;
wire n_12063;
wire n_7564;
wire n_628;
wire n_10396;
wire n_10646;
wire n_13471;
wire n_13021;
wire n_15589;
wire n_15322;
wire n_10955;
wire n_5863;
wire n_8185;
wire n_8313;
wire n_6633;
wire n_11382;
wire n_13062;
wire n_3790;
wire n_14298;
wire n_14931;
wire n_7775;
wire n_907;
wire n_7118;
wire n_9234;
wire n_16847;
wire n_13706;
wire n_7960;
wire n_14967;
wire n_6152;
wire n_9431;
wire n_5734;
wire n_15831;
wire n_10308;
wire n_10023;
wire n_8281;
wire n_12347;
wire n_847;
wire n_747;
wire n_12543;
wire n_1135;
wire n_2566;
wire n_12958;
wire n_11254;
wire n_5095;
wire n_3101;
wire n_10538;
wire n_14797;
wire n_3662;
wire n_6169;
wire n_5774;
wire n_12532;
wire n_15974;
wire n_7069;
wire n_11388;
wire n_5199;
wire n_13347;
wire n_6546;
wire n_15557;
wire n_14051;
wire n_4257;
wire n_15548;
wire n_4282;
wire n_11043;
wire n_7636;
wire n_4341;
wire n_10199;
wire n_1694;
wire n_10673;
wire n_6925;
wire n_7186;
wire n_593;
wire n_10467;
wire n_8766;
wire n_13976;
wire n_16823;
wire n_1695;
wire n_4027;
wire n_12334;
wire n_4650;
wire n_4309;
wire n_5480;
wire n_6428;
wire n_609;
wire n_6924;
wire n_12876;
wire n_16350;
wire n_3077;
wire n_4944;
wire n_8066;
wire n_11252;
wire n_9340;
wire n_12774;
wire n_12544;
wire n_13793;
wire n_9380;
wire n_7666;
wire n_15892;
wire n_12353;
wire n_6425;
wire n_12653;
wire n_11824;
wire n_10581;
wire n_14594;
wire n_15816;
wire n_3478;
wire n_14369;
wire n_3062;
wire n_1774;
wire n_9976;
wire n_4994;
wire n_10818;
wire n_10226;
wire n_7967;
wire n_14515;
wire n_519;
wire n_16052;
wire n_5977;
wire n_15998;
wire n_8314;
wire n_384;
wire n_16474;
wire n_3533;
wire n_5175;
wire n_7246;
wire n_1994;
wire n_11724;
wire n_3978;
wire n_12052;
wire n_11507;
wire n_3836;
wire n_11086;
wire n_10647;
wire n_13184;
wire n_9064;
wire n_3409;
wire n_15311;
wire n_4381;
wire n_8239;
wire n_9092;
wire n_14968;
wire n_14721;
wire n_3583;
wire n_16413;
wire n_11533;
wire n_4316;
wire n_15900;
wire n_7301;
wire n_11905;
wire n_14160;
wire n_4860;
wire n_4469;
wire n_16017;
wire n_9746;
wire n_12994;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_8497;
wire n_10637;
wire n_15824;
wire n_1157;
wire n_7262;
wire n_234;
wire n_5959;
wire n_15089;
wire n_13856;
wire n_16597;
wire n_8056;
wire n_8210;
wire n_3563;
wire n_10769;
wire n_5945;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_12215;
wire n_10519;
wire n_3689;
wire n_13218;
wire n_7584;
wire n_7748;
wire n_16409;
wire n_1789;
wire n_9066;
wire n_763;
wire n_14637;
wire n_6301;
wire n_14965;
wire n_15988;
wire n_2174;
wire n_13298;
wire n_540;
wire n_5668;
wire n_12535;
wire n_3442;
wire n_3972;
wire n_14248;
wire n_2315;
wire n_4209;
wire n_12582;
wire n_15175;
wire n_14982;
wire n_1687;
wire n_4703;
wire n_6282;
wire n_4934;
wire n_7686;
wire n_11800;
wire n_17082;
wire n_9870;
wire n_14391;
wire n_9817;
wire n_2638;
wire n_12505;
wire n_13396;
wire n_2046;
wire n_13988;
wire n_14648;
wire n_7059;
wire n_15349;
wire n_14947;
wire n_15725;
wire n_6985;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_5600;
wire n_13132;
wire n_395;
wire n_15546;
wire n_16364;
wire n_6737;
wire n_1587;
wire n_10723;
wire n_12875;
wire n_213;
wire n_2340;
wire n_9857;
wire n_13794;
wire n_4804;
wire n_8404;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_5767;
wire n_9455;
wire n_10056;
wire n_6459;
wire n_15126;
wire n_1427;
wire n_7670;
wire n_13400;
wire n_2977;
wire n_3991;
wire n_13813;
wire n_14307;
wire n_4936;
wire n_8505;
wire n_10653;
wire n_2199;
wire n_6384;
wire n_4669;
wire n_15345;
wire n_15509;
wire n_5228;
wire n_15571;
wire n_15678;
wire n_15777;
wire n_1100;
wire n_585;
wire n_9916;
wire n_1617;
wire n_10157;
wire n_2600;
wire n_8606;
wire n_13542;
wire n_7443;
wire n_10701;
wire n_10470;
wire n_10923;
wire n_12828;
wire n_3436;
wire n_5973;
wire n_7484;
wire n_1962;
wire n_12402;
wire n_14387;
wire n_3806;
wire n_9440;
wire n_4759;
wire n_10038;
wire n_9059;
wire n_11691;
wire n_9812;
wire n_14666;
wire n_5869;
wire n_5914;
wire n_2114;
wire n_6753;
wire n_9690;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_13879;
wire n_11594;
wire n_9912;
wire n_11687;
wire n_14793;
wire n_1175;
wire n_4887;
wire n_15913;
wire n_3751;
wire n_11513;
wire n_9002;
wire n_16057;
wire n_3402;
wire n_9620;
wire n_1621;
wire n_10619;
wire n_13522;
wire n_16901;
wire n_6448;
wire n_9229;
wire n_12524;
wire n_14535;
wire n_15051;
wire n_5186;
wire n_14196;
wire n_7930;
wire n_7487;
wire n_4585;
wire n_1785;
wire n_13403;
wire n_10454;
wire n_11655;
wire n_3406;
wire n_13241;
wire n_580;
wire n_3664;
wire n_4218;
wire n_9464;
wire n_11386;
wire n_434;
wire n_4687;
wire n_7077;
wire n_14060;
wire n_10656;
wire n_394;
wire n_10871;
wire n_1381;
wire n_15406;
wire n_3686;
wire n_1183;
wire n_8518;
wire n_11111;
wire n_4720;
wire n_2889;
wire n_13270;
wire n_11938;
wire n_15037;
wire n_6043;
wire n_6268;
wire n_12670;
wire n_9497;
wire n_2141;
wire n_14923;
wire n_1110;
wire n_1758;
wire n_14543;
wire n_5604;
wire n_3470;
wire n_243;
wire n_8350;
wire n_8741;
wire n_10444;
wire n_11833;
wire n_5221;
wire n_7024;
wire n_1407;
wire n_8148;
wire n_11866;
wire n_8408;
wire n_6145;
wire n_12308;
wire n_17020;
wire n_15523;
wire n_2865;
wire n_10846;
wire n_12659;
wire n_13934;
wire n_14854;
wire n_13024;
wire n_5925;
wire n_6529;
wire n_973;
wire n_5591;
wire n_4762;
wire n_13223;
wire n_3844;
wire n_3259;
wire n_8236;
wire n_14202;
wire n_11192;
wire n_15970;
wire n_11229;
wire n_7214;
wire n_11244;
wire n_16421;
wire n_8806;
wire n_14352;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_8295;
wire n_1176;
wire n_9587;
wire n_3677;
wire n_1054;
wire n_13888;
wire n_7977;
wire n_15370;
wire n_15166;
wire n_14719;
wire n_15260;
wire n_5387;
wire n_13529;
wire n_12452;
wire n_3292;
wire n_16340;
wire n_6311;
wire n_11848;
wire n_13530;
wire n_8377;
wire n_13591;
wire n_3989;
wire n_7652;
wire n_8167;
wire n_10558;
wire n_16518;
wire n_9783;
wire n_4644;
wire n_8956;
wire n_4752;
wire n_8673;
wire n_4746;
wire n_16957;
wire n_7566;
wire n_14631;
wire n_1057;
wire n_4131;
wire n_11876;
wire n_16120;
wire n_12667;
wire n_5449;
wire n_8760;
wire n_4215;
wire n_15032;
wire n_15121;
wire n_17161;
wire n_978;
wire n_12707;
wire n_2488;
wire n_1509;
wire n_828;
wire n_6134;
wire n_16246;
wire n_322;
wire n_4158;
wire n_10466;
wire n_14824;
wire n_6812;
wire n_3079;
wire n_10546;
wire n_10044;
wire n_12878;
wire n_14919;
wire n_5190;
wire n_15886;
wire n_6733;
wire n_11666;
wire n_3269;
wire n_558;
wire n_5325;
wire n_13354;
wire n_10527;
wire n_4231;
wire n_8960;
wire n_8957;
wire n_9008;
wire n_10143;
wire n_12361;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_10233;
wire n_653;
wire n_14856;
wire n_6262;
wire n_4926;
wire n_2050;
wire n_8207;
wire n_6938;
wire n_2197;
wire n_4872;
wire n_12709;
wire n_16734;
wire n_4778;
wire n_5876;
wire n_10461;
wire n_5344;
wire n_2550;
wire n_15827;
wire n_556;
wire n_170;
wire n_1536;
wire n_16428;
wire n_3177;
wire n_6160;
wire n_10186;
wire n_4667;
wire n_10113;
wire n_12721;
wire n_5813;
wire n_6235;
wire n_1471;
wire n_13023;
wire n_6212;
wire n_3440;
wire n_16150;
wire n_9381;
wire n_9194;
wire n_6816;
wire n_8904;
wire n_16772;
wire n_3658;
wire n_16725;
wire n_12264;
wire n_14683;
wire n_7374;
wire n_16839;
wire n_12464;
wire n_13268;
wire n_12753;
wire n_3404;
wire n_2291;
wire n_13887;
wire n_3346;
wire n_2816;
wire n_12968;
wire n_15107;
wire n_1620;
wire n_2542;
wire n_10120;
wire n_5892;
wire n_9549;
wire n_16809;
wire n_7678;
wire n_17076;
wire n_2165;
wire n_15402;
wire n_4837;
wire n_14848;
wire n_4210;
wire n_15539;
wire n_11248;
wire n_788;
wire n_13660;
wire n_7110;
wire n_15712;
wire n_5714;
wire n_17053;
wire n_12111;
wire n_2169;
wire n_6953;
wire n_9652;
wire n_9957;
wire n_7975;
wire n_13481;
wire n_15485;
wire n_12609;
wire n_13143;
wire n_12482;
wire n_8451;
wire n_17079;
wire n_6089;
wire n_591;
wire n_16363;
wire n_10591;
wire n_11780;
wire n_5634;
wire n_12966;
wire n_5133;
wire n_14607;
wire n_8527;
wire n_7553;
wire n_5990;
wire n_7086;
wire n_2175;
wire n_1625;
wire n_5305;
wire n_5689;
wire n_7732;
wire n_7891;
wire n_13419;
wire n_13383;
wire n_9089;
wire n_16332;
wire n_4578;
wire n_318;
wire n_8840;
wire n_11424;
wire n_16904;
wire n_11467;
wire n_5644;
wire n_9137;
wire n_9390;
wire n_3644;
wire n_11995;
wire n_12178;
wire n_8038;
wire n_8190;
wire n_9439;
wire n_11701;
wire n_2176;
wire n_15803;
wire n_1412;
wire n_15405;
wire n_3059;
wire n_6138;
wire n_528;
wire n_16333;
wire n_15621;
wire n_9080;
wire n_17141;
wire n_14773;
wire n_15706;
wire n_15878;
wire n_16752;
wire n_13351;
wire n_1922;
wire n_9296;
wire n_12997;
wire n_16169;
wire n_940;
wire n_10625;
wire n_13544;
wire n_16180;
wire n_1537;
wire n_4877;
wire n_15060;
wire n_14173;
wire n_9312;
wire n_10662;
wire n_2065;
wire n_12818;
wire n_9151;
wire n_16572;
wire n_8179;
wire n_7038;
wire n_7994;
wire n_4470;
wire n_4187;
wire n_9883;
wire n_13420;
wire n_14576;
wire n_10697;
wire n_8287;
wire n_14981;
wire n_1904;
wire n_16714;
wire n_8341;
wire n_8111;
wire n_13527;
wire n_16006;
wire n_8830;
wire n_13206;
wire n_13235;
wire n_16541;
wire n_4998;
wire n_10200;
wire n_14436;
wire n_5576;
wire n_13399;
wire n_16994;
wire n_2395;
wire n_2868;
wire n_10935;
wire n_7345;
wire n_9324;
wire n_13317;
wire n_9631;
wire n_8308;
wire n_10547;
wire n_1530;
wire n_4057;
wire n_6070;
wire n_15432;
wire n_5852;
wire n_5918;
wire n_631;
wire n_8021;
wire n_11092;
wire n_13622;
wire n_1170;
wire n_10933;
wire n_14790;
wire n_2724;
wire n_8965;
wire n_9736;
wire n_16635;
wire n_2258;
wire n_7041;
wire n_9365;
wire n_10632;
wire n_14651;
wire n_16083;
wire n_6717;
wire n_7593;
wire n_8265;
wire n_13564;
wire n_898;
wire n_11166;
wire n_6881;
wire n_10085;
wire n_14881;
wire n_3328;
wire n_17085;
wire n_2012;
wire n_9600;
wire n_3182;
wire n_6871;
wire n_15629;
wire n_2967;
wire n_9816;
wire n_5343;
wire n_9869;
wire n_6672;
wire n_16997;
wire n_7757;
wire n_1093;
wire n_13276;
wire n_8251;
wire n_7866;
wire n_6518;
wire n_7334;
wire n_9402;
wire n_4021;
wire n_6396;
wire n_7028;
wire n_3379;
wire n_4379;
wire n_8773;
wire n_12195;
wire n_14383;
wire n_16998;
wire n_14400;
wire n_5947;
wire n_6242;
wire n_14143;
wire n_336;
wire n_6601;
wire n_8570;
wire n_12536;
wire n_10645;
wire n_2268;
wire n_3469;
wire n_10041;
wire n_15392;
wire n_12168;
wire n_16373;
wire n_16868;
wire n_14858;
wire n_16544;
wire n_16505;
wire n_1452;
wire n_2835;
wire n_5835;
wire n_10096;
wire n_668;
wire n_12533;
wire n_8579;
wire n_15333;
wire n_2111;
wire n_3743;
wire n_15762;
wire n_8079;
wire n_5542;
wire n_9615;
wire n_11869;
wire n_14106;
wire n_2948;
wire n_5015;
wire n_13792;
wire n_3099;
wire n_12560;
wire n_16319;
wire n_5527;
wire n_2897;
wire n_9711;
wire n_9759;
wire n_4812;
wire n_8506;
wire n_8973;
wire n_13171;
wire n_4497;
wire n_6606;
wire n_2583;
wire n_13764;
wire n_8291;
wire n_3155;
wire n_14725;
wire n_4300;
wire n_16077;
wire n_2024;
wire n_11264;
wire n_10336;
wire n_16018;
wire n_9820;
wire n_1770;
wire n_701;
wire n_1003;
wire n_7758;
wire n_8320;
wire n_12477;
wire n_8635;
wire n_9703;
wire n_4472;
wire n_12516;
wire n_9819;
wire n_15422;
wire n_9118;
wire n_11060;
wire n_16922;
wire n_15722;
wire n_2699;
wire n_9321;
wire n_12523;
wire n_11493;
wire n_11562;
wire n_13698;
wire n_5819;
wire n_3901;
wire n_291;
wire n_5180;
wire n_1640;
wire n_8375;
wire n_10703;
wire n_11575;
wire n_2973;
wire n_10449;
wire n_13462;
wire n_14959;
wire n_16114;
wire n_14806;
wire n_16637;
wire n_10280;
wire n_9428;
wire n_8612;
wire n_10198;
wire n_8778;
wire n_16978;
wire n_11065;
wire n_5893;
wire n_9292;
wire n_11452;
wire n_15366;
wire n_2710;
wire n_7705;
wire n_16393;
wire n_6092;
wire n_12486;
wire n_6462;
wire n_2505;
wire n_15977;
wire n_11345;
wire n_4519;
wire n_15989;
wire n_9018;
wire n_16700;
wire n_13741;
wire n_5025;
wire n_2397;
wire n_8872;
wire n_12743;
wire n_240;
wire n_369;
wire n_10371;
wire n_7333;
wire n_3878;
wire n_12246;
wire n_4197;
wire n_12297;
wire n_13440;
wire n_6669;
wire n_8006;
wire n_11495;
wire n_9565;
wire n_2721;
wire n_13325;
wire n_1892;
wire n_6251;
wire n_2615;
wire n_4787;
wire n_8491;
wire n_8218;
wire n_1212;
wire n_13089;
wire n_13578;
wire n_7337;
wire n_4310;
wire n_5726;
wire n_3933;
wire n_4566;
wire n_7439;
wire n_4371;
wire n_12610;
wire n_14006;
wire n_14901;
wire n_16336;
wire n_14757;
wire n_10483;
wire n_188;
wire n_16422;
wire n_12771;
wire n_1902;
wire n_5828;
wire n_2784;
wire n_7210;
wire n_10346;
wire n_3898;
wire n_7744;
wire n_11864;
wire n_16426;
wire n_694;
wire n_6228;
wire n_15619;
wire n_16030;
wire n_10805;
wire n_14107;
wire n_6702;
wire n_7358;
wire n_8240;
wire n_10059;
wire n_9961;
wire n_15990;
wire n_4749;
wire n_12763;
wire n_16038;
wire n_7707;
wire n_5924;
wire n_1845;
wire n_7733;
wire n_13496;
wire n_921;
wire n_14536;
wire n_5545;
wire n_16174;
wire n_8458;
wire n_2104;
wire n_16678;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_8853;
wire n_9603;
wire n_11293;
wire n_14950;
wire n_5083;
wire n_15122;
wire n_15341;
wire n_15159;
wire n_7684;
wire n_14834;
wire n_16805;
wire n_10700;
wire n_11984;
wire n_3253;
wire n_16819;
wire n_17176;
wire n_11961;
wire n_8306;
wire n_2088;
wire n_11981;
wire n_1275;
wire n_14599;
wire n_6997;
wire n_9692;
wire n_4238;
wire n_6371;
wire n_13222;
wire n_904;
wire n_11559;
wire n_7673;
wire n_2005;
wire n_15391;
wire n_1696;
wire n_14642;
wire n_15674;
wire n_12172;
wire n_11942;
wire n_11207;
wire n_11686;
wire n_14809;
wire n_12280;
wire n_12883;
wire n_8013;
wire n_14897;
wire n_2108;
wire n_7187;
wire n_14476;
wire n_3824;
wire n_8342;
wire n_10502;
wire n_12064;
wire n_12480;
wire n_2246;
wire n_10974;
wire n_7313;
wire n_16212;
wire n_5899;
wire n_11239;
wire n_14221;
wire n_10511;
wire n_10250;
wire n_9012;
wire n_11482;
wire n_3846;
wire n_12682;
wire n_10831;
wire n_17180;
wire n_5122;
wire n_11992;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_12621;
wire n_15843;
wire n_4479;
wire n_13754;
wire n_10613;
wire n_16254;
wire n_6641;
wire n_3845;
wire n_12283;
wire n_10351;
wire n_10172;
wire n_3203;
wire n_13285;
wire n_383;
wire n_6463;
wire n_4986;
wire n_10333;
wire n_1316;
wire n_4668;
wire n_950;
wire n_9868;
wire n_711;
wire n_6264;
wire n_15789;
wire n_5782;
wire n_8119;
wire n_9264;
wire n_16460;
wire n_630;
wire n_4168;
wire n_1369;
wire n_8582;
wire n_11479;
wire n_11814;
wire n_4298;
wire n_10594;
wire n_7036;
wire n_7370;
wire n_7931;
wire n_4743;
wire n_13181;
wire n_11622;
wire n_8445;
wire n_12225;
wire n_1781;
wire n_9720;
wire n_4250;
wire n_15245;
wire n_13004;
wire n_11067;
wire n_3143;
wire n_8044;
wire n_13413;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_8363;
wire n_8464;
wire n_16784;
wire n_8921;
wire n_12208;
wire n_14072;
wire n_13608;
wire n_15858;
wire n_12126;
wire n_13397;
wire n_235;
wire n_2188;
wire n_15003;
wire n_11083;
wire n_14282;
wire n_10010;
wire n_10588;
wire n_11907;
wire n_2430;
wire n_2504;
wire n_12396;
wire n_12984;
wire n_17170;
wire n_11952;
wire n_4211;
wire n_6084;
wire n_3094;
wire n_741;
wire n_9646;
wire n_16109;
wire n_5637;
wire n_7480;
wire n_13997;
wire n_12158;
wire n_8843;
wire n_371;
wire n_13513;
wire n_5185;
wire n_16424;
wire n_8405;
wire n_13232;
wire n_2964;
wire n_13296;
wire n_13816;
wire n_14713;
wire n_8376;
wire n_308;
wire n_16414;
wire n_13859;
wire n_5032;
wire n_11506;
wire n_6990;
wire n_865;
wire n_5034;
wire n_3312;
wire n_7071;
wire n_1041;
wire n_2451;
wire n_10797;
wire n_8694;
wire n_16695;
wire n_2913;
wire n_8848;
wire n_6288;
wire n_993;
wire n_13989;
wire n_1862;
wire n_14573;
wire n_3752;
wire n_8752;
wire n_10643;
wire n_3672;
wire n_922;
wire n_1004;
wire n_8894;
wire n_8625;
wire n_7380;
wire n_14058;
wire n_2839;
wire n_16118;
wire n_8813;
wire n_3237;
wire n_7708;
wire n_12690;
wire n_12813;
wire n_16622;
wire n_11524;
wire n_10905;
wire n_9842;
wire n_11859;
wire n_4128;
wire n_11228;
wire n_16583;
wire n_12725;
wire n_4036;
wire n_9671;
wire n_5269;
wire n_15025;
wire n_8430;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_1764;
wire n_10784;
wire n_11035;
wire n_4807;
wire n_16949;
wire n_11023;
wire n_8770;
wire n_6277;
wire n_8426;
wire n_14009;
wire n_5115;
wire n_12474;
wire n_7376;
wire n_11174;
wire n_8411;
wire n_16992;
wire n_13759;
wire n_902;
wire n_8817;
wire n_8461;
wire n_10438;
wire n_1723;
wire n_15056;
wire n_3918;
wire n_14911;
wire n_10234;
wire n_17016;
wire n_10946;
wire n_11582;
wire n_9230;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_11705;
wire n_17093;
wire n_4391;
wire n_11796;
wire n_596;
wire n_12484;
wire n_9893;
wire n_6409;
wire n_4095;
wire n_8391;
wire n_17006;
wire n_8507;
wire n_1310;
wire n_12021;
wire n_5927;
wire n_11003;
wire n_9188;
wire n_8691;
wire n_4485;
wire n_9032;
wire n_7657;
wire n_6388;
wire n_16463;
wire n_10275;
wire n_574;
wire n_3593;
wire n_15279;
wire n_6839;
wire n_14284;
wire n_5163;
wire n_9614;
wire n_16852;
wire n_8967;
wire n_12990;
wire n_1229;
wire n_2582;
wire n_16872;
wire n_3327;
wire n_4356;
wire n_9628;
wire n_1896;
wire n_9231;
wire n_10854;
wire n_6864;
wire n_14309;
wire n_13652;
wire n_1516;
wire n_13207;
wire n_4890;
wire n_10204;
wire n_8084;
wire n_8856;
wire n_15963;
wire n_2485;
wire n_12685;
wire n_12778;
wire n_6679;
wire n_12862;
wire n_11528;
wire n_10734;
wire n_13442;
wire n_17008;
wire n_10201;
wire n_8631;
wire n_16144;
wire n_6051;
wire n_15128;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_8219;
wire n_16008;
wire n_9730;
wire n_5507;
wire n_15898;
wire n_10608;
wire n_16556;
wire n_195;
wire n_4573;
wire n_1328;
wire n_10746;
wire n_4943;
wire n_2875;
wire n_10676;
wire n_6599;
wire n_3519;
wire n_2209;
wire n_16609;
wire n_14423;
wire n_12177;
wire n_13128;
wire n_7504;
wire n_14086;
wire n_4042;
wire n_7099;
wire n_7586;
wire n_4244;
wire n_16554;
wire n_1928;
wire n_5642;
wire n_12672;
wire n_4708;
wire n_4883;
wire n_17122;
wire n_6227;
wire n_4553;
wire n_7052;
wire n_8428;
wire n_9172;
wire n_12141;
wire n_14665;
wire n_1634;
wire n_17057;
wire n_14342;
wire n_1203;
wire n_9926;
wire n_1699;
wire n_14634;
wire n_6738;
wire n_12665;
wire n_13719;
wire n_5226;
wire n_2081;
wire n_937;
wire n_1474;
wire n_11615;
wire n_11079;
wire n_8338;
wire n_14772;
wire n_1631;
wire n_7602;
wire n_9180;
wire n_12024;
wire n_12795;
wire n_156;
wire n_9017;
wire n_9269;
wire n_9026;
wire n_16540;
wire n_6566;
wire n_13453;
wire n_1794;
wire n_9462;
wire n_10900;
wire n_5696;
wire n_13370;
wire n_7998;
wire n_8666;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_7106;
wire n_6346;
wire n_204;
wire n_11438;
wire n_11700;
wire n_12940;
wire n_3772;
wire n_7408;
wire n_7557;
wire n_12555;
wire n_16123;
wire n_16551;
wire n_14539;
wire n_2891;
wire n_496;
wire n_4335;
wire n_10052;
wire n_3128;
wire n_7026;
wire n_16215;
wire n_13656;
wire n_11668;
wire n_15286;
wire n_6146;
wire n_13667;
wire n_5677;
wire n_13641;
wire n_4277;
wire n_12487;
wire n_16464;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_7394;
wire n_11387;
wire n_9515;
wire n_10560;
wire n_9502;
wire n_13103;
wire n_263;
wire n_4516;
wire n_5235;
wire n_360;
wire n_13183;
wire n_13720;
wire n_1129;
wire n_13971;
wire n_15650;
wire n_11099;
wire n_15929;
wire n_7627;
wire n_6436;
wire n_12305;
wire n_1464;
wire n_7719;
wire n_2798;
wire n_10773;
wire n_7450;
wire n_165;
wire n_9316;
wire n_3217;
wire n_11996;
wire n_15962;
wire n_8938;
wire n_6081;
wire n_13436;
wire n_14479;
wire n_16098;
wire n_10455;
wire n_1249;
wire n_14410;
wire n_16148;
wire n_329;
wire n_7852;
wire n_5724;
wire n_3821;
wire n_340;
wire n_12526;
wire n_3201;
wire n_12622;
wire n_12456;
wire n_7462;
wire n_7780;
wire n_3503;
wire n_10391;
wire n_8523;
wire n_12857;
wire n_5979;
wire n_10476;
wire n_10630;
wire n_10559;
wire n_13797;
wire n_6027;
wire n_13321;
wire n_1870;
wire n_10911;
wire n_11547;
wire n_10121;
wire n_11064;
wire n_12439;
wire n_4467;
wire n_15785;
wire n_177;
wire n_13809;
wire n_364;
wire n_258;
wire n_7582;
wire n_15522;
wire n_10540;
wire n_16304;
wire n_5521;
wire n_17135;
wire n_431;
wire n_15140;
wire n_2654;
wire n_3935;
wire n_7421;
wire n_13575;
wire n_16239;
wire n_1861;
wire n_11104;
wire n_9873;
wire n_1228;
wire n_2319;
wire n_10473;
wire n_15120;
wire n_15234;
wire n_12287;
wire n_10828;
wire n_12182;
wire n_13390;
wire n_8924;
wire n_2965;
wire n_12366;
wire n_7555;
wire n_4955;
wire n_11112;
wire n_16968;
wire n_14915;
wire n_10114;
wire n_17160;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_447;
wire n_2689;
wire n_6110;
wire n_12552;
wire n_14123;
wire n_1762;
wire n_10269;
wire n_14258;
wire n_6238;
wire n_7025;
wire n_3798;
wire n_3080;
wire n_8380;
wire n_13371;
wire n_12777;
wire n_16591;
wire n_9978;
wire n_5241;
wire n_16547;
wire n_12492;
wire n_10418;
wire n_4248;
wire n_1672;
wire n_16367;
wire n_2228;
wire n_4645;
wire n_15235;
wire n_16471;
wire n_17127;
wire n_13231;
wire n_5331;
wire n_7478;
wire n_3308;
wire n_6326;
wire n_841;
wire n_3204;
wire n_10672;
wire n_7451;
wire n_9494;
wire n_15918;
wire n_4134;
wire n_5018;
wire n_14601;
wire n_6917;
wire n_11850;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_12437;
wire n_2345;
wire n_1730;
wire n_6612;
wire n_10922;
wire n_5258;

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_3),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_5),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_29),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_128),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_12),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_110),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_126),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_8),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_18),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_67),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_0),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_95),
.Y(n_147)
);

BUFx10_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_13),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_51),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_106),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_52),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_17),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_60),
.Y(n_158)
);

BUFx10_ASAP7_75t_L g159 ( 
.A(n_47),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_61),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_39),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_14),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_74),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_35),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_31),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_71),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_100),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_87),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_97),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_116),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_11),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_105),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_83),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_15),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_33),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_76),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_36),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_41),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_54),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_131),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_24),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_38),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_130),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_91),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_101),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_3),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_113),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_98),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_85),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_6),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_49),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_2),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_10),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_81),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_72),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_28),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_124),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_56),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_20),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_132),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_55),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_79),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_107),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_19),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_46),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_50),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_68),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_77),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_45),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_43),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_80),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_30),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_0),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_59),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_114),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_92),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_112),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_118),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_58),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_23),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_64),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_4),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_2),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_22),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_7),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_21),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_4),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_123),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_127),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_134),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_133),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_108),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_65),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_42),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_78),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_125),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_25),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_122),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_16),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_63),
.Y(n_242)
);

CKINVDCx12_ASAP7_75t_R g243 ( 
.A(n_129),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_111),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_102),
.Y(n_245)
);

BUFx8_ASAP7_75t_SL g246 ( 
.A(n_73),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_57),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_26),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_62),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_27),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_103),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_86),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_1),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_99),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_93),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_89),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_70),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_69),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_48),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_32),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_109),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_117),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_66),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_88),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_53),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_104),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_40),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_44),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_37),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_215),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_139),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_229),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_154),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_236),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_148),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_144),
.B(n_1),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_246),
.Y(n_277)
);

BUFx8_ASAP7_75t_SL g278 ( 
.A(n_136),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_148),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_150),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_151),
.Y(n_281)
);

NOR2xp67_ASAP7_75t_L g282 ( 
.A(n_146),
.B(n_9),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_159),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_159),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_201),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_169),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_187),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_156),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_153),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_162),
.Y(n_290)
);

XNOR2x1_ASAP7_75t_L g291 ( 
.A(n_194),
.B(n_34),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_169),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_199),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_199),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_214),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_214),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_184),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_232),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_235),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_249),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_264),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_258),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_224),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_225),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_201),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_253),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_L g307 ( 
.A(n_155),
.B(n_82),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_137),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_160),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_264),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_171),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_177),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_287),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_270),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_309),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_272),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_288),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_297),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_285),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_296),
.B(n_164),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_174),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_271),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_280),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_290),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_298),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_292),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_281),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_289),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_299),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_300),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_311),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_312),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_285),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_303),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_275),
.B(n_181),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_277),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_285),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_305),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_305),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_302),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_278),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_301),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_305),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_304),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_306),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_279),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_276),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_283),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_276),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_273),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_274),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_R g352 ( 
.A(n_284),
.B(n_269),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_286),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_293),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_294),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_295),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_310),
.B(n_185),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_291),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_282),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_307),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_346),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_316),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_323),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_319),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_319),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_138),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_319),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_327),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_346),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_328),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_337),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_333),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_338),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_345),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_339),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_314),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_331),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_332),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_343),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_356),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_353),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_354),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_326),
.B(n_175),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_336),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_326),
.B(n_198),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_347),
.B(n_191),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_348),
.A2(n_212),
.B1(n_265),
.B2(n_227),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_320),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_342),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_355),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_335),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_350),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_317),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_351),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_318),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_349),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_315),
.B(n_210),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_360),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_321),
.B(n_140),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_357),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_315),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_359),
.Y(n_402)
);

OA21x2_ASAP7_75t_L g403 ( 
.A1(n_334),
.A2(n_268),
.B(n_266),
.Y(n_403)
);

AOI22x1_ASAP7_75t_SL g404 ( 
.A1(n_341),
.A2(n_261),
.B1(n_255),
.B2(n_239),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_313),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_352),
.B(n_325),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_329),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_358),
.A2(n_205),
.B1(n_233),
.B2(n_226),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_330),
.Y(n_409)
);

OA21x2_ASAP7_75t_L g410 ( 
.A1(n_340),
.A2(n_218),
.B(n_206),
.Y(n_410)
);

BUFx12f_ASAP7_75t_L g411 ( 
.A(n_322),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_324),
.B(n_197),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_347),
.B(n_141),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_316),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_348),
.A2(n_222),
.B1(n_216),
.B2(n_243),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_347),
.B(n_142),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_323),
.Y(n_417)
);

OA21x2_ASAP7_75t_L g418 ( 
.A1(n_335),
.A2(n_262),
.B(n_259),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_319),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_316),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_323),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_323),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_316),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_319),
.Y(n_424)
);

OA21x2_ASAP7_75t_L g425 ( 
.A1(n_335),
.A2(n_245),
.B(n_242),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_323),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_319),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_319),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_323),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_323),
.Y(n_430)
);

AOI22x1_ASAP7_75t_SL g431 ( 
.A1(n_341),
.A2(n_267),
.B1(n_263),
.B2(n_260),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_323),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_348),
.A2(n_196),
.B1(n_256),
.B2(n_252),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_331),
.B(n_240),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_323),
.Y(n_435)
);

OA21x2_ASAP7_75t_L g436 ( 
.A1(n_335),
.A2(n_238),
.B(n_157),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_323),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_316),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_326),
.B(n_149),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_319),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_346),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_316),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_326),
.B(n_195),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_323),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_326),
.B(n_193),
.Y(n_445)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_336),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_344),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_336),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_319),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_319),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_331),
.B(n_254),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_315),
.B(n_200),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_315),
.B(n_192),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_316),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_344),
.Y(n_455)
);

OA21x2_ASAP7_75t_L g456 ( 
.A1(n_335),
.A2(n_257),
.B(n_251),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_358),
.A2(n_190),
.B1(n_250),
.B2(n_248),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_323),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_322),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_313),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_326),
.B(n_183),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_323),
.Y(n_462)
);

OA21x2_ASAP7_75t_L g463 ( 
.A1(n_335),
.A2(n_189),
.B(n_247),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_323),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_316),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_316),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_326),
.B(n_182),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_326),
.B(n_180),
.Y(n_468)
);

NAND2xp33_ASAP7_75t_L g469 ( 
.A(n_344),
.B(n_244),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_323),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_323),
.Y(n_471)
);

NOR2x1_ASAP7_75t_L g472 ( 
.A(n_321),
.B(n_204),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_347),
.B(n_178),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_331),
.B(n_201),
.Y(n_474)
);

AND2x2_ASAP7_75t_SL g475 ( 
.A(n_320),
.B(n_254),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_315),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_336),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_347),
.B(n_179),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_319),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_316),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_313),
.Y(n_481)
);

OA21x2_ASAP7_75t_L g482 ( 
.A1(n_335),
.A2(n_202),
.B(n_241),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_316),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_323),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_323),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_344),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_316),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_323),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_319),
.Y(n_489)
);

OA21x2_ASAP7_75t_L g490 ( 
.A1(n_335),
.A2(n_173),
.B(n_237),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_323),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_316),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_394),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_362),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_376),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_401),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_477),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_406),
.B(n_176),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_414),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_420),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_378),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_423),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_438),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_459),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_442),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_454),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_391),
.B(n_172),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_455),
.A2(n_203),
.B1(n_234),
.B2(n_231),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_388),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_465),
.Y(n_510)
);

AND2x6_ASAP7_75t_L g511 ( 
.A(n_406),
.B(n_254),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_466),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_480),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_483),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_487),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_492),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_388),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_400),
.B(n_186),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_377),
.Y(n_519)
);

NAND2xp33_ASAP7_75t_L g520 ( 
.A(n_486),
.B(n_188),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_476),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_380),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_374),
.B(n_170),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_363),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_397),
.B(n_230),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_396),
.B(n_168),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_447),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_368),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_370),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_417),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_421),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_422),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_411),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_397),
.B(n_228),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_426),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_429),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_399),
.B(n_167),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_389),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_386),
.B(n_223),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_430),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_432),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_393),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_435),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_437),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_444),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_412),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_458),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_462),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_464),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_470),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_471),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_484),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_485),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_488),
.Y(n_554)
);

OAI21x1_ASAP7_75t_L g555 ( 
.A1(n_472),
.A2(n_418),
.B(n_425),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_384),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_491),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_395),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_446),
.B(n_448),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_475),
.B(n_166),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_395),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_384),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_407),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_382),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_373),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_390),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_460),
.Y(n_567)
);

BUFx6f_ASAP7_75t_SL g568 ( 
.A(n_407),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_371),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_452),
.B(n_221),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_481),
.B(n_165),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_381),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_451),
.Y(n_573)
);

NAND2x1p5_ASAP7_75t_L g574 ( 
.A(n_409),
.B(n_405),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_451),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_474),
.Y(n_576)
);

OA21x2_ASAP7_75t_L g577 ( 
.A1(n_413),
.A2(n_473),
.B(n_478),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_474),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_392),
.A2(n_220),
.B1(n_219),
.B2(n_217),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_379),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_372),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_434),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_409),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_434),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_372),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_416),
.A2(n_161),
.B1(n_211),
.B2(n_209),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_375),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_457),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_375),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_361),
.Y(n_590)
);

OAI21x1_ASAP7_75t_L g591 ( 
.A1(n_436),
.A2(n_188),
.B(n_213),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_461),
.B(n_152),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_364),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_369),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_441),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_453),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_364),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_439),
.B(n_158),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_365),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_365),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_443),
.B(n_147),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_367),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_367),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_419),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_402),
.B(n_163),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_419),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_424),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_424),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_427),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_445),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_427),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_433),
.B(n_145),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_428),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_428),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_SL g615 ( 
.A(n_467),
.B(n_208),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_440),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_440),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_449),
.Y(n_618)
);

NAND2xp33_ASAP7_75t_L g619 ( 
.A(n_387),
.B(n_188),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_SL g620 ( 
.A(n_408),
.B(n_143),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_449),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_450),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_450),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_479),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_479),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_489),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_468),
.B(n_207),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_489),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_383),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_398),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_385),
.B(n_188),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_403),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_415),
.B(n_204),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_456),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_410),
.Y(n_635)
);

OA21x2_ASAP7_75t_L g636 ( 
.A1(n_463),
.A2(n_188),
.B(n_204),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_482),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_490),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_431),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_404),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_366),
.B(n_84),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_469),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_362),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_475),
.B(n_96),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_477),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_394),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_391),
.A2(n_119),
.B1(n_386),
.B2(n_397),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_391),
.A2(n_386),
.B1(n_397),
.B2(n_392),
.Y(n_648)
);

CKINVDCx11_ASAP7_75t_R g649 ( 
.A(n_411),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_362),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_391),
.A2(n_386),
.B1(n_397),
.B2(n_392),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_394),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_477),
.Y(n_653)
);

OAI21x1_ASAP7_75t_L g654 ( 
.A1(n_472),
.A2(n_391),
.B(n_377),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_388),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_362),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_397),
.B(n_315),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_391),
.A2(n_386),
.B1(n_397),
.B2(n_392),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_411),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_394),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_406),
.B(n_344),
.Y(n_661)
);

OA21x2_ASAP7_75t_L g662 ( 
.A1(n_413),
.A2(n_473),
.B(n_416),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_477),
.Y(n_663)
);

OAI21x1_ASAP7_75t_L g664 ( 
.A1(n_472),
.A2(n_391),
.B(n_377),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_362),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_394),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_477),
.B(n_374),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_362),
.Y(n_668)
);

OA21x2_ASAP7_75t_L g669 ( 
.A1(n_413),
.A2(n_473),
.B(n_416),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_391),
.B(n_400),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_394),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_397),
.B(n_315),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_391),
.B(n_400),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_394),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_394),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_477),
.B(n_374),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_459),
.Y(n_677)
);

AND3x1_ASAP7_75t_L g678 ( 
.A(n_452),
.B(n_453),
.C(n_386),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_362),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_394),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_394),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_394),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_477),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_397),
.B(n_315),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_362),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_394),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_362),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_459),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_362),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_388),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_459),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_477),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_394),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_394),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_394),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_394),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_362),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_362),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_388),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_394),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_394),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_394),
.Y(n_702)
);

OA21x2_ASAP7_75t_L g703 ( 
.A1(n_413),
.A2(n_473),
.B(n_416),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_394),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_477),
.B(n_374),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_394),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_362),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_394),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_362),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_394),
.Y(n_710)
);

NAND3xp33_ASAP7_75t_L g711 ( 
.A(n_366),
.B(n_345),
.C(n_344),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_394),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_397),
.B(n_315),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_394),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_477),
.B(n_388),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_397),
.B(n_315),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_394),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_391),
.B(n_400),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_394),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_362),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_394),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_394),
.Y(n_722)
);

OA21x2_ASAP7_75t_L g723 ( 
.A1(n_413),
.A2(n_473),
.B(n_416),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_394),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_362),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_384),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_477),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_459),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_406),
.B(n_344),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_394),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_384),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_394),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_394),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_394),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_362),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_394),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_362),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_388),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_394),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_397),
.B(n_315),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_362),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_362),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_394),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_477),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_406),
.B(n_344),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_362),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_362),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_406),
.B(n_344),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_394),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_406),
.B(n_344),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_459),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_391),
.B(n_400),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_362),
.Y(n_753)
);

OA21x2_ASAP7_75t_L g754 ( 
.A1(n_413),
.A2(n_473),
.B(n_416),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_406),
.B(n_344),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_477),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_406),
.B(n_344),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_394),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_362),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_388),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_459),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_391),
.B(n_400),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_362),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_411),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_411),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_394),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_394),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_394),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_388),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_477),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_394),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_388),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_394),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_394),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_391),
.B(n_400),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_394),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_394),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_394),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_394),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_L g780 ( 
.A(n_455),
.B(n_344),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_394),
.Y(n_781)
);

OA21x2_ASAP7_75t_L g782 ( 
.A1(n_413),
.A2(n_473),
.B(n_416),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_388),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_394),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_362),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_391),
.B(n_400),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_394),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_362),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_394),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_477),
.B(n_374),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_477),
.B(n_374),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_391),
.B(n_400),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_394),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_459),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_394),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_362),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_394),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_394),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_394),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_394),
.Y(n_800)
);

XNOR2xp5_ASAP7_75t_L g801 ( 
.A(n_459),
.B(n_358),
.Y(n_801)
);

OAI21x1_ASAP7_75t_L g802 ( 
.A1(n_472),
.A2(n_391),
.B(n_377),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_497),
.B(n_645),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_495),
.Y(n_804)
);

NAND2xp33_ASAP7_75t_SL g805 ( 
.A(n_559),
.B(n_497),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_667),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_494),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_501),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_670),
.B(n_673),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_715),
.B(n_726),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_527),
.B(n_596),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_715),
.B(n_731),
.Y(n_812)
);

INVxp33_ASAP7_75t_L g813 ( 
.A(n_801),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_645),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_499),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_761),
.B(n_567),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_496),
.B(n_657),
.Y(n_817)
);

INVx8_ASAP7_75t_L g818 ( 
.A(n_568),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_542),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_672),
.B(n_684),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_500),
.Y(n_821)
);

AND2x6_ASAP7_75t_L g822 ( 
.A(n_644),
.B(n_642),
.Y(n_822)
);

INVxp33_ASAP7_75t_L g823 ( 
.A(n_801),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_648),
.B(n_651),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_502),
.Y(n_825)
);

OAI21xp33_ASAP7_75t_SL g826 ( 
.A1(n_658),
.A2(n_752),
.B(n_718),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_512),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_560),
.A2(n_633),
.B1(n_534),
.B2(n_525),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_653),
.Y(n_829)
);

INVx4_ASAP7_75t_L g830 ( 
.A(n_653),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_762),
.B(n_775),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_676),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_786),
.B(n_792),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_572),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_513),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_678),
.B(n_713),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_524),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_528),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_663),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_529),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_663),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_716),
.B(n_740),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_530),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_531),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_514),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_535),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_536),
.Y(n_847)
);

BUFx4f_ASAP7_75t_L g848 ( 
.A(n_705),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_540),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_570),
.B(n_582),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_543),
.Y(n_851)
);

AND3x2_ASAP7_75t_L g852 ( 
.A(n_659),
.B(n_764),
.C(n_538),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_584),
.B(n_539),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_790),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_515),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_504),
.B(n_677),
.Y(n_856)
);

BUFx6f_ASAP7_75t_SL g857 ( 
.A(n_791),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_643),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_647),
.B(n_711),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_544),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_547),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_650),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_683),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_549),
.Y(n_864)
);

NOR3xp33_ASAP7_75t_L g865 ( 
.A(n_780),
.B(n_508),
.C(n_661),
.Y(n_865)
);

INVx5_ASAP7_75t_L g866 ( 
.A(n_683),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_552),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_692),
.B(n_727),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_553),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_688),
.B(n_691),
.Y(n_870)
);

CKINVDCx16_ASAP7_75t_R g871 ( 
.A(n_765),
.Y(n_871)
);

INVx4_ASAP7_75t_L g872 ( 
.A(n_692),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_728),
.B(n_751),
.Y(n_873)
);

INVx6_ASAP7_75t_L g874 ( 
.A(n_727),
.Y(n_874)
);

INVxp33_ASAP7_75t_SL g875 ( 
.A(n_649),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_656),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_580),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_794),
.B(n_521),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_538),
.B(n_744),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_665),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_744),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_546),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_668),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_620),
.A2(n_541),
.B1(n_545),
.B2(n_532),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_756),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_679),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_685),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_756),
.B(n_770),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_770),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_556),
.B(n_562),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_548),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_518),
.B(n_573),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_687),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_659),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_689),
.Y(n_895)
);

BUFx6f_ASAP7_75t_SL g896 ( 
.A(n_556),
.Y(n_896)
);

INVx4_ASAP7_75t_L g897 ( 
.A(n_562),
.Y(n_897)
);

NOR2x1_ASAP7_75t_L g898 ( 
.A(n_729),
.B(n_745),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_550),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_571),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_697),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_698),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_563),
.B(n_610),
.Y(n_903)
);

INVxp33_ASAP7_75t_L g904 ( 
.A(n_563),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_707),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_709),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_507),
.B(n_523),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_629),
.B(n_598),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_558),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_551),
.Y(n_910)
);

BUFx10_ASAP7_75t_L g911 ( 
.A(n_511),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_629),
.B(n_605),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_554),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_509),
.B(n_517),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_593),
.B(n_606),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_655),
.B(n_690),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_593),
.B(n_606),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_557),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_699),
.B(n_738),
.Y(n_919)
);

BUFx10_ASAP7_75t_L g920 ( 
.A(n_511),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_493),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_720),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_607),
.Y(n_923)
);

AOI21x1_ASAP7_75t_L g924 ( 
.A1(n_637),
.A2(n_638),
.B(n_634),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_575),
.B(n_576),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_764),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_519),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_578),
.B(n_564),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_725),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_760),
.B(n_769),
.Y(n_930)
);

NAND2xp33_ASAP7_75t_SL g931 ( 
.A(n_748),
.B(n_750),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_561),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_566),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_607),
.B(n_614),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_646),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_652),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_583),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_619),
.A2(n_757),
.B1(n_755),
.B2(n_511),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_614),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_735),
.Y(n_940)
);

INVxp67_ASAP7_75t_SL g941 ( 
.A(n_772),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_660),
.Y(n_942)
);

NOR2x1p5_ASAP7_75t_L g943 ( 
.A(n_533),
.B(n_571),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_783),
.B(n_595),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_624),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_666),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_671),
.B(n_674),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_737),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_624),
.B(n_628),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_635),
.A2(n_682),
.B1(n_732),
.B2(n_730),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_675),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_680),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_681),
.B(n_686),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_741),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_628),
.Y(n_955)
);

INVx5_ASAP7_75t_L g956 ( 
.A(n_632),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_526),
.B(n_537),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_693),
.B(n_694),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_574),
.B(n_627),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_695),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_696),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_700),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_701),
.B(n_702),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_704),
.A2(n_768),
.B1(n_733),
.B2(n_724),
.Y(n_964)
);

INVx4_ASAP7_75t_L g965 ( 
.A(n_585),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_706),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_597),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_613),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_579),
.B(n_601),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_742),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_708),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_588),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_746),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_630),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_747),
.Y(n_975)
);

AND2x2_ASAP7_75t_SL g976 ( 
.A(n_520),
.B(n_639),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_616),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_710),
.B(n_712),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_714),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_615),
.B(n_590),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_594),
.B(n_498),
.Y(n_981)
);

AND2x6_ASAP7_75t_L g982 ( 
.A(n_632),
.B(n_717),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_753),
.Y(n_983)
);

NAND2xp33_ASAP7_75t_L g984 ( 
.A(n_592),
.B(n_641),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_640),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_719),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_721),
.B(n_722),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_577),
.B(n_662),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_577),
.B(n_662),
.Y(n_989)
);

INVx4_ASAP7_75t_L g990 ( 
.A(n_581),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_734),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_599),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_759),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_586),
.B(n_587),
.Y(n_994)
);

BUFx4f_ASAP7_75t_L g995 ( 
.A(n_600),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_763),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_736),
.A2(n_758),
.B1(n_749),
.B2(n_743),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_739),
.A2(n_781),
.B1(n_797),
.B2(n_766),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_669),
.B(n_703),
.Y(n_999)
);

BUFx10_ASAP7_75t_L g1000 ( 
.A(n_602),
.Y(n_1000)
);

OR2x6_ASAP7_75t_L g1001 ( 
.A(n_589),
.B(n_604),
.Y(n_1001)
);

OR2x6_ASAP7_75t_L g1002 ( 
.A(n_608),
.B(n_609),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_785),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_767),
.Y(n_1004)
);

AND2x2_ASAP7_75t_SL g1005 ( 
.A(n_669),
.B(n_782),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_771),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_773),
.A2(n_795),
.B1(n_793),
.B2(n_789),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_788),
.Y(n_1008)
);

NAND2xp33_ASAP7_75t_L g1009 ( 
.A(n_631),
.B(n_612),
.Y(n_1009)
);

INVxp67_ASAP7_75t_SL g1010 ( 
.A(n_611),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_774),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_776),
.A2(n_800),
.B1(n_784),
.B2(n_798),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_777),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_625),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_778),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_779),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_787),
.B(n_799),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_603),
.Y(n_1018)
);

INVxp67_ASAP7_75t_SL g1019 ( 
.A(n_617),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_618),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_621),
.B(n_623),
.Y(n_1021)
);

AND2x2_ASAP7_75t_SL g1022 ( 
.A(n_703),
.B(n_782),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_503),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_505),
.Y(n_1024)
);

NOR2x1p5_ASAP7_75t_L g1025 ( 
.A(n_622),
.B(n_626),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_723),
.B(n_754),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_506),
.Y(n_1027)
);

INVxp33_ASAP7_75t_L g1028 ( 
.A(n_796),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_565),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_569),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_510),
.B(n_516),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_522),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_723),
.B(n_754),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_636),
.A2(n_654),
.B1(n_664),
.B2(n_802),
.Y(n_1034)
);

OAI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_636),
.A2(n_620),
.B1(n_651),
.B2(n_648),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_555),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_591),
.A2(n_358),
.B1(n_644),
.B2(n_560),
.Y(n_1037)
);

NAND3xp33_ASAP7_75t_L g1038 ( 
.A(n_780),
.B(n_486),
.C(n_455),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_494),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_497),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_678),
.A2(n_647),
.B1(n_620),
.B2(n_596),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_497),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_527),
.B(n_288),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_495),
.Y(n_1044)
);

BUFx4f_ASAP7_75t_L g1045 ( 
.A(n_667),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_495),
.Y(n_1046)
);

BUFx4f_ASAP7_75t_L g1047 ( 
.A(n_667),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_494),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_495),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_494),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_495),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_644),
.A2(n_358),
.B1(n_560),
.B2(n_408),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_495),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_495),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_494),
.Y(n_1055)
);

INVxp67_ASAP7_75t_SL g1056 ( 
.A(n_504),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_495),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_648),
.B(n_651),
.Y(n_1058)
);

OR2x6_ASAP7_75t_L g1059 ( 
.A(n_497),
.B(n_645),
.Y(n_1059)
);

NAND2xp33_ASAP7_75t_SL g1060 ( 
.A(n_559),
.B(n_455),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_495),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_715),
.B(n_726),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_495),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_527),
.B(n_288),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_648),
.B(n_651),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_648),
.B(n_651),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_504),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_678),
.A2(n_647),
.B1(n_620),
.B2(n_596),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_648),
.B(n_651),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_527),
.B(n_288),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_494),
.Y(n_1071)
);

BUFx10_ASAP7_75t_L g1072 ( 
.A(n_568),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_494),
.Y(n_1073)
);

NAND2xp33_ASAP7_75t_SL g1074 ( 
.A(n_559),
.B(n_455),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_495),
.Y(n_1075)
);

AND2x6_ASAP7_75t_L g1076 ( 
.A(n_644),
.B(n_642),
.Y(n_1076)
);

NAND2xp33_ASAP7_75t_L g1077 ( 
.A(n_642),
.B(n_455),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_542),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_667),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_495),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_670),
.B(n_673),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_495),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_494),
.Y(n_1083)
);

BUFx10_ASAP7_75t_L g1084 ( 
.A(n_568),
.Y(n_1084)
);

OR2x6_ASAP7_75t_L g1085 ( 
.A(n_497),
.B(n_645),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_494),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_670),
.B(n_673),
.Y(n_1087)
);

BUFx4f_ASAP7_75t_L g1088 ( 
.A(n_667),
.Y(n_1088)
);

AO22x2_ASAP7_75t_L g1089 ( 
.A1(n_633),
.A2(n_408),
.B1(n_291),
.B2(n_459),
.Y(n_1089)
);

NAND3xp33_ASAP7_75t_L g1090 ( 
.A(n_780),
.B(n_486),
.C(n_455),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_670),
.B(n_673),
.Y(n_1091)
);

INVx4_ASAP7_75t_L g1092 ( 
.A(n_497),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_494),
.Y(n_1093)
);

INVxp67_ASAP7_75t_SL g1094 ( 
.A(n_504),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_495),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_670),
.B(n_673),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_495),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_761),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_527),
.B(n_288),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_527),
.B(n_288),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_495),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_670),
.B(n_673),
.Y(n_1102)
);

NAND2xp33_ASAP7_75t_SL g1103 ( 
.A(n_559),
.B(n_455),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_538),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_495),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_644),
.A2(n_358),
.B1(n_560),
.B2(n_408),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_527),
.B(n_288),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_495),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_495),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_539),
.A2(n_673),
.B1(n_718),
.B2(n_670),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_497),
.Y(n_1111)
);

INVx4_ASAP7_75t_L g1112 ( 
.A(n_497),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_494),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_495),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_670),
.B(n_673),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_494),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_542),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_497),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_648),
.B(n_651),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_527),
.B(n_288),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_648),
.B(n_651),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_648),
.B(n_651),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_657),
.B(n_459),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_761),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_495),
.Y(n_1125)
);

BUFx4f_ASAP7_75t_L g1126 ( 
.A(n_667),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_497),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_670),
.B(n_673),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_670),
.B(n_673),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_497),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_497),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_542),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_670),
.B(n_673),
.Y(n_1133)
);

INVx4_ASAP7_75t_L g1134 ( 
.A(n_497),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_542),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_495),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_542),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_495),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_657),
.B(n_459),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_497),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_497),
.Y(n_1141)
);

CKINVDCx20_ASAP7_75t_R g1142 ( 
.A(n_542),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_542),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_667),
.Y(n_1144)
);

NAND2xp33_ASAP7_75t_R g1145 ( 
.A(n_667),
.B(n_393),
.Y(n_1145)
);

CKINVDCx20_ASAP7_75t_R g1146 ( 
.A(n_542),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_670),
.B(n_673),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_657),
.B(n_672),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_494),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_497),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_678),
.A2(n_647),
.B1(n_620),
.B2(n_596),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_495),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_497),
.Y(n_1153)
);

AND2x6_ASAP7_75t_L g1154 ( 
.A(n_644),
.B(n_642),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_670),
.B(n_673),
.Y(n_1155)
);

INVx1_ASAP7_75t_SL g1156 ( 
.A(n_761),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_644),
.A2(n_358),
.B1(n_560),
.B2(n_408),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_542),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_497),
.Y(n_1159)
);

NAND2xp33_ASAP7_75t_L g1160 ( 
.A(n_642),
.B(n_455),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_504),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_670),
.B(n_673),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_494),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_678),
.A2(n_647),
.B1(n_620),
.B2(n_596),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_527),
.B(n_288),
.Y(n_1165)
);

INVx4_ASAP7_75t_L g1166 ( 
.A(n_497),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_542),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_542),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_495),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_494),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_495),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_667),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_497),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_497),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_542),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_497),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_527),
.B(n_288),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_657),
.B(n_459),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_495),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_495),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_667),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_495),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_497),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_497),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_780),
.B(n_486),
.C(n_455),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_670),
.B(n_673),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_497),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_761),
.Y(n_1188)
);

AND2x6_ASAP7_75t_L g1189 ( 
.A(n_644),
.B(n_642),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_657),
.B(n_672),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_494),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_670),
.B(n_673),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_527),
.B(n_288),
.Y(n_1193)
);

BUFx10_ASAP7_75t_L g1194 ( 
.A(n_568),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_495),
.Y(n_1195)
);

NAND2xp33_ASAP7_75t_SL g1196 ( 
.A(n_559),
.B(n_455),
.Y(n_1196)
);

NAND2xp33_ASAP7_75t_SL g1197 ( 
.A(n_559),
.B(n_455),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_495),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_495),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_495),
.Y(n_1200)
);

AND2x2_ASAP7_75t_SL g1201 ( 
.A(n_644),
.B(n_475),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_648),
.B(n_651),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_494),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_495),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_497),
.Y(n_1205)
);

INVx4_ASAP7_75t_L g1206 ( 
.A(n_497),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_495),
.Y(n_1207)
);

INVx2_ASAP7_75t_SL g1208 ( 
.A(n_667),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_542),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_539),
.A2(n_673),
.B1(n_718),
.B2(n_670),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_527),
.B(n_288),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_657),
.B(n_672),
.Y(n_1212)
);

OAI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_620),
.A2(n_651),
.B1(n_658),
.B2(n_648),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_648),
.B(n_651),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_494),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_495),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_494),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_495),
.Y(n_1218)
);

INVx4_ASAP7_75t_L g1219 ( 
.A(n_497),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_542),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_494),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_504),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_494),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_670),
.B(n_673),
.Y(n_1224)
);

BUFx4f_ASAP7_75t_L g1225 ( 
.A(n_667),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_497),
.Y(n_1226)
);

NAND3xp33_ASAP7_75t_L g1227 ( 
.A(n_780),
.B(n_486),
.C(n_455),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_648),
.B(n_651),
.Y(n_1228)
);

BUFx4f_ASAP7_75t_L g1229 ( 
.A(n_667),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_497),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_542),
.Y(n_1231)
);

INVx4_ASAP7_75t_L g1232 ( 
.A(n_497),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_657),
.B(n_672),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_495),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_678),
.A2(n_647),
.B1(n_620),
.B2(n_596),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_648),
.B(n_651),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_494),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_494),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_497),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_495),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_495),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_497),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_494),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_495),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_497),
.Y(n_1245)
);

BUFx4f_ASAP7_75t_L g1246 ( 
.A(n_667),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_539),
.A2(n_673),
.B1(n_718),
.B2(n_670),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_761),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_497),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1043),
.B(n_1064),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_820),
.B(n_809),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_816),
.A2(n_1052),
.B1(n_1157),
.B2(n_1106),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_831),
.B(n_833),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_1098),
.Y(n_1254)
);

NAND3xp33_ASAP7_75t_L g1255 ( 
.A(n_1070),
.B(n_1100),
.C(n_1099),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_826),
.A2(n_1068),
.B(n_1151),
.C(n_1041),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_817),
.B(n_811),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1123),
.B(n_1139),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_848),
.B(n_1045),
.Y(n_1259)
);

NAND2x1_ASAP7_75t_L g1260 ( 
.A(n_982),
.B(n_822),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1107),
.B(n_1120),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_804),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1047),
.B(n_1088),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1081),
.B(n_1087),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_889),
.Y(n_1265)
);

INVxp67_ASAP7_75t_L g1266 ( 
.A(n_856),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1032),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1091),
.B(n_1096),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_808),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_834),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_891),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1102),
.B(n_1115),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_SL g1273 ( 
.A(n_1126),
.B(n_1225),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1165),
.B(n_1177),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1229),
.B(n_1246),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_837),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1038),
.B(n_1090),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_899),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1185),
.B(n_1227),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1193),
.B(n_1211),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1164),
.A2(n_1235),
.B(n_859),
.C(n_1210),
.Y(n_1281)
);

OR2x6_ASAP7_75t_L g1282 ( 
.A(n_818),
.B(n_806),
.Y(n_1282)
);

NAND3xp33_ASAP7_75t_L g1283 ( 
.A(n_1110),
.B(n_1247),
.C(n_1160),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1128),
.B(n_1129),
.Y(n_1284)
);

NAND2xp33_ASAP7_75t_L g1285 ( 
.A(n_865),
.B(n_822),
.Y(n_1285)
);

XOR2x2_ASAP7_75t_L g1286 ( 
.A(n_1201),
.B(n_832),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_866),
.B(n_900),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1133),
.B(n_1147),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1148),
.B(n_1190),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1155),
.B(n_1162),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1186),
.B(n_1192),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_866),
.B(n_878),
.Y(n_1292)
);

BUFx8_ASAP7_75t_L g1293 ( 
.A(n_857),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_866),
.B(n_1104),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_910),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1224),
.B(n_1212),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1233),
.B(n_974),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1104),
.B(n_1178),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_813),
.B(n_823),
.Y(n_1299)
);

OR2x6_ASAP7_75t_L g1300 ( 
.A(n_818),
.B(n_854),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_913),
.Y(n_1301)
);

INVx3_ASAP7_75t_L g1302 ( 
.A(n_982),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_842),
.B(n_824),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1058),
.B(n_1065),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1066),
.B(n_1069),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1119),
.B(n_1121),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1122),
.B(n_1202),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1214),
.B(n_1228),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1236),
.B(n_828),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_810),
.B(n_812),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1213),
.B(n_836),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_810),
.B(n_812),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_870),
.B(n_873),
.Y(n_1313)
);

BUFx5_ASAP7_75t_L g1314 ( 
.A(n_982),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_853),
.B(n_850),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_838),
.B(n_840),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_889),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1067),
.B(n_1161),
.Y(n_1318)
);

NOR3xp33_ASAP7_75t_L g1319 ( 
.A(n_1060),
.B(n_1103),
.C(n_1074),
.Y(n_1319)
);

INVxp67_ASAP7_75t_L g1320 ( 
.A(n_1222),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1124),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_918),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1062),
.B(n_1111),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_1056),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_843),
.B(n_844),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_846),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1094),
.B(n_907),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1062),
.B(n_1111),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_847),
.B(n_849),
.Y(n_1329)
);

NAND2xp33_ASAP7_75t_SL g1330 ( 
.A(n_1145),
.B(n_892),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_882),
.B(n_1079),
.Y(n_1331)
);

OR2x6_ASAP7_75t_L g1332 ( 
.A(n_1144),
.B(n_1172),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_879),
.B(n_1181),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_851),
.B(n_860),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_957),
.A2(n_984),
.B(n_969),
.Y(n_1335)
);

NAND2xp33_ASAP7_75t_L g1336 ( 
.A(n_822),
.B(n_1076),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1208),
.B(n_926),
.Y(n_1337)
);

NOR2xp67_ASAP7_75t_L g1338 ( 
.A(n_1135),
.B(n_1158),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_861),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_864),
.Y(n_1340)
);

AOI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1196),
.A2(n_1197),
.B1(n_1077),
.B2(n_805),
.Y(n_1341)
);

INVxp67_ASAP7_75t_L g1342 ( 
.A(n_1156),
.Y(n_1342)
);

INVxp67_ASAP7_75t_L g1343 ( 
.A(n_1188),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1089),
.A2(n_877),
.B1(n_1037),
.B2(n_1076),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1017),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1248),
.B(n_904),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1118),
.B(n_1130),
.Y(n_1347)
);

BUFx2_ASAP7_75t_R g1348 ( 
.A(n_1209),
.Y(n_1348)
);

NAND2xp33_ASAP7_75t_SL g1349 ( 
.A(n_943),
.B(n_1132),
.Y(n_1349)
);

INVx3_ASAP7_75t_L g1350 ( 
.A(n_911),
.Y(n_1350)
);

AND2x2_ASAP7_75t_SL g1351 ( 
.A(n_871),
.B(n_976),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_867),
.B(n_869),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1089),
.A2(n_959),
.B1(n_1154),
.B2(n_1076),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1044),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1072),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_912),
.B(n_1020),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1118),
.B(n_1130),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1150),
.B(n_1159),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_807),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1150),
.B(n_1159),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_888),
.B(n_972),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1046),
.B(n_1049),
.Y(n_1362)
);

INVx4_ASAP7_75t_L g1363 ( 
.A(n_881),
.Y(n_1363)
);

INVxp33_ASAP7_75t_L g1364 ( 
.A(n_1173),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1051),
.Y(n_1365)
);

INVx8_ASAP7_75t_L g1366 ( 
.A(n_896),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1053),
.B(n_1054),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_819),
.Y(n_1368)
);

INVx2_ASAP7_75t_SL g1369 ( 
.A(n_1072),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_815),
.Y(n_1370)
);

BUFx4_ASAP7_75t_L g1371 ( 
.A(n_875),
.Y(n_1371)
);

INVxp67_ASAP7_75t_L g1372 ( 
.A(n_1078),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_803),
.B(n_1059),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_911),
.Y(n_1374)
);

AND2x6_ASAP7_75t_SL g1375 ( 
.A(n_803),
.B(n_1059),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1057),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1020),
.B(n_1023),
.Y(n_1377)
);

INVxp33_ASAP7_75t_L g1378 ( 
.A(n_1173),
.Y(n_1378)
);

NOR2x1p5_ASAP7_75t_L g1379 ( 
.A(n_1231),
.B(n_1117),
.Y(n_1379)
);

NOR3xp33_ASAP7_75t_L g1380 ( 
.A(n_931),
.B(n_898),
.C(n_980),
.Y(n_1380)
);

BUFx8_ASAP7_75t_L g1381 ( 
.A(n_1137),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1061),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1063),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1075),
.B(n_1080),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1084),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1082),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1174),
.B(n_1183),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1085),
.B(n_995),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_SL g1389 ( 
.A(n_1174),
.B(n_1183),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1095),
.B(n_1097),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1101),
.B(n_1105),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1108),
.B(n_1109),
.Y(n_1392)
);

NAND2xp33_ASAP7_75t_L g1393 ( 
.A(n_1154),
.B(n_1189),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_908),
.B(n_992),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1114),
.Y(n_1395)
);

BUFx5_ASAP7_75t_L g1396 ( 
.A(n_1036),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1125),
.B(n_1136),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1138),
.B(n_1152),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_821),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_825),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1169),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1014),
.B(n_1142),
.Y(n_1402)
);

NAND3xp33_ASAP7_75t_L g1403 ( 
.A(n_1009),
.B(n_994),
.C(n_938),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1184),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_827),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1085),
.B(n_1143),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1171),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_1184),
.B(n_1205),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1179),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1146),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1180),
.B(n_1182),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1195),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_1084),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1198),
.B(n_1199),
.Y(n_1414)
);

NAND2xp33_ASAP7_75t_L g1415 ( 
.A(n_1154),
.B(n_1189),
.Y(n_1415)
);

NAND3xp33_ASAP7_75t_SL g1416 ( 
.A(n_894),
.B(n_884),
.C(n_985),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1167),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1200),
.B(n_1204),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_SL g1419 ( 
.A(n_1194),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1207),
.B(n_1216),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1218),
.B(n_1234),
.Y(n_1421)
);

BUFx5_ASAP7_75t_L g1422 ( 
.A(n_1005),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1240),
.B(n_1241),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1205),
.B(n_1230),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1230),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1244),
.B(n_1189),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_835),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_845),
.Y(n_1428)
);

INVxp33_ASAP7_75t_L g1429 ( 
.A(n_939),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_928),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_939),
.B(n_945),
.Y(n_1431)
);

NAND2xp33_ASAP7_75t_L g1432 ( 
.A(n_945),
.B(n_925),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_855),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_897),
.B(n_830),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_944),
.B(n_981),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_990),
.B(n_941),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_916),
.B(n_909),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_SL g1438 ( 
.A(n_863),
.B(n_872),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_956),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1019),
.B(n_921),
.Y(n_1440)
);

INVx4_ASAP7_75t_L g1441 ( 
.A(n_1194),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_947),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_858),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_927),
.B(n_933),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_862),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_876),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_880),
.Y(n_1447)
);

NOR2xp67_ASAP7_75t_L g1448 ( 
.A(n_1092),
.B(n_1112),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_953),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_958),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_L g1451 ( 
.A(n_964),
.B(n_998),
.C(n_997),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_883),
.Y(n_1452)
);

INVx5_ASAP7_75t_L g1453 ( 
.A(n_874),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_SL g1454 ( 
.A(n_1131),
.B(n_1134),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1168),
.B(n_1175),
.Y(n_1455)
);

AND2x6_ASAP7_75t_SL g1456 ( 
.A(n_914),
.B(n_919),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_935),
.B(n_936),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_942),
.B(n_946),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1220),
.B(n_930),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_886),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_887),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_951),
.B(n_952),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_963),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1166),
.B(n_1206),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_923),
.B(n_955),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_932),
.B(n_874),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_978),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_841),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_893),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_960),
.B(n_961),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_814),
.B(n_829),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_962),
.B(n_966),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_839),
.B(n_885),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_987),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_971),
.B(n_979),
.Y(n_1475)
);

INVxp67_ASAP7_75t_L g1476 ( 
.A(n_937),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1026),
.A2(n_988),
.B(n_1033),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_895),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1040),
.B(n_1042),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_901),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_986),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1219),
.B(n_1226),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_902),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_991),
.B(n_1004),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1006),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1127),
.B(n_1140),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_956),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_956),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_905),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1141),
.B(n_1153),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1011),
.B(n_1013),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1025),
.B(n_1232),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1015),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1176),
.B(n_1187),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1239),
.B(n_1242),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_906),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_L g1497 ( 
.A(n_1007),
.B(n_1012),
.C(n_1021),
.Y(n_1497)
);

BUFx6f_ASAP7_75t_L g1498 ( 
.A(n_920),
.Y(n_1498)
);

INVxp67_ASAP7_75t_L g1499 ( 
.A(n_977),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_920),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1016),
.B(n_1024),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1027),
.B(n_1028),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_922),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_929),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_940),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1249),
.B(n_903),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_948),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_954),
.B(n_1029),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1001),
.B(n_1002),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_970),
.B(n_1008),
.Y(n_1510)
);

NOR3xp33_ASAP7_75t_L g1511 ( 
.A(n_965),
.B(n_890),
.C(n_967),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_973),
.B(n_1223),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_977),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1018),
.B(n_1245),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1031),
.B(n_868),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_915),
.B(n_917),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_975),
.B(n_1048),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_983),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_993),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_996),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_SL g1521 ( 
.A(n_1035),
.B(n_968),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1003),
.B(n_1071),
.Y(n_1522)
);

INVxp67_ASAP7_75t_L g1523 ( 
.A(n_934),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_949),
.A2(n_852),
.B1(n_1001),
.B2(n_1002),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1039),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1050),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1055),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1073),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1083),
.B(n_1116),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1243),
.B(n_1113),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1000),
.Y(n_1531)
);

NAND3xp33_ASAP7_75t_L g1532 ( 
.A(n_950),
.B(n_1034),
.C(n_989),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1086),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1000),
.B(n_1170),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1093),
.B(n_1191),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1149),
.B(n_1203),
.Y(n_1536)
);

NOR3xp33_ASAP7_75t_L g1537 ( 
.A(n_1163),
.B(n_1215),
.C(n_1237),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1217),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1221),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1238),
.B(n_1030),
.Y(n_1540)
);

CKINVDCx20_ASAP7_75t_R g1541 ( 
.A(n_999),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1010),
.B(n_1022),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_924),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_924),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1043),
.B(n_455),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_816),
.A2(n_486),
.B1(n_455),
.B2(n_393),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1098),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1032),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1043),
.B(n_455),
.Y(n_1549)
);

NOR3xp33_ASAP7_75t_L g1550 ( 
.A(n_1043),
.B(n_780),
.C(n_1064),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_817),
.B(n_395),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1032),
.Y(n_1552)
);

INVx2_ASAP7_75t_SL g1553 ( 
.A(n_848),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_SL g1554 ( 
.A(n_1132),
.B(n_455),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1032),
.Y(n_1555)
);

AO221x1_ASAP7_75t_L g1556 ( 
.A1(n_1213),
.A2(n_1089),
.B1(n_1035),
.B2(n_408),
.C(n_407),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_804),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1032),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_804),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_820),
.B(n_809),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_820),
.B(n_809),
.Y(n_1561)
);

INVx3_ASAP7_75t_L g1562 ( 
.A(n_982),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_820),
.B(n_809),
.Y(n_1563)
);

INVx2_ASAP7_75t_SL g1564 ( 
.A(n_848),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1032),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1032),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1032),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_817),
.B(n_395),
.Y(n_1568)
);

NAND2x1_ASAP7_75t_L g1569 ( 
.A(n_982),
.B(n_822),
.Y(n_1569)
);

INVxp67_ASAP7_75t_L g1570 ( 
.A(n_856),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_817),
.B(n_395),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_804),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_817),
.B(n_395),
.Y(n_1573)
);

NOR3xp33_ASAP7_75t_L g1574 ( 
.A(n_1043),
.B(n_780),
.C(n_1064),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1148),
.B(n_657),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_820),
.B(n_809),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1032),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_820),
.B(n_809),
.Y(n_1578)
);

INVx2_ASAP7_75t_SL g1579 ( 
.A(n_848),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_804),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1104),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_817),
.B(n_395),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1032),
.Y(n_1583)
);

INVxp67_ASAP7_75t_L g1584 ( 
.A(n_856),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_817),
.B(n_395),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_817),
.B(n_395),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1032),
.Y(n_1587)
);

NAND3xp33_ASAP7_75t_L g1588 ( 
.A(n_1052),
.B(n_1157),
.C(n_1106),
.Y(n_1588)
);

NOR2x1p5_ASAP7_75t_L g1589 ( 
.A(n_1135),
.B(n_477),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_817),
.B(n_395),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1032),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1098),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1043),
.B(n_455),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_804),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1032),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_804),
.Y(n_1596)
);

INVxp33_ASAP7_75t_L g1597 ( 
.A(n_816),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1032),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_889),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1043),
.B(n_455),
.Y(n_1600)
);

NOR2xp67_ASAP7_75t_L g1601 ( 
.A(n_1038),
.B(n_446),
.Y(n_1601)
);

NAND2xp33_ASAP7_75t_SL g1602 ( 
.A(n_1145),
.B(n_455),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1032),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1032),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_817),
.B(n_395),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1032),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_820),
.B(n_809),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1043),
.B(n_455),
.Y(n_1608)
);

AND2x6_ASAP7_75t_L g1609 ( 
.A(n_1041),
.B(n_644),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1032),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_804),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1052),
.A2(n_358),
.B1(n_1157),
.B2(n_1106),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1032),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_817),
.B(n_395),
.Y(n_1614)
);

NOR2xp67_ASAP7_75t_L g1615 ( 
.A(n_1038),
.B(n_446),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1148),
.B(n_657),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1135),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_820),
.B(n_809),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1043),
.B(n_455),
.Y(n_1619)
);

BUFx6f_ASAP7_75t_L g1620 ( 
.A(n_889),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_817),
.B(n_395),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1032),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_848),
.Y(n_1623)
);

INVx3_ASAP7_75t_L g1624 ( 
.A(n_982),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_817),
.B(n_395),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_820),
.B(n_809),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_817),
.B(n_395),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_820),
.B(n_809),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_820),
.B(n_809),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1032),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_820),
.B(n_809),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1032),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_820),
.B(n_809),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_820),
.B(n_809),
.Y(n_1634)
);

NOR3xp33_ASAP7_75t_L g1635 ( 
.A(n_1043),
.B(n_780),
.C(n_1064),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1032),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_804),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_820),
.B(n_809),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1032),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1043),
.B(n_455),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_820),
.B(n_809),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_817),
.B(n_395),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_804),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1032),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_804),
.Y(n_1645)
);

BUFx5_ASAP7_75t_L g1646 ( 
.A(n_982),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_820),
.B(n_809),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_804),
.Y(n_1648)
);

XOR2xp5_ASAP7_75t_L g1649 ( 
.A(n_1132),
.B(n_542),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_820),
.B(n_809),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1043),
.B(n_455),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_848),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_817),
.B(n_395),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1032),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1148),
.B(n_657),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1043),
.B(n_455),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_804),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1052),
.A2(n_358),
.B1(n_1157),
.B2(n_1106),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_817),
.B(n_395),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_804),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_820),
.B(n_809),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_804),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_804),
.Y(n_1663)
);

BUFx2_ASAP7_75t_L g1664 ( 
.A(n_1104),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1043),
.B(n_455),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_889),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1032),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_820),
.B(n_809),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_817),
.B(n_395),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_804),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_820),
.B(n_809),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_804),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_804),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1043),
.B(n_455),
.Y(n_1674)
);

BUFx6f_ASAP7_75t_L g1675 ( 
.A(n_889),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_820),
.B(n_809),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1032),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_804),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_SL g1679 ( 
.A(n_1072),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1043),
.B(n_455),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1032),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1032),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1032),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_848),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_804),
.Y(n_1685)
);

OR2x6_ASAP7_75t_L g1686 ( 
.A(n_818),
.B(n_806),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1104),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1043),
.B(n_455),
.Y(n_1688)
);

INVxp67_ASAP7_75t_L g1689 ( 
.A(n_856),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_817),
.B(n_395),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_820),
.B(n_809),
.Y(n_1691)
);

INVx3_ASAP7_75t_L g1692 ( 
.A(n_982),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_804),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_804),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_820),
.B(n_809),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1032),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_820),
.B(n_809),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_856),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_817),
.B(n_395),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_804),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1148),
.B(n_657),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1032),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_820),
.B(n_809),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1032),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_804),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_1135),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_817),
.B(n_395),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1043),
.B(n_455),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_856),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_820),
.B(n_809),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_820),
.B(n_809),
.Y(n_1711)
);

NOR3xp33_ASAP7_75t_L g1712 ( 
.A(n_1043),
.B(n_780),
.C(n_1064),
.Y(n_1712)
);

AND2x6_ASAP7_75t_L g1713 ( 
.A(n_1041),
.B(n_644),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_804),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_820),
.B(n_809),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_820),
.B(n_809),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_820),
.B(n_809),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_804),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_804),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_804),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1043),
.B(n_455),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_804),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_804),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_820),
.B(n_809),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1148),
.B(n_657),
.Y(n_1725)
);

INVx2_ASAP7_75t_SL g1726 ( 
.A(n_848),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_820),
.B(n_809),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_817),
.B(n_395),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_820),
.B(n_809),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1032),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_820),
.B(n_809),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_816),
.A2(n_486),
.B1(n_455),
.B2(n_393),
.Y(n_1732)
);

NAND2xp33_ASAP7_75t_L g1733 ( 
.A(n_865),
.B(n_455),
.Y(n_1733)
);

NAND3xp33_ASAP7_75t_L g1734 ( 
.A(n_1052),
.B(n_1157),
.C(n_1106),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_804),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1148),
.B(n_657),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_SL g1737 ( 
.A(n_817),
.B(n_395),
.Y(n_1737)
);

BUFx6f_ASAP7_75t_L g1738 ( 
.A(n_889),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_820),
.B(n_809),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1148),
.B(n_657),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_820),
.B(n_809),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_820),
.B(n_809),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_817),
.B(n_395),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1110),
.A2(n_1247),
.B(n_1210),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_820),
.B(n_809),
.Y(n_1745)
);

NOR2xp67_ASAP7_75t_L g1746 ( 
.A(n_1038),
.B(n_446),
.Y(n_1746)
);

CKINVDCx20_ASAP7_75t_R g1747 ( 
.A(n_1132),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1043),
.B(n_455),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_SL g1749 ( 
.A(n_817),
.B(n_395),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_820),
.B(n_809),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1032),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1043),
.B(n_455),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1032),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_804),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1032),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_820),
.B(n_809),
.Y(n_1756)
);

NOR2xp67_ASAP7_75t_L g1757 ( 
.A(n_1038),
.B(n_446),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1148),
.B(n_657),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_804),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_804),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1148),
.B(n_657),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_SL g1762 ( 
.A(n_1072),
.Y(n_1762)
);

INVxp67_ASAP7_75t_L g1763 ( 
.A(n_856),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1043),
.B(n_455),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1032),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_820),
.B(n_809),
.Y(n_1766)
);

NOR2xp67_ASAP7_75t_L g1767 ( 
.A(n_1038),
.B(n_446),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1043),
.B(n_455),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_816),
.A2(n_486),
.B1(n_455),
.B2(n_393),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_804),
.Y(n_1770)
);

INVx2_ASAP7_75t_SL g1771 ( 
.A(n_848),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1043),
.B(n_455),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_804),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1032),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_804),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1032),
.Y(n_1776)
);

BUFx3_ASAP7_75t_L g1777 ( 
.A(n_818),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1043),
.B(n_455),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_804),
.Y(n_1779)
);

INVxp67_ASAP7_75t_L g1780 ( 
.A(n_856),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_804),
.Y(n_1781)
);

INVxp67_ASAP7_75t_L g1782 ( 
.A(n_856),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_820),
.B(n_809),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_817),
.B(n_395),
.Y(n_1784)
);

NAND2xp33_ASAP7_75t_L g1785 ( 
.A(n_865),
.B(n_455),
.Y(n_1785)
);

NAND2x1_ASAP7_75t_L g1786 ( 
.A(n_982),
.B(n_822),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_SL g1787 ( 
.A(n_1132),
.B(n_455),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_817),
.B(n_395),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_804),
.Y(n_1789)
);

INVxp33_ASAP7_75t_L g1790 ( 
.A(n_816),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1043),
.B(n_455),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_810),
.B(n_812),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_820),
.B(n_809),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_804),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1043),
.B(n_455),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1043),
.B(n_455),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1032),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_820),
.B(n_809),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1032),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1032),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_804),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_817),
.B(n_395),
.Y(n_1802)
);

BUFx6f_ASAP7_75t_L g1803 ( 
.A(n_889),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_804),
.Y(n_1804)
);

OR2x6_ASAP7_75t_L g1805 ( 
.A(n_818),
.B(n_806),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_804),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_820),
.B(n_809),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_820),
.B(n_809),
.Y(n_1808)
);

INVxp67_ASAP7_75t_L g1809 ( 
.A(n_856),
.Y(n_1809)
);

BUFx5_ASAP7_75t_L g1810 ( 
.A(n_982),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1032),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_820),
.B(n_809),
.Y(n_1812)
);

INVx2_ASAP7_75t_SL g1813 ( 
.A(n_848),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1032),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1032),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1032),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_820),
.B(n_809),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1032),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_804),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_804),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1032),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_820),
.B(n_809),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_856),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1032),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_820),
.B(n_809),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_820),
.B(n_809),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_804),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1032),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_820),
.B(n_809),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_817),
.B(n_395),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_817),
.B(n_395),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1032),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_817),
.B(n_395),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_817),
.B(n_395),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_817),
.B(n_395),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_804),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_804),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1032),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_820),
.B(n_809),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_820),
.B(n_809),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1032),
.Y(n_1841)
);

NAND3xp33_ASAP7_75t_L g1842 ( 
.A(n_1052),
.B(n_1157),
.C(n_1106),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_817),
.B(n_395),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_820),
.B(n_809),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_889),
.Y(n_1845)
);

BUFx6f_ASAP7_75t_SL g1846 ( 
.A(n_1072),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_817),
.B(n_395),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_804),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_804),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1052),
.A2(n_358),
.B1(n_1157),
.B2(n_1106),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_820),
.B(n_809),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_820),
.B(n_809),
.Y(n_1852)
);

AOI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_816),
.A2(n_486),
.B1(n_455),
.B2(n_393),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_804),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_820),
.B(n_809),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_804),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_817),
.B(n_395),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_804),
.Y(n_1858)
);

INVxp67_ASAP7_75t_L g1859 ( 
.A(n_856),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1032),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_820),
.B(n_809),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_L g1862 ( 
.A(n_1043),
.B(n_455),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1032),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_804),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_820),
.B(n_809),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_SL g1866 ( 
.A(n_817),
.B(n_395),
.Y(n_1866)
);

NOR2xp67_ASAP7_75t_L g1867 ( 
.A(n_1038),
.B(n_446),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_820),
.B(n_809),
.Y(n_1868)
);

INVxp67_ASAP7_75t_L g1869 ( 
.A(n_856),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_820),
.B(n_809),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_820),
.B(n_809),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1043),
.B(n_455),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_820),
.B(n_809),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_820),
.B(n_809),
.Y(n_1874)
);

OAI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1052),
.A2(n_1106),
.B1(n_1157),
.B2(n_539),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_817),
.B(n_395),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_820),
.B(n_809),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_817),
.B(n_395),
.Y(n_1878)
);

NOR3xp33_ASAP7_75t_L g1879 ( 
.A(n_1043),
.B(n_780),
.C(n_1064),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_SL g1880 ( 
.A(n_817),
.B(n_395),
.Y(n_1880)
);

BUFx6f_ASAP7_75t_SL g1881 ( 
.A(n_1072),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1032),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1123),
.B(n_459),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_817),
.B(n_395),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_804),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_SL g1886 ( 
.A(n_817),
.B(n_395),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1052),
.A2(n_358),
.B1(n_1157),
.B2(n_1106),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1032),
.Y(n_1888)
);

NOR3xp33_ASAP7_75t_L g1889 ( 
.A(n_1043),
.B(n_780),
.C(n_1064),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_804),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_804),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_804),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1148),
.B(n_657),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_817),
.B(n_395),
.Y(n_1894)
);

INVx2_ASAP7_75t_SL g1895 ( 
.A(n_848),
.Y(n_1895)
);

INVx4_ASAP7_75t_L g1896 ( 
.A(n_818),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_810),
.B(n_812),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_820),
.B(n_809),
.Y(n_1898)
);

AO221x1_ASAP7_75t_L g1899 ( 
.A1(n_1213),
.A2(n_1089),
.B1(n_1035),
.B2(n_408),
.C(n_407),
.Y(n_1899)
);

NAND3xp33_ASAP7_75t_L g1900 ( 
.A(n_1052),
.B(n_1157),
.C(n_1106),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_820),
.B(n_809),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1032),
.Y(n_1902)
);

INVxp33_ASAP7_75t_L g1903 ( 
.A(n_816),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1032),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_1043),
.B(n_455),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_SL g1906 ( 
.A(n_817),
.B(n_395),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1043),
.B(n_455),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_804),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1032),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_820),
.B(n_809),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1043),
.B(n_455),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1032),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_804),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_820),
.B(n_809),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1052),
.A2(n_358),
.B1(n_1157),
.B2(n_1106),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_1135),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1043),
.B(n_455),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_817),
.B(n_395),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_820),
.B(n_809),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_SL g1920 ( 
.A(n_817),
.B(n_395),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1043),
.B(n_455),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_820),
.B(n_809),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1043),
.B(n_455),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1032),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1032),
.Y(n_1925)
);

BUFx5_ASAP7_75t_L g1926 ( 
.A(n_982),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1032),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1032),
.Y(n_1928)
);

OR2x6_ASAP7_75t_L g1929 ( 
.A(n_818),
.B(n_806),
.Y(n_1929)
);

NOR3xp33_ASAP7_75t_L g1930 ( 
.A(n_1043),
.B(n_780),
.C(n_1064),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1313),
.B(n_1251),
.Y(n_1931)
);

OAI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_1932)
);

AOI22xp33_ASAP7_75t_L g1933 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1734),
.B2(n_1842),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1560),
.B(n_1561),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1545),
.B(n_1549),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1543),
.Y(n_1936)
);

INVx3_ASAP7_75t_L g1937 ( 
.A(n_1260),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1563),
.B(n_1576),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1637),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1518),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1637),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1593),
.B(n_1600),
.Y(n_1942)
);

AOI22xp33_ASAP7_75t_L g1943 ( 
.A1(n_1588),
.A2(n_1900),
.B1(n_1850),
.B2(n_1658),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1311),
.B(n_1253),
.Y(n_1944)
);

HB1xp67_ASAP7_75t_L g1945 ( 
.A(n_1581),
.Y(n_1945)
);

AND2x4_ASAP7_75t_L g1946 ( 
.A(n_1792),
.B(n_1897),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1578),
.B(n_1607),
.Y(n_1947)
);

O2A1O1Ixp33_ASAP7_75t_L g1948 ( 
.A1(n_1875),
.A2(n_1744),
.B(n_1281),
.C(n_1255),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1518),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1618),
.B(n_1626),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1608),
.B(n_1619),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1453),
.Y(n_1952)
);

OAI22xp5_ASAP7_75t_SL g1953 ( 
.A1(n_1612),
.A2(n_1915),
.B1(n_1887),
.B2(n_1651),
.Y(n_1953)
);

AOI22xp33_ASAP7_75t_L g1954 ( 
.A1(n_1609),
.A2(n_1713),
.B1(n_1252),
.B2(n_1416),
.Y(n_1954)
);

O2A1O1Ixp33_ASAP7_75t_L g1955 ( 
.A1(n_1640),
.A2(n_1665),
.B(n_1674),
.C(n_1656),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1643),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1643),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1781),
.Y(n_1958)
);

AOI22xp33_ASAP7_75t_SL g1959 ( 
.A1(n_1609),
.A2(n_1713),
.B1(n_1309),
.B2(n_1435),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_SL g1960 ( 
.A(n_1628),
.B(n_1629),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1631),
.B(n_1633),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1634),
.B(n_1638),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1519),
.Y(n_1963)
);

OAI22xp5_ASAP7_75t_SL g1964 ( 
.A1(n_1680),
.A2(n_1721),
.B1(n_1748),
.B2(n_1688),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1264),
.B(n_1268),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1792),
.B(n_1897),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1272),
.B(n_1284),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_L g1968 ( 
.A(n_1708),
.B(n_1752),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1641),
.B(n_1647),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1747),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1283),
.A2(n_1661),
.B1(n_1668),
.B2(n_1650),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1304),
.B(n_1305),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1519),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1527),
.Y(n_1974)
);

AOI22xp33_ASAP7_75t_L g1975 ( 
.A1(n_1609),
.A2(n_1713),
.B1(n_1344),
.B2(n_1541),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1671),
.B(n_1676),
.Y(n_1976)
);

OAI22xp5_ASAP7_75t_SL g1977 ( 
.A1(n_1764),
.A2(n_1772),
.B1(n_1778),
.B2(n_1768),
.Y(n_1977)
);

AOI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1609),
.A2(n_1713),
.B1(n_1923),
.B2(n_1795),
.Y(n_1978)
);

NOR2xp33_ASAP7_75t_L g1979 ( 
.A(n_1791),
.B(n_1796),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1691),
.B(n_1695),
.Y(n_1980)
);

OAI22xp33_ASAP7_75t_L g1981 ( 
.A1(n_1697),
.A2(n_1703),
.B1(n_1711),
.B2(n_1710),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1781),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1862),
.B(n_1872),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1527),
.Y(n_1984)
);

AOI22xp33_ASAP7_75t_SL g1985 ( 
.A1(n_1351),
.A2(n_1285),
.B1(n_1451),
.B2(n_1905),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1306),
.Y(n_1986)
);

O2A1O1Ixp33_ASAP7_75t_L g1987 ( 
.A1(n_1907),
.A2(n_1917),
.B(n_1911),
.C(n_1921),
.Y(n_1987)
);

INVx1_ASAP7_75t_SL g1988 ( 
.A(n_1254),
.Y(n_1988)
);

AND2x6_ASAP7_75t_SL g1989 ( 
.A(n_1299),
.B(n_1402),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1715),
.B(n_1716),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1307),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1717),
.B(n_1724),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1308),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1481),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_L g1995 ( 
.A(n_1266),
.B(n_1570),
.Y(n_1995)
);

AO22x1_ASAP7_75t_L g1996 ( 
.A1(n_1550),
.A2(n_1574),
.B1(n_1712),
.B2(n_1635),
.Y(n_1996)
);

NOR2xp33_ASAP7_75t_L g1997 ( 
.A(n_1584),
.B(n_1689),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1288),
.B(n_1290),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1727),
.B(n_1729),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1731),
.B(n_1739),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1698),
.B(n_1709),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_SL g2002 ( 
.A(n_1741),
.B(n_1742),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1267),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_SL g2004 ( 
.A(n_1745),
.B(n_1750),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1548),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1756),
.B(n_1766),
.Y(n_2006)
);

INVx2_ASAP7_75t_SL g2007 ( 
.A(n_1453),
.Y(n_2007)
);

A2O1A1Ixp33_ASAP7_75t_SL g2008 ( 
.A1(n_1879),
.A2(n_1889),
.B(n_1930),
.C(n_1319),
.Y(n_2008)
);

A2O1A1Ixp33_ASAP7_75t_L g2009 ( 
.A1(n_1256),
.A2(n_1793),
.B(n_1798),
.C(n_1783),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1552),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1807),
.B(n_1808),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1812),
.B(n_1817),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1822),
.B(n_1825),
.Y(n_2013)
);

AOI22xp33_ASAP7_75t_L g2014 ( 
.A1(n_1497),
.A2(n_1852),
.B1(n_1901),
.B2(n_1826),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1555),
.Y(n_2015)
);

A2O1A1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_1829),
.A2(n_1840),
.B(n_1844),
.C(n_1839),
.Y(n_2016)
);

OR2x2_ASAP7_75t_L g2017 ( 
.A(n_1258),
.B(n_1664),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_R g2018 ( 
.A(n_1602),
.B(n_1410),
.Y(n_2018)
);

BUFx3_ASAP7_75t_L g2019 ( 
.A(n_1777),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1851),
.B(n_1855),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_L g2021 ( 
.A(n_1763),
.B(n_1780),
.Y(n_2021)
);

AOI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_1546),
.A2(n_1732),
.B1(n_1853),
.B2(n_1769),
.Y(n_2022)
);

OAI22xp5_ASAP7_75t_SL g2023 ( 
.A1(n_1649),
.A2(n_1782),
.B1(n_1823),
.B2(n_1809),
.Y(n_2023)
);

OAI22xp5_ASAP7_75t_SL g2024 ( 
.A1(n_1859),
.A2(n_1869),
.B1(n_1353),
.B2(n_1706),
.Y(n_2024)
);

OAI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_1861),
.A2(n_1865),
.B1(n_1870),
.B2(n_1868),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1485),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1558),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1871),
.B(n_1873),
.Y(n_2028)
);

NAND3xp33_ASAP7_75t_L g2029 ( 
.A(n_1403),
.B(n_1785),
.C(n_1733),
.Y(n_2029)
);

AOI21xp5_ASAP7_75t_L g2030 ( 
.A1(n_1291),
.A2(n_1877),
.B(n_1874),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1898),
.B(n_1910),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_SL g2032 ( 
.A(n_1914),
.B(n_1919),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1565),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1922),
.B(n_1296),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1493),
.Y(n_2035)
);

AOI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_1335),
.A2(n_1393),
.B(n_1336),
.Y(n_2036)
);

AND2x2_ASAP7_75t_SL g2037 ( 
.A(n_1415),
.B(n_1477),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1262),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1575),
.B(n_1616),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1655),
.B(n_1701),
.Y(n_2040)
);

O2A1O1Ixp33_ASAP7_75t_L g2041 ( 
.A1(n_1257),
.A2(n_1568),
.B(n_1571),
.C(n_1551),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1566),
.Y(n_2042)
);

AO221x1_ASAP7_75t_L g2043 ( 
.A1(n_1302),
.A2(n_1562),
.B1(n_1692),
.B2(n_1624),
.C(n_1324),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1567),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1725),
.B(n_1736),
.Y(n_2045)
);

INVx3_ASAP7_75t_L g2046 ( 
.A(n_1569),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1740),
.B(n_1758),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1577),
.Y(n_2048)
);

INVx2_ASAP7_75t_SL g2049 ( 
.A(n_1453),
.Y(n_2049)
);

AOI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_1597),
.A2(n_1790),
.B1(n_1903),
.B2(n_1883),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1761),
.B(n_1893),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1269),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1583),
.Y(n_2053)
);

AND2x6_ASAP7_75t_SL g2054 ( 
.A(n_1361),
.B(n_1282),
.Y(n_2054)
);

AOI22xp33_ASAP7_75t_L g2055 ( 
.A1(n_1330),
.A2(n_1345),
.B1(n_1591),
.B2(n_1587),
.Y(n_2055)
);

INVx1_ASAP7_75t_SL g2056 ( 
.A(n_1321),
.Y(n_2056)
);

INVx2_ASAP7_75t_SL g2057 ( 
.A(n_1366),
.Y(n_2057)
);

INVx4_ASAP7_75t_L g2058 ( 
.A(n_1439),
.Y(n_2058)
);

NAND3xp33_ASAP7_75t_L g2059 ( 
.A(n_1380),
.B(n_1341),
.C(n_1377),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1595),
.Y(n_2060)
);

A2O1A1Ixp33_ASAP7_75t_L g2061 ( 
.A1(n_1303),
.A2(n_1315),
.B(n_1426),
.C(n_1515),
.Y(n_2061)
);

AND2x4_ASAP7_75t_L g2062 ( 
.A(n_1310),
.B(n_1312),
.Y(n_2062)
);

AOI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_1554),
.A2(n_1787),
.B1(n_1298),
.B2(n_1327),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_1477),
.A2(n_1532),
.B(n_1325),
.Y(n_2064)
);

AOI22xp33_ASAP7_75t_L g2065 ( 
.A1(n_1598),
.A2(n_1604),
.B1(n_1606),
.B2(n_1603),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1289),
.B(n_1430),
.Y(n_2066)
);

INVx4_ASAP7_75t_L g2067 ( 
.A(n_1439),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1297),
.B(n_1442),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1449),
.B(n_1450),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1610),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1463),
.B(n_1467),
.Y(n_2071)
);

NAND3xp33_ASAP7_75t_L g2072 ( 
.A(n_1573),
.B(n_1585),
.C(n_1582),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1474),
.B(n_1318),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1270),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1687),
.B(n_1547),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1276),
.B(n_1326),
.Y(n_2076)
);

NOR2xp33_ASAP7_75t_R g2077 ( 
.A(n_1617),
.B(n_1916),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_L g2078 ( 
.A(n_1259),
.B(n_1263),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1592),
.B(n_1342),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1613),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1622),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1343),
.B(n_1333),
.Y(n_2082)
);

AND2x6_ASAP7_75t_L g2083 ( 
.A(n_1302),
.B(n_1562),
.Y(n_2083)
);

BUFx12f_ASAP7_75t_L g2084 ( 
.A(n_1293),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_1630),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1320),
.B(n_1337),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_L g2087 ( 
.A(n_1273),
.B(n_1275),
.Y(n_2087)
);

AOI22xp33_ASAP7_75t_L g2088 ( 
.A1(n_1632),
.A2(n_1639),
.B1(n_1644),
.B2(n_1636),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1654),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_1542),
.B(n_1316),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_SL g2091 ( 
.A(n_1439),
.B(n_1487),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1331),
.B(n_1437),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1346),
.B(n_1329),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1334),
.B(n_1352),
.Y(n_2094)
);

INVx1_ASAP7_75t_SL g2095 ( 
.A(n_1459),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1667),
.Y(n_2096)
);

AOI22xp33_ASAP7_75t_L g2097 ( 
.A1(n_1677),
.A2(n_1682),
.B1(n_1683),
.B2(n_1681),
.Y(n_2097)
);

AOI22xp33_ASAP7_75t_L g2098 ( 
.A1(n_1696),
.A2(n_1704),
.B1(n_1730),
.B2(n_1702),
.Y(n_2098)
);

A2O1A1Ixp33_ASAP7_75t_L g2099 ( 
.A1(n_1521),
.A2(n_1356),
.B(n_1516),
.C(n_1432),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_1339),
.B(n_1340),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1362),
.B(n_1367),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1354),
.Y(n_2102)
);

BUFx3_ASAP7_75t_L g2103 ( 
.A(n_1366),
.Y(n_2103)
);

BUFx8_ASAP7_75t_L g2104 ( 
.A(n_1419),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1384),
.B(n_1390),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_1365),
.B(n_1376),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1391),
.B(n_1392),
.Y(n_2107)
);

INVx8_ASAP7_75t_L g2108 ( 
.A(n_1375),
.Y(n_2108)
);

AOI22xp33_ASAP7_75t_L g2109 ( 
.A1(n_1751),
.A2(n_1755),
.B1(n_1765),
.B2(n_1753),
.Y(n_2109)
);

INVxp67_ASAP7_75t_L g2110 ( 
.A(n_1468),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_L g2111 ( 
.A(n_1586),
.B(n_1590),
.Y(n_2111)
);

NOR2x1_ASAP7_75t_R g2112 ( 
.A(n_1896),
.B(n_1363),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_1397),
.B(n_1398),
.Y(n_2113)
);

INVxp67_ASAP7_75t_SL g2114 ( 
.A(n_1440),
.Y(n_2114)
);

INVx2_ASAP7_75t_SL g2115 ( 
.A(n_1487),
.Y(n_2115)
);

INVx2_ASAP7_75t_SL g2116 ( 
.A(n_1487),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_1382),
.B(n_1383),
.Y(n_2117)
);

BUFx3_ASAP7_75t_L g2118 ( 
.A(n_1293),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1411),
.B(n_1414),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1418),
.B(n_1420),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1421),
.B(n_1423),
.Y(n_2121)
);

INVxp67_ASAP7_75t_L g2122 ( 
.A(n_1479),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_L g2123 ( 
.A(n_1605),
.B(n_1614),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1553),
.B(n_1564),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1579),
.B(n_1623),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1652),
.B(n_1684),
.Y(n_2126)
);

INVx4_ASAP7_75t_L g2127 ( 
.A(n_1488),
.Y(n_2127)
);

AND2x4_ASAP7_75t_L g2128 ( 
.A(n_1624),
.B(n_1692),
.Y(n_2128)
);

AOI21xp5_ASAP7_75t_L g2129 ( 
.A1(n_1786),
.A2(n_1279),
.B(n_1277),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_SL g2130 ( 
.A(n_1488),
.B(n_1292),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1726),
.B(n_1771),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_SL g2132 ( 
.A(n_1488),
.B(n_1436),
.Y(n_2132)
);

NAND2x1p5_ASAP7_75t_L g2133 ( 
.A(n_1350),
.B(n_1374),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_1386),
.B(n_1395),
.Y(n_2134)
);

INVx3_ASAP7_75t_L g2135 ( 
.A(n_1314),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1813),
.B(n_1895),
.Y(n_2136)
);

NOR2xp33_ASAP7_75t_L g2137 ( 
.A(n_1621),
.B(n_1625),
.Y(n_2137)
);

AOI22xp33_ASAP7_75t_L g2138 ( 
.A1(n_1774),
.A2(n_1797),
.B1(n_1799),
.B2(n_1776),
.Y(n_2138)
);

NOR2xp33_ASAP7_75t_SL g2139 ( 
.A(n_1348),
.B(n_1363),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_SL g2140 ( 
.A(n_1627),
.B(n_1642),
.Y(n_2140)
);

OR2x6_ASAP7_75t_L g2141 ( 
.A(n_1509),
.B(n_1492),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1388),
.B(n_1401),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1407),
.B(n_1409),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_1412),
.B(n_1557),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1559),
.B(n_1572),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1800),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_SL g2147 ( 
.A(n_1653),
.B(n_1659),
.Y(n_2147)
);

INVx2_ASAP7_75t_SL g2148 ( 
.A(n_1265),
.Y(n_2148)
);

AND2x6_ASAP7_75t_SL g2149 ( 
.A(n_1282),
.B(n_1300),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_L g2150 ( 
.A(n_1669),
.B(n_1690),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_SL g2151 ( 
.A(n_1699),
.B(n_1707),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1811),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1580),
.B(n_1594),
.Y(n_2153)
);

NOR2xp33_ASAP7_75t_L g2154 ( 
.A(n_1728),
.B(n_1737),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_SL g2155 ( 
.A(n_1743),
.B(n_1749),
.Y(n_2155)
);

AND2x4_ASAP7_75t_L g2156 ( 
.A(n_1350),
.B(n_1374),
.Y(n_2156)
);

O2A1O1Ixp33_ASAP7_75t_L g2157 ( 
.A1(n_1784),
.A2(n_1802),
.B(n_1830),
.C(n_1788),
.Y(n_2157)
);

INVx2_ASAP7_75t_SL g2158 ( 
.A(n_1265),
.Y(n_2158)
);

CKINVDCx20_ASAP7_75t_R g2159 ( 
.A(n_1381),
.Y(n_2159)
);

NAND3xp33_ASAP7_75t_SL g2160 ( 
.A(n_1831),
.B(n_1834),
.C(n_1833),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1596),
.B(n_1611),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_SL g2162 ( 
.A(n_1835),
.B(n_1843),
.Y(n_2162)
);

INVx2_ASAP7_75t_SL g2163 ( 
.A(n_1265),
.Y(n_2163)
);

INVxp67_ASAP7_75t_SL g2164 ( 
.A(n_1502),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1814),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1645),
.B(n_1648),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1657),
.Y(n_2167)
);

NOR2xp33_ASAP7_75t_L g2168 ( 
.A(n_1847),
.B(n_1857),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1660),
.B(n_1662),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1663),
.B(n_1670),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1672),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_SL g2172 ( 
.A(n_1866),
.B(n_1876),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_1878),
.B(n_1880),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1673),
.Y(n_2174)
);

NOR2xp33_ASAP7_75t_L g2175 ( 
.A(n_1884),
.B(n_1886),
.Y(n_2175)
);

NAND2xp33_ASAP7_75t_L g2176 ( 
.A(n_1396),
.B(n_1314),
.Y(n_2176)
);

AND2x4_ASAP7_75t_L g2177 ( 
.A(n_1373),
.B(n_1498),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_1894),
.B(n_1906),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_L g2179 ( 
.A(n_1918),
.B(n_1920),
.Y(n_2179)
);

AOI22xp33_ASAP7_75t_L g2180 ( 
.A1(n_1815),
.A2(n_1818),
.B1(n_1821),
.B2(n_1816),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_L g2181 ( 
.A(n_1368),
.B(n_1372),
.Y(n_2181)
);

AND2x6_ASAP7_75t_SL g2182 ( 
.A(n_1300),
.B(n_1686),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1678),
.B(n_1685),
.Y(n_2183)
);

OAI22xp33_ASAP7_75t_L g2184 ( 
.A1(n_1417),
.A2(n_1531),
.B1(n_1805),
.B2(n_1686),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1693),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_1694),
.B(n_1700),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1705),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1824),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1714),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_1718),
.B(n_1719),
.Y(n_2190)
);

NOR2xp33_ASAP7_75t_L g2191 ( 
.A(n_1364),
.B(n_1378),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1720),
.B(n_1722),
.Y(n_2192)
);

NAND3xp33_ASAP7_75t_SL g2193 ( 
.A(n_1511),
.B(n_1349),
.C(n_1287),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_1723),
.B(n_1735),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_1492),
.B(n_1317),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1828),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_SL g2197 ( 
.A(n_1317),
.B(n_1404),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1832),
.Y(n_2198)
);

AOI22xp5_ASAP7_75t_L g2199 ( 
.A1(n_1589),
.A2(n_1506),
.B1(n_1523),
.B2(n_1406),
.Y(n_2199)
);

NAND3xp33_ASAP7_75t_L g2200 ( 
.A(n_1394),
.B(n_1490),
.C(n_1486),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_1754),
.B(n_1759),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1838),
.Y(n_2202)
);

CKINVDCx5p33_ASAP7_75t_R g2203 ( 
.A(n_1381),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1760),
.B(n_1770),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1773),
.B(n_1775),
.Y(n_2205)
);

INVx2_ASAP7_75t_SL g2206 ( 
.A(n_1317),
.Y(n_2206)
);

AOI22xp5_ASAP7_75t_L g2207 ( 
.A1(n_1514),
.A2(n_1294),
.B1(n_1805),
.B2(n_1929),
.Y(n_2207)
);

AOI22xp33_ASAP7_75t_L g2208 ( 
.A1(n_1841),
.A2(n_1860),
.B1(n_1928),
.B2(n_1863),
.Y(n_2208)
);

O2A1O1Ixp5_ASAP7_75t_L g2209 ( 
.A1(n_1534),
.A2(n_1431),
.B(n_1424),
.C(n_1408),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1779),
.B(n_1789),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1794),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_1429),
.B(n_1455),
.Y(n_2212)
);

NAND2xp33_ASAP7_75t_L g2213 ( 
.A(n_1396),
.B(n_1314),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1801),
.B(n_1804),
.Y(n_2214)
);

NOR2xp33_ASAP7_75t_L g2215 ( 
.A(n_1404),
.B(n_1425),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1882),
.Y(n_2216)
);

AOI22xp33_ASAP7_75t_L g2217 ( 
.A1(n_1888),
.A2(n_1909),
.B1(n_1902),
.B2(n_1904),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_1806),
.B(n_1819),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1820),
.Y(n_2219)
);

NOR2xp33_ASAP7_75t_L g2220 ( 
.A(n_1404),
.B(n_1425),
.Y(n_2220)
);

NOR2xp33_ASAP7_75t_L g2221 ( 
.A(n_1425),
.B(n_1599),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_SL g2222 ( 
.A(n_1599),
.B(n_1620),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_1827),
.B(n_1836),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1912),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1837),
.B(n_1848),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_1849),
.B(n_1854),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1856),
.B(n_1858),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_1864),
.B(n_1885),
.Y(n_2228)
);

INVx3_ASAP7_75t_L g2229 ( 
.A(n_1314),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1890),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1891),
.Y(n_2231)
);

AOI22xp5_ASAP7_75t_L g2232 ( 
.A1(n_1929),
.A2(n_1286),
.B1(n_1466),
.B2(n_1338),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_SL g2233 ( 
.A(n_1599),
.B(n_1620),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1892),
.B(n_1908),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1913),
.Y(n_2235)
);

HB1xp67_ASAP7_75t_L g2236 ( 
.A(n_1465),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_SL g2237 ( 
.A(n_1620),
.B(n_1666),
.Y(n_2237)
);

INVx4_ASAP7_75t_L g2238 ( 
.A(n_1314),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_1444),
.B(n_1457),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_1271),
.B(n_1278),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_1458),
.B(n_1462),
.Y(n_2241)
);

AOI22xp5_ASAP7_75t_L g2242 ( 
.A1(n_1323),
.A2(n_1328),
.B1(n_1495),
.B2(n_1494),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1544),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1470),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_SL g2245 ( 
.A(n_1666),
.B(n_1675),
.Y(n_2245)
);

HB1xp67_ASAP7_75t_L g2246 ( 
.A(n_1332),
.Y(n_2246)
);

OAI22xp5_ASAP7_75t_L g2247 ( 
.A1(n_1601),
.A2(n_1757),
.B1(n_1615),
.B2(n_1746),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1472),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1475),
.Y(n_2249)
);

AOI22xp33_ASAP7_75t_L g2250 ( 
.A1(n_1924),
.A2(n_1927),
.B1(n_1925),
.B2(n_1489),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_1484),
.B(n_1491),
.Y(n_2251)
);

INVx8_ASAP7_75t_L g2252 ( 
.A(n_1419),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_1501),
.B(n_1295),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_1301),
.B(n_1322),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1471),
.B(n_1473),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_SL g2256 ( 
.A(n_1666),
.B(n_1675),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_1359),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_SL g2258 ( 
.A(n_1675),
.B(n_1738),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_SL g2259 ( 
.A(n_1738),
.B(n_1803),
.Y(n_2259)
);

NAND2xp33_ASAP7_75t_L g2260 ( 
.A(n_1396),
.B(n_1646),
.Y(n_2260)
);

AOI22xp5_ASAP7_75t_L g2261 ( 
.A1(n_1379),
.A2(n_1332),
.B1(n_1347),
.B2(n_1357),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_1738),
.B(n_1803),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1370),
.Y(n_2263)
);

AOI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_1358),
.A2(n_1387),
.B1(n_1360),
.B2(n_1389),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_1803),
.B(n_1845),
.Y(n_2265)
);

NOR2xp33_ASAP7_75t_L g2266 ( 
.A(n_1845),
.B(n_1499),
.Y(n_2266)
);

BUFx2_ASAP7_75t_L g2267 ( 
.A(n_1422),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_1845),
.B(n_1530),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_1399),
.B(n_1400),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_1405),
.B(n_1427),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_1513),
.B(n_1504),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_1513),
.B(n_1505),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_SL g2273 ( 
.A(n_1422),
.B(n_1867),
.Y(n_2273)
);

AND2x6_ASAP7_75t_SL g2274 ( 
.A(n_1371),
.B(n_1881),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_1513),
.B(n_1538),
.Y(n_2275)
);

HB1xp67_ASAP7_75t_L g2276 ( 
.A(n_1476),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1539),
.B(n_1461),
.Y(n_2277)
);

BUFx6f_ASAP7_75t_L g2278 ( 
.A(n_1498),
.Y(n_2278)
);

INVxp67_ASAP7_75t_L g2279 ( 
.A(n_1438),
.Y(n_2279)
);

NAND3xp33_ASAP7_75t_SL g2280 ( 
.A(n_1524),
.B(n_1896),
.C(n_1441),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1508),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_1428),
.B(n_1460),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_1433),
.B(n_1525),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_1443),
.B(n_1446),
.Y(n_2284)
);

INVx4_ASAP7_75t_L g2285 ( 
.A(n_1646),
.Y(n_2285)
);

NOR2xp33_ASAP7_75t_L g2286 ( 
.A(n_1456),
.B(n_1441),
.Y(n_2286)
);

INVx5_ASAP7_75t_L g2287 ( 
.A(n_1498),
.Y(n_2287)
);

AOI22xp33_ASAP7_75t_L g2288 ( 
.A1(n_1445),
.A2(n_1526),
.B1(n_1507),
.B2(n_1483),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_1447),
.B(n_1469),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_1452),
.B(n_1478),
.Y(n_2290)
);

AND2x6_ASAP7_75t_SL g2291 ( 
.A(n_1679),
.B(n_1881),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_1480),
.B(n_1520),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1510),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_1512),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1496),
.B(n_1528),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_1503),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_1533),
.B(n_1448),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_1500),
.B(n_1529),
.Y(n_2298)
);

AOI22xp33_ASAP7_75t_L g2299 ( 
.A1(n_1537),
.A2(n_1536),
.B1(n_1535),
.B2(n_1517),
.Y(n_2299)
);

AOI22xp33_ASAP7_75t_L g2300 ( 
.A1(n_1522),
.A2(n_1540),
.B1(n_1422),
.B2(n_1646),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_SL g2301 ( 
.A(n_1422),
.B(n_1767),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_1500),
.B(n_1464),
.Y(n_2302)
);

INVx2_ASAP7_75t_SL g2303 ( 
.A(n_1500),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_1454),
.B(n_1482),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_SL g2305 ( 
.A(n_1422),
.B(n_1646),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_1434),
.B(n_1355),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_SL g2307 ( 
.A(n_1646),
.B(n_1926),
.Y(n_2307)
);

AO22x1_ASAP7_75t_L g2308 ( 
.A1(n_1369),
.A2(n_1413),
.B1(n_1385),
.B2(n_1926),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_SL g2309 ( 
.A(n_1810),
.B(n_1926),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_1810),
.B(n_1926),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_1810),
.B(n_1926),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_SL g2312 ( 
.A(n_1810),
.B(n_1396),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_1396),
.Y(n_2313)
);

INVxp67_ASAP7_75t_L g2314 ( 
.A(n_1679),
.Y(n_2314)
);

NAND2x1_ASAP7_75t_L g2315 ( 
.A(n_1810),
.B(n_1762),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_1762),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_1846),
.B(n_1313),
.Y(n_2317)
);

BUFx3_ASAP7_75t_L g2318 ( 
.A(n_1846),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1543),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_1543),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_SL g2321 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2322)
);

NOR2xp33_ASAP7_75t_L g2323 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2323)
);

INVx2_ASAP7_75t_SL g2324 ( 
.A(n_1453),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2325)
);

BUFx3_ASAP7_75t_L g2326 ( 
.A(n_1777),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_1311),
.B(n_1253),
.Y(n_2327)
);

AND2x4_ASAP7_75t_SL g2328 ( 
.A(n_1896),
.B(n_1072),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1543),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2330)
);

BUFx3_ASAP7_75t_L g2331 ( 
.A(n_1777),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_1543),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2333)
);

OAI22xp33_ASAP7_75t_SL g2334 ( 
.A1(n_1252),
.A2(n_1875),
.B1(n_620),
.B2(n_1309),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_1543),
.Y(n_2335)
);

BUFx4f_ASAP7_75t_L g2336 ( 
.A(n_1439),
.Y(n_2336)
);

BUFx6f_ASAP7_75t_L g2337 ( 
.A(n_1439),
.Y(n_2337)
);

AOI22xp5_ASAP7_75t_L g2338 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2338)
);

BUFx6f_ASAP7_75t_L g2339 ( 
.A(n_1439),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2340)
);

INVxp33_ASAP7_75t_L g2341 ( 
.A(n_1313),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_SL g2342 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2342)
);

AOI21xp5_ASAP7_75t_L g2343 ( 
.A1(n_1744),
.A2(n_1283),
.B(n_1264),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_1543),
.Y(n_2344)
);

OAI22xp5_ASAP7_75t_L g2345 ( 
.A1(n_1250),
.A2(n_1274),
.B1(n_1280),
.B2(n_1261),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2346)
);

BUFx3_ASAP7_75t_L g2347 ( 
.A(n_1777),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2348)
);

NAND2x1_ASAP7_75t_L g2349 ( 
.A(n_1744),
.B(n_1283),
.Y(n_2349)
);

OAI21xp5_ASAP7_75t_L g2350 ( 
.A1(n_1744),
.A2(n_1261),
.B(n_1250),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2351)
);

NAND2xp33_ASAP7_75t_L g2352 ( 
.A(n_1744),
.B(n_1550),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_1543),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2354)
);

OR2x2_ASAP7_75t_L g2355 ( 
.A(n_1309),
.B(n_1304),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_SL g2356 ( 
.A(n_1348),
.B(n_542),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2357)
);

AND2x4_ASAP7_75t_SL g2358 ( 
.A(n_1896),
.B(n_1072),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_1543),
.Y(n_2359)
);

OAI21xp5_ASAP7_75t_L g2360 ( 
.A1(n_1744),
.A2(n_1261),
.B(n_1250),
.Y(n_2360)
);

INVxp67_ASAP7_75t_L g2361 ( 
.A(n_1318),
.Y(n_2361)
);

BUFx3_ASAP7_75t_L g2362 ( 
.A(n_1777),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_1543),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2364)
);

O2A1O1Ixp33_ASAP7_75t_L g2365 ( 
.A1(n_1250),
.A2(n_1274),
.B(n_1280),
.C(n_1261),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_1543),
.Y(n_2366)
);

INVx4_ASAP7_75t_L g2367 ( 
.A(n_1439),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_SL g2369 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2369)
);

CKINVDCx5p33_ASAP7_75t_R g2370 ( 
.A(n_1747),
.Y(n_2370)
);

NOR3x1_ASAP7_75t_L g2371 ( 
.A(n_1255),
.B(n_1734),
.C(n_1588),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2374)
);

BUFx8_ASAP7_75t_L g2375 ( 
.A(n_1419),
.Y(n_2375)
);

AOI22xp33_ASAP7_75t_L g2376 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_SL g2377 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2378)
);

AND2x6_ASAP7_75t_SL g2379 ( 
.A(n_1545),
.B(n_1549),
.Y(n_2379)
);

NOR2xp33_ASAP7_75t_L g2380 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2380)
);

NOR2xp33_ASAP7_75t_L g2381 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_1543),
.Y(n_2383)
);

AOI22xp33_ASAP7_75t_L g2384 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2384)
);

OAI22xp5_ASAP7_75t_SL g2385 ( 
.A1(n_1250),
.A2(n_1274),
.B1(n_1280),
.B2(n_1261),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1543),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_SL g2387 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2387)
);

INVxp67_ASAP7_75t_L g2388 ( 
.A(n_1318),
.Y(n_2388)
);

AOI22xp5_ASAP7_75t_L g2389 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2389)
);

CKINVDCx6p67_ASAP7_75t_R g2390 ( 
.A(n_1366),
.Y(n_2390)
);

INVxp67_ASAP7_75t_L g2391 ( 
.A(n_1318),
.Y(n_2391)
);

O2A1O1Ixp33_ASAP7_75t_L g2392 ( 
.A1(n_1250),
.A2(n_1274),
.B(n_1280),
.C(n_1261),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_1543),
.Y(n_2394)
);

AOI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2395)
);

NOR2xp67_ASAP7_75t_L g2396 ( 
.A(n_1283),
.B(n_1403),
.Y(n_2396)
);

AOI22xp5_ASAP7_75t_L g2397 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_1543),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_1543),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_SL g2401 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2401)
);

AOI21xp5_ASAP7_75t_L g2402 ( 
.A1(n_1744),
.A2(n_1283),
.B(n_1264),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2404)
);

AND2x4_ASAP7_75t_L g2405 ( 
.A(n_1792),
.B(n_1897),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_1543),
.Y(n_2407)
);

OAI22xp5_ASAP7_75t_L g2408 ( 
.A1(n_1250),
.A2(n_1274),
.B1(n_1280),
.B2(n_1261),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_1543),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_1543),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_1543),
.Y(n_2414)
);

NOR2xp33_ASAP7_75t_SL g2415 ( 
.A(n_1348),
.B(n_542),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2416)
);

INVx3_ASAP7_75t_L g2417 ( 
.A(n_1260),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_SL g2419 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2421)
);

BUFx6f_ASAP7_75t_L g2422 ( 
.A(n_1439),
.Y(n_2422)
);

AOI21xp5_ASAP7_75t_L g2423 ( 
.A1(n_1744),
.A2(n_1283),
.B(n_1264),
.Y(n_2423)
);

AOI21xp5_ASAP7_75t_L g2424 ( 
.A1(n_1744),
.A2(n_1283),
.B(n_1264),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2425)
);

AOI22xp33_ASAP7_75t_L g2426 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2426)
);

AOI22xp5_ASAP7_75t_L g2427 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2427)
);

INVx2_ASAP7_75t_SL g2428 ( 
.A(n_1453),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_1543),
.Y(n_2429)
);

OAI22xp33_ASAP7_75t_L g2430 ( 
.A1(n_1252),
.A2(n_1588),
.B1(n_1842),
.B2(n_1734),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2431)
);

AOI22xp5_ASAP7_75t_L g2432 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2432)
);

AOI22xp5_ASAP7_75t_L g2433 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_1543),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_1543),
.Y(n_2436)
);

NOR2xp33_ASAP7_75t_L g2437 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_SL g2438 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2439)
);

HB1xp67_ASAP7_75t_L g2440 ( 
.A(n_1581),
.Y(n_2440)
);

NAND2xp33_ASAP7_75t_L g2441 ( 
.A(n_1744),
.B(n_1550),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2442)
);

INVx8_ASAP7_75t_L g2443 ( 
.A(n_1366),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_1543),
.Y(n_2444)
);

NOR2xp33_ASAP7_75t_L g2445 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2445)
);

INVxp67_ASAP7_75t_L g2446 ( 
.A(n_1318),
.Y(n_2446)
);

AOI22xp33_ASAP7_75t_SL g2447 ( 
.A1(n_1588),
.A2(n_1201),
.B1(n_1089),
.B2(n_1734),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_1543),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2449)
);

INVxp67_ASAP7_75t_L g2450 ( 
.A(n_1318),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_SL g2451 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2451)
);

O2A1O1Ixp33_ASAP7_75t_L g2452 ( 
.A1(n_1250),
.A2(n_1274),
.B(n_1280),
.C(n_1261),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2453)
);

NOR2xp33_ASAP7_75t_L g2454 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_1543),
.Y(n_2457)
);

NOR2xp33_ASAP7_75t_L g2458 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2459)
);

AOI22xp33_ASAP7_75t_L g2460 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2460)
);

INVx8_ASAP7_75t_L g2461 ( 
.A(n_1366),
.Y(n_2461)
);

BUFx6f_ASAP7_75t_L g2462 ( 
.A(n_1439),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_SL g2463 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2463)
);

NAND2xp33_ASAP7_75t_SL g2464 ( 
.A(n_1744),
.B(n_1875),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_1543),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_SL g2466 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_1543),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2469)
);

INVx3_ASAP7_75t_L g2470 ( 
.A(n_1260),
.Y(n_2470)
);

AOI22xp5_ASAP7_75t_SL g2471 ( 
.A1(n_1609),
.A2(n_588),
.B1(n_1713),
.B2(n_1261),
.Y(n_2471)
);

INVx2_ASAP7_75t_SL g2472 ( 
.A(n_1453),
.Y(n_2472)
);

NOR2xp33_ASAP7_75t_L g2473 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_1543),
.Y(n_2474)
);

NOR2xp33_ASAP7_75t_L g2475 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2475)
);

INVx8_ASAP7_75t_L g2476 ( 
.A(n_1366),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_1543),
.Y(n_2477)
);

NOR2xp33_ASAP7_75t_L g2478 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_1543),
.Y(n_2480)
);

AOI22xp5_ASAP7_75t_L g2481 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2481)
);

AOI22xp33_ASAP7_75t_L g2482 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2482)
);

HB1xp67_ASAP7_75t_L g2483 ( 
.A(n_1581),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2484)
);

NOR2xp33_ASAP7_75t_L g2485 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2486)
);

OAI22xp5_ASAP7_75t_SL g2487 ( 
.A1(n_1250),
.A2(n_1274),
.B1(n_1280),
.B2(n_1261),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_1543),
.Y(n_2488)
);

INVx2_ASAP7_75t_SL g2489 ( 
.A(n_1453),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2490)
);

AOI22xp33_ASAP7_75t_L g2491 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_1543),
.Y(n_2492)
);

NOR2xp33_ASAP7_75t_SL g2493 ( 
.A(n_1348),
.B(n_542),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_1543),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_1543),
.Y(n_2497)
);

AOI22xp5_ASAP7_75t_L g2498 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2498)
);

OAI21xp5_ASAP7_75t_L g2499 ( 
.A1(n_1744),
.A2(n_1261),
.B(n_1250),
.Y(n_2499)
);

NAND3xp33_ASAP7_75t_L g2500 ( 
.A(n_1250),
.B(n_1274),
.C(n_1261),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_SL g2502 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_SL g2506 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_SL g2509 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2510)
);

INVx8_ASAP7_75t_L g2511 ( 
.A(n_1366),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_1543),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_SL g2513 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_SL g2514 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2514)
);

AOI22xp33_ASAP7_75t_SL g2515 ( 
.A1(n_1588),
.A2(n_1201),
.B1(n_1089),
.B2(n_1734),
.Y(n_2515)
);

OAI22xp33_ASAP7_75t_L g2516 ( 
.A1(n_1252),
.A2(n_1588),
.B1(n_1842),
.B2(n_1734),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_SL g2518 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_1311),
.B(n_1253),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2520)
);

INVx1_ASAP7_75t_SL g2521 ( 
.A(n_1747),
.Y(n_2521)
);

INVx2_ASAP7_75t_SL g2522 ( 
.A(n_1453),
.Y(n_2522)
);

OAI21xp5_ASAP7_75t_L g2523 ( 
.A1(n_1744),
.A2(n_1261),
.B(n_1250),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_SL g2524 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_SL g2525 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2526)
);

NOR2xp33_ASAP7_75t_L g2527 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_1543),
.Y(n_2528)
);

NOR3xp33_ASAP7_75t_L g2529 ( 
.A(n_1250),
.B(n_1274),
.C(n_1261),
.Y(n_2529)
);

NOR2xp33_ASAP7_75t_L g2530 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_1543),
.Y(n_2531)
);

AOI22xp5_ASAP7_75t_L g2532 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_SL g2533 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2533)
);

OAI21xp5_ASAP7_75t_L g2534 ( 
.A1(n_1744),
.A2(n_1261),
.B(n_1250),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_1543),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2536)
);

AOI22xp5_ASAP7_75t_L g2537 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_1543),
.Y(n_2538)
);

AND2x4_ASAP7_75t_L g2539 ( 
.A(n_1792),
.B(n_1897),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_1543),
.Y(n_2540)
);

AOI22xp5_ASAP7_75t_L g2541 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_1543),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_1543),
.Y(n_2544)
);

NOR2xp33_ASAP7_75t_L g2545 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_1543),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_1543),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_SL g2548 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2549)
);

NAND2x1p5_ASAP7_75t_L g2550 ( 
.A(n_1260),
.B(n_1569),
.Y(n_2550)
);

AOI21xp5_ASAP7_75t_L g2551 ( 
.A1(n_1744),
.A2(n_1283),
.B(n_1264),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_1543),
.Y(n_2553)
);

AOI22xp5_ASAP7_75t_L g2554 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2554)
);

INVx3_ASAP7_75t_L g2555 ( 
.A(n_1260),
.Y(n_2555)
);

A2O1A1Ixp33_ASAP7_75t_L g2556 ( 
.A1(n_1744),
.A2(n_1875),
.B(n_1311),
.C(n_1734),
.Y(n_2556)
);

AOI22xp33_ASAP7_75t_L g2557 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2557)
);

AOI22xp33_ASAP7_75t_L g2558 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2558)
);

INVx4_ASAP7_75t_L g2559 ( 
.A(n_1439),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2560)
);

INVx2_ASAP7_75t_SL g2561 ( 
.A(n_1453),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_1543),
.Y(n_2563)
);

AOI22xp33_ASAP7_75t_L g2564 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2564)
);

INVxp67_ASAP7_75t_SL g2565 ( 
.A(n_1324),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_SL g2566 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2566)
);

NOR2xp33_ASAP7_75t_L g2567 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_SL g2569 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2569)
);

AOI22xp5_ASAP7_75t_L g2570 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_1543),
.Y(n_2571)
);

AND2x2_ASAP7_75t_SL g2572 ( 
.A(n_1336),
.B(n_1201),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_1543),
.Y(n_2573)
);

NOR2xp67_ASAP7_75t_L g2574 ( 
.A(n_1283),
.B(n_1403),
.Y(n_2574)
);

NOR2x2_ASAP7_75t_L g2575 ( 
.A(n_1282),
.B(n_1300),
.Y(n_2575)
);

INVx3_ASAP7_75t_L g2576 ( 
.A(n_1260),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2578)
);

NOR2xp67_ASAP7_75t_L g2579 ( 
.A(n_1283),
.B(n_1403),
.Y(n_2579)
);

INVx8_ASAP7_75t_L g2580 ( 
.A(n_1366),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_1543),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_1543),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2585)
);

BUFx4f_ASAP7_75t_L g2586 ( 
.A(n_1439),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_1543),
.Y(n_2588)
);

NOR2xp33_ASAP7_75t_SL g2589 ( 
.A(n_1348),
.B(n_542),
.Y(n_2589)
);

AOI21xp5_ASAP7_75t_L g2590 ( 
.A1(n_1744),
.A2(n_1283),
.B(n_1264),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_SL g2591 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2591)
);

INVx3_ASAP7_75t_L g2592 ( 
.A(n_1260),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2593)
);

AOI22xp33_ASAP7_75t_L g2594 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2594)
);

AOI22xp33_ASAP7_75t_L g2595 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2595)
);

AND2x6_ASAP7_75t_L g2596 ( 
.A(n_1302),
.B(n_1562),
.Y(n_2596)
);

BUFx3_ASAP7_75t_L g2597 ( 
.A(n_1777),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2598)
);

INVx2_ASAP7_75t_SL g2599 ( 
.A(n_1453),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_1543),
.Y(n_2600)
);

INVx3_ASAP7_75t_L g2601 ( 
.A(n_1260),
.Y(n_2601)
);

BUFx2_ASAP7_75t_L g2602 ( 
.A(n_1664),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_1543),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_1543),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_SL g2606 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2607)
);

INVx3_ASAP7_75t_L g2608 ( 
.A(n_1260),
.Y(n_2608)
);

OAI22xp5_ASAP7_75t_L g2609 ( 
.A1(n_1250),
.A2(n_1274),
.B1(n_1280),
.B2(n_1261),
.Y(n_2609)
);

AOI22xp5_ASAP7_75t_L g2610 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_SL g2611 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2611)
);

A2O1A1Ixp33_ASAP7_75t_SL g2612 ( 
.A1(n_1250),
.A2(n_1274),
.B(n_1280),
.C(n_1261),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_1543),
.Y(n_2614)
);

NAND2x1_ASAP7_75t_L g2615 ( 
.A(n_1744),
.B(n_1283),
.Y(n_2615)
);

AOI22xp33_ASAP7_75t_L g2616 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_SL g2617 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2617)
);

BUFx6f_ASAP7_75t_L g2618 ( 
.A(n_1439),
.Y(n_2618)
);

INVx3_ASAP7_75t_L g2619 ( 
.A(n_1260),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2620)
);

NOR2xp33_ASAP7_75t_L g2621 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_SL g2622 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_1543),
.Y(n_2626)
);

BUFx3_ASAP7_75t_L g2627 ( 
.A(n_1777),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_1543),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_SL g2629 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2630)
);

AO22x1_ASAP7_75t_L g2631 ( 
.A1(n_1609),
.A2(n_1713),
.B1(n_1311),
.B2(n_1875),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2632)
);

AND3x1_ASAP7_75t_L g2633 ( 
.A(n_1554),
.B(n_1787),
.C(n_1261),
.Y(n_2633)
);

AND2x4_ASAP7_75t_L g2634 ( 
.A(n_1792),
.B(n_1897),
.Y(n_2634)
);

NOR2xp67_ASAP7_75t_L g2635 ( 
.A(n_1283),
.B(n_1403),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_1543),
.Y(n_2636)
);

CKINVDCx16_ASAP7_75t_R g2637 ( 
.A(n_1554),
.Y(n_2637)
);

AND2x6_ASAP7_75t_SL g2638 ( 
.A(n_1545),
.B(n_1549),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_SL g2639 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_SL g2640 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2640)
);

INVx2_ASAP7_75t_SL g2641 ( 
.A(n_1453),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_SL g2642 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2642)
);

AOI22xp5_ASAP7_75t_L g2643 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2644)
);

NAND2xp33_ASAP7_75t_SL g2645 ( 
.A(n_1744),
.B(n_1875),
.Y(n_2645)
);

INVxp33_ASAP7_75t_SL g2646 ( 
.A(n_1554),
.Y(n_2646)
);

CKINVDCx5p33_ASAP7_75t_R g2647 ( 
.A(n_1747),
.Y(n_2647)
);

OAI22xp33_ASAP7_75t_L g2648 ( 
.A1(n_1252),
.A2(n_1588),
.B1(n_1842),
.B2(n_1734),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2649)
);

AOI22xp5_ASAP7_75t_L g2650 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2650)
);

AOI22xp33_ASAP7_75t_L g2651 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2651)
);

O2A1O1Ixp5_ASAP7_75t_L g2652 ( 
.A1(n_1744),
.A2(n_1261),
.B(n_1274),
.C(n_1250),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2653)
);

BUFx3_ASAP7_75t_L g2654 ( 
.A(n_1777),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_SL g2655 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2655)
);

AOI22xp5_ASAP7_75t_L g2656 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2656)
);

AOI22xp33_ASAP7_75t_L g2657 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2657)
);

INVx2_ASAP7_75t_SL g2658 ( 
.A(n_1453),
.Y(n_2658)
);

NOR2xp33_ASAP7_75t_L g2659 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2659)
);

BUFx6f_ASAP7_75t_L g2660 ( 
.A(n_1439),
.Y(n_2660)
);

OR2x2_ASAP7_75t_L g2661 ( 
.A(n_1309),
.B(n_1304),
.Y(n_2661)
);

AOI22xp33_ASAP7_75t_L g2662 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2662)
);

NOR3xp33_ASAP7_75t_L g2663 ( 
.A(n_1250),
.B(n_1274),
.C(n_1261),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_1543),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_SL g2665 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_1543),
.Y(n_2666)
);

NOR2xp33_ASAP7_75t_L g2667 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_SL g2668 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2668)
);

INVx2_ASAP7_75t_L g2669 ( 
.A(n_1543),
.Y(n_2669)
);

INVx4_ASAP7_75t_L g2670 ( 
.A(n_1439),
.Y(n_2670)
);

NOR2xp33_ASAP7_75t_L g2671 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2672)
);

NOR2xp33_ASAP7_75t_SL g2673 ( 
.A(n_1348),
.B(n_542),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_1543),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2676)
);

OR2x2_ASAP7_75t_L g2677 ( 
.A(n_1309),
.B(n_1304),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2679)
);

INVxp67_ASAP7_75t_L g2680 ( 
.A(n_1318),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_1543),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_1543),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2686)
);

NOR2xp33_ASAP7_75t_L g2687 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_SL g2688 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_1543),
.Y(n_2690)
);

NOR2xp33_ASAP7_75t_L g2691 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_1543),
.Y(n_2693)
);

AOI221xp5_ASAP7_75t_L g2694 ( 
.A1(n_1875),
.A2(n_1658),
.B1(n_1887),
.B2(n_1850),
.C(n_1612),
.Y(n_2694)
);

HB1xp67_ASAP7_75t_L g2695 ( 
.A(n_1581),
.Y(n_2695)
);

NOR2x2_ASAP7_75t_L g2696 ( 
.A(n_1282),
.B(n_1300),
.Y(n_2696)
);

NOR2xp33_ASAP7_75t_L g2697 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_1543),
.Y(n_2698)
);

NOR2xp33_ASAP7_75t_L g2699 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2699)
);

NOR2xp33_ASAP7_75t_L g2700 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_SL g2701 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2702)
);

AOI22xp33_ASAP7_75t_L g2703 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2703)
);

NOR2xp33_ASAP7_75t_SL g2704 ( 
.A(n_1348),
.B(n_542),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_SL g2705 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2707)
);

AOI22xp33_ASAP7_75t_L g2708 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2708)
);

BUFx3_ASAP7_75t_L g2709 ( 
.A(n_1777),
.Y(n_2709)
);

AOI22xp33_ASAP7_75t_L g2710 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2711)
);

AND2x4_ASAP7_75t_L g2712 ( 
.A(n_1792),
.B(n_1897),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_SL g2713 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_SL g2714 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2714)
);

AOI22xp33_ASAP7_75t_L g2715 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2716)
);

NOR2xp33_ASAP7_75t_SL g2717 ( 
.A(n_1348),
.B(n_542),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2718)
);

NOR2xp33_ASAP7_75t_L g2719 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_1543),
.Y(n_2721)
);

AOI22xp33_ASAP7_75t_L g2722 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_1311),
.B(n_1253),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2724)
);

AND2x6_ASAP7_75t_SL g2725 ( 
.A(n_1545),
.B(n_1549),
.Y(n_2725)
);

AOI22xp33_ASAP7_75t_L g2726 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_1543),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2729)
);

AOI21xp5_ASAP7_75t_L g2730 ( 
.A1(n_1744),
.A2(n_1283),
.B(n_1264),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_1543),
.Y(n_2731)
);

OAI22xp5_ASAP7_75t_SL g2732 ( 
.A1(n_1250),
.A2(n_1274),
.B1(n_1280),
.B2(n_1261),
.Y(n_2732)
);

AOI22xp5_ASAP7_75t_L g2733 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_1543),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_1543),
.Y(n_2735)
);

AOI21xp5_ASAP7_75t_L g2736 ( 
.A1(n_1744),
.A2(n_1283),
.B(n_1264),
.Y(n_2736)
);

INVx2_ASAP7_75t_SL g2737 ( 
.A(n_1453),
.Y(n_2737)
);

CKINVDCx5p33_ASAP7_75t_R g2738 ( 
.A(n_1747),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2739)
);

AND2x2_ASAP7_75t_SL g2740 ( 
.A(n_1336),
.B(n_1201),
.Y(n_2740)
);

OR2x2_ASAP7_75t_L g2741 ( 
.A(n_1309),
.B(n_1304),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_1543),
.Y(n_2742)
);

NOR2xp33_ASAP7_75t_L g2743 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2743)
);

NOR2xp33_ASAP7_75t_L g2744 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2744)
);

CKINVDCx20_ASAP7_75t_R g2745 ( 
.A(n_1747),
.Y(n_2745)
);

INVx8_ASAP7_75t_L g2746 ( 
.A(n_1366),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_1543),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_SL g2750 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_1543),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_1543),
.Y(n_2753)
);

AND2x2_ASAP7_75t_L g2754 ( 
.A(n_1311),
.B(n_1253),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_SL g2755 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2755)
);

AND2x4_ASAP7_75t_L g2756 ( 
.A(n_1792),
.B(n_1897),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_L g2757 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2757)
);

NOR2xp67_ASAP7_75t_L g2758 ( 
.A(n_1283),
.B(n_1403),
.Y(n_2758)
);

AOI22xp33_ASAP7_75t_L g2759 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2759)
);

INVx2_ASAP7_75t_SL g2760 ( 
.A(n_1453),
.Y(n_2760)
);

NAND2xp33_ASAP7_75t_SL g2761 ( 
.A(n_1744),
.B(n_1875),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_1543),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_1543),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_1543),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_SL g2766 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2766)
);

NOR2xp33_ASAP7_75t_SL g2767 ( 
.A(n_1348),
.B(n_542),
.Y(n_2767)
);

OR2x6_ASAP7_75t_L g2768 ( 
.A(n_1260),
.B(n_1569),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2769)
);

AOI22xp33_ASAP7_75t_L g2770 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2770)
);

AOI22xp5_ASAP7_75t_L g2771 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_SL g2772 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2772)
);

INVx8_ASAP7_75t_L g2773 ( 
.A(n_1366),
.Y(n_2773)
);

AOI21xp5_ASAP7_75t_L g2774 ( 
.A1(n_1744),
.A2(n_1283),
.B(n_1264),
.Y(n_2774)
);

AND2x2_ASAP7_75t_L g2775 ( 
.A(n_1311),
.B(n_1253),
.Y(n_2775)
);

AOI22xp5_ASAP7_75t_L g2776 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2776)
);

BUFx6f_ASAP7_75t_L g2777 ( 
.A(n_1439),
.Y(n_2777)
);

NOR2xp33_ASAP7_75t_L g2778 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2778)
);

NOR2xp67_ASAP7_75t_L g2779 ( 
.A(n_1283),
.B(n_1403),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_1543),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_1543),
.Y(n_2781)
);

A2O1A1Ixp33_ASAP7_75t_L g2782 ( 
.A1(n_1744),
.A2(n_1875),
.B(n_1311),
.C(n_1734),
.Y(n_2782)
);

CKINVDCx5p33_ASAP7_75t_R g2783 ( 
.A(n_1747),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_1543),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2785)
);

NOR2xp33_ASAP7_75t_L g2786 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_SL g2787 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2788)
);

HB1xp67_ASAP7_75t_L g2789 ( 
.A(n_1581),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_1543),
.Y(n_2790)
);

NOR2xp33_ASAP7_75t_SL g2791 ( 
.A(n_1348),
.B(n_542),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2792)
);

O2A1O1Ixp33_ASAP7_75t_L g2793 ( 
.A1(n_1250),
.A2(n_1274),
.B(n_1280),
.C(n_1261),
.Y(n_2793)
);

NOR2xp33_ASAP7_75t_L g2794 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_SL g2795 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_1543),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_1543),
.Y(n_2797)
);

INVx3_ASAP7_75t_L g2798 ( 
.A(n_1260),
.Y(n_2798)
);

INVxp67_ASAP7_75t_L g2799 ( 
.A(n_1318),
.Y(n_2799)
);

CKINVDCx5p33_ASAP7_75t_R g2800 ( 
.A(n_1747),
.Y(n_2800)
);

AND2x2_ASAP7_75t_L g2801 ( 
.A(n_1311),
.B(n_1253),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_1543),
.Y(n_2802)
);

INVxp67_ASAP7_75t_SL g2803 ( 
.A(n_1324),
.Y(n_2803)
);

AOI22xp5_ASAP7_75t_L g2804 ( 
.A1(n_1588),
.A2(n_1734),
.B1(n_1900),
.B2(n_1842),
.Y(n_2804)
);

NOR2xp33_ASAP7_75t_SL g2805 ( 
.A(n_1348),
.B(n_542),
.Y(n_2805)
);

OAI22xp5_ASAP7_75t_SL g2806 ( 
.A1(n_1250),
.A2(n_1274),
.B1(n_1280),
.B2(n_1261),
.Y(n_2806)
);

AOI22xp33_ASAP7_75t_L g2807 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_1543),
.Y(n_2808)
);

AOI22xp5_ASAP7_75t_L g2809 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2810)
);

AOI22xp5_ASAP7_75t_L g2811 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2811)
);

INVx2_ASAP7_75t_SL g2812 ( 
.A(n_1453),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2813)
);

CKINVDCx11_ASAP7_75t_R g2814 ( 
.A(n_1747),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_1543),
.Y(n_2815)
);

INVx8_ASAP7_75t_L g2816 ( 
.A(n_1366),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_1543),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_SL g2819 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_1543),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_1543),
.Y(n_2821)
);

AOI22xp33_ASAP7_75t_L g2822 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2822)
);

NOR2xp33_ASAP7_75t_L g2823 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2823)
);

OAI22xp5_ASAP7_75t_SL g2824 ( 
.A1(n_1250),
.A2(n_1274),
.B1(n_1280),
.B2(n_1261),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_1543),
.Y(n_2827)
);

NOR2xp33_ASAP7_75t_L g2828 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2828)
);

OAI22xp5_ASAP7_75t_SL g2829 ( 
.A1(n_1250),
.A2(n_1274),
.B1(n_1280),
.B2(n_1261),
.Y(n_2829)
);

INVx2_ASAP7_75t_SL g2830 ( 
.A(n_1453),
.Y(n_2830)
);

NOR3xp33_ASAP7_75t_SL g2831 ( 
.A(n_1545),
.B(n_486),
.C(n_455),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_L g2832 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2833)
);

NOR2xp33_ASAP7_75t_L g2834 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2834)
);

AOI21xp5_ASAP7_75t_L g2835 ( 
.A1(n_1744),
.A2(n_1283),
.B(n_1264),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_1543),
.Y(n_2836)
);

AND2x6_ASAP7_75t_L g2837 ( 
.A(n_1302),
.B(n_1562),
.Y(n_2837)
);

INVxp33_ASAP7_75t_L g2838 ( 
.A(n_1313),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_SL g2839 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2839)
);

AND2x6_ASAP7_75t_SL g2840 ( 
.A(n_1545),
.B(n_1549),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2841)
);

AO22x1_ASAP7_75t_L g2842 ( 
.A1(n_1609),
.A2(n_1713),
.B1(n_1311),
.B2(n_1875),
.Y(n_2842)
);

HB1xp67_ASAP7_75t_L g2843 ( 
.A(n_1581),
.Y(n_2843)
);

INVx3_ASAP7_75t_L g2844 ( 
.A(n_1260),
.Y(n_2844)
);

OAI221xp5_ASAP7_75t_L g2845 ( 
.A1(n_1261),
.A2(n_1274),
.B1(n_1280),
.B2(n_1250),
.C(n_1612),
.Y(n_2845)
);

INVx2_ASAP7_75t_SL g2846 ( 
.A(n_1453),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_1543),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_SL g2849 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_SL g2852 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2852)
);

BUFx2_ASAP7_75t_L g2853 ( 
.A(n_1664),
.Y(n_2853)
);

NOR2xp33_ASAP7_75t_L g2854 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2855)
);

AOI22xp5_ASAP7_75t_L g2856 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2856)
);

AOI22xp33_ASAP7_75t_L g2857 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_1543),
.Y(n_2858)
);

INVx2_ASAP7_75t_SL g2859 ( 
.A(n_1453),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_SL g2860 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2860)
);

NOR2xp33_ASAP7_75t_L g2861 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_SL g2863 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2863)
);

NOR2xp33_ASAP7_75t_L g2864 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_1543),
.Y(n_2865)
);

INVx8_ASAP7_75t_L g2866 ( 
.A(n_1366),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_1543),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_SL g2868 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2868)
);

INVx4_ASAP7_75t_L g2869 ( 
.A(n_1439),
.Y(n_2869)
);

AND2x2_ASAP7_75t_L g2870 ( 
.A(n_1311),
.B(n_1253),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_SL g2871 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2871)
);

INVx4_ASAP7_75t_L g2872 ( 
.A(n_1439),
.Y(n_2872)
);

AND2x4_ASAP7_75t_L g2873 ( 
.A(n_1792),
.B(n_1897),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_1543),
.Y(n_2874)
);

O2A1O1Ixp33_ASAP7_75t_L g2875 ( 
.A1(n_1250),
.A2(n_1274),
.B(n_1280),
.C(n_1261),
.Y(n_2875)
);

AOI21xp5_ASAP7_75t_L g2876 ( 
.A1(n_1744),
.A2(n_1283),
.B(n_1264),
.Y(n_2876)
);

AND2x2_ASAP7_75t_L g2877 ( 
.A(n_1311),
.B(n_1253),
.Y(n_2877)
);

HB1xp67_ASAP7_75t_L g2878 ( 
.A(n_1581),
.Y(n_2878)
);

CKINVDCx11_ASAP7_75t_R g2879 ( 
.A(n_1747),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_SL g2881 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2881)
);

AOI22xp33_ASAP7_75t_L g2882 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2884)
);

NOR2x1_ASAP7_75t_R g2885 ( 
.A(n_1896),
.B(n_455),
.Y(n_2885)
);

INVx2_ASAP7_75t_SL g2886 ( 
.A(n_1453),
.Y(n_2886)
);

O2A1O1Ixp33_ASAP7_75t_L g2887 ( 
.A1(n_1250),
.A2(n_1274),
.B(n_1280),
.C(n_1261),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_1311),
.B(n_1253),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_1543),
.Y(n_2889)
);

A2O1A1Ixp33_ASAP7_75t_L g2890 ( 
.A1(n_1744),
.A2(n_1875),
.B(n_1311),
.C(n_1734),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_1543),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2895)
);

BUFx6f_ASAP7_75t_L g2896 ( 
.A(n_1439),
.Y(n_2896)
);

NOR2xp33_ASAP7_75t_L g2897 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2897)
);

OAI22xp5_ASAP7_75t_L g2898 ( 
.A1(n_1250),
.A2(n_1274),
.B1(n_1280),
.B2(n_1261),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2901)
);

HB1xp67_ASAP7_75t_L g2902 ( 
.A(n_1581),
.Y(n_2902)
);

INVx4_ASAP7_75t_L g2903 ( 
.A(n_1439),
.Y(n_2903)
);

NOR2xp33_ASAP7_75t_L g2904 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2905)
);

NOR2xp33_ASAP7_75t_L g2906 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2907)
);

BUFx3_ASAP7_75t_L g2908 ( 
.A(n_1777),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_1543),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_1543),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_1543),
.Y(n_2911)
);

OR2x2_ASAP7_75t_L g2912 ( 
.A(n_1309),
.B(n_1304),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_SL g2914 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2914)
);

OAI22xp5_ASAP7_75t_L g2915 ( 
.A1(n_1250),
.A2(n_1274),
.B1(n_1280),
.B2(n_1261),
.Y(n_2915)
);

NOR2xp33_ASAP7_75t_L g2916 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_SL g2917 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2917)
);

NOR2x1p5_ASAP7_75t_L g2918 ( 
.A(n_1588),
.B(n_1734),
.Y(n_2918)
);

NAND2x1_ASAP7_75t_L g2919 ( 
.A(n_1744),
.B(n_1283),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_SL g2920 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2920)
);

AND2x6_ASAP7_75t_SL g2921 ( 
.A(n_1545),
.B(n_1549),
.Y(n_2921)
);

BUFx3_ASAP7_75t_L g2922 ( 
.A(n_1777),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_1543),
.Y(n_2923)
);

AND2x4_ASAP7_75t_L g2924 ( 
.A(n_1792),
.B(n_1897),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_1543),
.Y(n_2925)
);

INVx8_ASAP7_75t_L g2926 ( 
.A(n_1366),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_SL g2928 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_1543),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2930)
);

AOI22xp5_ASAP7_75t_L g2931 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2931)
);

AOI22xp33_ASAP7_75t_SL g2932 ( 
.A1(n_1588),
.A2(n_1201),
.B1(n_1089),
.B2(n_1734),
.Y(n_2932)
);

BUFx6f_ASAP7_75t_L g2933 ( 
.A(n_1439),
.Y(n_2933)
);

O2A1O1Ixp5_ASAP7_75t_L g2934 ( 
.A1(n_1744),
.A2(n_1261),
.B(n_1274),
.C(n_1250),
.Y(n_2934)
);

AOI22xp5_ASAP7_75t_L g2935 ( 
.A1(n_1250),
.A2(n_1261),
.B1(n_1280),
.B2(n_1274),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_SL g2937 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_1543),
.Y(n_2938)
);

INVx2_ASAP7_75t_SL g2939 ( 
.A(n_1453),
.Y(n_2939)
);

INVx2_ASAP7_75t_L g2940 ( 
.A(n_1543),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_SL g2941 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2941)
);

INVx2_ASAP7_75t_L g2942 ( 
.A(n_1543),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_1543),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_1543),
.Y(n_2944)
);

INVx2_ASAP7_75t_SL g2945 ( 
.A(n_1453),
.Y(n_2945)
);

AND2x4_ASAP7_75t_SL g2946 ( 
.A(n_1896),
.B(n_1072),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_1543),
.Y(n_2947)
);

AND2x2_ASAP7_75t_L g2948 ( 
.A(n_1311),
.B(n_1253),
.Y(n_2948)
);

AOI21xp5_ASAP7_75t_L g2949 ( 
.A1(n_1744),
.A2(n_1283),
.B(n_1264),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_1543),
.Y(n_2950)
);

AOI22xp33_ASAP7_75t_L g2951 ( 
.A1(n_1556),
.A2(n_1899),
.B1(n_1089),
.B2(n_1201),
.Y(n_2951)
);

NOR3xp33_ASAP7_75t_L g2952 ( 
.A(n_1250),
.B(n_1274),
.C(n_1261),
.Y(n_2952)
);

AND2x2_ASAP7_75t_L g2953 ( 
.A(n_1311),
.B(n_1253),
.Y(n_2953)
);

NAND3xp33_ASAP7_75t_SL g2954 ( 
.A(n_1250),
.B(n_1274),
.C(n_1261),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_1313),
.B(n_1251),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_1543),
.Y(n_2956)
);

NOR2xp33_ASAP7_75t_L g2957 ( 
.A(n_1250),
.B(n_1261),
.Y(n_2957)
);

AND2x2_ASAP7_75t_L g2958 ( 
.A(n_1311),
.B(n_1253),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_SL g2959 ( 
.A(n_1313),
.B(n_1435),
.Y(n_2959)
);

AOI22xp33_ASAP7_75t_L g2960 ( 
.A1(n_2447),
.A2(n_2515),
.B1(n_2932),
.B2(n_1953),
.Y(n_2960)
);

INVx3_ASAP7_75t_L g2961 ( 
.A(n_2349),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_SL g2962 ( 
.A(n_2350),
.B(n_2360),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_1944),
.B(n_2327),
.Y(n_2963)
);

AOI21xp5_ASAP7_75t_L g2964 ( 
.A1(n_2499),
.A2(n_2534),
.B(n_2523),
.Y(n_2964)
);

AO21x1_ASAP7_75t_L g2965 ( 
.A1(n_2464),
.A2(n_2761),
.B(n_2645),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_1944),
.B(n_2327),
.Y(n_2966)
);

AOI21xp5_ASAP7_75t_L g2967 ( 
.A1(n_2464),
.A2(n_2761),
.B(n_2645),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2519),
.B(n_2723),
.Y(n_2968)
);

AOI21xp5_ASAP7_75t_L g2969 ( 
.A1(n_2352),
.A2(n_2441),
.B(n_2349),
.Y(n_2969)
);

A2O1A1Ixp33_ASAP7_75t_L g2970 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1948),
.C(n_2782),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2519),
.B(n_2723),
.Y(n_2971)
);

OAI21xp5_ASAP7_75t_L g2972 ( 
.A1(n_2556),
.A2(n_2890),
.B(n_2345),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_SL g2973 ( 
.A(n_2338),
.B(n_2389),
.Y(n_2973)
);

O2A1O1Ixp33_ASAP7_75t_L g2974 ( 
.A1(n_1932),
.A2(n_2609),
.B(n_2898),
.C(n_2408),
.Y(n_2974)
);

INVx4_ASAP7_75t_L g2975 ( 
.A(n_2768),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2754),
.B(n_2775),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2754),
.B(n_2775),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_SL g2978 ( 
.A(n_2395),
.B(n_2397),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_SL g2979 ( 
.A(n_2427),
.B(n_2432),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2319),
.Y(n_2980)
);

NOR2xp33_ASAP7_75t_L g2981 ( 
.A(n_2915),
.B(n_2385),
.Y(n_2981)
);

AOI21xp5_ASAP7_75t_L g2982 ( 
.A1(n_2352),
.A2(n_2441),
.B(n_2615),
.Y(n_2982)
);

OAI321xp33_ASAP7_75t_L g2983 ( 
.A1(n_2845),
.A2(n_2516),
.A3(n_2648),
.B1(n_2430),
.B2(n_2804),
.C(n_2694),
.Y(n_2983)
);

NOR2xp67_ASAP7_75t_R g2984 ( 
.A(n_2631),
.B(n_2842),
.Y(n_2984)
);

A2O1A1Ixp33_ASAP7_75t_L g2985 ( 
.A1(n_2365),
.A2(n_2452),
.B(n_2793),
.C(n_2392),
.Y(n_2985)
);

AOI21x1_ASAP7_75t_L g2986 ( 
.A1(n_1996),
.A2(n_2842),
.B(n_2631),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_SL g2987 ( 
.A(n_2433),
.B(n_2481),
.Y(n_2987)
);

AOI21xp5_ASAP7_75t_L g2988 ( 
.A1(n_2615),
.A2(n_2919),
.B(n_2402),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2801),
.B(n_2870),
.Y(n_2989)
);

NOR2xp33_ASAP7_75t_L g2990 ( 
.A(n_2487),
.B(n_2732),
.Y(n_2990)
);

OAI21xp5_ASAP7_75t_L g2991 ( 
.A1(n_2875),
.A2(n_2887),
.B(n_2532),
.Y(n_2991)
);

NOR2xp67_ASAP7_75t_L g2992 ( 
.A(n_2029),
.B(n_2129),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2801),
.B(n_2870),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2877),
.B(n_2888),
.Y(n_2994)
);

AND2x4_ASAP7_75t_L g2995 ( 
.A(n_2267),
.B(n_2768),
.Y(n_2995)
);

OR2x2_ASAP7_75t_L g2996 ( 
.A(n_2090),
.B(n_2948),
.Y(n_2996)
);

AOI21xp5_ASAP7_75t_L g2997 ( 
.A1(n_2919),
.A2(n_2423),
.B(n_2343),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2877),
.B(n_2888),
.Y(n_2998)
);

AOI21x1_ASAP7_75t_L g2999 ( 
.A1(n_1996),
.A2(n_2574),
.B(n_2396),
.Y(n_2999)
);

HB1xp67_ASAP7_75t_L g3000 ( 
.A(n_1945),
.Y(n_3000)
);

AOI21x1_ASAP7_75t_L g3001 ( 
.A1(n_2396),
.A2(n_2579),
.B(n_2574),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_SL g3002 ( 
.A(n_2498),
.B(n_2537),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2956),
.Y(n_3003)
);

OAI21xp5_ASAP7_75t_L g3004 ( 
.A1(n_2541),
.A2(n_2570),
.B(n_2554),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_SL g3005 ( 
.A(n_2610),
.B(n_2643),
.Y(n_3005)
);

AOI21xp5_ASAP7_75t_L g3006 ( 
.A1(n_2424),
.A2(n_2590),
.B(n_2551),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_SL g3007 ( 
.A(n_2650),
.B(n_2656),
.Y(n_3007)
);

AOI22xp5_ASAP7_75t_L g3008 ( 
.A1(n_2323),
.A2(n_2380),
.B1(n_2437),
.B2(n_2381),
.Y(n_3008)
);

BUFx6f_ASAP7_75t_L g3009 ( 
.A(n_2037),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2948),
.B(n_2953),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2953),
.B(n_2958),
.Y(n_3011)
);

O2A1O1Ixp33_ASAP7_75t_L g3012 ( 
.A1(n_2612),
.A2(n_2454),
.B(n_2458),
.C(n_2445),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_2958),
.B(n_2730),
.Y(n_3013)
);

CKINVDCx5p33_ASAP7_75t_R g3014 ( 
.A(n_2084),
.Y(n_3014)
);

AOI21xp5_ASAP7_75t_L g3015 ( 
.A1(n_2736),
.A2(n_2835),
.B(n_2774),
.Y(n_3015)
);

OAI21xp5_ASAP7_75t_L g3016 ( 
.A1(n_2733),
.A2(n_2776),
.B(n_2771),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2876),
.B(n_2949),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_SL g3018 ( 
.A(n_2809),
.B(n_2811),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2804),
.B(n_1965),
.Y(n_3019)
);

BUFx12f_ASAP7_75t_L g3020 ( 
.A(n_2814),
.Y(n_3020)
);

AOI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_2176),
.A2(n_2260),
.B(n_2213),
.Y(n_3021)
);

A2O1A1Ixp33_ASAP7_75t_L g3022 ( 
.A1(n_2471),
.A2(n_2475),
.B(n_2478),
.C(n_2473),
.Y(n_3022)
);

AOI21xp5_ASAP7_75t_L g3023 ( 
.A1(n_2176),
.A2(n_2260),
.B(n_2213),
.Y(n_3023)
);

A2O1A1Ixp33_ASAP7_75t_L g3024 ( 
.A1(n_2485),
.A2(n_2530),
.B(n_2567),
.C(n_2545),
.Y(n_3024)
);

O2A1O1Ixp33_ASAP7_75t_L g3025 ( 
.A1(n_2527),
.A2(n_2659),
.B(n_2667),
.C(n_2621),
.Y(n_3025)
);

AOI21x1_ASAP7_75t_L g3026 ( 
.A1(n_2579),
.A2(n_2758),
.B(n_2635),
.Y(n_3026)
);

BUFx6f_ASAP7_75t_L g3027 ( 
.A(n_2037),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_1965),
.B(n_1967),
.Y(n_3028)
);

AND2x2_ASAP7_75t_L g3029 ( 
.A(n_1939),
.B(n_1941),
.Y(n_3029)
);

AND2x4_ASAP7_75t_L g3030 ( 
.A(n_2267),
.B(n_2768),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_1967),
.B(n_1998),
.Y(n_3031)
);

O2A1O1Ixp5_ASAP7_75t_L g3032 ( 
.A1(n_2957),
.A2(n_2687),
.B(n_2691),
.C(n_2671),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2319),
.Y(n_3033)
);

AOI21xp5_ASAP7_75t_L g3034 ( 
.A1(n_1971),
.A2(n_2758),
.B(n_2635),
.Y(n_3034)
);

AOI21xp5_ASAP7_75t_L g3035 ( 
.A1(n_2779),
.A2(n_2829),
.B(n_2824),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_1998),
.B(n_2009),
.Y(n_3036)
);

A2O1A1Ixp33_ASAP7_75t_L g3037 ( 
.A1(n_2697),
.A2(n_2700),
.B(n_2719),
.C(n_2699),
.Y(n_3037)
);

AOI21xp5_ASAP7_75t_L g3038 ( 
.A1(n_2779),
.A2(n_2806),
.B(n_2036),
.Y(n_3038)
);

NOR2xp33_ASAP7_75t_L g3039 ( 
.A(n_2743),
.B(n_2744),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2918),
.B(n_1981),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2320),
.Y(n_3041)
);

OAI21xp5_ASAP7_75t_L g3042 ( 
.A1(n_2856),
.A2(n_2935),
.B(n_2931),
.Y(n_3042)
);

AOI21xp5_ASAP7_75t_L g3043 ( 
.A1(n_2030),
.A2(n_2313),
.B(n_2008),
.Y(n_3043)
);

AND2x2_ASAP7_75t_L g3044 ( 
.A(n_1939),
.B(n_1941),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2320),
.Y(n_3045)
);

AOI22xp5_ASAP7_75t_L g3046 ( 
.A1(n_2757),
.A2(n_2778),
.B1(n_2794),
.B2(n_2786),
.Y(n_3046)
);

AOI21xp5_ASAP7_75t_L g3047 ( 
.A1(n_2313),
.A2(n_2312),
.B(n_2823),
.Y(n_3047)
);

AOI21xp5_ASAP7_75t_L g3048 ( 
.A1(n_2828),
.A2(n_2854),
.B(n_2832),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2918),
.B(n_2025),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2329),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_1986),
.B(n_1991),
.Y(n_3051)
);

AOI22x1_ASAP7_75t_L g3052 ( 
.A1(n_2954),
.A2(n_2529),
.B1(n_2952),
.B2(n_2663),
.Y(n_3052)
);

NOR2xp33_ASAP7_75t_L g3053 ( 
.A(n_2834),
.B(n_2861),
.Y(n_3053)
);

O2A1O1Ixp33_ASAP7_75t_SL g3054 ( 
.A1(n_2864),
.A2(n_2897),
.B(n_2906),
.C(n_2904),
.Y(n_3054)
);

AOI21xp5_ASAP7_75t_L g3055 ( 
.A1(n_2916),
.A2(n_1978),
.B(n_2016),
.Y(n_3055)
);

AOI22xp33_ASAP7_75t_L g3056 ( 
.A1(n_2376),
.A2(n_2384),
.B1(n_2460),
.B2(n_2426),
.Y(n_3056)
);

AOI21xp5_ASAP7_75t_L g3057 ( 
.A1(n_2094),
.A2(n_2105),
.B(n_2101),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_SL g3058 ( 
.A(n_1959),
.B(n_1985),
.Y(n_3058)
);

OAI21xp5_ASAP7_75t_L g3059 ( 
.A1(n_2500),
.A2(n_1942),
.B(n_1935),
.Y(n_3059)
);

INVx2_ASAP7_75t_L g3060 ( 
.A(n_2942),
.Y(n_3060)
);

AOI21xp5_ASAP7_75t_L g3061 ( 
.A1(n_2107),
.A2(n_2120),
.B(n_2119),
.Y(n_3061)
);

OAI21xp5_ASAP7_75t_L g3062 ( 
.A1(n_1951),
.A2(n_1979),
.B(n_1968),
.Y(n_3062)
);

NOR3xp33_ASAP7_75t_L g3063 ( 
.A(n_1983),
.B(n_1977),
.C(n_1964),
.Y(n_3063)
);

OAI22xp5_ASAP7_75t_L g3064 ( 
.A1(n_1943),
.A2(n_2321),
.B1(n_2369),
.B2(n_2342),
.Y(n_3064)
);

OAI21xp5_ASAP7_75t_L g3065 ( 
.A1(n_1955),
.A2(n_1987),
.B(n_2377),
.Y(n_3065)
);

NOR2xp33_ASAP7_75t_L g3066 ( 
.A(n_2341),
.B(n_2838),
.Y(n_3066)
);

BUFx3_ASAP7_75t_L g3067 ( 
.A(n_2602),
.Y(n_3067)
);

AOI21xp5_ASAP7_75t_L g3068 ( 
.A1(n_2121),
.A2(n_2241),
.B(n_2239),
.Y(n_3068)
);

AOI21xp5_ASAP7_75t_L g3069 ( 
.A1(n_2251),
.A2(n_2064),
.B(n_2959),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2329),
.Y(n_3070)
);

OAI21xp5_ASAP7_75t_L g3071 ( 
.A1(n_2387),
.A2(n_2419),
.B(n_2401),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_1936),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_1986),
.B(n_1991),
.Y(n_3073)
);

NOR2xp33_ASAP7_75t_L g3074 ( 
.A(n_2341),
.B(n_2838),
.Y(n_3074)
);

NOR2xp67_ASAP7_75t_L g3075 ( 
.A(n_2059),
.B(n_1937),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_SL g3076 ( 
.A(n_2063),
.B(n_2633),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_SL g3077 ( 
.A(n_2014),
.B(n_2438),
.Y(n_3077)
);

BUFx6f_ASAP7_75t_L g3078 ( 
.A(n_2768),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_1993),
.B(n_2355),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_1993),
.B(n_2355),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2661),
.B(n_2677),
.Y(n_3081)
);

OAI21xp33_ASAP7_75t_L g3082 ( 
.A1(n_2451),
.A2(n_2466),
.B(n_2463),
.Y(n_3082)
);

OAI21xp5_ASAP7_75t_L g3083 ( 
.A1(n_2502),
.A2(n_2509),
.B(n_2506),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2940),
.Y(n_3084)
);

NAND3xp33_ASAP7_75t_L g3085 ( 
.A(n_2937),
.B(n_2514),
.C(n_2513),
.Y(n_3085)
);

AOI21xp5_ASAP7_75t_L g3086 ( 
.A1(n_2941),
.A2(n_2524),
.B(n_2518),
.Y(n_3086)
);

AOI21xp5_ASAP7_75t_L g3087 ( 
.A1(n_2525),
.A2(n_2548),
.B(n_2533),
.Y(n_3087)
);

BUFx8_ASAP7_75t_L g3088 ( 
.A(n_2084),
.Y(n_3088)
);

A2O1A1Ixp33_ASAP7_75t_L g3089 ( 
.A1(n_1954),
.A2(n_1975),
.B(n_1934),
.C(n_1947),
.Y(n_3089)
);

AOI21x1_ASAP7_75t_L g3090 ( 
.A1(n_2308),
.A2(n_2301),
.B(n_2273),
.Y(n_3090)
);

BUFx24_ASAP7_75t_L g3091 ( 
.A(n_2177),
.Y(n_3091)
);

BUFx3_ASAP7_75t_L g3092 ( 
.A(n_2602),
.Y(n_3092)
);

NOR2xp33_ASAP7_75t_L g3093 ( 
.A(n_2566),
.B(n_2569),
.Y(n_3093)
);

BUFx3_ASAP7_75t_L g3094 ( 
.A(n_2853),
.Y(n_3094)
);

AOI21xp5_ASAP7_75t_L g3095 ( 
.A1(n_2591),
.A2(n_2611),
.B(n_2606),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_SL g3096 ( 
.A(n_2617),
.B(n_2622),
.Y(n_3096)
);

BUFx4f_ASAP7_75t_L g3097 ( 
.A(n_2572),
.Y(n_3097)
);

AOI21xp5_ASAP7_75t_L g3098 ( 
.A1(n_2629),
.A2(n_2639),
.B(n_2630),
.Y(n_3098)
);

AND2x6_ASAP7_75t_L g3099 ( 
.A(n_2135),
.B(n_2229),
.Y(n_3099)
);

A2O1A1Ixp33_ASAP7_75t_L g3100 ( 
.A1(n_1938),
.A2(n_1962),
.B(n_1969),
.C(n_1950),
.Y(n_3100)
);

NOR2xp33_ASAP7_75t_L g3101 ( 
.A(n_2640),
.B(n_2642),
.Y(n_3101)
);

NOR2xp33_ASAP7_75t_L g3102 ( 
.A(n_2655),
.B(n_2665),
.Y(n_3102)
);

AOI33xp33_ASAP7_75t_L g3103 ( 
.A1(n_2022),
.A2(n_2066),
.A3(n_2491),
.B1(n_2558),
.B2(n_2557),
.B3(n_2482),
.Y(n_3103)
);

NOR2xp33_ASAP7_75t_L g3104 ( 
.A(n_2668),
.B(n_2688),
.Y(n_3104)
);

NOR2xp33_ASAP7_75t_L g3105 ( 
.A(n_2701),
.B(n_2705),
.Y(n_3105)
);

AOI22xp5_ASAP7_75t_L g3106 ( 
.A1(n_1931),
.A2(n_2325),
.B1(n_2330),
.B2(n_2322),
.Y(n_3106)
);

AOI22xp5_ASAP7_75t_L g3107 ( 
.A1(n_2333),
.A2(n_2346),
.B1(n_2348),
.B2(n_2340),
.Y(n_3107)
);

CKINVDCx10_ASAP7_75t_R g3108 ( 
.A(n_2637),
.Y(n_3108)
);

O2A1O1Ixp5_ASAP7_75t_L g3109 ( 
.A1(n_2713),
.A2(n_2750),
.B(n_2755),
.C(n_2714),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2335),
.Y(n_3110)
);

AND2x2_ASAP7_75t_L g3111 ( 
.A(n_1956),
.B(n_1957),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2661),
.B(n_2677),
.Y(n_3112)
);

BUFx8_ASAP7_75t_SL g3113 ( 
.A(n_2745),
.Y(n_3113)
);

AOI22xp33_ASAP7_75t_L g3114 ( 
.A1(n_2564),
.A2(n_2595),
.B1(n_2616),
.B2(n_2594),
.Y(n_3114)
);

AOI21xp5_ASAP7_75t_L g3115 ( 
.A1(n_2766),
.A2(n_2787),
.B(n_2772),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2741),
.B(n_2912),
.Y(n_3116)
);

O2A1O1Ixp33_ASAP7_75t_L g3117 ( 
.A1(n_2852),
.A2(n_2914),
.B(n_2863),
.C(n_2819),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_SL g3118 ( 
.A(n_2795),
.B(n_2839),
.Y(n_3118)
);

BUFx6f_ASAP7_75t_L g3119 ( 
.A(n_2285),
.Y(n_3119)
);

NOR2xp33_ASAP7_75t_L g3120 ( 
.A(n_2849),
.B(n_2860),
.Y(n_3120)
);

AOI21xp5_ASAP7_75t_L g3121 ( 
.A1(n_2351),
.A2(n_2364),
.B(n_2357),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_SL g3122 ( 
.A(n_2868),
.B(n_2871),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_SL g3123 ( 
.A(n_2881),
.B(n_2917),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2741),
.B(n_2912),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2244),
.B(n_2248),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2244),
.B(n_2248),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2249),
.B(n_2090),
.Y(n_3127)
);

OAI22xp5_ASAP7_75t_L g3128 ( 
.A1(n_2920),
.A2(n_2928),
.B1(n_2368),
.B2(n_2372),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2249),
.B(n_1972),
.Y(n_3129)
);

OAI21xp33_ASAP7_75t_L g3130 ( 
.A1(n_2354),
.A2(n_2374),
.B(n_2373),
.Y(n_3130)
);

OAI22xp5_ASAP7_75t_L g3131 ( 
.A1(n_2378),
.A2(n_2393),
.B1(n_2399),
.B2(n_2382),
.Y(n_3131)
);

NOR2xp33_ASAP7_75t_SL g3132 ( 
.A(n_2334),
.B(n_2572),
.Y(n_3132)
);

CKINVDCx8_ASAP7_75t_R g3133 ( 
.A(n_2274),
.Y(n_3133)
);

INVxp33_ASAP7_75t_SL g3134 ( 
.A(n_2356),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_1972),
.B(n_2113),
.Y(n_3135)
);

AOI21xp5_ASAP7_75t_L g3136 ( 
.A1(n_2403),
.A2(n_2406),
.B(n_2404),
.Y(n_3136)
);

OAI22xp5_ASAP7_75t_L g3137 ( 
.A1(n_2410),
.A2(n_2413),
.B1(n_2416),
.B2(n_2411),
.Y(n_3137)
);

AOI21xp33_ASAP7_75t_L g3138 ( 
.A1(n_1933),
.A2(n_2657),
.B(n_2651),
.Y(n_3138)
);

AOI21xp5_ASAP7_75t_L g3139 ( 
.A1(n_2418),
.A2(n_2425),
.B(n_2420),
.Y(n_3139)
);

HB1xp67_ASAP7_75t_L g3140 ( 
.A(n_2440),
.Y(n_3140)
);

AOI21xp5_ASAP7_75t_L g3141 ( 
.A1(n_2421),
.A2(n_2435),
.B(n_2431),
.Y(n_3141)
);

NOR2xp33_ASAP7_75t_L g3142 ( 
.A(n_2439),
.B(n_2442),
.Y(n_3142)
);

AOI21xp5_ASAP7_75t_L g3143 ( 
.A1(n_2453),
.A2(n_2456),
.B(n_2455),
.Y(n_3143)
);

NOR2xp33_ASAP7_75t_L g3144 ( 
.A(n_2449),
.B(n_2459),
.Y(n_3144)
);

INVx2_ASAP7_75t_L g3145 ( 
.A(n_2940),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_2943),
.Y(n_3146)
);

AND2x2_ASAP7_75t_L g3147 ( 
.A(n_1956),
.B(n_1957),
.Y(n_3147)
);

AOI21xp5_ASAP7_75t_L g3148 ( 
.A1(n_2467),
.A2(n_2479),
.B(n_2469),
.Y(n_3148)
);

NOR2xp33_ASAP7_75t_L g3149 ( 
.A(n_2484),
.B(n_2486),
.Y(n_3149)
);

AOI21xp33_ASAP7_75t_L g3150 ( 
.A1(n_2662),
.A2(n_2708),
.B(n_2703),
.Y(n_3150)
);

OAI321xp33_ASAP7_75t_L g3151 ( 
.A1(n_2710),
.A2(n_2759),
.A3(n_2722),
.B1(n_2770),
.B2(n_2726),
.C(n_2715),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2113),
.B(n_1976),
.Y(n_3152)
);

AOI21xp5_ASAP7_75t_L g3153 ( 
.A1(n_2490),
.A2(n_2496),
.B(n_2495),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_1980),
.B(n_1990),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_1992),
.B(n_1999),
.Y(n_3155)
);

BUFx2_ASAP7_75t_L g3156 ( 
.A(n_2243),
.Y(n_3156)
);

OAI21xp5_ASAP7_75t_L g3157 ( 
.A1(n_2061),
.A2(n_2503),
.B(n_2501),
.Y(n_3157)
);

INVx2_ASAP7_75t_SL g3158 ( 
.A(n_2337),
.Y(n_3158)
);

BUFx12f_ASAP7_75t_L g3159 ( 
.A(n_2814),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2000),
.B(n_2006),
.Y(n_3160)
);

OAI21xp5_ASAP7_75t_L g3161 ( 
.A1(n_2504),
.A2(n_2507),
.B(n_2505),
.Y(n_3161)
);

AO21x2_ASAP7_75t_L g3162 ( 
.A1(n_2243),
.A2(n_2344),
.B(n_2335),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_2011),
.B(n_2012),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_SL g3164 ( 
.A(n_2092),
.B(n_2740),
.Y(n_3164)
);

INVx4_ASAP7_75t_L g3165 ( 
.A(n_1937),
.Y(n_3165)
);

AOI21xp5_ASAP7_75t_L g3166 ( 
.A1(n_2508),
.A2(n_2517),
.B(n_2510),
.Y(n_3166)
);

BUFx2_ASAP7_75t_L g3167 ( 
.A(n_2344),
.Y(n_3167)
);

OAI21xp5_ASAP7_75t_L g3168 ( 
.A1(n_2520),
.A2(n_2536),
.B(n_2526),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2353),
.Y(n_3169)
);

NOR2xp33_ASAP7_75t_L g3170 ( 
.A(n_2543),
.B(n_2549),
.Y(n_3170)
);

NOR2x1_ASAP7_75t_L g3171 ( 
.A(n_1937),
.B(n_2046),
.Y(n_3171)
);

AOI21xp5_ASAP7_75t_L g3172 ( 
.A1(n_2552),
.A2(n_2562),
.B(n_2560),
.Y(n_3172)
);

OR2x2_ASAP7_75t_L g3173 ( 
.A(n_2017),
.B(n_2947),
.Y(n_3173)
);

A2O1A1Ixp33_ASAP7_75t_L g3174 ( 
.A1(n_2013),
.A2(n_2028),
.B(n_2020),
.C(n_2099),
.Y(n_3174)
);

AOI21xp5_ASAP7_75t_L g3175 ( 
.A1(n_2568),
.A2(n_2578),
.B(n_2577),
.Y(n_3175)
);

AOI21xp5_ASAP7_75t_L g3176 ( 
.A1(n_2581),
.A2(n_2585),
.B(n_2584),
.Y(n_3176)
);

OAI21xp33_ASAP7_75t_SL g3177 ( 
.A1(n_2043),
.A2(n_2740),
.B(n_1982),
.Y(n_3177)
);

AOI21xp5_ASAP7_75t_L g3178 ( 
.A1(n_2587),
.A2(n_2598),
.B(n_2593),
.Y(n_3178)
);

AOI21xp5_ASAP7_75t_L g3179 ( 
.A1(n_2605),
.A2(n_2613),
.B(n_2607),
.Y(n_3179)
);

AOI21xp5_ASAP7_75t_L g3180 ( 
.A1(n_2620),
.A2(n_2624),
.B(n_2623),
.Y(n_3180)
);

O2A1O1Ixp33_ASAP7_75t_L g3181 ( 
.A1(n_2625),
.A2(n_2644),
.B(n_2649),
.C(n_2632),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2353),
.Y(n_3182)
);

NOR2xp33_ASAP7_75t_SL g3183 ( 
.A(n_2637),
.B(n_2286),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_SL g3184 ( 
.A(n_2317),
.B(n_2675),
.Y(n_3184)
);

AOI21xp5_ASAP7_75t_L g3185 ( 
.A1(n_2653),
.A2(n_2676),
.B(n_2672),
.Y(n_3185)
);

AOI21xp5_ASAP7_75t_L g3186 ( 
.A1(n_2678),
.A2(n_2682),
.B(n_2679),
.Y(n_3186)
);

AOI21xp5_ASAP7_75t_L g3187 ( 
.A1(n_2683),
.A2(n_2686),
.B(n_2685),
.Y(n_3187)
);

AOI21xp5_ASAP7_75t_L g3188 ( 
.A1(n_2689),
.A2(n_2702),
.B(n_2692),
.Y(n_3188)
);

NOR2xp33_ASAP7_75t_SL g3189 ( 
.A(n_2415),
.B(n_2493),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2114),
.B(n_2034),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_L g3191 ( 
.A(n_2706),
.B(n_2707),
.Y(n_3191)
);

INVxp67_ASAP7_75t_L g3192 ( 
.A(n_1995),
.Y(n_3192)
);

AOI21xp5_ASAP7_75t_L g3193 ( 
.A1(n_2711),
.A2(n_2718),
.B(n_2716),
.Y(n_3193)
);

NOR2xp33_ASAP7_75t_L g3194 ( 
.A(n_2720),
.B(n_2724),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_SL g3195 ( 
.A(n_2769),
.B(n_2850),
.Y(n_3195)
);

AOI21xp5_ASAP7_75t_L g3196 ( 
.A1(n_2727),
.A2(n_2739),
.B(n_2729),
.Y(n_3196)
);

NOR2xp33_ASAP7_75t_L g3197 ( 
.A(n_2748),
.B(n_2749),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2751),
.B(n_2762),
.Y(n_3198)
);

BUFx2_ASAP7_75t_L g3199 ( 
.A(n_2359),
.Y(n_3199)
);

NOR2xp67_ASAP7_75t_L g3200 ( 
.A(n_2046),
.B(n_2417),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_2785),
.B(n_2788),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_2792),
.B(n_2810),
.Y(n_3202)
);

AOI21xp5_ASAP7_75t_L g3203 ( 
.A1(n_2813),
.A2(n_2825),
.B(n_2817),
.Y(n_3203)
);

O2A1O1Ixp33_ASAP7_75t_L g3204 ( 
.A1(n_2826),
.A2(n_2841),
.B(n_2848),
.C(n_2833),
.Y(n_3204)
);

AOI21xp5_ASAP7_75t_L g3205 ( 
.A1(n_2851),
.A2(n_2862),
.B(n_2855),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_SL g3206 ( 
.A(n_2895),
.B(n_2880),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2883),
.B(n_2884),
.Y(n_3207)
);

AOI21xp5_ASAP7_75t_L g3208 ( 
.A1(n_2892),
.A2(n_2894),
.B(n_2893),
.Y(n_3208)
);

O2A1O1Ixp33_ASAP7_75t_L g3209 ( 
.A1(n_2899),
.A2(n_2901),
.B(n_2905),
.C(n_2900),
.Y(n_3209)
);

BUFx2_ASAP7_75t_L g3210 ( 
.A(n_2359),
.Y(n_3210)
);

AOI21xp5_ASAP7_75t_L g3211 ( 
.A1(n_2907),
.A2(n_2927),
.B(n_2913),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2930),
.B(n_2936),
.Y(n_3212)
);

O2A1O1Ixp5_ASAP7_75t_L g3213 ( 
.A1(n_2140),
.A2(n_2151),
.B(n_2155),
.C(n_2147),
.Y(n_3213)
);

BUFx6f_ASAP7_75t_L g3214 ( 
.A(n_2315),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_SL g3215 ( 
.A(n_2955),
.B(n_2646),
.Y(n_3215)
);

BUFx2_ASAP7_75t_L g3216 ( 
.A(n_2363),
.Y(n_3216)
);

OAI21xp33_ASAP7_75t_L g3217 ( 
.A1(n_2646),
.A2(n_1961),
.B(n_1960),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_1958),
.B(n_1982),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2363),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2366),
.Y(n_3220)
);

NOR3xp33_ASAP7_75t_L g3221 ( 
.A(n_2193),
.B(n_2160),
.C(n_2024),
.Y(n_3221)
);

AOI21xp5_ASAP7_75t_L g3222 ( 
.A1(n_2002),
.A2(n_2031),
.B(n_2004),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_2366),
.Y(n_3223)
);

O2A1O1Ixp33_ASAP7_75t_L g3224 ( 
.A1(n_2032),
.A2(n_2041),
.B(n_2172),
.C(n_2162),
.Y(n_3224)
);

AND2x2_ASAP7_75t_L g3225 ( 
.A(n_1958),
.B(n_2076),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_SL g3226 ( 
.A(n_2184),
.B(n_2093),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_SL g3227 ( 
.A(n_2361),
.B(n_2388),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2383),
.Y(n_3228)
);

INVxp67_ASAP7_75t_L g3229 ( 
.A(n_1997),
.Y(n_3229)
);

AOI21xp5_ASAP7_75t_L g3230 ( 
.A1(n_2310),
.A2(n_2311),
.B(n_2069),
.Y(n_3230)
);

AOI21x1_ASAP7_75t_L g3231 ( 
.A1(n_2308),
.A2(n_2305),
.B(n_2307),
.Y(n_3231)
);

OR2x2_ASAP7_75t_L g3232 ( 
.A(n_2017),
.B(n_2332),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_2383),
.Y(n_3233)
);

NOR2xp33_ASAP7_75t_L g3234 ( 
.A(n_2023),
.B(n_2379),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_2071),
.B(n_2371),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_SL g3236 ( 
.A(n_2391),
.B(n_2446),
.Y(n_3236)
);

OAI21xp33_ASAP7_75t_SL g3237 ( 
.A1(n_2043),
.A2(n_2822),
.B(n_2807),
.Y(n_3237)
);

AOI21xp5_ASAP7_75t_L g3238 ( 
.A1(n_2309),
.A2(n_2253),
.B(n_2229),
.Y(n_3238)
);

AOI21x1_ASAP7_75t_L g3239 ( 
.A1(n_2386),
.A2(n_2412),
.B(n_2400),
.Y(n_3239)
);

AOI21xp5_ASAP7_75t_L g3240 ( 
.A1(n_2135),
.A2(n_2229),
.B(n_2145),
.Y(n_3240)
);

AND2x2_ASAP7_75t_SL g3241 ( 
.A(n_2371),
.B(n_2857),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_2071),
.B(n_1994),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2386),
.Y(n_3243)
);

OAI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_2072),
.A2(n_2073),
.B(n_2066),
.Y(n_3244)
);

AOI21xp5_ASAP7_75t_L g3245 ( 
.A1(n_2135),
.A2(n_2153),
.B(n_2143),
.Y(n_3245)
);

AOI21xp5_ASAP7_75t_L g3246 ( 
.A1(n_2161),
.A2(n_2169),
.B(n_2166),
.Y(n_3246)
);

OAI21xp5_ASAP7_75t_L g3247 ( 
.A1(n_2157),
.A2(n_2209),
.B(n_2178),
.Y(n_3247)
);

OAI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_2173),
.A2(n_2123),
.B(n_2111),
.Y(n_3248)
);

AND2x2_ASAP7_75t_L g3249 ( 
.A(n_2076),
.B(n_2100),
.Y(n_3249)
);

OAI21xp5_ASAP7_75t_L g3250 ( 
.A1(n_2137),
.A2(n_2154),
.B(n_2150),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_1994),
.B(n_2026),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_SL g3252 ( 
.A(n_2450),
.B(n_2680),
.Y(n_3252)
);

AOI21xp5_ASAP7_75t_L g3253 ( 
.A1(n_2170),
.A2(n_2186),
.B(n_2183),
.Y(n_3253)
);

AOI22x1_ASAP7_75t_L g3254 ( 
.A1(n_2133),
.A2(n_2725),
.B1(n_2840),
.B2(n_2638),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_2026),
.B(n_2035),
.Y(n_3255)
);

AOI21xp5_ASAP7_75t_L g3256 ( 
.A1(n_2190),
.A2(n_2201),
.B(n_2192),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_2035),
.B(n_2038),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_2038),
.B(n_2052),
.Y(n_3258)
);

BUFx6f_ASAP7_75t_L g3259 ( 
.A(n_2315),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_2400),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_2052),
.B(n_2074),
.Y(n_3261)
);

OAI22xp5_ASAP7_75t_L g3262 ( 
.A1(n_2882),
.A2(n_2951),
.B1(n_2799),
.B2(n_2040),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_2074),
.B(n_2102),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2412),
.Y(n_3264)
);

AOI22xp5_ASAP7_75t_L g3265 ( 
.A1(n_2062),
.A2(n_2045),
.B1(n_2047),
.B2(n_2039),
.Y(n_3265)
);

AOI21xp5_ASAP7_75t_L g3266 ( 
.A1(n_2204),
.A2(n_2210),
.B(n_2205),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_2950),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_2102),
.B(n_2167),
.Y(n_3268)
);

O2A1O1Ixp33_ASAP7_75t_L g3269 ( 
.A1(n_2001),
.A2(n_2021),
.B(n_2110),
.C(n_2087),
.Y(n_3269)
);

NAND3xp33_ASAP7_75t_L g3270 ( 
.A(n_2086),
.B(n_2175),
.C(n_2168),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_L g3271 ( 
.A(n_2167),
.B(n_2171),
.Y(n_3271)
);

OAI21xp5_ASAP7_75t_L g3272 ( 
.A1(n_2179),
.A2(n_2106),
.B(n_2100),
.Y(n_3272)
);

NAND2xp33_ASAP7_75t_L g3273 ( 
.A(n_2831),
.B(n_2018),
.Y(n_3273)
);

HB1xp67_ASAP7_75t_L g3274 ( 
.A(n_2483),
.Y(n_3274)
);

OAI21xp5_ASAP7_75t_L g3275 ( 
.A1(n_2106),
.A2(n_2134),
.B(n_2117),
.Y(n_3275)
);

AOI21xp33_ASAP7_75t_L g3276 ( 
.A1(n_2565),
.A2(n_2803),
.B(n_2055),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_2171),
.B(n_2174),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_2174),
.B(n_2185),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_2185),
.B(n_2187),
.Y(n_3279)
);

AND2x4_ASAP7_75t_L g3280 ( 
.A(n_2046),
.B(n_2417),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2187),
.B(n_2189),
.Y(n_3281)
);

AND2x2_ASAP7_75t_L g3282 ( 
.A(n_2117),
.B(n_2134),
.Y(n_3282)
);

AOI21xp5_ASAP7_75t_L g3283 ( 
.A1(n_2214),
.A2(n_2223),
.B(n_2218),
.Y(n_3283)
);

AOI21xp5_ASAP7_75t_L g3284 ( 
.A1(n_2225),
.A2(n_2228),
.B(n_2226),
.Y(n_3284)
);

NOR2xp67_ASAP7_75t_L g3285 ( 
.A(n_2417),
.B(n_2470),
.Y(n_3285)
);

AOI22xp5_ASAP7_75t_L g3286 ( 
.A1(n_2062),
.A2(n_2051),
.B1(n_2095),
.B2(n_2589),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_2189),
.B(n_2211),
.Y(n_3287)
);

BUFx6f_ASAP7_75t_L g3288 ( 
.A(n_2550),
.Y(n_3288)
);

OAI21xp5_ASAP7_75t_L g3289 ( 
.A1(n_2144),
.A2(n_2227),
.B(n_2194),
.Y(n_3289)
);

AND2x2_ASAP7_75t_L g3290 ( 
.A(n_2144),
.B(n_2194),
.Y(n_3290)
);

BUFx2_ASAP7_75t_L g3291 ( 
.A(n_2414),
.Y(n_3291)
);

A2O1A1Ixp33_ASAP7_75t_L g3292 ( 
.A1(n_2078),
.A2(n_2062),
.B(n_2242),
.C(n_2068),
.Y(n_3292)
);

AOI21xp5_ASAP7_75t_L g3293 ( 
.A1(n_2234),
.A2(n_2247),
.B(n_2470),
.Y(n_3293)
);

NOR2xp67_ASAP7_75t_L g3294 ( 
.A(n_2470),
.B(n_2555),
.Y(n_3294)
);

HB1xp67_ASAP7_75t_L g3295 ( 
.A(n_2695),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_2211),
.B(n_2219),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_2219),
.B(n_2230),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_2230),
.B(n_2231),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_2231),
.B(n_2235),
.Y(n_3299)
);

AOI21x1_ASAP7_75t_L g3300 ( 
.A1(n_2429),
.A2(n_2457),
.B(n_2448),
.Y(n_3300)
);

NOR2xp33_ASAP7_75t_L g3301 ( 
.A(n_2921),
.B(n_2521),
.Y(n_3301)
);

OR2x6_ASAP7_75t_L g3302 ( 
.A(n_2108),
.B(n_2550),
.Y(n_3302)
);

NOR2xp33_ASAP7_75t_L g3303 ( 
.A(n_2745),
.B(n_1970),
.Y(n_3303)
);

AND2x4_ASAP7_75t_L g3304 ( 
.A(n_2555),
.B(n_2576),
.Y(n_3304)
);

AO21x1_ASAP7_75t_L g3305 ( 
.A1(n_2235),
.A2(n_2448),
.B(n_2429),
.Y(n_3305)
);

O2A1O1Ixp33_ASAP7_75t_L g3306 ( 
.A1(n_2789),
.A2(n_2843),
.B(n_2902),
.C(n_2878),
.Y(n_3306)
);

AOI21xp5_ASAP7_75t_L g3307 ( 
.A1(n_2555),
.A2(n_2592),
.B(n_2576),
.Y(n_3307)
);

AND2x2_ASAP7_75t_L g3308 ( 
.A(n_2227),
.B(n_1940),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_1940),
.B(n_1949),
.Y(n_3309)
);

AOI21xp5_ASAP7_75t_L g3310 ( 
.A1(n_2576),
.A2(n_2601),
.B(n_2592),
.Y(n_3310)
);

OAI21xp5_ASAP7_75t_L g3311 ( 
.A1(n_2457),
.A2(n_2468),
.B(n_2465),
.Y(n_3311)
);

OAI22xp5_ASAP7_75t_L g3312 ( 
.A1(n_2853),
.A2(n_2232),
.B1(n_2199),
.B2(n_2261),
.Y(n_3312)
);

INVx2_ASAP7_75t_SL g3313 ( 
.A(n_2337),
.Y(n_3313)
);

NOR2xp33_ASAP7_75t_SL g3314 ( 
.A(n_2673),
.B(n_2704),
.Y(n_3314)
);

OAI22xp5_ASAP7_75t_L g3315 ( 
.A1(n_2075),
.A2(n_2133),
.B1(n_2200),
.B2(n_2207),
.Y(n_3315)
);

OAI21xp33_ASAP7_75t_L g3316 ( 
.A1(n_2717),
.A2(n_2791),
.B(n_2767),
.Y(n_3316)
);

NOR2xp33_ASAP7_75t_SL g3317 ( 
.A(n_2805),
.B(n_2139),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_1949),
.B(n_1963),
.Y(n_3318)
);

NOR2xp33_ASAP7_75t_L g3319 ( 
.A(n_1970),
.B(n_2370),
.Y(n_3319)
);

OAI21xp5_ASAP7_75t_L g3320 ( 
.A1(n_2465),
.A2(n_2477),
.B(n_2468),
.Y(n_3320)
);

O2A1O1Ixp33_ASAP7_75t_L g3321 ( 
.A1(n_2276),
.A2(n_2279),
.B(n_2255),
.C(n_2122),
.Y(n_3321)
);

AOI21xp5_ASAP7_75t_L g3322 ( 
.A1(n_2592),
.A2(n_2608),
.B(n_2601),
.Y(n_3322)
);

INVx3_ASAP7_75t_L g3323 ( 
.A(n_2601),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_1963),
.B(n_1973),
.Y(n_3324)
);

OAI21xp5_ASAP7_75t_L g3325 ( 
.A1(n_2477),
.A2(n_2494),
.B(n_2488),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_1973),
.B(n_1974),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_L g3327 ( 
.A(n_1974),
.B(n_1984),
.Y(n_3327)
);

AOI21xp5_ASAP7_75t_L g3328 ( 
.A1(n_2608),
.A2(n_2798),
.B(n_2619),
.Y(n_3328)
);

A2O1A1Ixp33_ASAP7_75t_L g3329 ( 
.A1(n_2264),
.A2(n_2268),
.B(n_2142),
.C(n_2298),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_L g3330 ( 
.A(n_1984),
.B(n_2281),
.Y(n_3330)
);

AOI21xp5_ASAP7_75t_L g3331 ( 
.A1(n_2608),
.A2(n_2798),
.B(n_2619),
.Y(n_3331)
);

AOI21xp5_ASAP7_75t_L g3332 ( 
.A1(n_2619),
.A2(n_2844),
.B(n_2798),
.Y(n_3332)
);

OAI22xp5_ASAP7_75t_L g3333 ( 
.A1(n_2133),
.A2(n_2050),
.B1(n_2156),
.B2(n_1966),
.Y(n_3333)
);

AOI21xp5_ASAP7_75t_L g3334 ( 
.A1(n_2844),
.A2(n_2494),
.B(n_2488),
.Y(n_3334)
);

AOI21xp5_ASAP7_75t_L g3335 ( 
.A1(n_2844),
.A2(n_2528),
.B(n_2512),
.Y(n_3335)
);

AOI21xp5_ASAP7_75t_L g3336 ( 
.A1(n_2512),
.A2(n_2531),
.B(n_2528),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_SL g3337 ( 
.A(n_2337),
.B(n_2339),
.Y(n_3337)
);

NOR2xp33_ASAP7_75t_L g3338 ( 
.A(n_2370),
.B(n_2647),
.Y(n_3338)
);

AOI21xp5_ASAP7_75t_L g3339 ( 
.A1(n_2531),
.A2(n_2547),
.B(n_2535),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_2535),
.Y(n_3340)
);

A2O1A1Ixp33_ASAP7_75t_L g3341 ( 
.A1(n_2164),
.A2(n_2220),
.B(n_2221),
.C(n_2215),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_SL g3342 ( 
.A(n_2337),
.B(n_2339),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_L g3343 ( 
.A(n_2281),
.B(n_2293),
.Y(n_3343)
);

NAND2x1p5_ASAP7_75t_L g3344 ( 
.A(n_2128),
.B(n_2547),
.Y(n_3344)
);

O2A1O1Ixp33_ASAP7_75t_L g3345 ( 
.A1(n_2304),
.A2(n_2280),
.B(n_2181),
.C(n_2132),
.Y(n_3345)
);

AOI21xp5_ASAP7_75t_L g3346 ( 
.A1(n_2553),
.A2(n_2582),
.B(n_2571),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_2293),
.B(n_2294),
.Y(n_3347)
);

AOI21xp5_ASAP7_75t_L g3348 ( 
.A1(n_2553),
.A2(n_2582),
.B(n_2571),
.Y(n_3348)
);

AOI21xp5_ASAP7_75t_L g3349 ( 
.A1(n_2583),
.A2(n_2603),
.B(n_2600),
.Y(n_3349)
);

AOI21xp5_ASAP7_75t_L g3350 ( 
.A1(n_2583),
.A2(n_2603),
.B(n_2600),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_2294),
.B(n_2240),
.Y(n_3351)
);

CKINVDCx5p33_ASAP7_75t_R g3352 ( 
.A(n_2077),
.Y(n_3352)
);

NOR2x1_ASAP7_75t_R g3353 ( 
.A(n_2879),
.B(n_2118),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_2240),
.B(n_2626),
.Y(n_3354)
);

OAI21xp5_ASAP7_75t_L g3355 ( 
.A1(n_2626),
.A2(n_2636),
.B(n_2628),
.Y(n_3355)
);

AOI21xp5_ASAP7_75t_L g3356 ( 
.A1(n_2628),
.A2(n_2664),
.B(n_2636),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_2664),
.Y(n_3357)
);

AOI21xp5_ASAP7_75t_L g3358 ( 
.A1(n_2681),
.A2(n_2693),
.B(n_2690),
.Y(n_3358)
);

A2O1A1Ixp33_ASAP7_75t_L g3359 ( 
.A1(n_2297),
.A2(n_2300),
.B(n_2272),
.C(n_2275),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_2681),
.B(n_2690),
.Y(n_3360)
);

AOI21x1_ASAP7_75t_L g3361 ( 
.A1(n_2693),
.A2(n_2721),
.B(n_2698),
.Y(n_3361)
);

A2O1A1Ixp33_ASAP7_75t_L g3362 ( 
.A1(n_2271),
.A2(n_2130),
.B(n_2128),
.C(n_2336),
.Y(n_3362)
);

AOI22xp5_ASAP7_75t_L g3363 ( 
.A1(n_1946),
.A2(n_2405),
.B1(n_2539),
.B2(n_1966),
.Y(n_3363)
);

O2A1O1Ixp33_ASAP7_75t_L g3364 ( 
.A1(n_2306),
.A2(n_2314),
.B(n_2195),
.C(n_2236),
.Y(n_3364)
);

AOI21xp5_ASAP7_75t_L g3365 ( 
.A1(n_2698),
.A2(n_2728),
.B(n_2721),
.Y(n_3365)
);

AOI21xp5_ASAP7_75t_L g3366 ( 
.A1(n_2728),
.A2(n_2735),
.B(n_2734),
.Y(n_3366)
);

A2O1A1Ixp33_ASAP7_75t_L g3367 ( 
.A1(n_2128),
.A2(n_2336),
.B(n_2586),
.C(n_2266),
.Y(n_3367)
);

OAI21xp5_ASAP7_75t_L g3368 ( 
.A1(n_2734),
.A2(n_2763),
.B(n_2735),
.Y(n_3368)
);

INVx3_ASAP7_75t_L g3369 ( 
.A(n_2550),
.Y(n_3369)
);

AOI21xp5_ASAP7_75t_L g3370 ( 
.A1(n_2763),
.A2(n_2784),
.B(n_2780),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_2780),
.B(n_2784),
.Y(n_3371)
);

AO21x1_ASAP7_75t_L g3372 ( 
.A1(n_2790),
.A2(n_2797),
.B(n_2796),
.Y(n_3372)
);

NOR2xp33_ASAP7_75t_L g3373 ( 
.A(n_2647),
.B(n_2738),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_SL g3374 ( 
.A(n_2337),
.B(n_2339),
.Y(n_3374)
);

BUFx2_ASAP7_75t_L g3375 ( 
.A(n_2790),
.Y(n_3375)
);

HB1xp67_ASAP7_75t_L g3376 ( 
.A(n_2246),
.Y(n_3376)
);

NOR2xp33_ASAP7_75t_L g3377 ( 
.A(n_2738),
.B(n_2783),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_2796),
.Y(n_3378)
);

NOR2xp33_ASAP7_75t_L g3379 ( 
.A(n_2783),
.B(n_2800),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_L g3380 ( 
.A(n_2797),
.B(n_2802),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_2802),
.B(n_2820),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_2820),
.B(n_2821),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2821),
.Y(n_3383)
);

OAI21x1_ASAP7_75t_L g3384 ( 
.A1(n_2827),
.A2(n_2865),
.B(n_2847),
.Y(n_3384)
);

INVx3_ASAP7_75t_L g3385 ( 
.A(n_2827),
.Y(n_3385)
);

AOI21xp5_ASAP7_75t_L g3386 ( 
.A1(n_2847),
.A2(n_2867),
.B(n_2865),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_2867),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_2874),
.B(n_2889),
.Y(n_3388)
);

HB1xp67_ASAP7_75t_L g3389 ( 
.A(n_2082),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_2874),
.B(n_2889),
.Y(n_3390)
);

NOR2xp33_ASAP7_75t_SL g3391 ( 
.A(n_2108),
.B(n_2885),
.Y(n_3391)
);

INVx5_ASAP7_75t_L g3392 ( 
.A(n_2083),
.Y(n_3392)
);

NOR2xp33_ASAP7_75t_L g3393 ( 
.A(n_2800),
.B(n_2879),
.Y(n_3393)
);

OAI21xp5_ASAP7_75t_L g3394 ( 
.A1(n_2891),
.A2(n_2923),
.B(n_2909),
.Y(n_3394)
);

AOI21xp33_ASAP7_75t_L g3395 ( 
.A1(n_2299),
.A2(n_2909),
.B(n_2891),
.Y(n_3395)
);

AOI21xp5_ASAP7_75t_L g3396 ( 
.A1(n_2923),
.A2(n_2938),
.B(n_2925),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_2925),
.B(n_2938),
.Y(n_3397)
);

O2A1O1Ixp5_ASAP7_75t_L g3398 ( 
.A1(n_2197),
.A2(n_2222),
.B(n_2237),
.C(n_2233),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_SL g3399 ( 
.A(n_2339),
.B(n_2422),
.Y(n_3399)
);

AOI21xp5_ASAP7_75t_L g3400 ( 
.A1(n_2944),
.A2(n_2398),
.B(n_2394),
.Y(n_3400)
);

AO21x1_ASAP7_75t_L g3401 ( 
.A1(n_2944),
.A2(n_2256),
.B(n_2245),
.Y(n_3401)
);

A2O1A1Ixp33_ASAP7_75t_L g3402 ( 
.A1(n_2336),
.A2(n_2586),
.B(n_2125),
.C(n_2126),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_2394),
.Y(n_3403)
);

AOI22xp5_ASAP7_75t_L g3404 ( 
.A1(n_1946),
.A2(n_2405),
.B1(n_2539),
.B2(n_1966),
.Y(n_3404)
);

AOI21xp5_ASAP7_75t_L g3405 ( 
.A1(n_2398),
.A2(n_2409),
.B(n_2407),
.Y(n_3405)
);

NOR2x1_ASAP7_75t_L g3406 ( 
.A(n_2316),
.B(n_2058),
.Y(n_3406)
);

NAND3xp33_ASAP7_75t_L g3407 ( 
.A(n_2104),
.B(n_2375),
.C(n_2287),
.Y(n_3407)
);

O2A1O1Ixp5_ASAP7_75t_L g3408 ( 
.A1(n_2258),
.A2(n_2259),
.B(n_2091),
.C(n_2302),
.Y(n_3408)
);

A2O1A1Ixp33_ASAP7_75t_L g3409 ( 
.A1(n_2586),
.A2(n_2131),
.B(n_2136),
.C(n_2124),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_2407),
.B(n_2409),
.Y(n_3410)
);

AOI21xp5_ASAP7_75t_L g3411 ( 
.A1(n_2434),
.A2(n_2444),
.B(n_2436),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_2434),
.B(n_2436),
.Y(n_3412)
);

INVx3_ASAP7_75t_L g3413 ( 
.A(n_2156),
.Y(n_3413)
);

OAI21xp33_ASAP7_75t_L g3414 ( 
.A1(n_2019),
.A2(n_2331),
.B(n_2326),
.Y(n_3414)
);

O2A1O1Ixp33_ASAP7_75t_L g3415 ( 
.A1(n_2057),
.A2(n_2316),
.B(n_2156),
.C(n_2007),
.Y(n_3415)
);

AOI21xp5_ASAP7_75t_L g3416 ( 
.A1(n_2474),
.A2(n_2492),
.B(n_2480),
.Y(n_3416)
);

AOI21xp5_ASAP7_75t_L g3417 ( 
.A1(n_2474),
.A2(n_2492),
.B(n_2480),
.Y(n_3417)
);

AOI21xp5_ASAP7_75t_L g3418 ( 
.A1(n_2497),
.A2(n_2540),
.B(n_2538),
.Y(n_3418)
);

NOR2xp33_ASAP7_75t_L g3419 ( 
.A(n_1989),
.B(n_2212),
.Y(n_3419)
);

OAI321xp33_ASAP7_75t_L g3420 ( 
.A1(n_2079),
.A2(n_2846),
.A3(n_1952),
.B1(n_2324),
.B2(n_2939),
.C(n_2658),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_2497),
.B(n_2538),
.Y(n_3421)
);

BUFx4f_ASAP7_75t_L g3422 ( 
.A(n_2083),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_2540),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_2542),
.B(n_2544),
.Y(n_3424)
);

AOI22xp5_ASAP7_75t_L g3425 ( 
.A1(n_1946),
.A2(n_2712),
.B1(n_2405),
.B2(n_2539),
.Y(n_3425)
);

O2A1O1Ixp33_ASAP7_75t_L g3426 ( 
.A1(n_2057),
.A2(n_1952),
.B(n_2945),
.C(n_2939),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_SL g3427 ( 
.A(n_2339),
.B(n_2422),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_2542),
.B(n_2544),
.Y(n_3428)
);

NOR2xp33_ASAP7_75t_L g3429 ( 
.A(n_2885),
.B(n_2191),
.Y(n_3429)
);

AOI21xp5_ASAP7_75t_L g3430 ( 
.A1(n_2546),
.A2(n_2573),
.B(n_2563),
.Y(n_3430)
);

AOI21xp5_ASAP7_75t_L g3431 ( 
.A1(n_2573),
.A2(n_2604),
.B(n_2588),
.Y(n_3431)
);

NOR2xp33_ASAP7_75t_L g3432 ( 
.A(n_2262),
.B(n_2265),
.Y(n_3432)
);

OAI22xp5_ASAP7_75t_L g3433 ( 
.A1(n_2634),
.A2(n_2756),
.B1(n_2924),
.B2(n_2873),
.Y(n_3433)
);

AOI21xp5_ASAP7_75t_L g3434 ( 
.A1(n_2588),
.A2(n_2614),
.B(n_2604),
.Y(n_3434)
);

AOI21xp5_ASAP7_75t_L g3435 ( 
.A1(n_2614),
.A2(n_2669),
.B(n_2666),
.Y(n_3435)
);

AOI21xp5_ASAP7_75t_L g3436 ( 
.A1(n_2666),
.A2(n_2674),
.B(n_2669),
.Y(n_3436)
);

INVx2_ASAP7_75t_SL g3437 ( 
.A(n_2422),
.Y(n_3437)
);

INVx2_ASAP7_75t_SL g3438 ( 
.A(n_2422),
.Y(n_3438)
);

A2O1A1Ixp33_ASAP7_75t_L g3439 ( 
.A1(n_2007),
.A2(n_2599),
.B(n_2561),
.C(n_2886),
.Y(n_3439)
);

OAI22xp5_ASAP7_75t_L g3440 ( 
.A1(n_2634),
.A2(n_2756),
.B1(n_2924),
.B2(n_2712),
.Y(n_3440)
);

AO21x1_ASAP7_75t_L g3441 ( 
.A1(n_2684),
.A2(n_2742),
.B(n_2731),
.Y(n_3441)
);

O2A1O1Ixp33_ASAP7_75t_L g3442 ( 
.A1(n_2049),
.A2(n_2641),
.B(n_2945),
.C(n_2324),
.Y(n_3442)
);

AOI21xp5_ASAP7_75t_L g3443 ( 
.A1(n_2684),
.A2(n_2742),
.B(n_2731),
.Y(n_3443)
);

AOI21xp5_ASAP7_75t_L g3444 ( 
.A1(n_2747),
.A2(n_2753),
.B(n_2752),
.Y(n_3444)
);

AOI21xp5_ASAP7_75t_L g3445 ( 
.A1(n_2747),
.A2(n_2753),
.B(n_2752),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_SL g3446 ( 
.A(n_2422),
.B(n_2462),
.Y(n_3446)
);

AOI22xp5_ASAP7_75t_L g3447 ( 
.A1(n_2634),
.A2(n_2873),
.B1(n_2712),
.B2(n_2756),
.Y(n_3447)
);

AOI21xp5_ASAP7_75t_L g3448 ( 
.A1(n_2764),
.A2(n_2781),
.B(n_2765),
.Y(n_3448)
);

OAI22xp5_ASAP7_75t_L g3449 ( 
.A1(n_2873),
.A2(n_2924),
.B1(n_2287),
.B2(n_2141),
.Y(n_3449)
);

AOI21xp5_ASAP7_75t_L g3450 ( 
.A1(n_2764),
.A2(n_2781),
.B(n_2765),
.Y(n_3450)
);

INVx2_ASAP7_75t_SL g3451 ( 
.A(n_2462),
.Y(n_3451)
);

AOI21xp5_ASAP7_75t_L g3452 ( 
.A1(n_2808),
.A2(n_2818),
.B(n_2815),
.Y(n_3452)
);

NOR3xp33_ASAP7_75t_L g3453 ( 
.A(n_2112),
.B(n_2067),
.C(n_2058),
.Y(n_3453)
);

OR2x2_ASAP7_75t_L g3454 ( 
.A(n_2815),
.B(n_2818),
.Y(n_3454)
);

INVx4_ASAP7_75t_L g3455 ( 
.A(n_2083),
.Y(n_3455)
);

NOR2xp67_ASAP7_75t_L g3456 ( 
.A(n_2836),
.B(n_2858),
.Y(n_3456)
);

AND2x2_ASAP7_75t_L g3457 ( 
.A(n_2910),
.B(n_2911),
.Y(n_3457)
);

AO21x1_ASAP7_75t_L g3458 ( 
.A1(n_2910),
.A2(n_2929),
.B(n_2911),
.Y(n_3458)
);

INVx1_ASAP7_75t_SL g3459 ( 
.A(n_2575),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_2254),
.B(n_2003),
.Y(n_3460)
);

AND2x2_ASAP7_75t_L g3461 ( 
.A(n_2269),
.B(n_2270),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_2003),
.Y(n_3462)
);

AND2x2_ASAP7_75t_L g3463 ( 
.A(n_2269),
.B(n_2270),
.Y(n_3463)
);

AOI21x1_ASAP7_75t_L g3464 ( 
.A1(n_2277),
.A2(n_2283),
.B(n_2282),
.Y(n_3464)
);

OAI21xp5_ASAP7_75t_L g3465 ( 
.A1(n_2148),
.A2(n_2163),
.B(n_2158),
.Y(n_3465)
);

OAI22xp5_ASAP7_75t_L g3466 ( 
.A1(n_2287),
.A2(n_2141),
.B1(n_2278),
.B2(n_2159),
.Y(n_3466)
);

OAI21xp5_ASAP7_75t_L g3467 ( 
.A1(n_2148),
.A2(n_2163),
.B(n_2158),
.Y(n_3467)
);

OAI21xp5_ASAP7_75t_L g3468 ( 
.A1(n_2206),
.A2(n_2303),
.B(n_2083),
.Y(n_3468)
);

INVx2_ASAP7_75t_L g3469 ( 
.A(n_2257),
.Y(n_3469)
);

AO21x1_ASAP7_75t_L g3470 ( 
.A1(n_2058),
.A2(n_2127),
.B(n_2067),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_2005),
.B(n_2010),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_2005),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_2010),
.Y(n_3473)
);

AOI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_2284),
.A2(n_2290),
.B(n_2289),
.Y(n_3474)
);

INVx2_ASAP7_75t_SL g3475 ( 
.A(n_2462),
.Y(n_3475)
);

AOI21x1_ASAP7_75t_L g3476 ( 
.A1(n_2292),
.A2(n_2295),
.B(n_2015),
.Y(n_3476)
);

AOI21xp5_ASAP7_75t_L g3477 ( 
.A1(n_2015),
.A2(n_2202),
.B(n_2216),
.Y(n_3477)
);

OAI21xp5_ASAP7_75t_L g3478 ( 
.A1(n_2206),
.A2(n_2303),
.B(n_2083),
.Y(n_3478)
);

O2A1O1Ixp33_ASAP7_75t_L g3479 ( 
.A1(n_2049),
.A2(n_2561),
.B(n_2846),
.C(n_2522),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_2027),
.Y(n_3480)
);

BUFx12f_ASAP7_75t_L g3481 ( 
.A(n_2291),
.Y(n_3481)
);

O2A1O1Ixp5_ASAP7_75t_L g3482 ( 
.A1(n_2067),
.A2(n_2903),
.B(n_2869),
.C(n_2127),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_2027),
.B(n_2033),
.Y(n_3483)
);

OAI21xp5_ASAP7_75t_L g3484 ( 
.A1(n_2083),
.A2(n_2837),
.B(n_2596),
.Y(n_3484)
);

AOI21xp5_ASAP7_75t_L g3485 ( 
.A1(n_2033),
.A2(n_2080),
.B(n_2152),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_2042),
.B(n_2044),
.Y(n_3486)
);

AOI21xp5_ASAP7_75t_L g3487 ( 
.A1(n_2042),
.A2(n_2165),
.B(n_2146),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_2044),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_2048),
.B(n_2053),
.Y(n_3489)
);

AOI21xp5_ASAP7_75t_L g3490 ( 
.A1(n_2048),
.A2(n_2202),
.B(n_2152),
.Y(n_3490)
);

AND2x2_ASAP7_75t_L g3491 ( 
.A(n_2053),
.B(n_2060),
.Y(n_3491)
);

AOI21xp33_ASAP7_75t_L g3492 ( 
.A1(n_2060),
.A2(n_2188),
.B(n_2224),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_2070),
.Y(n_3493)
);

BUFx2_ASAP7_75t_L g3494 ( 
.A(n_2575),
.Y(n_3494)
);

AOI21xp5_ASAP7_75t_L g3495 ( 
.A1(n_2070),
.A2(n_2224),
.B(n_2146),
.Y(n_3495)
);

INVx2_ASAP7_75t_L g3496 ( 
.A(n_2257),
.Y(n_3496)
);

O2A1O1Ixp33_ASAP7_75t_L g3497 ( 
.A1(n_2428),
.A2(n_2472),
.B(n_2489),
.C(n_2522),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_2080),
.B(n_2081),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_2263),
.Y(n_3499)
);

AOI22xp5_ASAP7_75t_L g3500 ( 
.A1(n_2159),
.A2(n_2596),
.B1(n_2837),
.B2(n_2177),
.Y(n_3500)
);

BUFx12f_ASAP7_75t_L g3501 ( 
.A(n_2203),
.Y(n_3501)
);

OAI321xp33_ASAP7_75t_L g3502 ( 
.A1(n_2428),
.A2(n_2859),
.A3(n_2886),
.B1(n_2599),
.B2(n_2658),
.C(n_2830),
.Y(n_3502)
);

O2A1O1Ixp5_ASAP7_75t_L g3503 ( 
.A1(n_2127),
.A2(n_2872),
.B(n_2559),
.C(n_2670),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_SL g3504 ( 
.A(n_2462),
.B(n_2618),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_2081),
.B(n_2085),
.Y(n_3505)
);

HB1xp67_ASAP7_75t_L g3506 ( 
.A(n_2462),
.Y(n_3506)
);

AOI22xp33_ASAP7_75t_L g3507 ( 
.A1(n_2108),
.A2(n_2198),
.B1(n_2188),
.B2(n_2196),
.Y(n_3507)
);

OAI21xp5_ASAP7_75t_L g3508 ( 
.A1(n_2596),
.A2(n_2837),
.B(n_2115),
.Y(n_3508)
);

AOI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_2085),
.A2(n_2216),
.B(n_2198),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_2089),
.B(n_2096),
.Y(n_3510)
);

O2A1O1Ixp33_ASAP7_75t_L g3511 ( 
.A1(n_2472),
.A2(n_2641),
.B(n_2489),
.C(n_2737),
.Y(n_3511)
);

NOR2xp33_ASAP7_75t_L g3512 ( 
.A(n_2019),
.B(n_2326),
.Y(n_3512)
);

AOI21xp5_ASAP7_75t_L g3513 ( 
.A1(n_2089),
.A2(n_2165),
.B(n_2196),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_2096),
.B(n_2263),
.Y(n_3514)
);

OAI22xp5_ASAP7_75t_L g3515 ( 
.A1(n_2287),
.A2(n_2141),
.B1(n_2278),
.B2(n_2390),
.Y(n_3515)
);

OAI21xp5_ASAP7_75t_L g3516 ( 
.A1(n_2596),
.A2(n_2837),
.B(n_2115),
.Y(n_3516)
);

A2O1A1Ixp33_ASAP7_75t_L g3517 ( 
.A1(n_2737),
.A2(n_2830),
.B(n_2859),
.C(n_2812),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_2296),
.Y(n_3518)
);

NOR2xp33_ASAP7_75t_L g3519 ( 
.A(n_2331),
.B(n_2347),
.Y(n_3519)
);

O2A1O1Ixp33_ASAP7_75t_L g3520 ( 
.A1(n_2760),
.A2(n_2812),
.B(n_2627),
.C(n_2362),
.Y(n_3520)
);

NOR3xp33_ASAP7_75t_L g3521 ( 
.A(n_2112),
.B(n_2367),
.C(n_2559),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_SL g3522 ( 
.A(n_2618),
.B(n_2660),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_2296),
.B(n_2596),
.Y(n_3523)
);

AOI21xp5_ASAP7_75t_L g3524 ( 
.A1(n_2618),
.A2(n_2660),
.B(n_2933),
.Y(n_3524)
);

OR2x6_ASAP7_75t_L g3525 ( 
.A(n_2108),
.B(n_2141),
.Y(n_3525)
);

INVx4_ASAP7_75t_L g3526 ( 
.A(n_2596),
.Y(n_3526)
);

NAND2x1p5_ASAP7_75t_L g3527 ( 
.A(n_2287),
.B(n_2933),
.Y(n_3527)
);

INVx11_ASAP7_75t_L g3528 ( 
.A(n_2104),
.Y(n_3528)
);

A2O1A1Ixp33_ASAP7_75t_L g3529 ( 
.A1(n_2760),
.A2(n_2116),
.B(n_2177),
.C(n_2278),
.Y(n_3529)
);

AOI21xp5_ASAP7_75t_L g3530 ( 
.A1(n_2618),
.A2(n_2660),
.B(n_2933),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_SL g3531 ( 
.A(n_2618),
.B(n_2660),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_SL g3532 ( 
.A(n_2660),
.B(n_2896),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_2065),
.Y(n_3533)
);

AND2x2_ASAP7_75t_L g3534 ( 
.A(n_2777),
.B(n_2896),
.Y(n_3534)
);

INVx3_ASAP7_75t_L g3535 ( 
.A(n_2278),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_2837),
.B(n_2217),
.Y(n_3536)
);

A2O1A1Ixp33_ASAP7_75t_L g3537 ( 
.A1(n_2116),
.A2(n_2278),
.B(n_2933),
.C(n_2896),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_L g3538 ( 
.A(n_2837),
.B(n_2208),
.Y(n_3538)
);

INVx2_ASAP7_75t_L g3539 ( 
.A(n_2777),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_2088),
.B(n_2138),
.Y(n_3540)
);

AOI21xp5_ASAP7_75t_L g3541 ( 
.A1(n_2777),
.A2(n_2933),
.B(n_2896),
.Y(n_3541)
);

OAI21xp33_ASAP7_75t_L g3542 ( 
.A1(n_2347),
.A2(n_2597),
.B(n_2922),
.Y(n_3542)
);

O2A1O1Ixp33_ASAP7_75t_SL g3543 ( 
.A1(n_1988),
.A2(n_2056),
.B(n_2252),
.C(n_2375),
.Y(n_3543)
);

AOI22xp5_ASAP7_75t_L g3544 ( 
.A1(n_2203),
.A2(n_2118),
.B1(n_2390),
.B2(n_2252),
.Y(n_3544)
);

OAI21xp5_ASAP7_75t_L g3545 ( 
.A1(n_2097),
.A2(n_2180),
.B(n_2098),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_2109),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_2777),
.B(n_2896),
.Y(n_3547)
);

O2A1O1Ixp33_ASAP7_75t_L g3548 ( 
.A1(n_2362),
.A2(n_2597),
.B(n_2627),
.C(n_2654),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_SL g3549 ( 
.A(n_2777),
.B(n_2559),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_2250),
.B(n_2288),
.Y(n_3550)
);

INVx2_ASAP7_75t_L g3551 ( 
.A(n_2696),
.Y(n_3551)
);

O2A1O1Ixp33_ASAP7_75t_L g3552 ( 
.A1(n_2654),
.A2(n_2709),
.B(n_2908),
.C(n_2922),
.Y(n_3552)
);

BUFx6f_ASAP7_75t_L g3553 ( 
.A(n_2149),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_2367),
.B(n_2872),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_SL g3555 ( 
.A(n_2367),
.B(n_2670),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_SL g3556 ( 
.A(n_2670),
.B(n_2869),
.Y(n_3556)
);

AND2x2_ASAP7_75t_L g3557 ( 
.A(n_2869),
.B(n_2872),
.Y(n_3557)
);

OAI21xp33_ASAP7_75t_L g3558 ( 
.A1(n_2709),
.A2(n_2908),
.B(n_2946),
.Y(n_3558)
);

OR2x6_ASAP7_75t_L g3559 ( 
.A(n_2252),
.B(n_2903),
.Y(n_3559)
);

AOI21x1_ASAP7_75t_L g3560 ( 
.A1(n_2696),
.A2(n_2903),
.B(n_2054),
.Y(n_3560)
);

INVx11_ASAP7_75t_L g3561 ( 
.A(n_2104),
.Y(n_3561)
);

AOI21xp5_ASAP7_75t_L g3562 ( 
.A1(n_2328),
.A2(n_2946),
.B(n_2358),
.Y(n_3562)
);

AND2x4_ASAP7_75t_L g3563 ( 
.A(n_2318),
.B(n_2103),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_2182),
.Y(n_3564)
);

AOI21xp5_ASAP7_75t_L g3565 ( 
.A1(n_2328),
.A2(n_2358),
.B(n_2252),
.Y(n_3565)
);

AOI22xp33_ASAP7_75t_L g3566 ( 
.A1(n_2318),
.A2(n_2103),
.B1(n_2580),
.B2(n_2443),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_2443),
.Y(n_3567)
);

AO21x1_ASAP7_75t_L g3568 ( 
.A1(n_2375),
.A2(n_2443),
.B(n_2461),
.Y(n_3568)
);

A2O1A1Ixp33_ASAP7_75t_L g3569 ( 
.A1(n_2443),
.A2(n_2461),
.B(n_2476),
.C(n_2511),
.Y(n_3569)
);

AOI21xp5_ASAP7_75t_L g3570 ( 
.A1(n_2926),
.A2(n_2461),
.B(n_2476),
.Y(n_3570)
);

AOI22xp5_ASAP7_75t_L g3571 ( 
.A1(n_2461),
.A2(n_2476),
.B1(n_2511),
.B2(n_2580),
.Y(n_3571)
);

BUFx6f_ASAP7_75t_L g3572 ( 
.A(n_2476),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_2511),
.B(n_2580),
.Y(n_3573)
);

AOI21xp5_ASAP7_75t_L g3574 ( 
.A1(n_2926),
.A2(n_2511),
.B(n_2580),
.Y(n_3574)
);

AOI21xp5_ASAP7_75t_L g3575 ( 
.A1(n_2926),
.A2(n_2746),
.B(n_2773),
.Y(n_3575)
);

A2O1A1Ixp33_ASAP7_75t_L g3576 ( 
.A1(n_2746),
.A2(n_2773),
.B(n_2816),
.C(n_2866),
.Y(n_3576)
);

O2A1O1Ixp33_ASAP7_75t_SL g3577 ( 
.A1(n_2746),
.A2(n_2773),
.B(n_2816),
.C(n_2866),
.Y(n_3577)
);

NOR2xp33_ASAP7_75t_L g3578 ( 
.A(n_2746),
.B(n_2773),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_SL g3579 ( 
.A(n_2816),
.B(n_2866),
.Y(n_3579)
);

AOI21xp5_ASAP7_75t_L g3580 ( 
.A1(n_2816),
.A2(n_2866),
.B(n_2926),
.Y(n_3580)
);

NOR2xp33_ASAP7_75t_L g3581 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_2319),
.Y(n_3582)
);

NOR2xp33_ASAP7_75t_L g3583 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3583)
);

HB1xp67_ASAP7_75t_L g3584 ( 
.A(n_1945),
.Y(n_3584)
);

OAI21xp5_ASAP7_75t_L g3585 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3585)
);

INVx3_ASAP7_75t_L g3586 ( 
.A(n_2349),
.Y(n_3586)
);

AOI21xp5_ASAP7_75t_L g3587 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3587)
);

OAI22xp5_ASAP7_75t_L g3588 ( 
.A1(n_2338),
.A2(n_2395),
.B1(n_2397),
.B2(n_2389),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_2319),
.Y(n_3589)
);

BUFx6f_ASAP7_75t_L g3590 ( 
.A(n_2037),
.Y(n_3590)
);

AOI21xp5_ASAP7_75t_L g3591 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3593)
);

O2A1O1Ixp33_ASAP7_75t_L g3594 ( 
.A1(n_1932),
.A2(n_2345),
.B(n_2609),
.C(n_2408),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3595)
);

AOI22xp33_ASAP7_75t_L g3596 ( 
.A1(n_2447),
.A2(n_1556),
.B1(n_1899),
.B2(n_2515),
.Y(n_3596)
);

O2A1O1Ixp33_ASAP7_75t_L g3597 ( 
.A1(n_1932),
.A2(n_2345),
.B(n_2609),
.C(n_2408),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_2319),
.Y(n_3598)
);

OAI21xp33_ASAP7_75t_L g3599 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3599)
);

INVxp67_ASAP7_75t_L g3600 ( 
.A(n_1995),
.Y(n_3600)
);

AOI21xp5_ASAP7_75t_L g3601 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_SL g3602 ( 
.A(n_2350),
.B(n_2360),
.Y(n_3602)
);

XOR2x2_ASAP7_75t_L g3603 ( 
.A(n_2471),
.B(n_2845),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3604)
);

AOI21xp5_ASAP7_75t_L g3605 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3605)
);

NOR2x1_ASAP7_75t_R g3606 ( 
.A(n_2084),
.B(n_649),
.Y(n_3606)
);

OR2x2_ASAP7_75t_L g3607 ( 
.A(n_2090),
.B(n_1944),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3608)
);

INVxp67_ASAP7_75t_L g3609 ( 
.A(n_1995),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_SL g3611 ( 
.A(n_2350),
.B(n_2360),
.Y(n_3611)
);

BUFx2_ASAP7_75t_L g3612 ( 
.A(n_2267),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3613)
);

HB1xp67_ASAP7_75t_L g3614 ( 
.A(n_1945),
.Y(n_3614)
);

AO22x1_ASAP7_75t_L g3615 ( 
.A1(n_2371),
.A2(n_1609),
.B1(n_1713),
.B2(n_2350),
.Y(n_3615)
);

AND2x4_ASAP7_75t_L g3616 ( 
.A(n_2267),
.B(n_2768),
.Y(n_3616)
);

AND2x2_ASAP7_75t_L g3617 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_L g3618 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_2319),
.Y(n_3619)
);

INVx2_ASAP7_75t_SL g3620 ( 
.A(n_2337),
.Y(n_3620)
);

A2O1A1Ixp33_ASAP7_75t_L g3621 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1588),
.C(n_1842),
.Y(n_3621)
);

AOI21xp5_ASAP7_75t_L g3622 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3622)
);

AOI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3623)
);

OR2x2_ASAP7_75t_L g3624 ( 
.A(n_2090),
.B(n_1944),
.Y(n_3624)
);

AOI21xp5_ASAP7_75t_L g3625 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3625)
);

HB1xp67_ASAP7_75t_L g3626 ( 
.A(n_1945),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3627)
);

AOI22xp5_ASAP7_75t_L g3628 ( 
.A1(n_1953),
.A2(n_1734),
.B1(n_1842),
.B2(n_1588),
.Y(n_3628)
);

AOI22xp5_ASAP7_75t_L g3629 ( 
.A1(n_1953),
.A2(n_1734),
.B1(n_1842),
.B2(n_1588),
.Y(n_3629)
);

AND2x2_ASAP7_75t_L g3630 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3630)
);

AOI21xp5_ASAP7_75t_L g3631 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3631)
);

AOI21xp5_ASAP7_75t_L g3632 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3633)
);

INVx2_ASAP7_75t_SL g3634 ( 
.A(n_2337),
.Y(n_3634)
);

AND2x2_ASAP7_75t_L g3635 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3635)
);

AO21x1_ASAP7_75t_L g3636 ( 
.A1(n_2464),
.A2(n_2761),
.B(n_2645),
.Y(n_3636)
);

OAI21xp5_ASAP7_75t_L g3637 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_L g3639 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3639)
);

OR2x2_ASAP7_75t_L g3640 ( 
.A(n_2090),
.B(n_1944),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_L g3641 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3641)
);

AOI21xp5_ASAP7_75t_L g3642 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3642)
);

INVx2_ASAP7_75t_SL g3643 ( 
.A(n_2337),
.Y(n_3643)
);

NOR2xp33_ASAP7_75t_L g3644 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3644)
);

HB1xp67_ASAP7_75t_L g3645 ( 
.A(n_1945),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3646)
);

BUFx3_ASAP7_75t_L g3647 ( 
.A(n_2602),
.Y(n_3647)
);

AND2x2_ASAP7_75t_L g3648 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3648)
);

AOI21xp5_ASAP7_75t_L g3649 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3649)
);

AND2x4_ASAP7_75t_L g3650 ( 
.A(n_2267),
.B(n_2768),
.Y(n_3650)
);

AOI21xp5_ASAP7_75t_L g3651 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3651)
);

O2A1O1Ixp33_ASAP7_75t_L g3652 ( 
.A1(n_1932),
.A2(n_2345),
.B(n_2609),
.C(n_2408),
.Y(n_3652)
);

OAI21x1_ASAP7_75t_L g3653 ( 
.A1(n_2349),
.A2(n_2919),
.B(n_2615),
.Y(n_3653)
);

AOI22xp33_ASAP7_75t_L g3654 ( 
.A1(n_2447),
.A2(n_1556),
.B1(n_1899),
.B2(n_2515),
.Y(n_3654)
);

AOI21xp5_ASAP7_75t_L g3655 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_2319),
.Y(n_3656)
);

BUFx6f_ASAP7_75t_L g3657 ( 
.A(n_2037),
.Y(n_3657)
);

INVx3_ASAP7_75t_L g3658 ( 
.A(n_2349),
.Y(n_3658)
);

BUFx6f_ASAP7_75t_L g3659 ( 
.A(n_2037),
.Y(n_3659)
);

AOI21xp5_ASAP7_75t_L g3660 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3660)
);

AOI21xp5_ASAP7_75t_L g3661 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3661)
);

A2O1A1Ixp33_ASAP7_75t_L g3662 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1588),
.C(n_1842),
.Y(n_3662)
);

AOI21xp5_ASAP7_75t_L g3663 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3663)
);

AOI22xp5_ASAP7_75t_L g3664 ( 
.A1(n_1953),
.A2(n_1734),
.B1(n_1842),
.B2(n_1588),
.Y(n_3664)
);

AOI21xp5_ASAP7_75t_L g3665 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3665)
);

AND2x2_ASAP7_75t_L g3666 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3666)
);

AOI21xp5_ASAP7_75t_L g3667 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3667)
);

O2A1O1Ixp5_ASAP7_75t_SL g3668 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2523),
.C(n_2360),
.Y(n_3668)
);

INVx2_ASAP7_75t_SL g3669 ( 
.A(n_2337),
.Y(n_3669)
);

HB1xp67_ASAP7_75t_L g3670 ( 
.A(n_1945),
.Y(n_3670)
);

OAI22xp5_ASAP7_75t_L g3671 ( 
.A1(n_2338),
.A2(n_2395),
.B1(n_2397),
.B2(n_2389),
.Y(n_3671)
);

AOI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3672)
);

OAI21xp5_ASAP7_75t_L g3673 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3673)
);

AOI21xp5_ASAP7_75t_L g3674 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3674)
);

AO21x1_ASAP7_75t_L g3675 ( 
.A1(n_2464),
.A2(n_2761),
.B(n_2645),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_SL g3676 ( 
.A(n_2350),
.B(n_2360),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_2319),
.Y(n_3677)
);

O2A1O1Ixp33_ASAP7_75t_SL g3678 ( 
.A1(n_2612),
.A2(n_1932),
.B(n_2408),
.C(n_2345),
.Y(n_3678)
);

INVxp67_ASAP7_75t_L g3679 ( 
.A(n_1995),
.Y(n_3679)
);

AOI33xp33_ASAP7_75t_L g3680 ( 
.A1(n_2338),
.A2(n_2427),
.A3(n_2395),
.B1(n_2432),
.B2(n_2397),
.B3(n_2389),
.Y(n_3680)
);

INVx2_ASAP7_75t_SL g3681 ( 
.A(n_2337),
.Y(n_3681)
);

AOI21xp5_ASAP7_75t_L g3682 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_2319),
.Y(n_3683)
);

BUFx3_ASAP7_75t_L g3684 ( 
.A(n_2602),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_L g3685 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_SL g3686 ( 
.A(n_2350),
.B(n_2360),
.Y(n_3686)
);

AOI21xp5_ASAP7_75t_L g3687 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3687)
);

OAI21xp5_ASAP7_75t_L g3688 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3688)
);

AOI21xp5_ASAP7_75t_L g3689 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3689)
);

INVx3_ASAP7_75t_L g3690 ( 
.A(n_2349),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_L g3691 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3692)
);

BUFx3_ASAP7_75t_L g3693 ( 
.A(n_2602),
.Y(n_3693)
);

BUFx4f_ASAP7_75t_L g3694 ( 
.A(n_2572),
.Y(n_3694)
);

AOI21x1_ASAP7_75t_L g3695 ( 
.A1(n_1996),
.A2(n_2842),
.B(n_2631),
.Y(n_3695)
);

O2A1O1Ixp5_ASAP7_75t_L g3696 ( 
.A1(n_1932),
.A2(n_2345),
.B(n_2609),
.C(n_2408),
.Y(n_3696)
);

OAI22xp5_ASAP7_75t_L g3697 ( 
.A1(n_2338),
.A2(n_2395),
.B1(n_2397),
.B2(n_2389),
.Y(n_3697)
);

AOI21xp5_ASAP7_75t_L g3698 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3698)
);

AOI21xp5_ASAP7_75t_L g3699 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3699)
);

INVx2_ASAP7_75t_SL g3700 ( 
.A(n_2337),
.Y(n_3700)
);

O2A1O1Ixp33_ASAP7_75t_L g3701 ( 
.A1(n_1932),
.A2(n_2345),
.B(n_2609),
.C(n_2408),
.Y(n_3701)
);

OAI21xp5_ASAP7_75t_L g3702 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3703)
);

OAI21xp5_ASAP7_75t_L g3704 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3704)
);

AOI21xp5_ASAP7_75t_L g3705 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3705)
);

AOI21xp5_ASAP7_75t_L g3706 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3706)
);

NOR2xp33_ASAP7_75t_L g3707 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3707)
);

BUFx6f_ASAP7_75t_L g3708 ( 
.A(n_2037),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_2319),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3712)
);

AOI21xp5_ASAP7_75t_L g3713 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3713)
);

AOI22xp5_ASAP7_75t_L g3714 ( 
.A1(n_1953),
.A2(n_1734),
.B1(n_1842),
.B2(n_1588),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3716)
);

AOI22xp5_ASAP7_75t_L g3717 ( 
.A1(n_1953),
.A2(n_1734),
.B1(n_1842),
.B2(n_1588),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3718)
);

OAI22xp5_ASAP7_75t_L g3719 ( 
.A1(n_2338),
.A2(n_2395),
.B1(n_2397),
.B2(n_2389),
.Y(n_3719)
);

AOI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3720)
);

AOI21xp5_ASAP7_75t_L g3721 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3721)
);

OAI21xp5_ASAP7_75t_L g3722 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3722)
);

NOR2xp33_ASAP7_75t_L g3723 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3723)
);

A2O1A1Ixp33_ASAP7_75t_L g3724 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1588),
.C(n_1842),
.Y(n_3724)
);

INVx3_ASAP7_75t_L g3725 ( 
.A(n_2349),
.Y(n_3725)
);

AOI21xp5_ASAP7_75t_L g3726 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3726)
);

AOI21xp5_ASAP7_75t_L g3727 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3727)
);

O2A1O1Ixp33_ASAP7_75t_SL g3728 ( 
.A1(n_2612),
.A2(n_1932),
.B(n_2408),
.C(n_2345),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3729)
);

AND2x4_ASAP7_75t_L g3730 ( 
.A(n_2267),
.B(n_2768),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_2319),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3733)
);

OAI21xp5_ASAP7_75t_L g3734 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3734)
);

NAND3xp33_ASAP7_75t_SL g3735 ( 
.A(n_2338),
.B(n_2395),
.C(n_2389),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_SL g3736 ( 
.A(n_2350),
.B(n_2360),
.Y(n_3736)
);

AOI21xp5_ASAP7_75t_L g3737 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_L g3738 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3738)
);

NOR2xp33_ASAP7_75t_L g3739 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3739)
);

AOI21xp5_ASAP7_75t_L g3740 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3740)
);

BUFx12f_ASAP7_75t_L g3741 ( 
.A(n_2814),
.Y(n_3741)
);

AOI21xp5_ASAP7_75t_L g3742 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3742)
);

OAI21xp5_ASAP7_75t_L g3743 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3743)
);

A2O1A1Ixp33_ASAP7_75t_L g3744 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1588),
.C(n_1842),
.Y(n_3744)
);

AOI21xp5_ASAP7_75t_L g3745 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3745)
);

BUFx8_ASAP7_75t_SL g3746 ( 
.A(n_2084),
.Y(n_3746)
);

BUFx6f_ASAP7_75t_L g3747 ( 
.A(n_2037),
.Y(n_3747)
);

AND2x2_ASAP7_75t_L g3748 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_2319),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_2319),
.Y(n_3750)
);

AO21x1_ASAP7_75t_L g3751 ( 
.A1(n_2464),
.A2(n_2761),
.B(n_2645),
.Y(n_3751)
);

AOI22xp5_ASAP7_75t_L g3752 ( 
.A1(n_1953),
.A2(n_1734),
.B1(n_1842),
.B2(n_1588),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_L g3753 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3753)
);

AOI21xp5_ASAP7_75t_L g3754 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3754)
);

INVx4_ASAP7_75t_L g3755 ( 
.A(n_2768),
.Y(n_3755)
);

O2A1O1Ixp33_ASAP7_75t_L g3756 ( 
.A1(n_1932),
.A2(n_2345),
.B(n_2609),
.C(n_2408),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_L g3757 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_2319),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3760)
);

NOR2xp33_ASAP7_75t_L g3761 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3761)
);

HB1xp67_ASAP7_75t_L g3762 ( 
.A(n_1945),
.Y(n_3762)
);

AOI21xp5_ASAP7_75t_L g3763 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_SL g3764 ( 
.A(n_2350),
.B(n_2360),
.Y(n_3764)
);

AND2x4_ASAP7_75t_L g3765 ( 
.A(n_2267),
.B(n_2768),
.Y(n_3765)
);

AOI21x1_ASAP7_75t_L g3766 ( 
.A1(n_1996),
.A2(n_2842),
.B(n_2631),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3767)
);

OAI21xp5_ASAP7_75t_L g3768 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3768)
);

NOR3xp33_ASAP7_75t_L g3769 ( 
.A(n_1932),
.B(n_2408),
.C(n_2345),
.Y(n_3769)
);

NOR2xp33_ASAP7_75t_L g3770 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3770)
);

OAI21xp5_ASAP7_75t_L g3771 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3771)
);

INVx3_ASAP7_75t_L g3772 ( 
.A(n_2349),
.Y(n_3772)
);

INVx3_ASAP7_75t_L g3773 ( 
.A(n_2349),
.Y(n_3773)
);

INVx4_ASAP7_75t_L g3774 ( 
.A(n_2768),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3776)
);

AOI21xp5_ASAP7_75t_L g3777 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3777)
);

BUFx2_ASAP7_75t_L g3778 ( 
.A(n_2267),
.Y(n_3778)
);

AOI22xp5_ASAP7_75t_L g3779 ( 
.A1(n_1953),
.A2(n_1734),
.B1(n_1842),
.B2(n_1588),
.Y(n_3779)
);

AOI22xp33_ASAP7_75t_L g3780 ( 
.A1(n_2447),
.A2(n_1556),
.B1(n_1899),
.B2(n_2515),
.Y(n_3780)
);

AOI21xp5_ASAP7_75t_L g3781 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3781)
);

A2O1A1Ixp33_ASAP7_75t_L g3782 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1588),
.C(n_1842),
.Y(n_3782)
);

AOI21xp5_ASAP7_75t_L g3783 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3783)
);

INVx2_ASAP7_75t_SL g3784 ( 
.A(n_2337),
.Y(n_3784)
);

AOI22xp5_ASAP7_75t_L g3785 ( 
.A1(n_1953),
.A2(n_1734),
.B1(n_1842),
.B2(n_1588),
.Y(n_3785)
);

AOI21x1_ASAP7_75t_L g3786 ( 
.A1(n_1996),
.A2(n_2842),
.B(n_2631),
.Y(n_3786)
);

AOI21xp5_ASAP7_75t_L g3787 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3787)
);

CKINVDCx5p33_ASAP7_75t_R g3788 ( 
.A(n_2084),
.Y(n_3788)
);

AOI21xp5_ASAP7_75t_L g3789 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_2319),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_2319),
.Y(n_3791)
);

NOR2xp67_ASAP7_75t_L g3792 ( 
.A(n_2029),
.B(n_1283),
.Y(n_3792)
);

AOI21xp5_ASAP7_75t_L g3793 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3793)
);

AO21x1_ASAP7_75t_L g3794 ( 
.A1(n_2464),
.A2(n_2761),
.B(n_2645),
.Y(n_3794)
);

NOR2xp67_ASAP7_75t_L g3795 ( 
.A(n_2029),
.B(n_1283),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_L g3796 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3796)
);

NOR2xp33_ASAP7_75t_L g3797 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3799)
);

O2A1O1Ixp33_ASAP7_75t_L g3800 ( 
.A1(n_1932),
.A2(n_2345),
.B(n_2609),
.C(n_2408),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_2319),
.Y(n_3801)
);

AOI21xp5_ASAP7_75t_L g3802 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3802)
);

OAI21xp33_ASAP7_75t_L g3803 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3803)
);

AOI21xp5_ASAP7_75t_L g3804 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3804)
);

AOI21xp5_ASAP7_75t_L g3805 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3805)
);

NOR3xp33_ASAP7_75t_L g3806 ( 
.A(n_1932),
.B(n_2408),
.C(n_2345),
.Y(n_3806)
);

AOI22xp5_ASAP7_75t_L g3807 ( 
.A1(n_1953),
.A2(n_1734),
.B1(n_1842),
.B2(n_1588),
.Y(n_3807)
);

CKINVDCx10_ASAP7_75t_R g3808 ( 
.A(n_2637),
.Y(n_3808)
);

CKINVDCx8_ASAP7_75t_R g3809 ( 
.A(n_2274),
.Y(n_3809)
);

NAND2x1p5_ASAP7_75t_L g3810 ( 
.A(n_2238),
.B(n_1260),
.Y(n_3810)
);

AOI21xp5_ASAP7_75t_L g3811 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3811)
);

AOI21xp5_ASAP7_75t_L g3812 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3812)
);

INVx11_ASAP7_75t_L g3813 ( 
.A(n_2084),
.Y(n_3813)
);

INVxp67_ASAP7_75t_L g3814 ( 
.A(n_1995),
.Y(n_3814)
);

AOI21xp5_ASAP7_75t_L g3815 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3815)
);

AOI21x1_ASAP7_75t_L g3816 ( 
.A1(n_1996),
.A2(n_2842),
.B(n_2631),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3817)
);

AND2x4_ASAP7_75t_L g3818 ( 
.A(n_2267),
.B(n_2768),
.Y(n_3818)
);

INVx5_ASAP7_75t_L g3819 ( 
.A(n_2768),
.Y(n_3819)
);

A2O1A1Ixp33_ASAP7_75t_L g3820 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1588),
.C(n_1842),
.Y(n_3820)
);

A2O1A1Ixp33_ASAP7_75t_L g3821 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1588),
.C(n_1842),
.Y(n_3821)
);

AOI22xp5_ASAP7_75t_L g3822 ( 
.A1(n_1953),
.A2(n_1734),
.B1(n_1842),
.B2(n_1588),
.Y(n_3822)
);

OAI22xp5_ASAP7_75t_L g3823 ( 
.A1(n_2338),
.A2(n_2395),
.B1(n_2397),
.B2(n_2389),
.Y(n_3823)
);

OAI21xp5_ASAP7_75t_L g3824 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3825)
);

BUFx6f_ASAP7_75t_L g3826 ( 
.A(n_2037),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3827)
);

AOI21xp5_ASAP7_75t_L g3828 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3828)
);

OAI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3829)
);

NOR2xp33_ASAP7_75t_L g3830 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3830)
);

AOI21xp5_ASAP7_75t_L g3831 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3831)
);

OAI21xp5_ASAP7_75t_L g3832 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3832)
);

NOR2xp33_ASAP7_75t_SL g3833 ( 
.A(n_2556),
.B(n_2782),
.Y(n_3833)
);

AOI21xp5_ASAP7_75t_L g3834 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3834)
);

NOR2xp33_ASAP7_75t_L g3835 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3835)
);

AOI21xp33_ASAP7_75t_L g3836 ( 
.A1(n_1948),
.A2(n_1744),
.B(n_2430),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3837)
);

AOI21xp5_ASAP7_75t_L g3838 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3838)
);

BUFx2_ASAP7_75t_L g3839 ( 
.A(n_2267),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_2319),
.Y(n_3840)
);

AOI21xp5_ASAP7_75t_L g3841 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3841)
);

INVx1_ASAP7_75t_L g3842 ( 
.A(n_2319),
.Y(n_3842)
);

AOI21xp5_ASAP7_75t_L g3843 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_SL g3844 ( 
.A(n_2350),
.B(n_2360),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_2319),
.Y(n_3845)
);

BUFx2_ASAP7_75t_L g3846 ( 
.A(n_2267),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3847)
);

BUFx12f_ASAP7_75t_L g3848 ( 
.A(n_2814),
.Y(n_3848)
);

O2A1O1Ixp33_ASAP7_75t_L g3849 ( 
.A1(n_1932),
.A2(n_2345),
.B(n_2609),
.C(n_2408),
.Y(n_3849)
);

BUFx6f_ASAP7_75t_L g3850 ( 
.A(n_2037),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_SL g3851 ( 
.A(n_2350),
.B(n_2360),
.Y(n_3851)
);

OAI21xp5_ASAP7_75t_L g3852 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3852)
);

NAND2x1p5_ASAP7_75t_L g3853 ( 
.A(n_2238),
.B(n_1260),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_L g3854 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3854)
);

A2O1A1Ixp33_ASAP7_75t_L g3855 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1588),
.C(n_1842),
.Y(n_3855)
);

INVxp67_ASAP7_75t_L g3856 ( 
.A(n_1995),
.Y(n_3856)
);

OAI21xp5_ASAP7_75t_L g3857 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3857)
);

AOI21xp5_ASAP7_75t_L g3858 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3858)
);

BUFx6f_ASAP7_75t_L g3859 ( 
.A(n_2037),
.Y(n_3859)
);

AOI21xp5_ASAP7_75t_L g3860 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3860)
);

AOI21xp5_ASAP7_75t_L g3861 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3862)
);

OAI21xp5_ASAP7_75t_L g3863 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3864)
);

NOR2xp33_ASAP7_75t_L g3865 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3866)
);

INVx4_ASAP7_75t_L g3867 ( 
.A(n_2768),
.Y(n_3867)
);

O2A1O1Ixp33_ASAP7_75t_L g3868 ( 
.A1(n_1932),
.A2(n_2345),
.B(n_2609),
.C(n_2408),
.Y(n_3868)
);

OR2x2_ASAP7_75t_L g3869 ( 
.A(n_2090),
.B(n_1944),
.Y(n_3869)
);

INVx3_ASAP7_75t_L g3870 ( 
.A(n_2349),
.Y(n_3870)
);

NOR2xp33_ASAP7_75t_L g3871 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3871)
);

HB1xp67_ASAP7_75t_L g3872 ( 
.A(n_1945),
.Y(n_3872)
);

AND2x2_ASAP7_75t_L g3873 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3873)
);

OAI21xp5_ASAP7_75t_L g3874 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3874)
);

NOR2xp67_ASAP7_75t_L g3875 ( 
.A(n_2029),
.B(n_1283),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_SL g3876 ( 
.A(n_2350),
.B(n_2360),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_2319),
.Y(n_3878)
);

BUFx3_ASAP7_75t_L g3879 ( 
.A(n_2602),
.Y(n_3879)
);

AOI21xp5_ASAP7_75t_L g3880 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_2319),
.Y(n_3881)
);

NOR2xp33_ASAP7_75t_SL g3882 ( 
.A(n_2556),
.B(n_2782),
.Y(n_3882)
);

AOI21xp5_ASAP7_75t_L g3883 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3883)
);

INVx3_ASAP7_75t_L g3884 ( 
.A(n_2349),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_SL g3885 ( 
.A(n_2350),
.B(n_2360),
.Y(n_3885)
);

OAI22xp5_ASAP7_75t_L g3886 ( 
.A1(n_2338),
.A2(n_2395),
.B1(n_2397),
.B2(n_2389),
.Y(n_3886)
);

AOI21xp5_ASAP7_75t_L g3887 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3887)
);

AOI21xp5_ASAP7_75t_L g3888 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_L g3889 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3889)
);

AOI21xp5_ASAP7_75t_L g3890 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3890)
);

AOI21xp5_ASAP7_75t_L g3891 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3891)
);

NOR2xp33_ASAP7_75t_L g3892 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3892)
);

AOI21xp5_ASAP7_75t_L g3893 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3893)
);

AOI21xp33_ASAP7_75t_L g3894 ( 
.A1(n_1948),
.A2(n_1744),
.B(n_2430),
.Y(n_3894)
);

AOI21xp5_ASAP7_75t_L g3895 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_SL g3896 ( 
.A(n_2350),
.B(n_2360),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_2319),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3898)
);

HB1xp67_ASAP7_75t_L g3899 ( 
.A(n_1945),
.Y(n_3899)
);

NOR2xp33_ASAP7_75t_L g3900 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3900)
);

OAI22xp5_ASAP7_75t_L g3901 ( 
.A1(n_2338),
.A2(n_2395),
.B1(n_2397),
.B2(n_2389),
.Y(n_3901)
);

INVx4_ASAP7_75t_L g3902 ( 
.A(n_2768),
.Y(n_3902)
);

AOI21xp5_ASAP7_75t_L g3903 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3903)
);

AO21x1_ASAP7_75t_L g3904 ( 
.A1(n_2464),
.A2(n_2761),
.B(n_2645),
.Y(n_3904)
);

BUFx6f_ASAP7_75t_L g3905 ( 
.A(n_2037),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_SL g3908 ( 
.A(n_2350),
.B(n_2360),
.Y(n_3908)
);

BUFx4f_ASAP7_75t_L g3909 ( 
.A(n_2572),
.Y(n_3909)
);

AND2x2_ASAP7_75t_L g3910 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3910)
);

AND2x4_ASAP7_75t_L g3911 ( 
.A(n_2267),
.B(n_2768),
.Y(n_3911)
);

BUFx6f_ASAP7_75t_L g3912 ( 
.A(n_2037),
.Y(n_3912)
);

INVx4_ASAP7_75t_L g3913 ( 
.A(n_2768),
.Y(n_3913)
);

AOI21xp5_ASAP7_75t_L g3914 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3914)
);

AOI21xp5_ASAP7_75t_L g3915 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3915)
);

A2O1A1Ixp33_ASAP7_75t_L g3916 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1588),
.C(n_1842),
.Y(n_3916)
);

AOI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3917)
);

AOI21xp5_ASAP7_75t_L g3918 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3918)
);

HB1xp67_ASAP7_75t_L g3919 ( 
.A(n_1945),
.Y(n_3919)
);

NOR2xp33_ASAP7_75t_L g3920 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3920)
);

OAI321xp33_ASAP7_75t_L g3921 ( 
.A1(n_2350),
.A2(n_1744),
.A3(n_2499),
.B1(n_2534),
.B2(n_2523),
.C(n_2360),
.Y(n_3921)
);

NOR2xp33_ASAP7_75t_L g3922 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3922)
);

AOI21xp5_ASAP7_75t_L g3923 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3923)
);

OAI21xp5_ASAP7_75t_L g3924 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3924)
);

HB1xp67_ASAP7_75t_L g3925 ( 
.A(n_1945),
.Y(n_3925)
);

BUFx2_ASAP7_75t_SL g3926 ( 
.A(n_2396),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_L g3927 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3927)
);

BUFx12f_ASAP7_75t_L g3928 ( 
.A(n_2814),
.Y(n_3928)
);

OR2x2_ASAP7_75t_L g3929 ( 
.A(n_2090),
.B(n_1944),
.Y(n_3929)
);

NOR2x1_ASAP7_75t_L g3930 ( 
.A(n_2396),
.B(n_1283),
.Y(n_3930)
);

NOR2xp33_ASAP7_75t_L g3931 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3931)
);

BUFx4f_ASAP7_75t_L g3932 ( 
.A(n_2572),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3933)
);

AOI21xp5_ASAP7_75t_L g3934 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3934)
);

AOI21xp5_ASAP7_75t_L g3935 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3935)
);

A2O1A1Ixp33_ASAP7_75t_L g3936 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1588),
.C(n_1842),
.Y(n_3936)
);

AOI21xp5_ASAP7_75t_L g3937 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3937)
);

AO22x1_ASAP7_75t_L g3938 ( 
.A1(n_2371),
.A2(n_1609),
.B1(n_1713),
.B2(n_2350),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_L g3939 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3939)
);

NOR2xp67_ASAP7_75t_SL g3940 ( 
.A(n_2350),
.B(n_1744),
.Y(n_3940)
);

O2A1O1Ixp33_ASAP7_75t_L g3941 ( 
.A1(n_1932),
.A2(n_2345),
.B(n_2609),
.C(n_2408),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3942)
);

AOI21xp5_ASAP7_75t_L g3943 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3943)
);

AOI21xp5_ASAP7_75t_L g3944 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_L g3945 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_2319),
.Y(n_3946)
);

INVx3_ASAP7_75t_L g3947 ( 
.A(n_2349),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3950)
);

AND2x2_ASAP7_75t_L g3951 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3951)
);

AOI21xp5_ASAP7_75t_L g3952 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_SL g3953 ( 
.A(n_2350),
.B(n_2360),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_L g3954 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3954)
);

AOI22xp33_ASAP7_75t_L g3955 ( 
.A1(n_2447),
.A2(n_1556),
.B1(n_1899),
.B2(n_2515),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3956)
);

HB1xp67_ASAP7_75t_L g3957 ( 
.A(n_1945),
.Y(n_3957)
);

OAI21xp5_ASAP7_75t_L g3958 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3958)
);

AOI21xp5_ASAP7_75t_L g3959 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3959)
);

AOI21x1_ASAP7_75t_L g3960 ( 
.A1(n_1996),
.A2(n_2842),
.B(n_2631),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3962)
);

NOR2xp33_ASAP7_75t_L g3963 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3963)
);

AOI21xp5_ASAP7_75t_L g3964 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3965)
);

NOR2xp33_ASAP7_75t_L g3966 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3966)
);

NOR2xp33_ASAP7_75t_L g3967 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_L g3968 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3968)
);

BUFx8_ASAP7_75t_L g3969 ( 
.A(n_2084),
.Y(n_3969)
);

AOI21xp5_ASAP7_75t_L g3970 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_L g3971 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_2319),
.Y(n_3972)
);

INVx3_ASAP7_75t_L g3973 ( 
.A(n_2349),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3974)
);

O2A1O1Ixp33_ASAP7_75t_L g3975 ( 
.A1(n_1932),
.A2(n_2345),
.B(n_2609),
.C(n_2408),
.Y(n_3975)
);

AOI21xp5_ASAP7_75t_L g3976 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3976)
);

AOI22xp5_ASAP7_75t_L g3977 ( 
.A1(n_1953),
.A2(n_1734),
.B1(n_1842),
.B2(n_1588),
.Y(n_3977)
);

INVx2_ASAP7_75t_SL g3978 ( 
.A(n_2337),
.Y(n_3978)
);

OAI22xp5_ASAP7_75t_L g3979 ( 
.A1(n_2338),
.A2(n_2395),
.B1(n_2397),
.B2(n_2389),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3980)
);

BUFx3_ASAP7_75t_L g3981 ( 
.A(n_2602),
.Y(n_3981)
);

AOI21x1_ASAP7_75t_L g3982 ( 
.A1(n_1996),
.A2(n_2842),
.B(n_2631),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3983)
);

AOI33xp33_ASAP7_75t_L g3984 ( 
.A1(n_2338),
.A2(n_2427),
.A3(n_2395),
.B1(n_2432),
.B2(n_2397),
.B3(n_2389),
.Y(n_3984)
);

NOR2xp33_ASAP7_75t_L g3985 ( 
.A(n_1932),
.B(n_2345),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3986)
);

OAI22xp5_ASAP7_75t_L g3987 ( 
.A1(n_2338),
.A2(n_2395),
.B1(n_2397),
.B2(n_2389),
.Y(n_3987)
);

OAI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_3988)
);

O2A1O1Ixp33_ASAP7_75t_L g3989 ( 
.A1(n_1932),
.A2(n_2345),
.B(n_2609),
.C(n_2408),
.Y(n_3989)
);

HB1xp67_ASAP7_75t_L g3990 ( 
.A(n_1945),
.Y(n_3990)
);

AOI21xp5_ASAP7_75t_L g3991 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3991)
);

OR2x6_ASAP7_75t_L g3992 ( 
.A(n_2631),
.B(n_2842),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_2319),
.Y(n_3993)
);

AOI21xp5_ASAP7_75t_L g3994 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3995)
);

O2A1O1Ixp33_ASAP7_75t_SL g3996 ( 
.A1(n_2612),
.A2(n_1932),
.B(n_2408),
.C(n_2345),
.Y(n_3996)
);

A2O1A1Ixp33_ASAP7_75t_L g3997 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1588),
.C(n_1842),
.Y(n_3997)
);

BUFx8_ASAP7_75t_SL g3998 ( 
.A(n_2084),
.Y(n_3998)
);

AND2x2_ASAP7_75t_L g3999 ( 
.A(n_1944),
.B(n_2327),
.Y(n_3999)
);

INVx4_ASAP7_75t_L g4000 ( 
.A(n_2768),
.Y(n_4000)
);

AO21x1_ASAP7_75t_L g4001 ( 
.A1(n_2464),
.A2(n_2761),
.B(n_2645),
.Y(n_4001)
);

NOR2xp33_ASAP7_75t_L g4002 ( 
.A(n_1932),
.B(n_2345),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_SL g4003 ( 
.A(n_2350),
.B(n_2360),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_SL g4004 ( 
.A(n_2350),
.B(n_2360),
.Y(n_4004)
);

AND2x4_ASAP7_75t_L g4005 ( 
.A(n_2267),
.B(n_2768),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_L g4006 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_L g4007 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4007)
);

AOI21xp5_ASAP7_75t_L g4008 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4008)
);

NOR3xp33_ASAP7_75t_L g4009 ( 
.A(n_1932),
.B(n_2408),
.C(n_2345),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_2319),
.Y(n_4010)
);

BUFx3_ASAP7_75t_L g4011 ( 
.A(n_2602),
.Y(n_4011)
);

NOR2xp33_ASAP7_75t_L g4012 ( 
.A(n_1932),
.B(n_2345),
.Y(n_4012)
);

NOR2xp33_ASAP7_75t_L g4013 ( 
.A(n_1932),
.B(n_2345),
.Y(n_4013)
);

OAI22xp5_ASAP7_75t_L g4014 ( 
.A1(n_2338),
.A2(n_2395),
.B1(n_2397),
.B2(n_2389),
.Y(n_4014)
);

AOI21x1_ASAP7_75t_L g4015 ( 
.A1(n_1996),
.A2(n_2842),
.B(n_2631),
.Y(n_4015)
);

BUFx3_ASAP7_75t_L g4016 ( 
.A(n_2602),
.Y(n_4016)
);

INVx3_ASAP7_75t_L g4017 ( 
.A(n_2349),
.Y(n_4017)
);

A2O1A1Ixp33_ASAP7_75t_L g4018 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1588),
.C(n_1842),
.Y(n_4018)
);

A2O1A1Ixp33_ASAP7_75t_L g4019 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1588),
.C(n_1842),
.Y(n_4019)
);

BUFx6f_ASAP7_75t_L g4020 ( 
.A(n_2037),
.Y(n_4020)
);

A2O1A1Ixp33_ASAP7_75t_L g4021 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1588),
.C(n_1842),
.Y(n_4021)
);

AOI21xp5_ASAP7_75t_L g4022 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4022)
);

AOI21xp5_ASAP7_75t_L g4023 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4024)
);

INVx1_ASAP7_75t_SL g4025 ( 
.A(n_2602),
.Y(n_4025)
);

NAND2xp33_ASAP7_75t_L g4026 ( 
.A(n_2529),
.B(n_2663),
.Y(n_4026)
);

AND2x4_ASAP7_75t_L g4027 ( 
.A(n_2267),
.B(n_2768),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_2319),
.Y(n_4028)
);

AOI33xp33_ASAP7_75t_L g4029 ( 
.A1(n_2338),
.A2(n_2427),
.A3(n_2395),
.B1(n_2432),
.B2(n_2397),
.B3(n_2389),
.Y(n_4029)
);

NOR2x1_ASAP7_75t_L g4030 ( 
.A(n_2396),
.B(n_1283),
.Y(n_4030)
);

INVxp67_ASAP7_75t_L g4031 ( 
.A(n_1995),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4032)
);

NOR2xp33_ASAP7_75t_L g4033 ( 
.A(n_1932),
.B(n_2345),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4034)
);

AOI21xp5_ASAP7_75t_L g4035 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4035)
);

INVx2_ASAP7_75t_L g4036 ( 
.A(n_2947),
.Y(n_4036)
);

AND2x4_ASAP7_75t_L g4037 ( 
.A(n_2267),
.B(n_2768),
.Y(n_4037)
);

INVx2_ASAP7_75t_L g4038 ( 
.A(n_2947),
.Y(n_4038)
);

OAI321xp33_ASAP7_75t_L g4039 ( 
.A1(n_2350),
.A2(n_1744),
.A3(n_2499),
.B1(n_2534),
.B2(n_2523),
.C(n_2360),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4040)
);

INVxp67_ASAP7_75t_SL g4041 ( 
.A(n_2114),
.Y(n_4041)
);

INVx2_ASAP7_75t_L g4042 ( 
.A(n_2947),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4043)
);

INVx2_ASAP7_75t_L g4044 ( 
.A(n_2947),
.Y(n_4044)
);

A2O1A1Ixp33_ASAP7_75t_L g4045 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1588),
.C(n_1842),
.Y(n_4045)
);

INVx2_ASAP7_75t_L g4046 ( 
.A(n_2947),
.Y(n_4046)
);

AOI22xp33_ASAP7_75t_L g4047 ( 
.A1(n_2447),
.A2(n_1556),
.B1(n_1899),
.B2(n_2515),
.Y(n_4047)
);

OAI21xp5_ASAP7_75t_L g4048 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_4048)
);

HB1xp67_ASAP7_75t_L g4049 ( 
.A(n_1945),
.Y(n_4049)
);

AOI21xp5_ASAP7_75t_L g4050 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_L g4051 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4051)
);

AND2x6_ASAP7_75t_SL g4052 ( 
.A(n_1935),
.B(n_1942),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_2319),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_2319),
.Y(n_4054)
);

AOI21xp5_ASAP7_75t_L g4055 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4055)
);

AOI21xp5_ASAP7_75t_L g4056 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_L g4058 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_SL g4059 ( 
.A(n_2350),
.B(n_2360),
.Y(n_4059)
);

A2O1A1Ixp33_ASAP7_75t_L g4060 ( 
.A1(n_2652),
.A2(n_2934),
.B(n_1588),
.C(n_1842),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_2947),
.Y(n_4061)
);

CKINVDCx10_ASAP7_75t_R g4062 ( 
.A(n_2637),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_2319),
.Y(n_4063)
);

INVx2_ASAP7_75t_L g4064 ( 
.A(n_2947),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_2947),
.Y(n_4065)
);

INVx2_ASAP7_75t_L g4066 ( 
.A(n_2947),
.Y(n_4066)
);

NOR2xp67_ASAP7_75t_L g4067 ( 
.A(n_2029),
.B(n_1283),
.Y(n_4067)
);

INVx2_ASAP7_75t_L g4068 ( 
.A(n_2947),
.Y(n_4068)
);

O2A1O1Ixp5_ASAP7_75t_L g4069 ( 
.A1(n_1932),
.A2(n_2345),
.B(n_2609),
.C(n_2408),
.Y(n_4069)
);

INVx2_ASAP7_75t_L g4070 ( 
.A(n_2947),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_SL g4071 ( 
.A(n_2350),
.B(n_2360),
.Y(n_4071)
);

AOI21xp5_ASAP7_75t_L g4072 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4072)
);

AOI21xp5_ASAP7_75t_L g4073 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4073)
);

BUFx6f_ASAP7_75t_L g4074 ( 
.A(n_2037),
.Y(n_4074)
);

OAI21xp5_ASAP7_75t_L g4075 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_4075)
);

AOI21xp5_ASAP7_75t_L g4076 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4076)
);

BUFx10_ASAP7_75t_L g4077 ( 
.A(n_2274),
.Y(n_4077)
);

AOI21xp5_ASAP7_75t_L g4078 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4078)
);

NOR2xp33_ASAP7_75t_L g4079 ( 
.A(n_1932),
.B(n_2345),
.Y(n_4079)
);

AOI21xp5_ASAP7_75t_L g4080 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4080)
);

AOI21xp5_ASAP7_75t_L g4081 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4081)
);

AOI21xp5_ASAP7_75t_L g4082 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_L g4083 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4083)
);

AOI21xp5_ASAP7_75t_L g4084 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4084)
);

AOI21xp5_ASAP7_75t_L g4085 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4085)
);

AOI21xp5_ASAP7_75t_L g4086 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4086)
);

BUFx6f_ASAP7_75t_L g4087 ( 
.A(n_2037),
.Y(n_4087)
);

AND2x2_ASAP7_75t_L g4088 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4088)
);

INVx2_ASAP7_75t_L g4089 ( 
.A(n_2947),
.Y(n_4089)
);

AOI21x1_ASAP7_75t_L g4090 ( 
.A1(n_1996),
.A2(n_2842),
.B(n_2631),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_SL g4092 ( 
.A(n_2350),
.B(n_2360),
.Y(n_4092)
);

AOI21xp5_ASAP7_75t_L g4093 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4094)
);

NOR2xp33_ASAP7_75t_L g4095 ( 
.A(n_1932),
.B(n_2345),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_L g4096 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_2319),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4100)
);

BUFx3_ASAP7_75t_L g4101 ( 
.A(n_2602),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_2319),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_L g4103 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4103)
);

OAI21xp5_ASAP7_75t_L g4104 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_4104)
);

NOR3xp33_ASAP7_75t_L g4105 ( 
.A(n_1932),
.B(n_2408),
.C(n_2345),
.Y(n_4105)
);

AOI21xp5_ASAP7_75t_L g4106 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4106)
);

NOR2xp67_ASAP7_75t_L g4107 ( 
.A(n_2029),
.B(n_1283),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_SL g4108 ( 
.A(n_2350),
.B(n_2360),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4109)
);

AOI21xp5_ASAP7_75t_L g4110 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4110)
);

INVx4_ASAP7_75t_L g4111 ( 
.A(n_2768),
.Y(n_4111)
);

AOI21xp5_ASAP7_75t_L g4112 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4112)
);

OAI21xp5_ASAP7_75t_L g4113 ( 
.A1(n_2350),
.A2(n_2499),
.B(n_2360),
.Y(n_4113)
);

AOI21x1_ASAP7_75t_L g4114 ( 
.A1(n_1996),
.A2(n_2842),
.B(n_2631),
.Y(n_4114)
);

AOI21xp5_ASAP7_75t_L g4115 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_SL g4116 ( 
.A(n_2350),
.B(n_2360),
.Y(n_4116)
);

AOI21xp5_ASAP7_75t_L g4117 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4117)
);

AOI21xp5_ASAP7_75t_L g4118 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_SL g4119 ( 
.A(n_2350),
.B(n_2360),
.Y(n_4119)
);

AOI21xp5_ASAP7_75t_L g4120 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_2319),
.Y(n_4121)
);

AOI21xp5_ASAP7_75t_L g4122 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_L g4123 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4123)
);

AND2x2_ASAP7_75t_L g4124 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4124)
);

AO21x2_ASAP7_75t_L g4125 ( 
.A1(n_2064),
.A2(n_1744),
.B(n_1026),
.Y(n_4125)
);

O2A1O1Ixp33_ASAP7_75t_L g4126 ( 
.A1(n_1932),
.A2(n_2345),
.B(n_2609),
.C(n_2408),
.Y(n_4126)
);

AOI21xp5_ASAP7_75t_L g4127 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_L g4128 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_L g4129 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4129)
);

NAND2xp5_ASAP7_75t_SL g4130 ( 
.A(n_2350),
.B(n_2360),
.Y(n_4130)
);

O2A1O1Ixp33_ASAP7_75t_SL g4131 ( 
.A1(n_2612),
.A2(n_1932),
.B(n_2408),
.C(n_2345),
.Y(n_4131)
);

NOR2xp33_ASAP7_75t_L g4132 ( 
.A(n_1932),
.B(n_2345),
.Y(n_4132)
);

INVx1_ASAP7_75t_SL g4133 ( 
.A(n_2602),
.Y(n_4133)
);

O2A1O1Ixp33_ASAP7_75t_L g4134 ( 
.A1(n_1932),
.A2(n_2345),
.B(n_2609),
.C(n_2408),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_SL g4135 ( 
.A(n_2350),
.B(n_2360),
.Y(n_4135)
);

AOI21xp5_ASAP7_75t_L g4136 ( 
.A1(n_2350),
.A2(n_1744),
.B(n_2360),
.Y(n_4136)
);

OAI22xp5_ASAP7_75t_L g4137 ( 
.A1(n_2338),
.A2(n_2395),
.B1(n_2397),
.B2(n_2389),
.Y(n_4137)
);

AOI22x1_ASAP7_75t_L g4138 ( 
.A1(n_2350),
.A2(n_2360),
.B1(n_2523),
.B2(n_2499),
.Y(n_4138)
);

BUFx2_ASAP7_75t_L g4139 ( 
.A(n_2267),
.Y(n_4139)
);

OAI22xp5_ASAP7_75t_L g4140 ( 
.A1(n_2338),
.A2(n_2395),
.B1(n_2397),
.B2(n_2389),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_L g4141 ( 
.A(n_1944),
.B(n_2327),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_3013),
.B(n_3019),
.Y(n_4142)
);

INVx2_ASAP7_75t_SL g4143 ( 
.A(n_2995),
.Y(n_4143)
);

INVx4_ASAP7_75t_L g4144 ( 
.A(n_3392),
.Y(n_4144)
);

INVx3_ASAP7_75t_L g4145 ( 
.A(n_2961),
.Y(n_4145)
);

NAND2xp5_ASAP7_75t_L g4146 ( 
.A(n_3013),
.B(n_3019),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_L g4147 ( 
.A(n_3057),
.B(n_3061),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_SL g4148 ( 
.A(n_2965),
.B(n_3636),
.Y(n_4148)
);

A2O1A1Ixp33_ASAP7_75t_L g4149 ( 
.A1(n_3034),
.A2(n_2983),
.B(n_2972),
.C(n_3833),
.Y(n_4149)
);

AND2x2_ASAP7_75t_L g4150 ( 
.A(n_3249),
.B(n_3282),
.Y(n_4150)
);

BUFx2_ASAP7_75t_L g4151 ( 
.A(n_3612),
.Y(n_4151)
);

BUFx6f_ASAP7_75t_L g4152 ( 
.A(n_3653),
.Y(n_4152)
);

CKINVDCx5p33_ASAP7_75t_R g4153 ( 
.A(n_3113),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_3239),
.Y(n_4154)
);

OA22x2_ASAP7_75t_L g4155 ( 
.A1(n_3628),
.A2(n_3629),
.B1(n_3714),
.B2(n_3664),
.Y(n_4155)
);

HB1xp67_ASAP7_75t_L g4156 ( 
.A(n_3156),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3239),
.Y(n_4157)
);

BUFx6f_ASAP7_75t_L g4158 ( 
.A(n_3653),
.Y(n_4158)
);

CKINVDCx5p33_ASAP7_75t_R g4159 ( 
.A(n_3528),
.Y(n_4159)
);

AO22x1_ASAP7_75t_L g4160 ( 
.A1(n_2972),
.A2(n_3040),
.B1(n_3049),
.B2(n_3819),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_3057),
.B(n_3061),
.Y(n_4161)
);

AOI22xp33_ASAP7_75t_L g4162 ( 
.A1(n_3603),
.A2(n_3833),
.B1(n_3882),
.B2(n_3241),
.Y(n_4162)
);

INVx2_ASAP7_75t_L g4163 ( 
.A(n_3384),
.Y(n_4163)
);

CKINVDCx5p33_ASAP7_75t_R g4164 ( 
.A(n_3528),
.Y(n_4164)
);

INVx2_ASAP7_75t_L g4165 ( 
.A(n_3384),
.Y(n_4165)
);

INVx2_ASAP7_75t_L g4166 ( 
.A(n_3384),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_3300),
.Y(n_4167)
);

NAND2xp5_ASAP7_75t_L g4168 ( 
.A(n_3068),
.B(n_3587),
.Y(n_4168)
);

NAND2xp5_ASAP7_75t_L g4169 ( 
.A(n_3068),
.B(n_3587),
.Y(n_4169)
);

INVx2_ASAP7_75t_SL g4170 ( 
.A(n_2995),
.Y(n_4170)
);

INVx2_ASAP7_75t_L g4171 ( 
.A(n_3300),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_L g4172 ( 
.A(n_3591),
.B(n_3601),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_3361),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_3361),
.Y(n_4174)
);

CKINVDCx5p33_ASAP7_75t_R g4175 ( 
.A(n_3561),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_SL g4176 ( 
.A(n_2965),
.B(n_3636),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_3372),
.Y(n_4177)
);

INVx3_ASAP7_75t_L g4178 ( 
.A(n_2961),
.Y(n_4178)
);

OAI22xp5_ASAP7_75t_L g4179 ( 
.A1(n_3581),
.A2(n_3583),
.B1(n_3707),
.B2(n_3644),
.Y(n_4179)
);

AND2x2_ASAP7_75t_L g4180 ( 
.A(n_3249),
.B(n_3282),
.Y(n_4180)
);

HB1xp67_ASAP7_75t_L g4181 ( 
.A(n_3156),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_3372),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_3305),
.Y(n_4183)
);

AOI22xp5_ASAP7_75t_L g4184 ( 
.A1(n_3882),
.A2(n_3603),
.B1(n_3040),
.B2(n_3241),
.Y(n_4184)
);

OAI22xp33_ASAP7_75t_L g4185 ( 
.A1(n_2983),
.A2(n_3049),
.B1(n_3629),
.B2(n_3628),
.Y(n_4185)
);

INVxp67_ASAP7_75t_L g4186 ( 
.A(n_3167),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_L g4187 ( 
.A(n_3591),
.B(n_3601),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_3605),
.B(n_3622),
.Y(n_4188)
);

OR2x2_ASAP7_75t_L g4189 ( 
.A(n_3167),
.B(n_3199),
.Y(n_4189)
);

BUFx4f_ASAP7_75t_SL g4190 ( 
.A(n_3020),
.Y(n_4190)
);

NOR2xp33_ASAP7_75t_L g4191 ( 
.A(n_2981),
.B(n_3723),
.Y(n_4191)
);

HB1xp67_ASAP7_75t_L g4192 ( 
.A(n_3162),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_3605),
.B(n_3622),
.Y(n_4193)
);

NAND2xp5_ASAP7_75t_L g4194 ( 
.A(n_3623),
.B(n_3625),
.Y(n_4194)
);

OR2x6_ASAP7_75t_L g4195 ( 
.A(n_3992),
.B(n_3023),
.Y(n_4195)
);

AND2x2_ASAP7_75t_L g4196 ( 
.A(n_3290),
.B(n_3385),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_3623),
.B(n_3625),
.Y(n_4197)
);

BUFx6f_ASAP7_75t_L g4198 ( 
.A(n_3653),
.Y(n_4198)
);

BUFx6f_ASAP7_75t_L g4199 ( 
.A(n_2986),
.Y(n_4199)
);

OAI22xp5_ASAP7_75t_L g4200 ( 
.A1(n_3739),
.A2(n_3770),
.B1(n_3797),
.B2(n_3761),
.Y(n_4200)
);

NOR2xp33_ASAP7_75t_L g4201 ( 
.A(n_3830),
.B(n_3835),
.Y(n_4201)
);

INVx2_ASAP7_75t_SL g4202 ( 
.A(n_2995),
.Y(n_4202)
);

BUFx6f_ASAP7_75t_L g4203 ( 
.A(n_2986),
.Y(n_4203)
);

INVx2_ASAP7_75t_SL g4204 ( 
.A(n_2995),
.Y(n_4204)
);

CKINVDCx20_ASAP7_75t_R g4205 ( 
.A(n_3746),
.Y(n_4205)
);

OR2x2_ASAP7_75t_L g4206 ( 
.A(n_3199),
.B(n_3210),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_3305),
.Y(n_4207)
);

BUFx6f_ASAP7_75t_L g4208 ( 
.A(n_3695),
.Y(n_4208)
);

INVx2_ASAP7_75t_L g4209 ( 
.A(n_3003),
.Y(n_4209)
);

BUFx2_ASAP7_75t_L g4210 ( 
.A(n_3612),
.Y(n_4210)
);

BUFx6f_ASAP7_75t_L g4211 ( 
.A(n_3695),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_3631),
.B(n_3632),
.Y(n_4212)
);

INVx3_ASAP7_75t_L g4213 ( 
.A(n_2961),
.Y(n_4213)
);

INVx2_ASAP7_75t_L g4214 ( 
.A(n_3003),
.Y(n_4214)
);

AND3x1_ASAP7_75t_L g4215 ( 
.A(n_3063),
.B(n_3806),
.C(n_3769),
.Y(n_4215)
);

AOI21xp5_ASAP7_75t_L g4216 ( 
.A1(n_2967),
.A2(n_3023),
.B(n_3021),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_SL g4217 ( 
.A(n_3675),
.B(n_3751),
.Y(n_4217)
);

NAND2xp5_ASAP7_75t_L g4218 ( 
.A(n_3631),
.B(n_3632),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_SL g4219 ( 
.A(n_3675),
.B(n_3751),
.Y(n_4219)
);

AND2x2_ASAP7_75t_L g4220 ( 
.A(n_3290),
.B(n_3385),
.Y(n_4220)
);

INVx2_ASAP7_75t_L g4221 ( 
.A(n_3003),
.Y(n_4221)
);

AND2x4_ASAP7_75t_L g4222 ( 
.A(n_3021),
.B(n_3030),
.Y(n_4222)
);

INVx2_ASAP7_75t_L g4223 ( 
.A(n_3060),
.Y(n_4223)
);

NAND2xp5_ASAP7_75t_L g4224 ( 
.A(n_3642),
.B(n_3649),
.Y(n_4224)
);

INVx4_ASAP7_75t_L g4225 ( 
.A(n_3392),
.Y(n_4225)
);

CKINVDCx5p33_ASAP7_75t_R g4226 ( 
.A(n_3561),
.Y(n_4226)
);

NAND2xp33_ASAP7_75t_SL g4227 ( 
.A(n_3940),
.B(n_3680),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_3642),
.B(n_3649),
.Y(n_4228)
);

INVx4_ASAP7_75t_L g4229 ( 
.A(n_3392),
.Y(n_4229)
);

BUFx6f_ASAP7_75t_L g4230 ( 
.A(n_3766),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_L g4231 ( 
.A(n_3651),
.B(n_3777),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_3162),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_L g4233 ( 
.A(n_3651),
.B(n_3777),
.Y(n_4233)
);

INVx2_ASAP7_75t_L g4234 ( 
.A(n_3060),
.Y(n_4234)
);

BUFx6f_ASAP7_75t_L g4235 ( 
.A(n_3766),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_SL g4236 ( 
.A(n_3794),
.B(n_3904),
.Y(n_4236)
);

CKINVDCx5p33_ASAP7_75t_R g4237 ( 
.A(n_3813),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_L g4238 ( 
.A(n_3781),
.B(n_3783),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_L g4239 ( 
.A(n_3781),
.B(n_3783),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_L g4240 ( 
.A(n_3787),
.B(n_3789),
.Y(n_4240)
);

BUFx6f_ASAP7_75t_L g4241 ( 
.A(n_3786),
.Y(n_4241)
);

CKINVDCx5p33_ASAP7_75t_R g4242 ( 
.A(n_3813),
.Y(n_4242)
);

AND2x2_ASAP7_75t_L g4243 ( 
.A(n_3385),
.B(n_3225),
.Y(n_4243)
);

INVx2_ASAP7_75t_L g4244 ( 
.A(n_3072),
.Y(n_4244)
);

NOR2xp33_ASAP7_75t_L g4245 ( 
.A(n_3865),
.B(n_3871),
.Y(n_4245)
);

OR2x6_ASAP7_75t_L g4246 ( 
.A(n_3992),
.B(n_3484),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_3162),
.Y(n_4247)
);

NOR2xp33_ASAP7_75t_L g4248 ( 
.A(n_3892),
.B(n_3900),
.Y(n_4248)
);

INVx2_ASAP7_75t_L g4249 ( 
.A(n_3072),
.Y(n_4249)
);

BUFx6f_ASAP7_75t_L g4250 ( 
.A(n_3786),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_SL g4251 ( 
.A(n_3794),
.B(n_3904),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_L g4252 ( 
.A(n_3787),
.B(n_3789),
.Y(n_4252)
);

CKINVDCx5p33_ASAP7_75t_R g4253 ( 
.A(n_3108),
.Y(n_4253)
);

BUFx2_ASAP7_75t_L g4254 ( 
.A(n_3778),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_SL g4255 ( 
.A(n_4001),
.B(n_3921),
.Y(n_4255)
);

NAND2x1p5_ASAP7_75t_L g4256 ( 
.A(n_3392),
.B(n_3819),
.Y(n_4256)
);

BUFx2_ASAP7_75t_L g4257 ( 
.A(n_3778),
.Y(n_4257)
);

BUFx6f_ASAP7_75t_L g4258 ( 
.A(n_3816),
.Y(n_4258)
);

INVx3_ASAP7_75t_L g4259 ( 
.A(n_2961),
.Y(n_4259)
);

BUFx4f_ASAP7_75t_SL g4260 ( 
.A(n_3020),
.Y(n_4260)
);

AND2x2_ASAP7_75t_L g4261 ( 
.A(n_3385),
.B(n_3225),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_3162),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_L g4263 ( 
.A(n_3793),
.B(n_3802),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_L g4264 ( 
.A(n_3793),
.B(n_3802),
.Y(n_4264)
);

BUFx4f_ASAP7_75t_SL g4265 ( 
.A(n_3020),
.Y(n_4265)
);

INVx1_ASAP7_75t_L g4266 ( 
.A(n_2980),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_3804),
.B(n_3805),
.Y(n_4267)
);

NOR2xp67_ASAP7_75t_L g4268 ( 
.A(n_2969),
.B(n_3392),
.Y(n_4268)
);

AND2x2_ASAP7_75t_L g4269 ( 
.A(n_2980),
.B(n_3033),
.Y(n_4269)
);

AOI22xp33_ASAP7_75t_L g4270 ( 
.A1(n_3603),
.A2(n_3241),
.B1(n_2960),
.B2(n_3664),
.Y(n_4270)
);

HB1xp67_ASAP7_75t_L g4271 ( 
.A(n_3210),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_3033),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_3041),
.Y(n_4273)
);

INVx6_ASAP7_75t_L g4274 ( 
.A(n_3392),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_SL g4275 ( 
.A(n_4001),
.B(n_3921),
.Y(n_4275)
);

INVx4_ASAP7_75t_L g4276 ( 
.A(n_3392),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_3041),
.Y(n_4277)
);

BUFx3_ASAP7_75t_L g4278 ( 
.A(n_3078),
.Y(n_4278)
);

INVx1_ASAP7_75t_SL g4279 ( 
.A(n_3926),
.Y(n_4279)
);

AOI22xp5_ASAP7_75t_L g4280 ( 
.A1(n_3714),
.A2(n_3752),
.B1(n_3779),
.B2(n_3717),
.Y(n_4280)
);

AOI21x1_ASAP7_75t_L g4281 ( 
.A1(n_3006),
.A2(n_3015),
.B(n_2997),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_L g4282 ( 
.A(n_3804),
.B(n_3805),
.Y(n_4282)
);

BUFx2_ASAP7_75t_L g4283 ( 
.A(n_3839),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_3045),
.Y(n_4284)
);

NOR2xp33_ASAP7_75t_L g4285 ( 
.A(n_3920),
.B(n_3922),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_SL g4286 ( 
.A(n_4039),
.B(n_3034),
.Y(n_4286)
);

AO22x1_ASAP7_75t_L g4287 ( 
.A1(n_3819),
.A2(n_4030),
.B1(n_3930),
.B2(n_3484),
.Y(n_4287)
);

INVx3_ASAP7_75t_SL g4288 ( 
.A(n_3992),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_3045),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_L g4290 ( 
.A(n_3811),
.B(n_3812),
.Y(n_4290)
);

AOI22xp5_ASAP7_75t_L g4291 ( 
.A1(n_3717),
.A2(n_3779),
.B1(n_3785),
.B2(n_3752),
.Y(n_4291)
);

BUFx2_ASAP7_75t_SL g4292 ( 
.A(n_3819),
.Y(n_4292)
);

AOI22xp33_ASAP7_75t_L g4293 ( 
.A1(n_3785),
.A2(n_3822),
.B1(n_3977),
.B2(n_3807),
.Y(n_4293)
);

INVxp67_ASAP7_75t_L g4294 ( 
.A(n_3216),
.Y(n_4294)
);

INVx2_ASAP7_75t_L g4295 ( 
.A(n_3072),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_3050),
.Y(n_4296)
);

CKINVDCx5p33_ASAP7_75t_R g4297 ( 
.A(n_3108),
.Y(n_4297)
);

BUFx2_ASAP7_75t_L g4298 ( 
.A(n_3839),
.Y(n_4298)
);

NAND3xp33_ASAP7_75t_SL g4299 ( 
.A(n_3062),
.B(n_3046),
.C(n_3008),
.Y(n_4299)
);

BUFx10_ASAP7_75t_L g4300 ( 
.A(n_3931),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_3811),
.B(n_3812),
.Y(n_4301)
);

INVx2_ASAP7_75t_SL g4302 ( 
.A(n_3030),
.Y(n_4302)
);

BUFx3_ASAP7_75t_L g4303 ( 
.A(n_3078),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_L g4304 ( 
.A(n_3815),
.B(n_3828),
.Y(n_4304)
);

INVx1_ASAP7_75t_SL g4305 ( 
.A(n_3926),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_3050),
.Y(n_4306)
);

AOI22xp5_ASAP7_75t_L g4307 ( 
.A1(n_3807),
.A2(n_3977),
.B1(n_3822),
.B2(n_3966),
.Y(n_4307)
);

BUFx3_ASAP7_75t_L g4308 ( 
.A(n_3078),
.Y(n_4308)
);

INVx2_ASAP7_75t_L g4309 ( 
.A(n_3084),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_L g4310 ( 
.A(n_3815),
.B(n_3828),
.Y(n_4310)
);

AOI22xp5_ASAP7_75t_L g4311 ( 
.A1(n_3963),
.A2(n_3985),
.B1(n_4002),
.B2(n_3967),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_L g4312 ( 
.A(n_3831),
.B(n_3834),
.Y(n_4312)
);

INVx2_ASAP7_75t_L g4313 ( 
.A(n_3084),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_3831),
.B(n_3834),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_SL g4315 ( 
.A(n_4039),
.B(n_4012),
.Y(n_4315)
);

BUFx4f_ASAP7_75t_L g4316 ( 
.A(n_3992),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_SL g4317 ( 
.A(n_4013),
.B(n_4033),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_3070),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_L g4319 ( 
.A(n_3838),
.B(n_3841),
.Y(n_4319)
);

BUFx3_ASAP7_75t_L g4320 ( 
.A(n_3078),
.Y(n_4320)
);

BUFx6f_ASAP7_75t_L g4321 ( 
.A(n_3816),
.Y(n_4321)
);

OAI22xp5_ASAP7_75t_SL g4322 ( 
.A1(n_2990),
.A2(n_4095),
.B1(n_4132),
.B2(n_4079),
.Y(n_4322)
);

NOR2xp33_ASAP7_75t_L g4323 ( 
.A(n_3588),
.B(n_3671),
.Y(n_4323)
);

BUFx3_ASAP7_75t_L g4324 ( 
.A(n_3078),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_3838),
.B(n_3841),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_SL g4326 ( 
.A(n_3655),
.B(n_3660),
.Y(n_4326)
);

BUFx2_ASAP7_75t_L g4327 ( 
.A(n_3846),
.Y(n_4327)
);

NOR2xp67_ASAP7_75t_L g4328 ( 
.A(n_2982),
.B(n_3043),
.Y(n_4328)
);

A2O1A1Ixp33_ASAP7_75t_L g4329 ( 
.A1(n_3836),
.A2(n_3894),
.B(n_3055),
.C(n_3663),
.Y(n_4329)
);

AND2x2_ASAP7_75t_L g4330 ( 
.A(n_3070),
.B(n_3110),
.Y(n_4330)
);

HB1xp67_ASAP7_75t_L g4331 ( 
.A(n_3216),
.Y(n_4331)
);

INVx2_ASAP7_75t_SL g4332 ( 
.A(n_3030),
.Y(n_4332)
);

AND2x2_ASAP7_75t_L g4333 ( 
.A(n_3110),
.B(n_3169),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_L g4334 ( 
.A(n_3843),
.B(n_3858),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_3843),
.B(n_3858),
.Y(n_4335)
);

HB1xp67_ASAP7_75t_L g4336 ( 
.A(n_3291),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_L g4337 ( 
.A(n_3860),
.B(n_3861),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_3169),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_3182),
.Y(n_4339)
);

CKINVDCx8_ASAP7_75t_R g4340 ( 
.A(n_3819),
.Y(n_4340)
);

AOI22xp33_ASAP7_75t_L g4341 ( 
.A1(n_3836),
.A2(n_3894),
.B1(n_3735),
.B2(n_4009),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_L g4342 ( 
.A(n_3860),
.B(n_3861),
.Y(n_4342)
);

OAI221xp5_ASAP7_75t_L g4343 ( 
.A1(n_3004),
.A2(n_3016),
.B1(n_3042),
.B2(n_3035),
.C(n_2991),
.Y(n_4343)
);

NAND2xp5_ASAP7_75t_L g4344 ( 
.A(n_3880),
.B(n_3883),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_L g4345 ( 
.A(n_3880),
.B(n_3883),
.Y(n_4345)
);

BUFx2_ASAP7_75t_L g4346 ( 
.A(n_3846),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_3182),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_3887),
.B(n_3888),
.Y(n_4348)
);

BUFx6f_ASAP7_75t_L g4349 ( 
.A(n_3960),
.Y(n_4349)
);

HB1xp67_ASAP7_75t_L g4350 ( 
.A(n_3291),
.Y(n_4350)
);

OR2x6_ASAP7_75t_L g4351 ( 
.A(n_3992),
.B(n_3009),
.Y(n_4351)
);

BUFx6f_ASAP7_75t_L g4352 ( 
.A(n_3960),
.Y(n_4352)
);

NOR2xp33_ASAP7_75t_L g4353 ( 
.A(n_3588),
.B(n_3671),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_3219),
.Y(n_4354)
);

NAND2xp5_ASAP7_75t_L g4355 ( 
.A(n_3887),
.B(n_3888),
.Y(n_4355)
);

NAND2xp5_ASAP7_75t_L g4356 ( 
.A(n_3890),
.B(n_3891),
.Y(n_4356)
);

AOI22xp5_ASAP7_75t_L g4357 ( 
.A1(n_3039),
.A2(n_3053),
.B1(n_4140),
.B2(n_4137),
.Y(n_4357)
);

NAND2xp5_ASAP7_75t_L g4358 ( 
.A(n_3890),
.B(n_3891),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_3893),
.B(n_3895),
.Y(n_4359)
);

BUFx6f_ASAP7_75t_L g4360 ( 
.A(n_3982),
.Y(n_4360)
);

AND2x4_ASAP7_75t_L g4361 ( 
.A(n_3030),
.B(n_3616),
.Y(n_4361)
);

NAND2xp5_ASAP7_75t_SL g4362 ( 
.A(n_3661),
.B(n_3665),
.Y(n_4362)
);

BUFx6f_ASAP7_75t_L g4363 ( 
.A(n_3982),
.Y(n_4363)
);

CKINVDCx5p33_ASAP7_75t_R g4364 ( 
.A(n_3808),
.Y(n_4364)
);

INVx2_ASAP7_75t_L g4365 ( 
.A(n_3145),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_3893),
.B(n_3895),
.Y(n_4366)
);

INVx2_ASAP7_75t_L g4367 ( 
.A(n_3146),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_3219),
.Y(n_4368)
);

INVx2_ASAP7_75t_L g4369 ( 
.A(n_3146),
.Y(n_4369)
);

INVxp67_ASAP7_75t_L g4370 ( 
.A(n_3375),
.Y(n_4370)
);

BUFx4f_ASAP7_75t_SL g4371 ( 
.A(n_3159),
.Y(n_4371)
);

AND2x2_ASAP7_75t_L g4372 ( 
.A(n_3220),
.B(n_3223),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_3220),
.Y(n_4373)
);

INVx1_ASAP7_75t_L g4374 ( 
.A(n_3223),
.Y(n_4374)
);

HB1xp67_ASAP7_75t_L g4375 ( 
.A(n_3375),
.Y(n_4375)
);

CKINVDCx5p33_ASAP7_75t_R g4376 ( 
.A(n_3808),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_3228),
.Y(n_4377)
);

NAND2xp5_ASAP7_75t_L g4378 ( 
.A(n_3903),
.B(n_3914),
.Y(n_4378)
);

AOI22xp33_ASAP7_75t_L g4379 ( 
.A1(n_4105),
.A2(n_3058),
.B1(n_2973),
.B2(n_2979),
.Y(n_4379)
);

BUFx8_ASAP7_75t_L g4380 ( 
.A(n_3494),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_3228),
.Y(n_4381)
);

AND2x4_ASAP7_75t_L g4382 ( 
.A(n_3616),
.B(n_3650),
.Y(n_4382)
);

AND2x4_ASAP7_75t_L g4383 ( 
.A(n_3616),
.B(n_3650),
.Y(n_4383)
);

OAI21xp5_ASAP7_75t_L g4384 ( 
.A1(n_3696),
.A2(n_4069),
.B(n_3048),
.Y(n_4384)
);

AND2x4_ASAP7_75t_L g4385 ( 
.A(n_3616),
.B(n_3650),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_3233),
.Y(n_4386)
);

BUFx2_ASAP7_75t_L g4387 ( 
.A(n_4139),
.Y(n_4387)
);

AND2x2_ASAP7_75t_L g4388 ( 
.A(n_3233),
.B(n_3243),
.Y(n_4388)
);

NAND2xp5_ASAP7_75t_SL g4389 ( 
.A(n_3667),
.B(n_3672),
.Y(n_4389)
);

NAND2xp5_ASAP7_75t_L g4390 ( 
.A(n_3903),
.B(n_3914),
.Y(n_4390)
);

CKINVDCx20_ASAP7_75t_R g4391 ( 
.A(n_3998),
.Y(n_4391)
);

BUFx6f_ASAP7_75t_L g4392 ( 
.A(n_4015),
.Y(n_4392)
);

AOI21xp5_ASAP7_75t_L g4393 ( 
.A1(n_3674),
.A2(n_3687),
.B(n_3682),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_3243),
.Y(n_4394)
);

AOI221xp5_ASAP7_75t_L g4395 ( 
.A1(n_4137),
.A2(n_4140),
.B1(n_3823),
.B2(n_3886),
.C(n_3719),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_3260),
.Y(n_4396)
);

NAND2xp5_ASAP7_75t_L g4397 ( 
.A(n_3915),
.B(n_3917),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_3260),
.Y(n_4398)
);

HB1xp67_ASAP7_75t_L g4399 ( 
.A(n_3311),
.Y(n_4399)
);

HB1xp67_ASAP7_75t_L g4400 ( 
.A(n_3311),
.Y(n_4400)
);

AOI21xp5_ASAP7_75t_L g4401 ( 
.A1(n_3689),
.A2(n_3699),
.B(n_3698),
.Y(n_4401)
);

INVxp67_ASAP7_75t_L g4402 ( 
.A(n_3067),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_L g4403 ( 
.A(n_3915),
.B(n_3917),
.Y(n_4403)
);

HB1xp67_ASAP7_75t_L g4404 ( 
.A(n_3320),
.Y(n_4404)
);

HB1xp67_ASAP7_75t_L g4405 ( 
.A(n_3320),
.Y(n_4405)
);

CKINVDCx5p33_ASAP7_75t_R g4406 ( 
.A(n_4062),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_SL g4407 ( 
.A(n_3705),
.B(n_3706),
.Y(n_4407)
);

HB1xp67_ASAP7_75t_L g4408 ( 
.A(n_3325),
.Y(n_4408)
);

AOI22xp33_ASAP7_75t_L g4409 ( 
.A1(n_2978),
.A2(n_2987),
.B1(n_3005),
.B2(n_3002),
.Y(n_4409)
);

AND2x2_ASAP7_75t_L g4410 ( 
.A(n_3264),
.B(n_3267),
.Y(n_4410)
);

NAND2xp5_ASAP7_75t_SL g4411 ( 
.A(n_3713),
.B(n_3720),
.Y(n_4411)
);

NOR2xp33_ASAP7_75t_L g4412 ( 
.A(n_3697),
.B(n_3719),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_L g4413 ( 
.A(n_3918),
.B(n_3923),
.Y(n_4413)
);

AND3x1_ASAP7_75t_SL g4414 ( 
.A(n_4052),
.B(n_3035),
.C(n_3678),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_L g4415 ( 
.A(n_3918),
.B(n_3923),
.Y(n_4415)
);

INVx5_ASAP7_75t_L g4416 ( 
.A(n_3455),
.Y(n_4416)
);

INVx4_ASAP7_75t_L g4417 ( 
.A(n_3422),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_L g4418 ( 
.A(n_3934),
.B(n_3935),
.Y(n_4418)
);

BUFx2_ASAP7_75t_L g4419 ( 
.A(n_4139),
.Y(n_4419)
);

BUFx3_ASAP7_75t_L g4420 ( 
.A(n_3009),
.Y(n_4420)
);

OAI21x1_ASAP7_75t_L g4421 ( 
.A1(n_3006),
.A2(n_3015),
.B(n_2997),
.Y(n_4421)
);

AND2x6_ASAP7_75t_SL g4422 ( 
.A(n_3234),
.B(n_3393),
.Y(n_4422)
);

CKINVDCx5p33_ASAP7_75t_R g4423 ( 
.A(n_4062),
.Y(n_4423)
);

AND2x4_ASAP7_75t_L g4424 ( 
.A(n_3650),
.B(n_3730),
.Y(n_4424)
);

NOR2xp33_ASAP7_75t_L g4425 ( 
.A(n_3697),
.B(n_3823),
.Y(n_4425)
);

NOR2xp33_ASAP7_75t_L g4426 ( 
.A(n_3886),
.B(n_3901),
.Y(n_4426)
);

BUFx2_ASAP7_75t_L g4427 ( 
.A(n_3586),
.Y(n_4427)
);

NOR2xp67_ASAP7_75t_L g4428 ( 
.A(n_2982),
.B(n_3043),
.Y(n_4428)
);

BUFx3_ASAP7_75t_L g4429 ( 
.A(n_3009),
.Y(n_4429)
);

CKINVDCx5p33_ASAP7_75t_R g4430 ( 
.A(n_3481),
.Y(n_4430)
);

AOI22xp33_ASAP7_75t_L g4431 ( 
.A1(n_3007),
.A2(n_3018),
.B1(n_3076),
.B2(n_3016),
.Y(n_4431)
);

AND2x4_ASAP7_75t_L g4432 ( 
.A(n_3730),
.B(n_3765),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_3340),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_3340),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_3357),
.Y(n_4435)
);

NOR2xp33_ASAP7_75t_L g4436 ( 
.A(n_3901),
.B(n_3979),
.Y(n_4436)
);

NAND2x1p5_ASAP7_75t_L g4437 ( 
.A(n_3819),
.B(n_3422),
.Y(n_4437)
);

INVxp67_ASAP7_75t_L g4438 ( 
.A(n_3067),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_3934),
.B(n_3935),
.Y(n_4439)
);

BUFx6f_ASAP7_75t_L g4440 ( 
.A(n_4015),
.Y(n_4440)
);

NAND2xp5_ASAP7_75t_L g4441 ( 
.A(n_3937),
.B(n_3943),
.Y(n_4441)
);

AOI21xp5_ASAP7_75t_L g4442 ( 
.A1(n_3721),
.A2(n_3727),
.B(n_3726),
.Y(n_4442)
);

CKINVDCx5p33_ASAP7_75t_R g4443 ( 
.A(n_3481),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_3357),
.Y(n_4444)
);

AND2x2_ASAP7_75t_L g4445 ( 
.A(n_3378),
.B(n_3383),
.Y(n_4445)
);

INVx2_ASAP7_75t_SL g4446 ( 
.A(n_3730),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_3937),
.B(n_3943),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_3378),
.Y(n_4448)
);

BUFx2_ASAP7_75t_L g4449 ( 
.A(n_3658),
.Y(n_4449)
);

HB1xp67_ASAP7_75t_L g4450 ( 
.A(n_3325),
.Y(n_4450)
);

BUFx4f_ASAP7_75t_L g4451 ( 
.A(n_3527),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_3944),
.B(n_3952),
.Y(n_4452)
);

CKINVDCx16_ASAP7_75t_R g4453 ( 
.A(n_3500),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_L g4454 ( 
.A(n_3944),
.B(n_3952),
.Y(n_4454)
);

BUFx2_ASAP7_75t_L g4455 ( 
.A(n_3658),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_3383),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_3387),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_L g4458 ( 
.A(n_3959),
.B(n_3964),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_L g4459 ( 
.A(n_3959),
.B(n_3964),
.Y(n_4459)
);

BUFx2_ASAP7_75t_L g4460 ( 
.A(n_3658),
.Y(n_4460)
);

BUFx4f_ASAP7_75t_L g4461 ( 
.A(n_3527),
.Y(n_4461)
);

INVx4_ASAP7_75t_L g4462 ( 
.A(n_3422),
.Y(n_4462)
);

NAND2xp5_ASAP7_75t_SL g4463 ( 
.A(n_3737),
.B(n_3740),
.Y(n_4463)
);

AND2x2_ASAP7_75t_L g4464 ( 
.A(n_3582),
.B(n_3589),
.Y(n_4464)
);

HB1xp67_ASAP7_75t_L g4465 ( 
.A(n_3355),
.Y(n_4465)
);

NOR2xp33_ASAP7_75t_L g4466 ( 
.A(n_3979),
.B(n_3987),
.Y(n_4466)
);

NOR2xp33_ASAP7_75t_L g4467 ( 
.A(n_3987),
.B(n_4014),
.Y(n_4467)
);

BUFx2_ASAP7_75t_L g4468 ( 
.A(n_3658),
.Y(n_4468)
);

AND2x2_ASAP7_75t_L g4469 ( 
.A(n_3589),
.B(n_3598),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_L g4470 ( 
.A(n_3970),
.B(n_3976),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_SL g4471 ( 
.A(n_3742),
.B(n_3745),
.Y(n_4471)
);

AND2x4_ASAP7_75t_L g4472 ( 
.A(n_3730),
.B(n_3765),
.Y(n_4472)
);

NAND2x1p5_ASAP7_75t_L g4473 ( 
.A(n_3819),
.B(n_3422),
.Y(n_4473)
);

NAND2xp5_ASAP7_75t_L g4474 ( 
.A(n_3970),
.B(n_3976),
.Y(n_4474)
);

INVx1_ASAP7_75t_SL g4475 ( 
.A(n_4025),
.Y(n_4475)
);

NOR2xp33_ASAP7_75t_SL g4476 ( 
.A(n_3455),
.B(n_3526),
.Y(n_4476)
);

AOI22xp33_ASAP7_75t_L g4477 ( 
.A1(n_3004),
.A2(n_3042),
.B1(n_4014),
.B2(n_4138),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_L g4478 ( 
.A(n_3991),
.B(n_3994),
.Y(n_4478)
);

BUFx6f_ASAP7_75t_L g4479 ( 
.A(n_4090),
.Y(n_4479)
);

BUFx12f_ASAP7_75t_L g4480 ( 
.A(n_3088),
.Y(n_4480)
);

NAND2xp5_ASAP7_75t_L g4481 ( 
.A(n_3991),
.B(n_3994),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_L g4482 ( 
.A(n_4008),
.B(n_4022),
.Y(n_4482)
);

OR2x2_ASAP7_75t_SL g4483 ( 
.A(n_3551),
.B(n_3407),
.Y(n_4483)
);

INVx1_ASAP7_75t_SL g4484 ( 
.A(n_4025),
.Y(n_4484)
);

AND2x4_ASAP7_75t_L g4485 ( 
.A(n_3765),
.B(n_3818),
.Y(n_4485)
);

AND2x4_ASAP7_75t_L g4486 ( 
.A(n_3765),
.B(n_3818),
.Y(n_4486)
);

AND2x4_ASAP7_75t_L g4487 ( 
.A(n_3818),
.B(n_3911),
.Y(n_4487)
);

AND2x2_ASAP7_75t_L g4488 ( 
.A(n_3619),
.B(n_3656),
.Y(n_4488)
);

NAND2xp5_ASAP7_75t_L g4489 ( 
.A(n_4008),
.B(n_4022),
.Y(n_4489)
);

INVx5_ASAP7_75t_L g4490 ( 
.A(n_3455),
.Y(n_4490)
);

HB1xp67_ASAP7_75t_L g4491 ( 
.A(n_3355),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_4023),
.B(n_4035),
.Y(n_4492)
);

INVxp67_ASAP7_75t_L g4493 ( 
.A(n_3067),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_L g4494 ( 
.A(n_4023),
.B(n_4035),
.Y(n_4494)
);

NAND2xp5_ASAP7_75t_L g4495 ( 
.A(n_4050),
.B(n_4055),
.Y(n_4495)
);

AOI22xp33_ASAP7_75t_L g4496 ( 
.A1(n_4138),
.A2(n_3599),
.B1(n_3803),
.B2(n_3654),
.Y(n_4496)
);

HB1xp67_ASAP7_75t_L g4497 ( 
.A(n_3368),
.Y(n_4497)
);

NAND2xp5_ASAP7_75t_L g4498 ( 
.A(n_4050),
.B(n_4055),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_4056),
.B(n_4072),
.Y(n_4499)
);

NAND2xp5_ASAP7_75t_SL g4500 ( 
.A(n_3754),
.B(n_3763),
.Y(n_4500)
);

OR2x6_ASAP7_75t_L g4501 ( 
.A(n_3027),
.B(n_3590),
.Y(n_4501)
);

AND2x2_ASAP7_75t_L g4502 ( 
.A(n_3677),
.B(n_3683),
.Y(n_4502)
);

AND2x2_ASAP7_75t_L g4503 ( 
.A(n_3677),
.B(n_3683),
.Y(n_4503)
);

HB1xp67_ASAP7_75t_L g4504 ( 
.A(n_3368),
.Y(n_4504)
);

CKINVDCx5p33_ASAP7_75t_R g4505 ( 
.A(n_3481),
.Y(n_4505)
);

NAND2xp5_ASAP7_75t_SL g4506 ( 
.A(n_4106),
.B(n_4110),
.Y(n_4506)
);

AND2x4_ASAP7_75t_L g4507 ( 
.A(n_3818),
.B(n_3911),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_L g4508 ( 
.A(n_4056),
.B(n_4072),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_L g4509 ( 
.A(n_4073),
.B(n_4076),
.Y(n_4509)
);

NAND2xp5_ASAP7_75t_L g4510 ( 
.A(n_4073),
.B(n_4076),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_3709),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_L g4512 ( 
.A(n_4078),
.B(n_4080),
.Y(n_4512)
);

HB1xp67_ASAP7_75t_L g4513 ( 
.A(n_3394),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_SL g4514 ( 
.A(n_4112),
.B(n_4115),
.Y(n_4514)
);

BUFx6f_ASAP7_75t_L g4515 ( 
.A(n_4090),
.Y(n_4515)
);

OAI22xp5_ASAP7_75t_L g4516 ( 
.A1(n_3008),
.A2(n_3046),
.B1(n_3594),
.B2(n_2974),
.Y(n_4516)
);

CKINVDCx5p33_ASAP7_75t_R g4517 ( 
.A(n_3088),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_3732),
.Y(n_4518)
);

CKINVDCx11_ASAP7_75t_R g4519 ( 
.A(n_3133),
.Y(n_4519)
);

INVx5_ASAP7_75t_L g4520 ( 
.A(n_3455),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_3732),
.Y(n_4521)
);

INVx1_ASAP7_75t_L g4522 ( 
.A(n_3749),
.Y(n_4522)
);

INVx5_ASAP7_75t_L g4523 ( 
.A(n_3526),
.Y(n_4523)
);

NAND2xp5_ASAP7_75t_L g4524 ( 
.A(n_4078),
.B(n_4080),
.Y(n_4524)
);

NOR2xp33_ASAP7_75t_L g4525 ( 
.A(n_3062),
.B(n_4052),
.Y(n_4525)
);

HB1xp67_ASAP7_75t_L g4526 ( 
.A(n_3394),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_3749),
.Y(n_4527)
);

AO22x1_ASAP7_75t_L g4528 ( 
.A1(n_3930),
.A2(n_4030),
.B1(n_4041),
.B2(n_3585),
.Y(n_4528)
);

OR2x6_ASAP7_75t_L g4529 ( 
.A(n_3027),
.B(n_3590),
.Y(n_4529)
);

BUFx6f_ASAP7_75t_L g4530 ( 
.A(n_4114),
.Y(n_4530)
);

HB1xp67_ASAP7_75t_L g4531 ( 
.A(n_4125),
.Y(n_4531)
);

AND2x2_ASAP7_75t_L g4532 ( 
.A(n_3750),
.B(n_3759),
.Y(n_4532)
);

BUFx2_ASAP7_75t_L g4533 ( 
.A(n_3690),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_L g4534 ( 
.A(n_4081),
.B(n_4082),
.Y(n_4534)
);

BUFx6f_ASAP7_75t_L g4535 ( 
.A(n_4114),
.Y(n_4535)
);

AND3x1_ASAP7_75t_L g4536 ( 
.A(n_3391),
.B(n_4029),
.C(n_3984),
.Y(n_4536)
);

AND2x6_ASAP7_75t_L g4537 ( 
.A(n_3500),
.B(n_3091),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_3750),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_4081),
.B(n_4082),
.Y(n_4539)
);

NAND2xp5_ASAP7_75t_L g4540 ( 
.A(n_4084),
.B(n_4085),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_L g4541 ( 
.A(n_4084),
.B(n_4085),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_SL g4542 ( 
.A(n_4117),
.B(n_4118),
.Y(n_4542)
);

CKINVDCx5p33_ASAP7_75t_R g4543 ( 
.A(n_3088),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_3759),
.Y(n_4544)
);

OR2x2_ASAP7_75t_L g4545 ( 
.A(n_3173),
.B(n_3232),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_SL g4546 ( 
.A(n_4120),
.B(n_4122),
.Y(n_4546)
);

NAND2xp33_ASAP7_75t_L g4547 ( 
.A(n_3599),
.B(n_3803),
.Y(n_4547)
);

NOR2xp33_ASAP7_75t_L g4548 ( 
.A(n_4126),
.B(n_4134),
.Y(n_4548)
);

NAND2xp5_ASAP7_75t_L g4549 ( 
.A(n_4086),
.B(n_4093),
.Y(n_4549)
);

NAND2xp5_ASAP7_75t_L g4550 ( 
.A(n_4086),
.B(n_4093),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_3790),
.Y(n_4551)
);

OR2x2_ASAP7_75t_L g4552 ( 
.A(n_3173),
.B(n_3232),
.Y(n_4552)
);

INVxp67_ASAP7_75t_L g4553 ( 
.A(n_3092),
.Y(n_4553)
);

HB1xp67_ASAP7_75t_L g4554 ( 
.A(n_4125),
.Y(n_4554)
);

NAND2x1_ASAP7_75t_L g4555 ( 
.A(n_3099),
.B(n_3690),
.Y(n_4555)
);

NAND2xp5_ASAP7_75t_L g4556 ( 
.A(n_4127),
.B(n_4136),
.Y(n_4556)
);

AND3x1_ASAP7_75t_SL g4557 ( 
.A(n_3728),
.B(n_4131),
.C(n_3996),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_3790),
.Y(n_4558)
);

INVx4_ASAP7_75t_L g4559 ( 
.A(n_3526),
.Y(n_4559)
);

AND2x6_ASAP7_75t_L g4560 ( 
.A(n_3363),
.B(n_3404),
.Y(n_4560)
);

AND2x2_ASAP7_75t_L g4561 ( 
.A(n_3791),
.B(n_3801),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_3791),
.Y(n_4562)
);

BUFx6f_ASAP7_75t_L g4563 ( 
.A(n_3119),
.Y(n_4563)
);

BUFx2_ASAP7_75t_L g4564 ( 
.A(n_3725),
.Y(n_4564)
);

HB1xp67_ASAP7_75t_L g4565 ( 
.A(n_4125),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_3801),
.Y(n_4566)
);

NAND2xp5_ASAP7_75t_L g4567 ( 
.A(n_3190),
.B(n_2964),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_3840),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_3840),
.Y(n_4569)
);

NAND2xp5_ASAP7_75t_L g4570 ( 
.A(n_3190),
.B(n_3079),
.Y(n_4570)
);

HB1xp67_ASAP7_75t_L g4571 ( 
.A(n_4125),
.Y(n_4571)
);

NAND2xp5_ASAP7_75t_SL g4572 ( 
.A(n_3597),
.B(n_3652),
.Y(n_4572)
);

AND2x2_ASAP7_75t_L g4573 ( 
.A(n_3842),
.B(n_3845),
.Y(n_4573)
);

NOR2xp33_ASAP7_75t_L g4574 ( 
.A(n_3701),
.B(n_3756),
.Y(n_4574)
);

NOR2xp33_ASAP7_75t_SL g4575 ( 
.A(n_3526),
.B(n_3097),
.Y(n_4575)
);

NAND2xp5_ASAP7_75t_L g4576 ( 
.A(n_3079),
.B(n_3080),
.Y(n_4576)
);

AND3x1_ASAP7_75t_L g4577 ( 
.A(n_3391),
.B(n_3022),
.C(n_3317),
.Y(n_4577)
);

INVx4_ASAP7_75t_L g4578 ( 
.A(n_3725),
.Y(n_4578)
);

NAND2xp5_ASAP7_75t_L g4579 ( 
.A(n_3080),
.B(n_3246),
.Y(n_4579)
);

NAND2xp5_ASAP7_75t_SL g4580 ( 
.A(n_3800),
.B(n_3849),
.Y(n_4580)
);

AOI221xp5_ASAP7_75t_L g4581 ( 
.A1(n_3131),
.A2(n_3137),
.B1(n_3064),
.B2(n_3157),
.C(n_3868),
.Y(n_4581)
);

AND2x2_ASAP7_75t_L g4582 ( 
.A(n_3842),
.B(n_3845),
.Y(n_4582)
);

OR2x6_ASAP7_75t_L g4583 ( 
.A(n_3590),
.B(n_3657),
.Y(n_4583)
);

BUFx4f_ASAP7_75t_L g4584 ( 
.A(n_3527),
.Y(n_4584)
);

NAND2xp5_ASAP7_75t_L g4585 ( 
.A(n_3246),
.B(n_3253),
.Y(n_4585)
);

NOR2x1_ASAP7_75t_R g4586 ( 
.A(n_3159),
.B(n_3741),
.Y(n_4586)
);

INVx4_ASAP7_75t_L g4587 ( 
.A(n_3725),
.Y(n_4587)
);

AOI22xp33_ASAP7_75t_L g4588 ( 
.A1(n_3596),
.A2(n_3955),
.B1(n_4047),
.B2(n_3780),
.Y(n_4588)
);

OAI22xp5_ASAP7_75t_L g4589 ( 
.A1(n_3941),
.A2(n_3989),
.B1(n_3975),
.B2(n_3037),
.Y(n_4589)
);

BUFx6f_ASAP7_75t_L g4590 ( 
.A(n_3119),
.Y(n_4590)
);

OAI22xp5_ASAP7_75t_L g4591 ( 
.A1(n_3024),
.A2(n_3673),
.B1(n_3688),
.B2(n_3585),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_3878),
.Y(n_4592)
);

BUFx2_ASAP7_75t_L g4593 ( 
.A(n_3725),
.Y(n_4593)
);

NOR2x2_ASAP7_75t_L g4594 ( 
.A(n_3559),
.B(n_3302),
.Y(n_4594)
);

OR2x6_ASAP7_75t_L g4595 ( 
.A(n_3590),
.B(n_3657),
.Y(n_4595)
);

NAND2xp5_ASAP7_75t_L g4596 ( 
.A(n_3253),
.B(n_3256),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_3878),
.Y(n_4597)
);

INVx2_ASAP7_75t_SL g4598 ( 
.A(n_3911),
.Y(n_4598)
);

NAND2xp5_ASAP7_75t_L g4599 ( 
.A(n_3256),
.B(n_3266),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_3881),
.Y(n_4600)
);

OR2x2_ASAP7_75t_SL g4601 ( 
.A(n_3551),
.B(n_3407),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_L g4602 ( 
.A(n_3266),
.B(n_3283),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_3881),
.Y(n_4603)
);

INVx1_ASAP7_75t_L g4604 ( 
.A(n_3897),
.Y(n_4604)
);

AOI22xp33_ASAP7_75t_L g4605 ( 
.A1(n_2991),
.A2(n_3077),
.B1(n_3940),
.B2(n_3064),
.Y(n_4605)
);

NOR2xp33_ASAP7_75t_L g4606 ( 
.A(n_3048),
.B(n_3615),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_3283),
.B(n_3284),
.Y(n_4607)
);

NOR2xp33_ASAP7_75t_R g4608 ( 
.A(n_2999),
.B(n_3001),
.Y(n_4608)
);

INVx2_ASAP7_75t_SL g4609 ( 
.A(n_3911),
.Y(n_4609)
);

NAND2xp5_ASAP7_75t_L g4610 ( 
.A(n_3284),
.B(n_3129),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_L g4611 ( 
.A(n_3129),
.B(n_3081),
.Y(n_4611)
);

AND2x2_ASAP7_75t_L g4612 ( 
.A(n_3897),
.B(n_3946),
.Y(n_4612)
);

NAND2xp5_ASAP7_75t_L g4613 ( 
.A(n_3081),
.B(n_3112),
.Y(n_4613)
);

BUFx4f_ASAP7_75t_SL g4614 ( 
.A(n_3159),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_3946),
.Y(n_4615)
);

AND2x2_ASAP7_75t_L g4616 ( 
.A(n_3972),
.B(n_3993),
.Y(n_4616)
);

BUFx2_ASAP7_75t_L g4617 ( 
.A(n_3772),
.Y(n_4617)
);

NOR2xp33_ASAP7_75t_L g4618 ( 
.A(n_3615),
.B(n_3938),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_3972),
.Y(n_4619)
);

OAI21xp5_ASAP7_75t_L g4620 ( 
.A1(n_3032),
.A2(n_3795),
.B(n_3792),
.Y(n_4620)
);

OR2x6_ASAP7_75t_L g4621 ( 
.A(n_3657),
.B(n_3659),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_3993),
.Y(n_4622)
);

INVx5_ASAP7_75t_L g4623 ( 
.A(n_2975),
.Y(n_4623)
);

AOI22xp5_ASAP7_75t_L g4624 ( 
.A1(n_3938),
.A2(n_3144),
.B1(n_3149),
.B2(n_3142),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4010),
.Y(n_4625)
);

AND2x2_ASAP7_75t_L g4626 ( 
.A(n_4010),
.B(n_4028),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_L g4627 ( 
.A(n_3112),
.B(n_3116),
.Y(n_4627)
);

OR2x2_ASAP7_75t_L g4628 ( 
.A(n_4028),
.B(n_4053),
.Y(n_4628)
);

A2O1A1Ixp33_ASAP7_75t_L g4629 ( 
.A1(n_3055),
.A2(n_3038),
.B(n_3089),
.C(n_2970),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_4053),
.Y(n_4630)
);

NAND2xp5_ASAP7_75t_SL g4631 ( 
.A(n_3637),
.B(n_3673),
.Y(n_4631)
);

CKINVDCx5p33_ASAP7_75t_R g4632 ( 
.A(n_3088),
.Y(n_4632)
);

AND2x2_ASAP7_75t_L g4633 ( 
.A(n_4054),
.B(n_4063),
.Y(n_4633)
);

NAND2xp5_ASAP7_75t_L g4634 ( 
.A(n_3116),
.B(n_3124),
.Y(n_4634)
);

NAND2xp5_ASAP7_75t_L g4635 ( 
.A(n_3124),
.B(n_3637),
.Y(n_4635)
);

NAND2xp5_ASAP7_75t_L g4636 ( 
.A(n_3688),
.B(n_3702),
.Y(n_4636)
);

NAND2x1p5_ASAP7_75t_L g4637 ( 
.A(n_2975),
.B(n_3755),
.Y(n_4637)
);

HB1xp67_ASAP7_75t_L g4638 ( 
.A(n_4054),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_SL g4639 ( 
.A(n_3702),
.B(n_3704),
.Y(n_4639)
);

NAND2xp5_ASAP7_75t_L g4640 ( 
.A(n_3704),
.B(n_3722),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4063),
.Y(n_4641)
);

INVx3_ASAP7_75t_SL g4642 ( 
.A(n_3302),
.Y(n_4642)
);

NAND2xp5_ASAP7_75t_L g4643 ( 
.A(n_4113),
.B(n_3722),
.Y(n_4643)
);

AND2x2_ASAP7_75t_L g4644 ( 
.A(n_4099),
.B(n_4102),
.Y(n_4644)
);

AND3x1_ASAP7_75t_L g4645 ( 
.A(n_3317),
.B(n_3065),
.C(n_2985),
.Y(n_4645)
);

AND2x2_ASAP7_75t_L g4646 ( 
.A(n_4099),
.B(n_4102),
.Y(n_4646)
);

NAND2xp5_ASAP7_75t_L g4647 ( 
.A(n_3734),
.B(n_3743),
.Y(n_4647)
);

NOR2xp33_ASAP7_75t_L g4648 ( 
.A(n_3054),
.B(n_2999),
.Y(n_4648)
);

CKINVDCx5p33_ASAP7_75t_R g4649 ( 
.A(n_3969),
.Y(n_4649)
);

AND2x2_ASAP7_75t_L g4650 ( 
.A(n_4121),
.B(n_3029),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_SL g4651 ( 
.A(n_3734),
.B(n_3743),
.Y(n_4651)
);

AOI22xp33_ASAP7_75t_L g4652 ( 
.A1(n_3150),
.A2(n_3771),
.B1(n_3824),
.B2(n_3768),
.Y(n_4652)
);

NAND2xp5_ASAP7_75t_L g4653 ( 
.A(n_3768),
.B(n_3771),
.Y(n_4653)
);

AND2x2_ASAP7_75t_L g4654 ( 
.A(n_4121),
.B(n_3029),
.Y(n_4654)
);

NAND2xp5_ASAP7_75t_L g4655 ( 
.A(n_3824),
.B(n_3829),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_3360),
.Y(n_4656)
);

AOI22xp33_ASAP7_75t_L g4657 ( 
.A1(n_3150),
.A2(n_3832),
.B1(n_3852),
.B2(n_3829),
.Y(n_4657)
);

NAND2xp5_ASAP7_75t_L g4658 ( 
.A(n_4113),
.B(n_3832),
.Y(n_4658)
);

AND2x4_ASAP7_75t_L g4659 ( 
.A(n_4005),
.B(n_4027),
.Y(n_4659)
);

BUFx2_ASAP7_75t_L g4660 ( 
.A(n_3773),
.Y(n_4660)
);

HB1xp67_ASAP7_75t_L g4661 ( 
.A(n_3044),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_3360),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_3371),
.Y(n_4663)
);

AOI22xp5_ASAP7_75t_L g4664 ( 
.A1(n_3170),
.A2(n_3197),
.B1(n_3194),
.B2(n_3137),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_3371),
.Y(n_4665)
);

BUFx8_ASAP7_75t_L g4666 ( 
.A(n_3494),
.Y(n_4666)
);

NAND2xp5_ASAP7_75t_L g4667 ( 
.A(n_3852),
.B(n_3857),
.Y(n_4667)
);

AOI22xp33_ASAP7_75t_L g4668 ( 
.A1(n_3857),
.A2(n_3874),
.B1(n_3924),
.B2(n_3863),
.Y(n_4668)
);

AOI22xp33_ASAP7_75t_L g4669 ( 
.A1(n_3863),
.A2(n_3924),
.B1(n_3958),
.B2(n_3874),
.Y(n_4669)
);

CKINVDCx5p33_ASAP7_75t_R g4670 ( 
.A(n_3969),
.Y(n_4670)
);

NAND2xp5_ASAP7_75t_L g4671 ( 
.A(n_3958),
.B(n_3988),
.Y(n_4671)
);

NAND2xp5_ASAP7_75t_L g4672 ( 
.A(n_3988),
.B(n_4048),
.Y(n_4672)
);

BUFx2_ASAP7_75t_L g4673 ( 
.A(n_3773),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_3380),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_3380),
.Y(n_4675)
);

AND2x4_ASAP7_75t_L g4676 ( 
.A(n_4005),
.B(n_4027),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_L g4677 ( 
.A(n_4048),
.B(n_4075),
.Y(n_4677)
);

NOR2xp33_ASAP7_75t_L g4678 ( 
.A(n_3025),
.B(n_3131),
.Y(n_4678)
);

OAI22xp5_ASAP7_75t_L g4679 ( 
.A1(n_4104),
.A2(n_4075),
.B1(n_4135),
.B2(n_4130),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_3381),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_3381),
.Y(n_4681)
);

CKINVDCx5p33_ASAP7_75t_R g4682 ( 
.A(n_3969),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_L g4683 ( 
.A(n_4104),
.B(n_3127),
.Y(n_4683)
);

NAND2xp5_ASAP7_75t_L g4684 ( 
.A(n_3127),
.B(n_3172),
.Y(n_4684)
);

NAND2xp5_ASAP7_75t_L g4685 ( 
.A(n_3172),
.B(n_3175),
.Y(n_4685)
);

AND2x4_ASAP7_75t_L g4686 ( 
.A(n_4005),
.B(n_4027),
.Y(n_4686)
);

BUFx2_ASAP7_75t_L g4687 ( 
.A(n_3870),
.Y(n_4687)
);

OR2x2_ASAP7_75t_L g4688 ( 
.A(n_3275),
.B(n_3289),
.Y(n_4688)
);

NOR2xp33_ASAP7_75t_L g4689 ( 
.A(n_3217),
.B(n_3001),
.Y(n_4689)
);

AOI22xp5_ASAP7_75t_L g4690 ( 
.A1(n_3235),
.A2(n_3265),
.B1(n_3130),
.B2(n_2962),
.Y(n_4690)
);

NAND2xp5_ASAP7_75t_SL g4691 ( 
.A(n_3038),
.B(n_3792),
.Y(n_4691)
);

NAND2xp5_ASAP7_75t_SL g4692 ( 
.A(n_3795),
.B(n_3875),
.Y(n_4692)
);

BUFx2_ASAP7_75t_L g4693 ( 
.A(n_3870),
.Y(n_4693)
);

INVx4_ASAP7_75t_L g4694 ( 
.A(n_3870),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_3382),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_SL g4696 ( 
.A(n_3875),
.B(n_4067),
.Y(n_4696)
);

NOR2xp33_ASAP7_75t_L g4697 ( 
.A(n_3217),
.B(n_3026),
.Y(n_4697)
);

AOI21xp5_ASAP7_75t_L g4698 ( 
.A1(n_2988),
.A2(n_3017),
.B(n_3602),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_3382),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_L g4700 ( 
.A(n_3175),
.B(n_3176),
.Y(n_4700)
);

AND2x2_ASAP7_75t_L g4701 ( 
.A(n_3044),
.B(n_3111),
.Y(n_4701)
);

O2A1O1Ixp33_ASAP7_75t_L g4702 ( 
.A1(n_4026),
.A2(n_3012),
.B(n_3059),
.C(n_3065),
.Y(n_4702)
);

NAND2xp5_ASAP7_75t_L g4703 ( 
.A(n_3176),
.B(n_3178),
.Y(n_4703)
);

BUFx2_ASAP7_75t_L g4704 ( 
.A(n_3870),
.Y(n_4704)
);

NAND2xp5_ASAP7_75t_SL g4705 ( 
.A(n_4067),
.B(n_4107),
.Y(n_4705)
);

CKINVDCx5p33_ASAP7_75t_R g4706 ( 
.A(n_3969),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_L g4707 ( 
.A(n_3178),
.B(n_3179),
.Y(n_4707)
);

INVx4_ASAP7_75t_L g4708 ( 
.A(n_3884),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_3388),
.Y(n_4709)
);

INVx1_ASAP7_75t_L g4710 ( 
.A(n_3388),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_3179),
.B(n_3180),
.Y(n_4711)
);

HB1xp67_ASAP7_75t_L g4712 ( 
.A(n_3111),
.Y(n_4712)
);

INVx2_ASAP7_75t_SL g4713 ( 
.A(n_4005),
.Y(n_4713)
);

HB1xp67_ASAP7_75t_L g4714 ( 
.A(n_3147),
.Y(n_4714)
);

NAND2xp5_ASAP7_75t_L g4715 ( 
.A(n_3180),
.B(n_3185),
.Y(n_4715)
);

AND3x1_ASAP7_75t_L g4716 ( 
.A(n_3059),
.B(n_3314),
.C(n_3189),
.Y(n_4716)
);

BUFx2_ASAP7_75t_L g4717 ( 
.A(n_3884),
.Y(n_4717)
);

INVx1_ASAP7_75t_L g4718 ( 
.A(n_3390),
.Y(n_4718)
);

CKINVDCx5p33_ASAP7_75t_R g4719 ( 
.A(n_3501),
.Y(n_4719)
);

NAND2xp5_ASAP7_75t_L g4720 ( 
.A(n_3185),
.B(n_3186),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_3390),
.Y(n_4721)
);

NAND2xp5_ASAP7_75t_L g4722 ( 
.A(n_3186),
.B(n_3187),
.Y(n_4722)
);

INVx1_ASAP7_75t_L g4723 ( 
.A(n_3397),
.Y(n_4723)
);

CKINVDCx20_ASAP7_75t_R g4724 ( 
.A(n_3133),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_SL g4725 ( 
.A(n_4107),
.B(n_3075),
.Y(n_4725)
);

NAND2xp5_ASAP7_75t_SL g4726 ( 
.A(n_3075),
.B(n_3026),
.Y(n_4726)
);

NAND3xp33_ASAP7_75t_SL g4727 ( 
.A(n_3221),
.B(n_3668),
.C(n_3157),
.Y(n_4727)
);

HB1xp67_ASAP7_75t_L g4728 ( 
.A(n_3147),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_L g4729 ( 
.A(n_3187),
.B(n_3188),
.Y(n_4729)
);

NAND2xp5_ASAP7_75t_L g4730 ( 
.A(n_3188),
.B(n_3193),
.Y(n_4730)
);

AND2x2_ASAP7_75t_L g4731 ( 
.A(n_3275),
.B(n_3289),
.Y(n_4731)
);

BUFx2_ASAP7_75t_L g4732 ( 
.A(n_3947),
.Y(n_4732)
);

AND2x4_ASAP7_75t_L g4733 ( 
.A(n_4027),
.B(n_4037),
.Y(n_4733)
);

NAND2xp5_ASAP7_75t_L g4734 ( 
.A(n_3193),
.B(n_3196),
.Y(n_4734)
);

CKINVDCx5p33_ASAP7_75t_R g4735 ( 
.A(n_3501),
.Y(n_4735)
);

INVx1_ASAP7_75t_L g4736 ( 
.A(n_3397),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_3441),
.Y(n_4737)
);

NOR2xp33_ASAP7_75t_L g4738 ( 
.A(n_3611),
.B(n_3676),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_3441),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_3458),
.Y(n_4740)
);

NAND2xp5_ASAP7_75t_L g4741 ( 
.A(n_3196),
.B(n_3203),
.Y(n_4741)
);

BUFx4f_ASAP7_75t_SL g4742 ( 
.A(n_3741),
.Y(n_4742)
);

NOR2xp33_ASAP7_75t_L g4743 ( 
.A(n_3686),
.B(n_3736),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_3458),
.Y(n_4744)
);

INVx1_ASAP7_75t_L g4745 ( 
.A(n_3358),
.Y(n_4745)
);

INVxp67_ASAP7_75t_SL g4746 ( 
.A(n_3017),
.Y(n_4746)
);

INVx5_ASAP7_75t_L g4747 ( 
.A(n_2975),
.Y(n_4747)
);

NOR2xp33_ASAP7_75t_L g4748 ( 
.A(n_3764),
.B(n_3844),
.Y(n_4748)
);

HB1xp67_ASAP7_75t_L g4749 ( 
.A(n_3218),
.Y(n_4749)
);

NAND2xp5_ASAP7_75t_L g4750 ( 
.A(n_3203),
.B(n_3205),
.Y(n_4750)
);

OAI21xp5_ASAP7_75t_L g4751 ( 
.A1(n_3668),
.A2(n_3662),
.B(n_3621),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_3358),
.Y(n_4752)
);

OR2x6_ASAP7_75t_L g4753 ( 
.A(n_3657),
.B(n_3659),
.Y(n_4753)
);

AND2x2_ASAP7_75t_L g4754 ( 
.A(n_3617),
.B(n_3630),
.Y(n_4754)
);

INVx4_ASAP7_75t_L g4755 ( 
.A(n_3947),
.Y(n_4755)
);

AND2x2_ASAP7_75t_L g4756 ( 
.A(n_3617),
.B(n_3630),
.Y(n_4756)
);

NOR2xp33_ASAP7_75t_SL g4757 ( 
.A(n_3097),
.B(n_3694),
.Y(n_4757)
);

NOR2x2_ASAP7_75t_L g4758 ( 
.A(n_3559),
.B(n_3302),
.Y(n_4758)
);

NAND2xp33_ASAP7_75t_L g4759 ( 
.A(n_3052),
.B(n_3724),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_3365),
.Y(n_4760)
);

CKINVDCx20_ASAP7_75t_R g4761 ( 
.A(n_3809),
.Y(n_4761)
);

INVx1_ASAP7_75t_SL g4762 ( 
.A(n_4133),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_3365),
.Y(n_4763)
);

NAND2xp5_ASAP7_75t_SL g4764 ( 
.A(n_2992),
.B(n_2988),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_3366),
.Y(n_4765)
);

NAND2xp5_ASAP7_75t_SL g4766 ( 
.A(n_2992),
.B(n_3097),
.Y(n_4766)
);

NOR2xp33_ASAP7_75t_L g4767 ( 
.A(n_3851),
.B(n_3876),
.Y(n_4767)
);

NOR2xp33_ASAP7_75t_L g4768 ( 
.A(n_3885),
.B(n_3896),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_3366),
.Y(n_4769)
);

NOR2xp33_ASAP7_75t_L g4770 ( 
.A(n_3908),
.B(n_3953),
.Y(n_4770)
);

OAI21x1_ASAP7_75t_L g4771 ( 
.A1(n_3307),
.A2(n_3322),
.B(n_3310),
.Y(n_4771)
);

BUFx8_ASAP7_75t_L g4772 ( 
.A(n_3659),
.Y(n_4772)
);

NAND2xp5_ASAP7_75t_L g4773 ( 
.A(n_3205),
.B(n_3208),
.Y(n_4773)
);

HB1xp67_ASAP7_75t_L g4774 ( 
.A(n_3218),
.Y(n_4774)
);

INVx1_ASAP7_75t_L g4775 ( 
.A(n_3370),
.Y(n_4775)
);

AND2x2_ASAP7_75t_L g4776 ( 
.A(n_3635),
.B(n_3648),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_3370),
.Y(n_4777)
);

NAND2xp5_ASAP7_75t_L g4778 ( 
.A(n_3208),
.B(n_3211),
.Y(n_4778)
);

OAI21xp5_ASAP7_75t_L g4779 ( 
.A1(n_3744),
.A2(n_3820),
.B(n_3782),
.Y(n_4779)
);

INVx1_ASAP7_75t_L g4780 ( 
.A(n_3386),
.Y(n_4780)
);

HB1xp67_ASAP7_75t_L g4781 ( 
.A(n_3251),
.Y(n_4781)
);

OR2x2_ASAP7_75t_L g4782 ( 
.A(n_3235),
.B(n_3272),
.Y(n_4782)
);

NAND2xp5_ASAP7_75t_L g4783 ( 
.A(n_3211),
.B(n_3125),
.Y(n_4783)
);

INVx1_ASAP7_75t_L g4784 ( 
.A(n_3386),
.Y(n_4784)
);

AND2x4_ASAP7_75t_L g4785 ( 
.A(n_4037),
.B(n_3755),
.Y(n_4785)
);

AOI22xp33_ASAP7_75t_L g4786 ( 
.A1(n_3138),
.A2(n_4004),
.B1(n_4059),
.B2(n_4003),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_L g4787 ( 
.A(n_3125),
.B(n_3126),
.Y(n_4787)
);

NAND2xp5_ASAP7_75t_L g4788 ( 
.A(n_3126),
.B(n_3135),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_L g4789 ( 
.A(n_3135),
.B(n_3051),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_3396),
.Y(n_4790)
);

NAND2xp5_ASAP7_75t_L g4791 ( 
.A(n_3051),
.B(n_3073),
.Y(n_4791)
);

AOI22xp33_ASAP7_75t_L g4792 ( 
.A1(n_3138),
.A2(n_4092),
.B1(n_4108),
.B2(n_4071),
.Y(n_4792)
);

INVx1_ASAP7_75t_SL g4793 ( 
.A(n_4133),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_3396),
.Y(n_4794)
);

INVx5_ASAP7_75t_L g4795 ( 
.A(n_3755),
.Y(n_4795)
);

AOI22xp5_ASAP7_75t_L g4796 ( 
.A1(n_3265),
.A2(n_3130),
.B1(n_4119),
.B2(n_4116),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_L g4797 ( 
.A(n_3073),
.B(n_3174),
.Y(n_4797)
);

AOI22x1_ASAP7_75t_L g4798 ( 
.A1(n_3086),
.A2(n_3087),
.B1(n_3098),
.B2(n_3095),
.Y(n_4798)
);

NAND2xp5_ASAP7_75t_SL g4799 ( 
.A(n_3097),
.B(n_3694),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_3403),
.Y(n_4800)
);

OR2x6_ASAP7_75t_L g4801 ( 
.A(n_3708),
.B(n_3747),
.Y(n_4801)
);

AND2x2_ASAP7_75t_L g4802 ( 
.A(n_3635),
.B(n_3648),
.Y(n_4802)
);

AND3x2_ASAP7_75t_SL g4803 ( 
.A(n_2984),
.B(n_3551),
.C(n_3132),
.Y(n_4803)
);

NAND2xp5_ASAP7_75t_L g4804 ( 
.A(n_3036),
.B(n_3152),
.Y(n_4804)
);

INVxp33_ASAP7_75t_L g4805 ( 
.A(n_3512),
.Y(n_4805)
);

INVx1_ASAP7_75t_L g4806 ( 
.A(n_3403),
.Y(n_4806)
);

NAND2xp5_ASAP7_75t_L g4807 ( 
.A(n_3036),
.B(n_3152),
.Y(n_4807)
);

NAND2xp5_ASAP7_75t_L g4808 ( 
.A(n_3069),
.B(n_3343),
.Y(n_4808)
);

INVx5_ASAP7_75t_L g4809 ( 
.A(n_3774),
.Y(n_4809)
);

NAND2xp5_ASAP7_75t_SL g4810 ( 
.A(n_3694),
.B(n_3909),
.Y(n_4810)
);

NOR2xp33_ASAP7_75t_L g4811 ( 
.A(n_3164),
.B(n_3226),
.Y(n_4811)
);

CKINVDCx5p33_ASAP7_75t_R g4812 ( 
.A(n_3501),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_3423),
.Y(n_4813)
);

NAND2xp5_ASAP7_75t_SL g4814 ( 
.A(n_3694),
.B(n_3909),
.Y(n_4814)
);

INVx4_ASAP7_75t_L g4815 ( 
.A(n_3973),
.Y(n_4815)
);

AND3x1_ASAP7_75t_SL g4816 ( 
.A(n_3052),
.B(n_3353),
.C(n_3254),
.Y(n_4816)
);

BUFx12f_ASAP7_75t_L g4817 ( 
.A(n_4077),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_L g4818 ( 
.A(n_3069),
.B(n_3343),
.Y(n_4818)
);

NAND2xp5_ASAP7_75t_L g4819 ( 
.A(n_3347),
.B(n_3666),
.Y(n_4819)
);

AOI22xp5_ASAP7_75t_L g4820 ( 
.A1(n_3106),
.A2(n_3107),
.B1(n_3132),
.B2(n_4124),
.Y(n_4820)
);

NAND2xp5_ASAP7_75t_L g4821 ( 
.A(n_3347),
.B(n_3666),
.Y(n_4821)
);

NAND2xp5_ASAP7_75t_L g4822 ( 
.A(n_3748),
.B(n_3873),
.Y(n_4822)
);

AOI22xp5_ASAP7_75t_L g4823 ( 
.A1(n_3106),
.A2(n_3107),
.B1(n_4124),
.B2(n_3873),
.Y(n_4823)
);

INVx1_ASAP7_75t_L g4824 ( 
.A(n_3410),
.Y(n_4824)
);

AOI22xp33_ASAP7_75t_L g4825 ( 
.A1(n_3056),
.A2(n_3114),
.B1(n_3262),
.B2(n_3748),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_3410),
.Y(n_4826)
);

HB1xp67_ASAP7_75t_L g4827 ( 
.A(n_3251),
.Y(n_4827)
);

NAND2xp5_ASAP7_75t_L g4828 ( 
.A(n_3910),
.B(n_3951),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_3412),
.Y(n_4829)
);

AND2x2_ASAP7_75t_L g4830 ( 
.A(n_3910),
.B(n_3951),
.Y(n_4830)
);

NOR2xp33_ASAP7_75t_L g4831 ( 
.A(n_3082),
.B(n_3128),
.Y(n_4831)
);

HB1xp67_ASAP7_75t_L g4832 ( 
.A(n_3255),
.Y(n_4832)
);

NAND2xp5_ASAP7_75t_L g4833 ( 
.A(n_3980),
.B(n_3999),
.Y(n_4833)
);

NAND2xp5_ASAP7_75t_SL g4834 ( 
.A(n_3909),
.B(n_3932),
.Y(n_4834)
);

NAND2xp5_ASAP7_75t_L g4835 ( 
.A(n_3980),
.B(n_3999),
.Y(n_4835)
);

CKINVDCx5p33_ASAP7_75t_R g4836 ( 
.A(n_3352),
.Y(n_4836)
);

CKINVDCx5p33_ASAP7_75t_R g4837 ( 
.A(n_3741),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_3412),
.Y(n_4838)
);

AND2x4_ASAP7_75t_L g4839 ( 
.A(n_4037),
.B(n_3774),
.Y(n_4839)
);

NOR3xp33_ASAP7_75t_L g4840 ( 
.A(n_3821),
.B(n_3916),
.C(n_3855),
.Y(n_4840)
);

NAND2xp5_ASAP7_75t_L g4841 ( 
.A(n_4088),
.B(n_3308),
.Y(n_4841)
);

INVxp67_ASAP7_75t_L g4842 ( 
.A(n_3092),
.Y(n_4842)
);

NAND2xp5_ASAP7_75t_L g4843 ( 
.A(n_4088),
.B(n_3308),
.Y(n_4843)
);

CKINVDCx20_ASAP7_75t_R g4844 ( 
.A(n_3809),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_3421),
.Y(n_4845)
);

HB1xp67_ASAP7_75t_L g4846 ( 
.A(n_3255),
.Y(n_4846)
);

AND2x2_ASAP7_75t_L g4847 ( 
.A(n_3457),
.B(n_3272),
.Y(n_4847)
);

OAI221xp5_ASAP7_75t_L g4848 ( 
.A1(n_3936),
.A2(n_3997),
.B1(n_4021),
.B2(n_4019),
.C(n_4018),
.Y(n_4848)
);

NAND2xp5_ASAP7_75t_SL g4849 ( 
.A(n_3909),
.B(n_3932),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_L g4850 ( 
.A(n_3121),
.B(n_3136),
.Y(n_4850)
);

HB1xp67_ASAP7_75t_L g4851 ( 
.A(n_3257),
.Y(n_4851)
);

NOR2xp33_ASAP7_75t_L g4852 ( 
.A(n_3082),
.B(n_3128),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_3421),
.Y(n_4853)
);

NAND2xp5_ASAP7_75t_SL g4854 ( 
.A(n_3932),
.B(n_3177),
.Y(n_4854)
);

AOI22xp33_ASAP7_75t_L g4855 ( 
.A1(n_3262),
.A2(n_3254),
.B1(n_3932),
.B2(n_2968),
.Y(n_4855)
);

NAND2xp5_ASAP7_75t_L g4856 ( 
.A(n_3139),
.B(n_3141),
.Y(n_4856)
);

HB1xp67_ASAP7_75t_L g4857 ( 
.A(n_3257),
.Y(n_4857)
);

AOI22xp33_ASAP7_75t_L g4858 ( 
.A1(n_2963),
.A2(n_2971),
.B1(n_2966),
.B2(n_2968),
.Y(n_4858)
);

NOR2xp33_ASAP7_75t_L g4859 ( 
.A(n_3085),
.B(n_3215),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_3424),
.Y(n_4860)
);

OAI22xp5_ASAP7_75t_L g4861 ( 
.A1(n_4045),
.A2(n_4060),
.B1(n_3085),
.B2(n_3198),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_3143),
.B(n_3148),
.Y(n_4862)
);

OAI221xp5_ASAP7_75t_L g4863 ( 
.A1(n_3161),
.A2(n_3168),
.B1(n_3166),
.B2(n_3153),
.C(n_3181),
.Y(n_4863)
);

INVxp67_ASAP7_75t_SL g4864 ( 
.A(n_3456),
.Y(n_4864)
);

OAI21xp5_ASAP7_75t_L g4865 ( 
.A1(n_3109),
.A2(n_3100),
.B(n_3204),
.Y(n_4865)
);

HB1xp67_ASAP7_75t_L g4866 ( 
.A(n_3258),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_3424),
.Y(n_4867)
);

CKINVDCx11_ASAP7_75t_R g4868 ( 
.A(n_3848),
.Y(n_4868)
);

NOR2xp33_ASAP7_75t_L g4869 ( 
.A(n_3270),
.B(n_3315),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_3428),
.Y(n_4870)
);

INVx1_ASAP7_75t_L g4871 ( 
.A(n_3428),
.Y(n_4871)
);

NAND2xp5_ASAP7_75t_SL g4872 ( 
.A(n_3177),
.B(n_4017),
.Y(n_4872)
);

NAND2xp5_ASAP7_75t_L g4873 ( 
.A(n_3242),
.B(n_2996),
.Y(n_4873)
);

CKINVDCx5p33_ASAP7_75t_R g4874 ( 
.A(n_3848),
.Y(n_4874)
);

NAND2xp5_ASAP7_75t_L g4875 ( 
.A(n_3242),
.B(n_2996),
.Y(n_4875)
);

OR2x2_ASAP7_75t_L g4876 ( 
.A(n_3607),
.B(n_3624),
.Y(n_4876)
);

NAND2xp5_ASAP7_75t_L g4877 ( 
.A(n_3607),
.B(n_3624),
.Y(n_4877)
);

NAND2xp5_ASAP7_75t_L g4878 ( 
.A(n_3640),
.B(n_3869),
.Y(n_4878)
);

BUFx2_ASAP7_75t_R g4879 ( 
.A(n_3014),
.Y(n_4879)
);

NAND2xp5_ASAP7_75t_L g4880 ( 
.A(n_3640),
.B(n_3869),
.Y(n_4880)
);

AND2x4_ASAP7_75t_L g4881 ( 
.A(n_4037),
.B(n_3774),
.Y(n_4881)
);

INVxp67_ASAP7_75t_L g4882 ( 
.A(n_3092),
.Y(n_4882)
);

NAND2xp5_ASAP7_75t_L g4883 ( 
.A(n_3929),
.B(n_2963),
.Y(n_4883)
);

NAND2xp5_ASAP7_75t_SL g4884 ( 
.A(n_4017),
.B(n_3420),
.Y(n_4884)
);

NAND2xp5_ASAP7_75t_L g4885 ( 
.A(n_3929),
.B(n_2966),
.Y(n_4885)
);

BUFx2_ASAP7_75t_L g4886 ( 
.A(n_3094),
.Y(n_4886)
);

NAND2xp5_ASAP7_75t_L g4887 ( 
.A(n_2971),
.B(n_2976),
.Y(n_4887)
);

BUFx2_ASAP7_75t_L g4888 ( 
.A(n_3094),
.Y(n_4888)
);

NAND2xp5_ASAP7_75t_L g4889 ( 
.A(n_2976),
.B(n_2977),
.Y(n_4889)
);

NOR2xp33_ASAP7_75t_R g4890 ( 
.A(n_3189),
.B(n_3314),
.Y(n_4890)
);

A2O1A1Ixp33_ASAP7_75t_L g4891 ( 
.A1(n_3237),
.A2(n_3103),
.B(n_3292),
.C(n_3151),
.Y(n_4891)
);

NOR2xp33_ASAP7_75t_L g4892 ( 
.A(n_3270),
.B(n_3315),
.Y(n_4892)
);

NAND2xp5_ASAP7_75t_L g4893 ( 
.A(n_2977),
.B(n_2989),
.Y(n_4893)
);

INVx5_ASAP7_75t_L g4894 ( 
.A(n_3774),
.Y(n_4894)
);

HB1xp67_ASAP7_75t_L g4895 ( 
.A(n_3258),
.Y(n_4895)
);

CKINVDCx11_ASAP7_75t_R g4896 ( 
.A(n_3848),
.Y(n_4896)
);

BUFx2_ASAP7_75t_L g4897 ( 
.A(n_3094),
.Y(n_4897)
);

NAND2xp5_ASAP7_75t_SL g4898 ( 
.A(n_3420),
.B(n_3293),
.Y(n_4898)
);

AND2x2_ASAP7_75t_SL g4899 ( 
.A(n_3867),
.B(n_3902),
.Y(n_4899)
);

HB1xp67_ASAP7_75t_L g4900 ( 
.A(n_3261),
.Y(n_4900)
);

OR2x6_ASAP7_75t_L g4901 ( 
.A(n_3747),
.B(n_3826),
.Y(n_4901)
);

NOR2xp67_ASAP7_75t_L g4902 ( 
.A(n_3047),
.B(n_3867),
.Y(n_4902)
);

NAND2xp5_ASAP7_75t_L g4903 ( 
.A(n_2989),
.B(n_2993),
.Y(n_4903)
);

NAND2xp5_ASAP7_75t_L g4904 ( 
.A(n_2993),
.B(n_2994),
.Y(n_4904)
);

AOI21xp5_ASAP7_75t_L g4905 ( 
.A1(n_2984),
.A2(n_3240),
.B(n_3047),
.Y(n_4905)
);

NAND2xp5_ASAP7_75t_L g4906 ( 
.A(n_2994),
.B(n_2998),
.Y(n_4906)
);

BUFx12f_ASAP7_75t_L g4907 ( 
.A(n_4077),
.Y(n_4907)
);

HB1xp67_ASAP7_75t_L g4908 ( 
.A(n_3261),
.Y(n_4908)
);

AOI22xp33_ASAP7_75t_L g4909 ( 
.A1(n_2998),
.A2(n_3011),
.B1(n_3592),
.B2(n_3010),
.Y(n_4909)
);

NOR2xp33_ASAP7_75t_L g4910 ( 
.A(n_3184),
.B(n_3191),
.Y(n_4910)
);

OR2x6_ASAP7_75t_L g4911 ( 
.A(n_3747),
.B(n_3826),
.Y(n_4911)
);

BUFx4f_ASAP7_75t_L g4912 ( 
.A(n_3302),
.Y(n_4912)
);

NAND2xp5_ASAP7_75t_L g4913 ( 
.A(n_3010),
.B(n_3011),
.Y(n_4913)
);

BUFx2_ASAP7_75t_SL g4914 ( 
.A(n_3401),
.Y(n_4914)
);

OR2x2_ASAP7_75t_SL g4915 ( 
.A(n_3826),
.B(n_3850),
.Y(n_4915)
);

BUFx2_ASAP7_75t_L g4916 ( 
.A(n_3647),
.Y(n_4916)
);

A2O1A1Ixp33_ASAP7_75t_L g4917 ( 
.A1(n_3237),
.A2(n_3151),
.B(n_3209),
.C(n_3224),
.Y(n_4917)
);

NAND2xp5_ASAP7_75t_L g4918 ( 
.A(n_3592),
.B(n_3593),
.Y(n_4918)
);

NAND2xp5_ASAP7_75t_L g4919 ( 
.A(n_3593),
.B(n_3595),
.Y(n_4919)
);

HB1xp67_ASAP7_75t_L g4920 ( 
.A(n_3263),
.Y(n_4920)
);

NOR2xp33_ASAP7_75t_L g4921 ( 
.A(n_3191),
.B(n_3198),
.Y(n_4921)
);

AOI22xp33_ASAP7_75t_L g4922 ( 
.A1(n_3595),
.A2(n_3604),
.B1(n_3610),
.B2(n_3608),
.Y(n_4922)
);

NAND2xp5_ASAP7_75t_L g4923 ( 
.A(n_3604),
.B(n_3608),
.Y(n_4923)
);

INVxp67_ASAP7_75t_SL g4924 ( 
.A(n_3456),
.Y(n_4924)
);

NOR2xp33_ASAP7_75t_L g4925 ( 
.A(n_3201),
.B(n_3202),
.Y(n_4925)
);

NAND2xp5_ASAP7_75t_L g4926 ( 
.A(n_3610),
.B(n_3613),
.Y(n_4926)
);

NAND2xp5_ASAP7_75t_L g4927 ( 
.A(n_3613),
.B(n_3618),
.Y(n_4927)
);

OR2x2_ASAP7_75t_L g4928 ( 
.A(n_3618),
.B(n_3627),
.Y(n_4928)
);

INVxp67_ASAP7_75t_SL g4929 ( 
.A(n_3401),
.Y(n_4929)
);

BUFx4f_ASAP7_75t_L g4930 ( 
.A(n_3302),
.Y(n_4930)
);

AOI22xp5_ASAP7_75t_L g4931 ( 
.A1(n_3627),
.A2(n_3638),
.B1(n_3639),
.B2(n_3633),
.Y(n_4931)
);

BUFx2_ASAP7_75t_L g4932 ( 
.A(n_3647),
.Y(n_4932)
);

O2A1O1Ixp33_ASAP7_75t_L g4933 ( 
.A1(n_3096),
.A2(n_3118),
.B(n_3123),
.C(n_3122),
.Y(n_4933)
);

BUFx2_ASAP7_75t_L g4934 ( 
.A(n_3647),
.Y(n_4934)
);

INVx1_ASAP7_75t_L g4935 ( 
.A(n_3400),
.Y(n_4935)
);

CKINVDCx5p33_ASAP7_75t_R g4936 ( 
.A(n_3928),
.Y(n_4936)
);

CKINVDCx5p33_ASAP7_75t_R g4937 ( 
.A(n_3928),
.Y(n_4937)
);

NOR2xp33_ASAP7_75t_L g4938 ( 
.A(n_3201),
.B(n_3202),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_3400),
.Y(n_4939)
);

OR2x2_ASAP7_75t_L g4940 ( 
.A(n_3633),
.B(n_3638),
.Y(n_4940)
);

NAND2xp5_ASAP7_75t_SL g4941 ( 
.A(n_3244),
.B(n_3345),
.Y(n_4941)
);

AND2x4_ASAP7_75t_L g4942 ( 
.A(n_3867),
.B(n_3902),
.Y(n_4942)
);

NAND2xp5_ASAP7_75t_L g4943 ( 
.A(n_3639),
.B(n_3641),
.Y(n_4943)
);

NOR2xp33_ASAP7_75t_L g4944 ( 
.A(n_3207),
.B(n_3212),
.Y(n_4944)
);

INVx4_ASAP7_75t_L g4945 ( 
.A(n_3902),
.Y(n_4945)
);

AOI22x1_ASAP7_75t_L g4946 ( 
.A1(n_3086),
.A2(n_3095),
.B1(n_3098),
.B2(n_3087),
.Y(n_4946)
);

INVx2_ASAP7_75t_SL g4947 ( 
.A(n_3214),
.Y(n_4947)
);

BUFx2_ASAP7_75t_L g4948 ( 
.A(n_3684),
.Y(n_4948)
);

NAND2xp5_ASAP7_75t_L g4949 ( 
.A(n_3641),
.B(n_3646),
.Y(n_4949)
);

OR2x2_ASAP7_75t_L g4950 ( 
.A(n_3646),
.B(n_3685),
.Y(n_4950)
);

NAND2xp5_ASAP7_75t_L g4951 ( 
.A(n_3685),
.B(n_3691),
.Y(n_4951)
);

NAND2xp5_ASAP7_75t_SL g4952 ( 
.A(n_3244),
.B(n_3502),
.Y(n_4952)
);

NAND2xp5_ASAP7_75t_L g4953 ( 
.A(n_3691),
.B(n_3692),
.Y(n_4953)
);

INVxp67_ASAP7_75t_SL g4954 ( 
.A(n_3336),
.Y(n_4954)
);

INVx5_ASAP7_75t_L g4955 ( 
.A(n_3913),
.Y(n_4955)
);

NAND2xp5_ASAP7_75t_L g4956 ( 
.A(n_3692),
.B(n_3703),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_3703),
.B(n_3710),
.Y(n_4957)
);

HB1xp67_ASAP7_75t_L g4958 ( 
.A(n_3263),
.Y(n_4958)
);

NOR2x1p5_ASAP7_75t_L g4959 ( 
.A(n_3913),
.B(n_4000),
.Y(n_4959)
);

NAND2xp5_ASAP7_75t_L g4960 ( 
.A(n_3710),
.B(n_3711),
.Y(n_4960)
);

BUFx4f_ASAP7_75t_L g4961 ( 
.A(n_3288),
.Y(n_4961)
);

BUFx2_ASAP7_75t_L g4962 ( 
.A(n_3684),
.Y(n_4962)
);

NAND2xp5_ASAP7_75t_SL g4963 ( 
.A(n_3502),
.B(n_3250),
.Y(n_4963)
);

CKINVDCx5p33_ASAP7_75t_R g4964 ( 
.A(n_3928),
.Y(n_4964)
);

BUFx4f_ASAP7_75t_L g4965 ( 
.A(n_3288),
.Y(n_4965)
);

NAND2xp5_ASAP7_75t_L g4966 ( 
.A(n_3711),
.B(n_3712),
.Y(n_4966)
);

NAND2xp5_ASAP7_75t_L g4967 ( 
.A(n_3712),
.B(n_3715),
.Y(n_4967)
);

AOI22xp33_ASAP7_75t_L g4968 ( 
.A1(n_3715),
.A2(n_3716),
.B1(n_3729),
.B2(n_3718),
.Y(n_4968)
);

NAND2xp5_ASAP7_75t_SL g4969 ( 
.A(n_3250),
.B(n_3247),
.Y(n_4969)
);

NAND2xp5_ASAP7_75t_L g4970 ( 
.A(n_3716),
.B(n_3718),
.Y(n_4970)
);

NAND2xp5_ASAP7_75t_L g4971 ( 
.A(n_3729),
.B(n_3731),
.Y(n_4971)
);

A2O1A1Ixp33_ASAP7_75t_L g4972 ( 
.A1(n_3222),
.A2(n_3161),
.B(n_3168),
.C(n_3247),
.Y(n_4972)
);

NAND2xp5_ASAP7_75t_L g4973 ( 
.A(n_3731),
.B(n_3733),
.Y(n_4973)
);

HB1xp67_ASAP7_75t_L g4974 ( 
.A(n_3268),
.Y(n_4974)
);

CKINVDCx5p33_ASAP7_75t_R g4975 ( 
.A(n_3788),
.Y(n_4975)
);

NAND2xp5_ASAP7_75t_L g4976 ( 
.A(n_3733),
.B(n_3738),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_L g4977 ( 
.A(n_3738),
.B(n_3753),
.Y(n_4977)
);

CKINVDCx14_ASAP7_75t_R g4978 ( 
.A(n_4077),
.Y(n_4978)
);

NOR2xp33_ASAP7_75t_L g4979 ( 
.A(n_3207),
.B(n_3212),
.Y(n_4979)
);

NAND2xp5_ASAP7_75t_L g4980 ( 
.A(n_3753),
.B(n_3757),
.Y(n_4980)
);

INVx3_ASAP7_75t_SL g4981 ( 
.A(n_3559),
.Y(n_4981)
);

OR2x6_ASAP7_75t_SL g4982 ( 
.A(n_3466),
.B(n_3449),
.Y(n_4982)
);

NOR2xp33_ASAP7_75t_L g4983 ( 
.A(n_3192),
.B(n_3229),
.Y(n_4983)
);

NAND2xp5_ASAP7_75t_L g4984 ( 
.A(n_3757),
.B(n_3758),
.Y(n_4984)
);

AOI22x1_ASAP7_75t_L g4985 ( 
.A1(n_3115),
.A2(n_3071),
.B1(n_3083),
.B2(n_3165),
.Y(n_4985)
);

HB1xp67_ASAP7_75t_L g4986 ( 
.A(n_3268),
.Y(n_4986)
);

HB1xp67_ASAP7_75t_L g4987 ( 
.A(n_3271),
.Y(n_4987)
);

OR2x2_ASAP7_75t_SL g4988 ( 
.A(n_3850),
.B(n_3859),
.Y(n_4988)
);

OR2x2_ASAP7_75t_L g4989 ( 
.A(n_3758),
.B(n_3760),
.Y(n_4989)
);

NAND2xp5_ASAP7_75t_L g4990 ( 
.A(n_3760),
.B(n_3767),
.Y(n_4990)
);

OR2x2_ASAP7_75t_L g4991 ( 
.A(n_3767),
.B(n_3775),
.Y(n_4991)
);

NAND2xp5_ASAP7_75t_SL g4992 ( 
.A(n_3321),
.B(n_3333),
.Y(n_4992)
);

BUFx12f_ASAP7_75t_L g4993 ( 
.A(n_4077),
.Y(n_4993)
);

NAND2xp5_ASAP7_75t_L g4994 ( 
.A(n_3775),
.B(n_3776),
.Y(n_4994)
);

INVxp67_ASAP7_75t_L g4995 ( 
.A(n_3684),
.Y(n_4995)
);

NOR2xp33_ASAP7_75t_L g4996 ( 
.A(n_3600),
.B(n_3609),
.Y(n_4996)
);

HB1xp67_ASAP7_75t_L g4997 ( 
.A(n_3271),
.Y(n_4997)
);

NAND2xp5_ASAP7_75t_L g4998 ( 
.A(n_3776),
.B(n_3796),
.Y(n_4998)
);

AOI22xp33_ASAP7_75t_L g4999 ( 
.A1(n_3796),
.A2(n_3798),
.B1(n_3817),
.B2(n_3799),
.Y(n_4999)
);

BUFx2_ASAP7_75t_L g5000 ( 
.A(n_3693),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_L g5001 ( 
.A(n_3798),
.B(n_3799),
.Y(n_5001)
);

INVxp67_ASAP7_75t_L g5002 ( 
.A(n_3693),
.Y(n_5002)
);

INVxp67_ASAP7_75t_L g5003 ( 
.A(n_3693),
.Y(n_5003)
);

AOI22xp5_ASAP7_75t_L g5004 ( 
.A1(n_3817),
.A2(n_3827),
.B1(n_3837),
.B2(n_3825),
.Y(n_5004)
);

NAND2xp5_ASAP7_75t_SL g5005 ( 
.A(n_3333),
.B(n_3306),
.Y(n_5005)
);

INVxp67_ASAP7_75t_L g5006 ( 
.A(n_3879),
.Y(n_5006)
);

INVxp67_ASAP7_75t_SL g5007 ( 
.A(n_3339),
.Y(n_5007)
);

AND3x1_ASAP7_75t_L g5008 ( 
.A(n_3316),
.B(n_3544),
.C(n_3569),
.Y(n_5008)
);

INVx4_ASAP7_75t_L g5009 ( 
.A(n_4000),
.Y(n_5009)
);

BUFx6f_ASAP7_75t_L g5010 ( 
.A(n_3214),
.Y(n_5010)
);

CKINVDCx20_ASAP7_75t_R g5011 ( 
.A(n_3303),
.Y(n_5011)
);

NAND2xp5_ASAP7_75t_L g5012 ( 
.A(n_3825),
.B(n_3827),
.Y(n_5012)
);

NAND2xp5_ASAP7_75t_L g5013 ( 
.A(n_3837),
.B(n_3847),
.Y(n_5013)
);

HB1xp67_ASAP7_75t_L g5014 ( 
.A(n_3277),
.Y(n_5014)
);

NAND2xp5_ASAP7_75t_SL g5015 ( 
.A(n_3312),
.B(n_3414),
.Y(n_5015)
);

BUFx2_ASAP7_75t_L g5016 ( 
.A(n_3879),
.Y(n_5016)
);

NAND2xp5_ASAP7_75t_L g5017 ( 
.A(n_3847),
.B(n_3854),
.Y(n_5017)
);

NAND2xp5_ASAP7_75t_L g5018 ( 
.A(n_3854),
.B(n_3862),
.Y(n_5018)
);

NAND2xp5_ASAP7_75t_L g5019 ( 
.A(n_3862),
.B(n_3864),
.Y(n_5019)
);

INVx2_ASAP7_75t_SL g5020 ( 
.A(n_3214),
.Y(n_5020)
);

BUFx2_ASAP7_75t_L g5021 ( 
.A(n_3879),
.Y(n_5021)
);

BUFx2_ASAP7_75t_L g5022 ( 
.A(n_3981),
.Y(n_5022)
);

AND2x4_ASAP7_75t_L g5023 ( 
.A(n_4111),
.B(n_3859),
.Y(n_5023)
);

BUFx6f_ASAP7_75t_L g5024 ( 
.A(n_3214),
.Y(n_5024)
);

A2O1A1Ixp33_ASAP7_75t_L g5025 ( 
.A1(n_3222),
.A2(n_3115),
.B(n_3155),
.C(n_3154),
.Y(n_5025)
);

CKINVDCx5p33_ASAP7_75t_R g5026 ( 
.A(n_3134),
.Y(n_5026)
);

NAND2xp5_ASAP7_75t_L g5027 ( 
.A(n_3864),
.B(n_3866),
.Y(n_5027)
);

NAND2xp5_ASAP7_75t_L g5028 ( 
.A(n_3866),
.B(n_3877),
.Y(n_5028)
);

CKINVDCx5p33_ASAP7_75t_R g5029 ( 
.A(n_3544),
.Y(n_5029)
);

NOR2xp33_ASAP7_75t_L g5030 ( 
.A(n_3679),
.B(n_3814),
.Y(n_5030)
);

BUFx6f_ASAP7_75t_L g5031 ( 
.A(n_3214),
.Y(n_5031)
);

NAND2xp5_ASAP7_75t_L g5032 ( 
.A(n_3877),
.B(n_3889),
.Y(n_5032)
);

AOI221xp5_ASAP7_75t_L g5033 ( 
.A1(n_3195),
.A2(n_3206),
.B1(n_3312),
.B2(n_3160),
.C(n_3163),
.Y(n_5033)
);

NAND2xp5_ASAP7_75t_L g5034 ( 
.A(n_3889),
.B(n_3898),
.Y(n_5034)
);

NAND2xp5_ASAP7_75t_L g5035 ( 
.A(n_3898),
.B(n_3906),
.Y(n_5035)
);

NAND2xp5_ASAP7_75t_L g5036 ( 
.A(n_3906),
.B(n_3907),
.Y(n_5036)
);

BUFx2_ASAP7_75t_L g5037 ( 
.A(n_3981),
.Y(n_5037)
);

BUFx4f_ASAP7_75t_L g5038 ( 
.A(n_3259),
.Y(n_5038)
);

NAND2xp5_ASAP7_75t_L g5039 ( 
.A(n_3907),
.B(n_3927),
.Y(n_5039)
);

INVxp33_ASAP7_75t_SL g5040 ( 
.A(n_3353),
.Y(n_5040)
);

AOI22xp5_ASAP7_75t_L g5041 ( 
.A1(n_3927),
.A2(n_3933),
.B1(n_3942),
.B2(n_3939),
.Y(n_5041)
);

CKINVDCx5p33_ASAP7_75t_R g5042 ( 
.A(n_3319),
.Y(n_5042)
);

NAND2xp5_ASAP7_75t_L g5043 ( 
.A(n_3933),
.B(n_3939),
.Y(n_5043)
);

AND3x1_ASAP7_75t_SL g5044 ( 
.A(n_3567),
.B(n_3568),
.C(n_3273),
.Y(n_5044)
);

INVx2_ASAP7_75t_SL g5045 ( 
.A(n_3259),
.Y(n_5045)
);

NAND2xp5_ASAP7_75t_L g5046 ( 
.A(n_3942),
.B(n_3945),
.Y(n_5046)
);

OR2x6_ASAP7_75t_L g5047 ( 
.A(n_3859),
.B(n_3905),
.Y(n_5047)
);

CKINVDCx5p33_ASAP7_75t_R g5048 ( 
.A(n_3338),
.Y(n_5048)
);

NAND2xp5_ASAP7_75t_SL g5049 ( 
.A(n_3414),
.B(n_3542),
.Y(n_5049)
);

AOI22xp33_ASAP7_75t_L g5050 ( 
.A1(n_3945),
.A2(n_3948),
.B1(n_3950),
.B2(n_3949),
.Y(n_5050)
);

NAND2xp5_ASAP7_75t_L g5051 ( 
.A(n_3948),
.B(n_3949),
.Y(n_5051)
);

INVx3_ASAP7_75t_L g5052 ( 
.A(n_3099),
.Y(n_5052)
);

OR2x2_ASAP7_75t_L g5053 ( 
.A(n_3950),
.B(n_3954),
.Y(n_5053)
);

BUFx2_ASAP7_75t_L g5054 ( 
.A(n_3981),
.Y(n_5054)
);

INVx2_ASAP7_75t_SL g5055 ( 
.A(n_3259),
.Y(n_5055)
);

BUFx2_ASAP7_75t_L g5056 ( 
.A(n_4011),
.Y(n_5056)
);

NAND2xp5_ASAP7_75t_L g5057 ( 
.A(n_3954),
.B(n_3956),
.Y(n_5057)
);

HB1xp67_ASAP7_75t_L g5058 ( 
.A(n_3277),
.Y(n_5058)
);

CKINVDCx5p33_ASAP7_75t_R g5059 ( 
.A(n_3373),
.Y(n_5059)
);

CKINVDCx5p33_ASAP7_75t_R g5060 ( 
.A(n_3377),
.Y(n_5060)
);

INVx1_ASAP7_75t_SL g5061 ( 
.A(n_4011),
.Y(n_5061)
);

BUFx4f_ASAP7_75t_L g5062 ( 
.A(n_3810),
.Y(n_5062)
);

AOI22xp33_ASAP7_75t_L g5063 ( 
.A1(n_3956),
.A2(n_3961),
.B1(n_3965),
.B2(n_3962),
.Y(n_5063)
);

NAND2xp5_ASAP7_75t_SL g5064 ( 
.A(n_3542),
.B(n_3961),
.Y(n_5064)
);

O2A1O1Ixp33_ASAP7_75t_L g5065 ( 
.A1(n_3117),
.A2(n_3071),
.B(n_3083),
.C(n_3227),
.Y(n_5065)
);

HB1xp67_ASAP7_75t_L g5066 ( 
.A(n_3278),
.Y(n_5066)
);

CKINVDCx5p33_ASAP7_75t_R g5067 ( 
.A(n_3379),
.Y(n_5067)
);

INVx1_ASAP7_75t_SL g5068 ( 
.A(n_4016),
.Y(n_5068)
);

OAI22xp5_ASAP7_75t_L g5069 ( 
.A1(n_3962),
.A2(n_3968),
.B1(n_3971),
.B2(n_3965),
.Y(n_5069)
);

NAND2xp5_ASAP7_75t_L g5070 ( 
.A(n_3968),
.B(n_3971),
.Y(n_5070)
);

HB1xp67_ASAP7_75t_L g5071 ( 
.A(n_3278),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_L g5072 ( 
.A(n_3974),
.B(n_3983),
.Y(n_5072)
);

BUFx6f_ASAP7_75t_L g5073 ( 
.A(n_3099),
.Y(n_5073)
);

BUFx2_ASAP7_75t_SL g5074 ( 
.A(n_4111),
.Y(n_5074)
);

NAND2xp5_ASAP7_75t_L g5075 ( 
.A(n_3974),
.B(n_3983),
.Y(n_5075)
);

AOI22xp33_ASAP7_75t_L g5076 ( 
.A1(n_3986),
.A2(n_3995),
.B1(n_4007),
.B2(n_4006),
.Y(n_5076)
);

BUFx12f_ASAP7_75t_L g5077 ( 
.A(n_3572),
.Y(n_5077)
);

NAND2xp5_ASAP7_75t_SL g5078 ( 
.A(n_3986),
.B(n_3995),
.Y(n_5078)
);

A2O1A1Ixp33_ASAP7_75t_L g5079 ( 
.A1(n_3154),
.A2(n_3160),
.B(n_3163),
.C(n_3155),
.Y(n_5079)
);

NAND2xp5_ASAP7_75t_L g5080 ( 
.A(n_4006),
.B(n_4007),
.Y(n_5080)
);

NAND2xp5_ASAP7_75t_L g5081 ( 
.A(n_4024),
.B(n_4032),
.Y(n_5081)
);

NAND2xp5_ASAP7_75t_L g5082 ( 
.A(n_4024),
.B(n_4032),
.Y(n_5082)
);

OR2x2_ASAP7_75t_L g5083 ( 
.A(n_4034),
.B(n_4040),
.Y(n_5083)
);

AND2x4_ASAP7_75t_L g5084 ( 
.A(n_4111),
.B(n_3859),
.Y(n_5084)
);

AOI22xp33_ASAP7_75t_L g5085 ( 
.A1(n_4034),
.A2(n_4040),
.B1(n_4051),
.B2(n_4043),
.Y(n_5085)
);

NOR2xp67_ASAP7_75t_L g5086 ( 
.A(n_4111),
.B(n_3524),
.Y(n_5086)
);

NAND2xp5_ASAP7_75t_L g5087 ( 
.A(n_4043),
.B(n_4051),
.Y(n_5087)
);

NAND2xp5_ASAP7_75t_L g5088 ( 
.A(n_4057),
.B(n_4058),
.Y(n_5088)
);

NAND2xp5_ASAP7_75t_L g5089 ( 
.A(n_4057),
.B(n_4058),
.Y(n_5089)
);

NAND2xp5_ASAP7_75t_L g5090 ( 
.A(n_4083),
.B(n_4091),
.Y(n_5090)
);

INVx3_ASAP7_75t_L g5091 ( 
.A(n_3099),
.Y(n_5091)
);

NAND2xp5_ASAP7_75t_L g5092 ( 
.A(n_4083),
.B(n_4091),
.Y(n_5092)
);

AND3x1_ASAP7_75t_SL g5093 ( 
.A(n_3567),
.B(n_3568),
.C(n_3606),
.Y(n_5093)
);

NAND2xp5_ASAP7_75t_L g5094 ( 
.A(n_4094),
.B(n_4096),
.Y(n_5094)
);

AND2x4_ASAP7_75t_L g5095 ( 
.A(n_3905),
.B(n_3912),
.Y(n_5095)
);

CKINVDCx8_ASAP7_75t_R g5096 ( 
.A(n_3905),
.Y(n_5096)
);

NOR2xp33_ASAP7_75t_L g5097 ( 
.A(n_3856),
.B(n_4031),
.Y(n_5097)
);

NOR2xp33_ASAP7_75t_L g5098 ( 
.A(n_3093),
.B(n_3101),
.Y(n_5098)
);

AOI22xp5_ASAP7_75t_L g5099 ( 
.A1(n_4094),
.A2(n_4096),
.B1(n_4098),
.B2(n_4097),
.Y(n_5099)
);

NAND2xp5_ASAP7_75t_L g5100 ( 
.A(n_4097),
.B(n_4098),
.Y(n_5100)
);

AOI22xp5_ASAP7_75t_L g5101 ( 
.A1(n_4100),
.A2(n_4103),
.B1(n_4123),
.B2(n_4109),
.Y(n_5101)
);

BUFx6f_ASAP7_75t_L g5102 ( 
.A(n_3099),
.Y(n_5102)
);

NAND2xp5_ASAP7_75t_L g5103 ( 
.A(n_4100),
.B(n_4103),
.Y(n_5103)
);

NAND2xp5_ASAP7_75t_SL g5104 ( 
.A(n_4109),
.B(n_4123),
.Y(n_5104)
);

INVx2_ASAP7_75t_SL g5105 ( 
.A(n_5010),
.Y(n_5105)
);

BUFx8_ASAP7_75t_L g5106 ( 
.A(n_5073),
.Y(n_5106)
);

BUFx3_ASAP7_75t_L g5107 ( 
.A(n_4151),
.Y(n_5107)
);

OAI22xp5_ASAP7_75t_L g5108 ( 
.A1(n_4307),
.A2(n_4129),
.B1(n_4141),
.B2(n_4128),
.Y(n_5108)
);

HB1xp67_ASAP7_75t_L g5109 ( 
.A(n_4271),
.Y(n_5109)
);

OAI22xp5_ASAP7_75t_L g5110 ( 
.A1(n_4307),
.A2(n_4129),
.B1(n_4141),
.B2(n_4128),
.Y(n_5110)
);

AOI22xp33_ASAP7_75t_L g5111 ( 
.A1(n_4155),
.A2(n_3419),
.B1(n_3301),
.B2(n_3286),
.Y(n_5111)
);

AND2x4_ASAP7_75t_L g5112 ( 
.A(n_4222),
.B(n_3905),
.Y(n_5112)
);

INVx1_ASAP7_75t_L g5113 ( 
.A(n_4266),
.Y(n_5113)
);

INVx2_ASAP7_75t_L g5114 ( 
.A(n_4163),
.Y(n_5114)
);

BUFx6f_ASAP7_75t_L g5115 ( 
.A(n_4152),
.Y(n_5115)
);

AOI21xp5_ASAP7_75t_L g5116 ( 
.A1(n_4216),
.A2(n_3245),
.B(n_3240),
.Y(n_5116)
);

INVx3_ASAP7_75t_L g5117 ( 
.A(n_4152),
.Y(n_5117)
);

BUFx4f_ASAP7_75t_L g5118 ( 
.A(n_4537),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_4266),
.Y(n_5119)
);

OAI21xp33_ASAP7_75t_L g5120 ( 
.A1(n_4315),
.A2(n_3104),
.B(n_3102),
.Y(n_5120)
);

INVx2_ASAP7_75t_L g5121 ( 
.A(n_4163),
.Y(n_5121)
);

O2A1O1Ixp33_ASAP7_75t_L g5122 ( 
.A1(n_4149),
.A2(n_3269),
.B(n_3248),
.C(n_3120),
.Y(n_5122)
);

AOI21xp5_ASAP7_75t_L g5123 ( 
.A1(n_4216),
.A2(n_3245),
.B(n_3328),
.Y(n_5123)
);

AOI22xp33_ASAP7_75t_L g5124 ( 
.A1(n_4155),
.A2(n_3286),
.B1(n_3031),
.B2(n_3028),
.Y(n_5124)
);

BUFx2_ASAP7_75t_L g5125 ( 
.A(n_4151),
.Y(n_5125)
);

INVx1_ASAP7_75t_L g5126 ( 
.A(n_4266),
.Y(n_5126)
);

BUFx8_ASAP7_75t_L g5127 ( 
.A(n_5073),
.Y(n_5127)
);

BUFx3_ASAP7_75t_L g5128 ( 
.A(n_4151),
.Y(n_5128)
);

BUFx6f_ASAP7_75t_L g5129 ( 
.A(n_4152),
.Y(n_5129)
);

INVx1_ASAP7_75t_L g5130 ( 
.A(n_4272),
.Y(n_5130)
);

NAND2xp5_ASAP7_75t_L g5131 ( 
.A(n_4567),
.B(n_3354),
.Y(n_5131)
);

NAND2xp5_ASAP7_75t_SL g5132 ( 
.A(n_4311),
.B(n_3558),
.Y(n_5132)
);

AOI222xp33_ASAP7_75t_L g5133 ( 
.A1(n_4293),
.A2(n_3316),
.B1(n_3028),
.B2(n_3031),
.C1(n_3606),
.C2(n_3105),
.Y(n_5133)
);

A2O1A1Ixp33_ASAP7_75t_L g5134 ( 
.A1(n_4280),
.A2(n_3558),
.B(n_3183),
.C(n_3276),
.Y(n_5134)
);

BUFx6f_ASAP7_75t_L g5135 ( 
.A(n_4152),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_4272),
.Y(n_5136)
);

INVx3_ASAP7_75t_L g5137 ( 
.A(n_4152),
.Y(n_5137)
);

INVx5_ASAP7_75t_L g5138 ( 
.A(n_4195),
.Y(n_5138)
);

NAND2xp5_ASAP7_75t_L g5139 ( 
.A(n_4567),
.B(n_3354),
.Y(n_5139)
);

BUFx6f_ASAP7_75t_L g5140 ( 
.A(n_4152),
.Y(n_5140)
);

AOI22xp5_ASAP7_75t_L g5141 ( 
.A1(n_4155),
.A2(n_3440),
.B1(n_3433),
.B2(n_3074),
.Y(n_5141)
);

NAND2xp5_ASAP7_75t_L g5142 ( 
.A(n_4684),
.B(n_3279),
.Y(n_5142)
);

OAI22xp5_ASAP7_75t_L g5143 ( 
.A1(n_4311),
.A2(n_3066),
.B1(n_3140),
.B2(n_3000),
.Y(n_5143)
);

AND2x4_ASAP7_75t_L g5144 ( 
.A(n_4222),
.B(n_3905),
.Y(n_5144)
);

AOI22xp5_ASAP7_75t_L g5145 ( 
.A1(n_4155),
.A2(n_3440),
.B1(n_3433),
.B2(n_3183),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_4272),
.Y(n_5146)
);

A2O1A1Ixp33_ASAP7_75t_L g5147 ( 
.A1(n_4280),
.A2(n_3276),
.B(n_3415),
.C(n_3548),
.Y(n_5147)
);

INVx2_ASAP7_75t_SL g5148 ( 
.A(n_5010),
.Y(n_5148)
);

BUFx6f_ASAP7_75t_L g5149 ( 
.A(n_4152),
.Y(n_5149)
);

INVx5_ASAP7_75t_L g5150 ( 
.A(n_4195),
.Y(n_5150)
);

AOI22xp33_ASAP7_75t_L g5151 ( 
.A1(n_4155),
.A2(n_3461),
.B1(n_3463),
.B2(n_3459),
.Y(n_5151)
);

INVx1_ASAP7_75t_SL g5152 ( 
.A(n_4279),
.Y(n_5152)
);

BUFx6f_ASAP7_75t_L g5153 ( 
.A(n_4152),
.Y(n_5153)
);

INVx2_ASAP7_75t_L g5154 ( 
.A(n_4163),
.Y(n_5154)
);

BUFx6f_ASAP7_75t_L g5155 ( 
.A(n_4152),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_4273),
.Y(n_5156)
);

CKINVDCx5p33_ASAP7_75t_R g5157 ( 
.A(n_4519),
.Y(n_5157)
);

NAND2x2_ASAP7_75t_L g5158 ( 
.A(n_4636),
.B(n_4016),
.Y(n_5158)
);

NAND2xp5_ASAP7_75t_L g5159 ( 
.A(n_4684),
.B(n_3279),
.Y(n_5159)
);

AND2x4_ASAP7_75t_L g5160 ( 
.A(n_4222),
.B(n_3912),
.Y(n_5160)
);

INVx1_ASAP7_75t_SL g5161 ( 
.A(n_4279),
.Y(n_5161)
);

AOI21xp5_ASAP7_75t_L g5162 ( 
.A1(n_4148),
.A2(n_3332),
.B(n_3331),
.Y(n_5162)
);

INVxp67_ASAP7_75t_SL g5163 ( 
.A(n_4954),
.Y(n_5163)
);

NAND2xp33_ASAP7_75t_L g5164 ( 
.A(n_4322),
.B(n_3453),
.Y(n_5164)
);

NOR2xp33_ASAP7_75t_L g5165 ( 
.A(n_4322),
.B(n_4101),
.Y(n_5165)
);

BUFx2_ASAP7_75t_L g5166 ( 
.A(n_4210),
.Y(n_5166)
);

NAND2xp5_ASAP7_75t_L g5167 ( 
.A(n_4685),
.B(n_3281),
.Y(n_5167)
);

NAND2xp5_ASAP7_75t_SL g5168 ( 
.A(n_4179),
.B(n_3520),
.Y(n_5168)
);

BUFx6f_ASAP7_75t_L g5169 ( 
.A(n_4158),
.Y(n_5169)
);

NOR2xp33_ASAP7_75t_L g5170 ( 
.A(n_4191),
.B(n_4201),
.Y(n_5170)
);

AND2x2_ASAP7_75t_L g5171 ( 
.A(n_4701),
.B(n_3912),
.Y(n_5171)
);

AOI22xp33_ASAP7_75t_SL g5172 ( 
.A1(n_4343),
.A2(n_3459),
.B1(n_3553),
.B2(n_3912),
.Y(n_5172)
);

BUFx6f_ASAP7_75t_L g5173 ( 
.A(n_4158),
.Y(n_5173)
);

AND2x4_ASAP7_75t_L g5174 ( 
.A(n_4222),
.B(n_5052),
.Y(n_5174)
);

AO22x1_ASAP7_75t_L g5175 ( 
.A1(n_4869),
.A2(n_3553),
.B1(n_3466),
.B2(n_3564),
.Y(n_5175)
);

INVxp67_ASAP7_75t_L g5176 ( 
.A(n_4914),
.Y(n_5176)
);

AOI21xp5_ASAP7_75t_L g5177 ( 
.A1(n_4148),
.A2(n_3478),
.B(n_3468),
.Y(n_5177)
);

NAND2xp5_ASAP7_75t_L g5178 ( 
.A(n_4685),
.B(n_3281),
.Y(n_5178)
);

INVx1_ASAP7_75t_L g5179 ( 
.A(n_4273),
.Y(n_5179)
);

OAI22xp5_ASAP7_75t_L g5180 ( 
.A1(n_4293),
.A2(n_3295),
.B1(n_3584),
.B2(n_3274),
.Y(n_5180)
);

NAND2xp5_ASAP7_75t_L g5181 ( 
.A(n_4700),
.B(n_3287),
.Y(n_5181)
);

BUFx3_ASAP7_75t_L g5182 ( 
.A(n_4210),
.Y(n_5182)
);

BUFx2_ASAP7_75t_L g5183 ( 
.A(n_4210),
.Y(n_5183)
);

AOI21xp5_ASAP7_75t_L g5184 ( 
.A1(n_4176),
.A2(n_3478),
.B(n_3468),
.Y(n_5184)
);

INVx2_ASAP7_75t_SL g5185 ( 
.A(n_5010),
.Y(n_5185)
);

AOI221xp5_ASAP7_75t_L g5186 ( 
.A1(n_4185),
.A2(n_3395),
.B1(n_3248),
.B2(n_3389),
.C(n_3236),
.Y(n_5186)
);

INVx6_ASAP7_75t_L g5187 ( 
.A(n_4772),
.Y(n_5187)
);

BUFx8_ASAP7_75t_L g5188 ( 
.A(n_5073),
.Y(n_5188)
);

INVx1_ASAP7_75t_L g5189 ( 
.A(n_4273),
.Y(n_5189)
);

INVx1_ASAP7_75t_L g5190 ( 
.A(n_4277),
.Y(n_5190)
);

INVx2_ASAP7_75t_L g5191 ( 
.A(n_4163),
.Y(n_5191)
);

NAND2xp5_ASAP7_75t_L g5192 ( 
.A(n_4700),
.B(n_3287),
.Y(n_5192)
);

INVxp67_ASAP7_75t_L g5193 ( 
.A(n_4914),
.Y(n_5193)
);

INVx1_ASAP7_75t_L g5194 ( 
.A(n_4277),
.Y(n_5194)
);

INVx2_ASAP7_75t_L g5195 ( 
.A(n_4165),
.Y(n_5195)
);

BUFx3_ASAP7_75t_L g5196 ( 
.A(n_4254),
.Y(n_5196)
);

OAI22xp5_ASAP7_75t_L g5197 ( 
.A1(n_4291),
.A2(n_4395),
.B1(n_4357),
.B2(n_4353),
.Y(n_5197)
);

INVx8_ASAP7_75t_L g5198 ( 
.A(n_4537),
.Y(n_5198)
);

BUFx2_ASAP7_75t_L g5199 ( 
.A(n_4254),
.Y(n_5199)
);

BUFx3_ASAP7_75t_L g5200 ( 
.A(n_4254),
.Y(n_5200)
);

NAND2xp5_ASAP7_75t_L g5201 ( 
.A(n_4703),
.B(n_3296),
.Y(n_5201)
);

OAI22xp5_ASAP7_75t_L g5202 ( 
.A1(n_4291),
.A2(n_3626),
.B1(n_3645),
.B2(n_3614),
.Y(n_5202)
);

A2O1A1Ixp33_ASAP7_75t_L g5203 ( 
.A1(n_4149),
.A2(n_3552),
.B(n_3564),
.C(n_3364),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_4277),
.Y(n_5204)
);

OR2x2_ASAP7_75t_L g5205 ( 
.A(n_4661),
.B(n_4101),
.Y(n_5205)
);

BUFx6f_ASAP7_75t_L g5206 ( 
.A(n_4158),
.Y(n_5206)
);

AOI21xp5_ASAP7_75t_L g5207 ( 
.A1(n_4176),
.A2(n_3516),
.B(n_3508),
.Y(n_5207)
);

OAI22xp5_ASAP7_75t_L g5208 ( 
.A1(n_4395),
.A2(n_3762),
.B1(n_3872),
.B2(n_3670),
.Y(n_5208)
);

BUFx2_ASAP7_75t_L g5209 ( 
.A(n_4257),
.Y(n_5209)
);

INVx2_ASAP7_75t_L g5210 ( 
.A(n_4165),
.Y(n_5210)
);

INVx3_ASAP7_75t_L g5211 ( 
.A(n_4158),
.Y(n_5211)
);

NOR2xp33_ASAP7_75t_L g5212 ( 
.A(n_4191),
.B(n_4101),
.Y(n_5212)
);

OR2x2_ASAP7_75t_L g5213 ( 
.A(n_4661),
.B(n_3899),
.Y(n_5213)
);

INVx1_ASAP7_75t_L g5214 ( 
.A(n_4284),
.Y(n_5214)
);

BUFx6f_ASAP7_75t_L g5215 ( 
.A(n_4158),
.Y(n_5215)
);

AO22x1_ASAP7_75t_L g5216 ( 
.A1(n_4869),
.A2(n_3553),
.B1(n_3564),
.B2(n_3449),
.Y(n_5216)
);

INVx1_ASAP7_75t_SL g5217 ( 
.A(n_4305),
.Y(n_5217)
);

INVx2_ASAP7_75t_L g5218 ( 
.A(n_4165),
.Y(n_5218)
);

INVx3_ASAP7_75t_L g5219 ( 
.A(n_4158),
.Y(n_5219)
);

NAND2xp5_ASAP7_75t_SL g5220 ( 
.A(n_4179),
.B(n_3553),
.Y(n_5220)
);

NOR2xp33_ASAP7_75t_SL g5221 ( 
.A(n_4343),
.B(n_3515),
.Y(n_5221)
);

BUFx4f_ASAP7_75t_SL g5222 ( 
.A(n_4205),
.Y(n_5222)
);

OAI22xp33_ASAP7_75t_L g5223 ( 
.A1(n_4184),
.A2(n_3404),
.B1(n_3425),
.B2(n_3363),
.Y(n_5223)
);

NAND2xp5_ASAP7_75t_L g5224 ( 
.A(n_4703),
.B(n_3296),
.Y(n_5224)
);

INVx3_ASAP7_75t_L g5225 ( 
.A(n_4158),
.Y(n_5225)
);

OAI22xp5_ASAP7_75t_L g5226 ( 
.A1(n_4357),
.A2(n_3925),
.B1(n_3957),
.B2(n_3919),
.Y(n_5226)
);

BUFx2_ASAP7_75t_L g5227 ( 
.A(n_4257),
.Y(n_5227)
);

INVx2_ASAP7_75t_L g5228 ( 
.A(n_4165),
.Y(n_5228)
);

CKINVDCx20_ASAP7_75t_R g5229 ( 
.A(n_4205),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_4284),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_L g5231 ( 
.A(n_4707),
.B(n_3297),
.Y(n_5231)
);

INVx3_ASAP7_75t_L g5232 ( 
.A(n_4158),
.Y(n_5232)
);

NAND2xp5_ASAP7_75t_L g5233 ( 
.A(n_4707),
.B(n_3297),
.Y(n_5233)
);

AOI22xp33_ASAP7_75t_SL g5234 ( 
.A1(n_4323),
.A2(n_3553),
.B1(n_4020),
.B2(n_3912),
.Y(n_5234)
);

AOI22xp33_ASAP7_75t_SL g5235 ( 
.A1(n_4323),
.A2(n_3553),
.B1(n_4020),
.B2(n_3912),
.Y(n_5235)
);

OR2x2_ASAP7_75t_L g5236 ( 
.A(n_4712),
.B(n_3990),
.Y(n_5236)
);

OAI21xp5_ASAP7_75t_L g5237 ( 
.A1(n_4315),
.A2(n_3213),
.B(n_3329),
.Y(n_5237)
);

NAND2xp5_ASAP7_75t_L g5238 ( 
.A(n_4711),
.B(n_4715),
.Y(n_5238)
);

NAND2xp5_ASAP7_75t_L g5239 ( 
.A(n_4711),
.B(n_3298),
.Y(n_5239)
);

INVx2_ASAP7_75t_L g5240 ( 
.A(n_4166),
.Y(n_5240)
);

INVx2_ASAP7_75t_L g5241 ( 
.A(n_4166),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_4284),
.Y(n_5242)
);

INVx1_ASAP7_75t_SL g5243 ( 
.A(n_4305),
.Y(n_5243)
);

A2O1A1Ixp33_ASAP7_75t_L g5244 ( 
.A1(n_4917),
.A2(n_3565),
.B(n_3426),
.C(n_3562),
.Y(n_5244)
);

AND2x2_ASAP7_75t_L g5245 ( 
.A(n_4701),
.B(n_4020),
.Y(n_5245)
);

BUFx2_ASAP7_75t_L g5246 ( 
.A(n_4283),
.Y(n_5246)
);

O2A1O1Ixp33_ASAP7_75t_L g5247 ( 
.A1(n_4759),
.A2(n_4702),
.B(n_4353),
.C(n_4425),
.Y(n_5247)
);

NOR2xp33_ASAP7_75t_L g5248 ( 
.A(n_4201),
.B(n_3252),
.Y(n_5248)
);

NOR2xp33_ASAP7_75t_L g5249 ( 
.A(n_4245),
.B(n_4049),
.Y(n_5249)
);

INVx3_ASAP7_75t_L g5250 ( 
.A(n_4198),
.Y(n_5250)
);

HB1xp67_ASAP7_75t_L g5251 ( 
.A(n_4271),
.Y(n_5251)
);

INVx1_ASAP7_75t_L g5252 ( 
.A(n_4289),
.Y(n_5252)
);

NOR2xp33_ASAP7_75t_L g5253 ( 
.A(n_4245),
.B(n_3413),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_4289),
.Y(n_5254)
);

A2O1A1Ixp33_ASAP7_75t_L g5255 ( 
.A1(n_4917),
.A2(n_3565),
.B(n_3562),
.C(n_3429),
.Y(n_5255)
);

INVx1_ASAP7_75t_L g5256 ( 
.A(n_4289),
.Y(n_5256)
);

AOI222xp33_ASAP7_75t_L g5257 ( 
.A1(n_4162),
.A2(n_3463),
.B1(n_3461),
.B2(n_3351),
.C1(n_3298),
.C2(n_3299),
.Y(n_5257)
);

INVx1_ASAP7_75t_L g5258 ( 
.A(n_4296),
.Y(n_5258)
);

BUFx6f_ASAP7_75t_L g5259 ( 
.A(n_4198),
.Y(n_5259)
);

AOI21xp5_ASAP7_75t_L g5260 ( 
.A1(n_4217),
.A2(n_3516),
.B(n_3508),
.Y(n_5260)
);

INVx1_ASAP7_75t_L g5261 ( 
.A(n_4296),
.Y(n_5261)
);

CKINVDCx5p33_ASAP7_75t_R g5262 ( 
.A(n_4519),
.Y(n_5262)
);

INVx1_ASAP7_75t_L g5263 ( 
.A(n_4296),
.Y(n_5263)
);

OR2x6_ASAP7_75t_L g5264 ( 
.A(n_4160),
.B(n_4020),
.Y(n_5264)
);

AOI21xp5_ASAP7_75t_L g5265 ( 
.A1(n_4217),
.A2(n_3530),
.B(n_3524),
.Y(n_5265)
);

BUFx2_ASAP7_75t_L g5266 ( 
.A(n_4298),
.Y(n_5266)
);

NAND2xp5_ASAP7_75t_L g5267 ( 
.A(n_4715),
.B(n_3299),
.Y(n_5267)
);

INVx1_ASAP7_75t_L g5268 ( 
.A(n_4306),
.Y(n_5268)
);

O2A1O1Ixp33_ASAP7_75t_L g5269 ( 
.A1(n_4759),
.A2(n_3409),
.B(n_3402),
.C(n_3376),
.Y(n_5269)
);

NAND2xp5_ASAP7_75t_SL g5270 ( 
.A(n_4200),
.B(n_4248),
.Y(n_5270)
);

O2A1O1Ixp5_ASAP7_75t_L g5271 ( 
.A1(n_4255),
.A2(n_3395),
.B(n_3230),
.C(n_3238),
.Y(n_5271)
);

NAND2xp5_ASAP7_75t_L g5272 ( 
.A(n_4720),
.B(n_3346),
.Y(n_5272)
);

NAND2xp5_ASAP7_75t_L g5273 ( 
.A(n_4720),
.B(n_3348),
.Y(n_5273)
);

BUFx2_ASAP7_75t_L g5274 ( 
.A(n_4298),
.Y(n_5274)
);

NOR2xp33_ASAP7_75t_L g5275 ( 
.A(n_4248),
.B(n_3413),
.Y(n_5275)
);

AND2x4_ASAP7_75t_L g5276 ( 
.A(n_4222),
.B(n_4020),
.Y(n_5276)
);

AOI21xp5_ASAP7_75t_L g5277 ( 
.A1(n_4219),
.A2(n_3541),
.B(n_3530),
.Y(n_5277)
);

A2O1A1Ixp33_ASAP7_75t_L g5278 ( 
.A1(n_4270),
.A2(n_3442),
.B(n_3479),
.C(n_3497),
.Y(n_5278)
);

AND2x2_ASAP7_75t_L g5279 ( 
.A(n_4701),
.B(n_4020),
.Y(n_5279)
);

NAND2xp5_ASAP7_75t_L g5280 ( 
.A(n_4722),
.B(n_3349),
.Y(n_5280)
);

AND2x2_ASAP7_75t_SL g5281 ( 
.A(n_4316),
.B(n_4074),
.Y(n_5281)
);

NOR2x1p5_ASAP7_75t_SL g5282 ( 
.A(n_4281),
.B(n_3231),
.Y(n_5282)
);

NOR2x1_ASAP7_75t_L g5283 ( 
.A(n_4850),
.B(n_3171),
.Y(n_5283)
);

INVx3_ASAP7_75t_L g5284 ( 
.A(n_4198),
.Y(n_5284)
);

AO32x2_ASAP7_75t_L g5285 ( 
.A1(n_5069),
.A2(n_3515),
.A3(n_3451),
.B1(n_3158),
.B2(n_3438),
.Y(n_5285)
);

BUFx2_ASAP7_75t_L g5286 ( 
.A(n_4327),
.Y(n_5286)
);

AOI21x1_ASAP7_75t_L g5287 ( 
.A1(n_4528),
.A2(n_3090),
.B(n_3231),
.Y(n_5287)
);

AND2x2_ASAP7_75t_L g5288 ( 
.A(n_4196),
.B(n_4074),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_4306),
.Y(n_5289)
);

NOR2xp33_ASAP7_75t_L g5290 ( 
.A(n_4285),
.B(n_3413),
.Y(n_5290)
);

AOI21x1_ASAP7_75t_L g5291 ( 
.A1(n_4528),
.A2(n_3090),
.B(n_3541),
.Y(n_5291)
);

AND2x4_ASAP7_75t_L g5292 ( 
.A(n_4222),
.B(n_4074),
.Y(n_5292)
);

HB1xp67_ASAP7_75t_L g5293 ( 
.A(n_4331),
.Y(n_5293)
);

OAI22xp33_ASAP7_75t_L g5294 ( 
.A1(n_4184),
.A2(n_3447),
.B1(n_3425),
.B2(n_3525),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_4306),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_4318),
.Y(n_5296)
);

NAND3xp33_ASAP7_75t_L g5297 ( 
.A(n_4581),
.B(n_3408),
.C(n_3359),
.Y(n_5297)
);

AND2x6_ASAP7_75t_L g5298 ( 
.A(n_5073),
.B(n_4074),
.Y(n_5298)
);

INVx1_ASAP7_75t_SL g5299 ( 
.A(n_4475),
.Y(n_5299)
);

BUFx4_ASAP7_75t_SL g5300 ( 
.A(n_4391),
.Y(n_5300)
);

OR2x6_ASAP7_75t_L g5301 ( 
.A(n_4160),
.B(n_4074),
.Y(n_5301)
);

AOI21xp5_ASAP7_75t_L g5302 ( 
.A1(n_4219),
.A2(n_3335),
.B(n_3334),
.Y(n_5302)
);

HB1xp67_ASAP7_75t_L g5303 ( 
.A(n_4331),
.Y(n_5303)
);

INVx1_ASAP7_75t_L g5304 ( 
.A(n_4318),
.Y(n_5304)
);

INVx2_ASAP7_75t_SL g5305 ( 
.A(n_5010),
.Y(n_5305)
);

AOI21xp5_ASAP7_75t_L g5306 ( 
.A1(n_4236),
.A2(n_3230),
.B(n_3171),
.Y(n_5306)
);

AND2x2_ASAP7_75t_L g5307 ( 
.A(n_4196),
.B(n_4087),
.Y(n_5307)
);

AOI21xp5_ASAP7_75t_L g5308 ( 
.A1(n_4236),
.A2(n_3537),
.B(n_3342),
.Y(n_5308)
);

INVx1_ASAP7_75t_L g5309 ( 
.A(n_4318),
.Y(n_5309)
);

NAND2xp5_ASAP7_75t_L g5310 ( 
.A(n_4722),
.B(n_3350),
.Y(n_5310)
);

AOI22xp33_ASAP7_75t_L g5311 ( 
.A1(n_4270),
.A2(n_3525),
.B1(n_3545),
.B2(n_3546),
.Y(n_5311)
);

OAI22xp5_ASAP7_75t_L g5312 ( 
.A1(n_4412),
.A2(n_3447),
.B1(n_3413),
.B2(n_3525),
.Y(n_5312)
);

INVx5_ASAP7_75t_L g5313 ( 
.A(n_4195),
.Y(n_5313)
);

AOI22xp33_ASAP7_75t_L g5314 ( 
.A1(n_4162),
.A2(n_3525),
.B1(n_3545),
.B2(n_3546),
.Y(n_5314)
);

NOR2x1_ASAP7_75t_L g5315 ( 
.A(n_4850),
.B(n_3200),
.Y(n_5315)
);

AOI22xp33_ASAP7_75t_L g5316 ( 
.A1(n_4185),
.A2(n_3525),
.B1(n_3533),
.B2(n_3351),
.Y(n_5316)
);

INVx1_ASAP7_75t_L g5317 ( 
.A(n_4338),
.Y(n_5317)
);

BUFx2_ASAP7_75t_L g5318 ( 
.A(n_4346),
.Y(n_5318)
);

OR2x6_ASAP7_75t_L g5319 ( 
.A(n_4160),
.B(n_4087),
.Y(n_5319)
);

INVx3_ASAP7_75t_L g5320 ( 
.A(n_4555),
.Y(n_5320)
);

HB1xp67_ASAP7_75t_L g5321 ( 
.A(n_4336),
.Y(n_5321)
);

INVx1_ASAP7_75t_L g5322 ( 
.A(n_4338),
.Y(n_5322)
);

AOI22xp33_ASAP7_75t_L g5323 ( 
.A1(n_4588),
.A2(n_3533),
.B1(n_4087),
.B2(n_3536),
.Y(n_5323)
);

NAND2xp5_ASAP7_75t_L g5324 ( 
.A(n_4729),
.B(n_3356),
.Y(n_5324)
);

AND2x2_ASAP7_75t_L g5325 ( 
.A(n_4196),
.B(n_4087),
.Y(n_5325)
);

INVx1_ASAP7_75t_SL g5326 ( 
.A(n_4475),
.Y(n_5326)
);

INVx1_ASAP7_75t_L g5327 ( 
.A(n_4338),
.Y(n_5327)
);

INVx3_ASAP7_75t_L g5328 ( 
.A(n_4555),
.Y(n_5328)
);

HB1xp67_ASAP7_75t_L g5329 ( 
.A(n_4336),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_4339),
.Y(n_5330)
);

A2O1A1Ixp33_ASAP7_75t_L g5331 ( 
.A1(n_4629),
.A2(n_3511),
.B(n_3519),
.C(n_3362),
.Y(n_5331)
);

INVx1_ASAP7_75t_SL g5332 ( 
.A(n_4484),
.Y(n_5332)
);

BUFx6f_ASAP7_75t_L g5333 ( 
.A(n_5010),
.Y(n_5333)
);

NAND2xp5_ASAP7_75t_L g5334 ( 
.A(n_4729),
.B(n_3405),
.Y(n_5334)
);

INVx3_ASAP7_75t_L g5335 ( 
.A(n_5010),
.Y(n_5335)
);

INVx2_ASAP7_75t_SL g5336 ( 
.A(n_5010),
.Y(n_5336)
);

OAI22xp33_ASAP7_75t_L g5337 ( 
.A1(n_4848),
.A2(n_3559),
.B1(n_4087),
.B2(n_3560),
.Y(n_5337)
);

INVx1_ASAP7_75t_SL g5338 ( 
.A(n_4484),
.Y(n_5338)
);

NAND2xp5_ASAP7_75t_SL g5339 ( 
.A(n_4200),
.B(n_3563),
.Y(n_5339)
);

INVx1_ASAP7_75t_L g5340 ( 
.A(n_4339),
.Y(n_5340)
);

INVxp67_ASAP7_75t_SL g5341 ( 
.A(n_4954),
.Y(n_5341)
);

CKINVDCx5p33_ASAP7_75t_R g5342 ( 
.A(n_4836),
.Y(n_5342)
);

INVx1_ASAP7_75t_SL g5343 ( 
.A(n_4762),
.Y(n_5343)
);

INVx5_ASAP7_75t_L g5344 ( 
.A(n_4195),
.Y(n_5344)
);

INVx4_ASAP7_75t_L g5345 ( 
.A(n_5102),
.Y(n_5345)
);

OAI22xp5_ASAP7_75t_L g5346 ( 
.A1(n_4412),
.A2(n_3571),
.B1(n_3344),
.B2(n_3559),
.Y(n_5346)
);

CKINVDCx5p33_ASAP7_75t_R g5347 ( 
.A(n_4836),
.Y(n_5347)
);

AOI222xp33_ASAP7_75t_L g5348 ( 
.A1(n_4581),
.A2(n_3330),
.B1(n_3550),
.B2(n_3540),
.C1(n_3563),
.C2(n_3536),
.Y(n_5348)
);

AOI21xp5_ASAP7_75t_L g5349 ( 
.A1(n_4251),
.A2(n_3374),
.B(n_3337),
.Y(n_5349)
);

AOI21xp5_ASAP7_75t_L g5350 ( 
.A1(n_4251),
.A2(n_3427),
.B(n_3399),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_4339),
.Y(n_5351)
);

NOR2xp33_ASAP7_75t_SL g5352 ( 
.A(n_4629),
.B(n_3563),
.Y(n_5352)
);

OAI22xp5_ASAP7_75t_L g5353 ( 
.A1(n_4425),
.A2(n_3571),
.B1(n_3344),
.B2(n_3576),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_4347),
.Y(n_5354)
);

INVx1_ASAP7_75t_L g5355 ( 
.A(n_4347),
.Y(n_5355)
);

AND2x2_ASAP7_75t_L g5356 ( 
.A(n_4220),
.B(n_4243),
.Y(n_5356)
);

CKINVDCx20_ASAP7_75t_R g5357 ( 
.A(n_4391),
.Y(n_5357)
);

BUFx2_ASAP7_75t_L g5358 ( 
.A(n_4387),
.Y(n_5358)
);

AOI221xp5_ASAP7_75t_L g5359 ( 
.A1(n_4848),
.A2(n_3543),
.B1(n_3563),
.B2(n_3432),
.C(n_3577),
.Y(n_5359)
);

NOR2xp67_ASAP7_75t_L g5360 ( 
.A(n_4856),
.B(n_3535),
.Y(n_5360)
);

BUFx12f_ASAP7_75t_L g5361 ( 
.A(n_4868),
.Y(n_5361)
);

BUFx4_ASAP7_75t_SL g5362 ( 
.A(n_4153),
.Y(n_5362)
);

BUFx2_ASAP7_75t_L g5363 ( 
.A(n_4387),
.Y(n_5363)
);

NAND2xp5_ASAP7_75t_L g5364 ( 
.A(n_4730),
.B(n_3405),
.Y(n_5364)
);

INVx4_ASAP7_75t_L g5365 ( 
.A(n_5073),
.Y(n_5365)
);

INVx3_ASAP7_75t_L g5366 ( 
.A(n_4578),
.Y(n_5366)
);

NAND2xp5_ASAP7_75t_SL g5367 ( 
.A(n_4285),
.B(n_3341),
.Y(n_5367)
);

HB1xp67_ASAP7_75t_L g5368 ( 
.A(n_4350),
.Y(n_5368)
);

AND2x2_ASAP7_75t_L g5369 ( 
.A(n_4220),
.B(n_4243),
.Y(n_5369)
);

INVx3_ASAP7_75t_SL g5370 ( 
.A(n_4691),
.Y(n_5370)
);

OAI22xp5_ASAP7_75t_L g5371 ( 
.A1(n_4426),
.A2(n_3344),
.B1(n_3566),
.B2(n_3560),
.Y(n_5371)
);

INVx1_ASAP7_75t_L g5372 ( 
.A(n_4347),
.Y(n_5372)
);

NAND2xp5_ASAP7_75t_L g5373 ( 
.A(n_4730),
.B(n_3411),
.Y(n_5373)
);

NAND2xp5_ASAP7_75t_L g5374 ( 
.A(n_4734),
.B(n_3411),
.Y(n_5374)
);

INVx1_ASAP7_75t_L g5375 ( 
.A(n_4354),
.Y(n_5375)
);

NOR2xp33_ASAP7_75t_L g5376 ( 
.A(n_4317),
.B(n_3554),
.Y(n_5376)
);

AOI21xp5_ASAP7_75t_L g5377 ( 
.A1(n_4393),
.A2(n_3504),
.B(n_3446),
.Y(n_5377)
);

INVx1_ASAP7_75t_L g5378 ( 
.A(n_4354),
.Y(n_5378)
);

INVx1_ASAP7_75t_L g5379 ( 
.A(n_4354),
.Y(n_5379)
);

BUFx2_ASAP7_75t_L g5380 ( 
.A(n_4387),
.Y(n_5380)
);

OAI21xp5_ASAP7_75t_L g5381 ( 
.A1(n_4426),
.A2(n_3238),
.B(n_3398),
.Y(n_5381)
);

AOI22xp33_ASAP7_75t_L g5382 ( 
.A1(n_4588),
.A2(n_3538),
.B1(n_3540),
.B2(n_3550),
.Y(n_5382)
);

HB1xp67_ASAP7_75t_L g5383 ( 
.A(n_4350),
.Y(n_5383)
);

INVx5_ASAP7_75t_L g5384 ( 
.A(n_4195),
.Y(n_5384)
);

AND2x2_ASAP7_75t_L g5385 ( 
.A(n_4243),
.B(n_4261),
.Y(n_5385)
);

A2O1A1Ixp33_ASAP7_75t_SL g5386 ( 
.A1(n_4751),
.A2(n_3578),
.B(n_3535),
.C(n_3521),
.Y(n_5386)
);

INVx1_ASAP7_75t_L g5387 ( 
.A(n_4368),
.Y(n_5387)
);

AND2x2_ASAP7_75t_SL g5388 ( 
.A(n_4316),
.B(n_3280),
.Y(n_5388)
);

INVx4_ASAP7_75t_L g5389 ( 
.A(n_5102),
.Y(n_5389)
);

INVxp67_ASAP7_75t_L g5390 ( 
.A(n_4914),
.Y(n_5390)
);

OAI22xp33_ASAP7_75t_L g5391 ( 
.A1(n_4624),
.A2(n_3538),
.B1(n_3369),
.B2(n_3330),
.Y(n_5391)
);

AOI222xp33_ASAP7_75t_L g5392 ( 
.A1(n_4436),
.A2(n_3579),
.B1(n_3327),
.B2(n_3326),
.C1(n_3324),
.C2(n_3309),
.Y(n_5392)
);

AOI22xp5_ASAP7_75t_L g5393 ( 
.A1(n_4645),
.A2(n_3406),
.B1(n_3507),
.B2(n_3523),
.Y(n_5393)
);

INVx4_ASAP7_75t_L g5394 ( 
.A(n_5073),
.Y(n_5394)
);

NAND2xp5_ASAP7_75t_L g5395 ( 
.A(n_4734),
.B(n_3416),
.Y(n_5395)
);

INVx1_ASAP7_75t_L g5396 ( 
.A(n_4368),
.Y(n_5396)
);

INVxp67_ASAP7_75t_L g5397 ( 
.A(n_4689),
.Y(n_5397)
);

NAND3xp33_ASAP7_75t_L g5398 ( 
.A(n_4605),
.B(n_3517),
.C(n_3439),
.Y(n_5398)
);

INVx4_ASAP7_75t_L g5399 ( 
.A(n_5073),
.Y(n_5399)
);

INVx1_ASAP7_75t_SL g5400 ( 
.A(n_4762),
.Y(n_5400)
);

AOI22xp33_ASAP7_75t_L g5401 ( 
.A1(n_4436),
.A2(n_4089),
.B1(n_4070),
.B2(n_4068),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_4368),
.Y(n_5402)
);

OR2x6_ASAP7_75t_L g5403 ( 
.A(n_4292),
.B(n_3416),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_4373),
.Y(n_5404)
);

AOI21xp5_ASAP7_75t_L g5405 ( 
.A1(n_4393),
.A2(n_3522),
.B(n_3531),
.Y(n_5405)
);

NOR2xp33_ASAP7_75t_L g5406 ( 
.A(n_4317),
.B(n_3554),
.Y(n_5406)
);

NAND2xp5_ASAP7_75t_L g5407 ( 
.A(n_4741),
.B(n_3417),
.Y(n_5407)
);

A2O1A1Ixp33_ASAP7_75t_L g5408 ( 
.A1(n_4891),
.A2(n_3367),
.B(n_3574),
.C(n_3575),
.Y(n_5408)
);

HB1xp67_ASAP7_75t_L g5409 ( 
.A(n_4375),
.Y(n_5409)
);

NAND2xp5_ASAP7_75t_L g5410 ( 
.A(n_4741),
.B(n_3417),
.Y(n_5410)
);

AOI21xp5_ASAP7_75t_L g5411 ( 
.A1(n_4401),
.A2(n_3532),
.B(n_3200),
.Y(n_5411)
);

OR2x2_ASAP7_75t_L g5412 ( 
.A(n_4712),
.B(n_3454),
.Y(n_5412)
);

BUFx2_ASAP7_75t_L g5413 ( 
.A(n_4419),
.Y(n_5413)
);

OAI22xp33_ASAP7_75t_L g5414 ( 
.A1(n_4624),
.A2(n_3369),
.B1(n_3572),
.B2(n_3523),
.Y(n_5414)
);

AND2x6_ASAP7_75t_SL g5415 ( 
.A(n_4525),
.B(n_3573),
.Y(n_5415)
);

AOI21xp5_ASAP7_75t_L g5416 ( 
.A1(n_4401),
.A2(n_3285),
.B(n_3294),
.Y(n_5416)
);

INVx1_ASAP7_75t_SL g5417 ( 
.A(n_4793),
.Y(n_5417)
);

INVx3_ASAP7_75t_L g5418 ( 
.A(n_4578),
.Y(n_5418)
);

NAND2x1p5_ASAP7_75t_L g5419 ( 
.A(n_4316),
.B(n_3369),
.Y(n_5419)
);

INVx2_ASAP7_75t_SL g5420 ( 
.A(n_5024),
.Y(n_5420)
);

INVx1_ASAP7_75t_L g5421 ( 
.A(n_4373),
.Y(n_5421)
);

O2A1O1Ixp33_ASAP7_75t_L g5422 ( 
.A1(n_4702),
.A2(n_3555),
.B(n_3556),
.C(n_3549),
.Y(n_5422)
);

INVx3_ASAP7_75t_L g5423 ( 
.A(n_5024),
.Y(n_5423)
);

AOI22xp5_ASAP7_75t_L g5424 ( 
.A1(n_4645),
.A2(n_3406),
.B1(n_3369),
.B2(n_3280),
.Y(n_5424)
);

O2A1O1Ixp33_ASAP7_75t_L g5425 ( 
.A1(n_4466),
.A2(n_3482),
.B(n_3503),
.C(n_3547),
.Y(n_5425)
);

AOI211xp5_ASAP7_75t_L g5426 ( 
.A1(n_4779),
.A2(n_3574),
.B(n_3570),
.C(n_3575),
.Y(n_5426)
);

OAI22xp5_ASAP7_75t_L g5427 ( 
.A1(n_4466),
.A2(n_3572),
.B1(n_3323),
.B2(n_3285),
.Y(n_5427)
);

NAND2xp5_ASAP7_75t_SL g5428 ( 
.A(n_4467),
.B(n_3470),
.Y(n_5428)
);

O2A1O1Ixp33_ASAP7_75t_L g5429 ( 
.A1(n_4467),
.A2(n_3547),
.B(n_3573),
.C(n_3570),
.Y(n_5429)
);

INVx1_ASAP7_75t_L g5430 ( 
.A(n_4373),
.Y(n_5430)
);

AOI21xp5_ASAP7_75t_L g5431 ( 
.A1(n_4442),
.A2(n_3294),
.B(n_3304),
.Y(n_5431)
);

NOR2x1_ASAP7_75t_L g5432 ( 
.A(n_4856),
.B(n_4862),
.Y(n_5432)
);

NOR2xp33_ASAP7_75t_L g5433 ( 
.A(n_4299),
.B(n_3557),
.Y(n_5433)
);

NAND2xp5_ASAP7_75t_L g5434 ( 
.A(n_4750),
.B(n_4773),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_4374),
.Y(n_5435)
);

AND2x2_ASAP7_75t_L g5436 ( 
.A(n_4261),
.B(n_4731),
.Y(n_5436)
);

NAND2xp5_ASAP7_75t_L g5437 ( 
.A(n_4750),
.B(n_3418),
.Y(n_5437)
);

CKINVDCx8_ASAP7_75t_R g5438 ( 
.A(n_4292),
.Y(n_5438)
);

O2A1O1Ixp5_ASAP7_75t_SL g5439 ( 
.A1(n_4286),
.A2(n_3506),
.B(n_3323),
.C(n_3535),
.Y(n_5439)
);

NOR2xp33_ASAP7_75t_L g5440 ( 
.A(n_4299),
.B(n_3557),
.Y(n_5440)
);

INVx1_ASAP7_75t_L g5441 ( 
.A(n_4374),
.Y(n_5441)
);

INVx1_ASAP7_75t_L g5442 ( 
.A(n_4374),
.Y(n_5442)
);

AOI21xp5_ASAP7_75t_L g5443 ( 
.A1(n_4442),
.A2(n_3304),
.B(n_3452),
.Y(n_5443)
);

AND2x2_ASAP7_75t_SL g5444 ( 
.A(n_4316),
.B(n_3304),
.Y(n_5444)
);

NOR2xp33_ASAP7_75t_L g5445 ( 
.A(n_4678),
.B(n_3535),
.Y(n_5445)
);

HB1xp67_ASAP7_75t_L g5446 ( 
.A(n_4375),
.Y(n_5446)
);

INVx3_ASAP7_75t_L g5447 ( 
.A(n_5024),
.Y(n_5447)
);

INVx3_ASAP7_75t_L g5448 ( 
.A(n_4578),
.Y(n_5448)
);

O2A1O1Ixp33_ASAP7_75t_L g5449 ( 
.A1(n_4589),
.A2(n_3580),
.B(n_3529),
.C(n_3465),
.Y(n_5449)
);

CKINVDCx20_ASAP7_75t_R g5450 ( 
.A(n_4724),
.Y(n_5450)
);

NOR2xp33_ASAP7_75t_L g5451 ( 
.A(n_4678),
.B(n_3470),
.Y(n_5451)
);

OAI22xp5_ASAP7_75t_L g5452 ( 
.A1(n_4477),
.A2(n_3572),
.B1(n_3323),
.B2(n_3580),
.Y(n_5452)
);

AOI22xp5_ASAP7_75t_L g5453 ( 
.A1(n_4431),
.A2(n_3572),
.B1(n_3534),
.B2(n_3467),
.Y(n_5453)
);

INVx1_ASAP7_75t_L g5454 ( 
.A(n_4377),
.Y(n_5454)
);

HB1xp67_ASAP7_75t_L g5455 ( 
.A(n_4156),
.Y(n_5455)
);

BUFx4f_ASAP7_75t_SL g5456 ( 
.A(n_4480),
.Y(n_5456)
);

AOI21x1_ASAP7_75t_L g5457 ( 
.A1(n_4528),
.A2(n_4275),
.B(n_4255),
.Y(n_5457)
);

O2A1O1Ixp33_ASAP7_75t_L g5458 ( 
.A1(n_4589),
.A2(n_3465),
.B(n_3467),
.C(n_3539),
.Y(n_5458)
);

INVx1_ASAP7_75t_L g5459 ( 
.A(n_4377),
.Y(n_5459)
);

INVx1_ASAP7_75t_L g5460 ( 
.A(n_4377),
.Y(n_5460)
);

AOI22xp33_ASAP7_75t_L g5461 ( 
.A1(n_4840),
.A2(n_4089),
.B1(n_4070),
.B2(n_4068),
.Y(n_5461)
);

AND2x4_ASAP7_75t_L g5462 ( 
.A(n_5091),
.B(n_5073),
.Y(n_5462)
);

BUFx12f_ASAP7_75t_L g5463 ( 
.A(n_4868),
.Y(n_5463)
);

INVx3_ASAP7_75t_L g5464 ( 
.A(n_4578),
.Y(n_5464)
);

OR2x2_ASAP7_75t_L g5465 ( 
.A(n_4714),
.B(n_3454),
.Y(n_5465)
);

AOI221xp5_ASAP7_75t_L g5466 ( 
.A1(n_4840),
.A2(n_3430),
.B1(n_3444),
.B2(n_3443),
.C(n_3448),
.Y(n_5466)
);

NAND2xp5_ASAP7_75t_L g5467 ( 
.A(n_4773),
.B(n_3418),
.Y(n_5467)
);

BUFx2_ASAP7_75t_L g5468 ( 
.A(n_4886),
.Y(n_5468)
);

INVx1_ASAP7_75t_L g5469 ( 
.A(n_4381),
.Y(n_5469)
);

AOI21xp5_ASAP7_75t_L g5470 ( 
.A1(n_4286),
.A2(n_3436),
.B(n_3452),
.Y(n_5470)
);

INVx2_ASAP7_75t_L g5471 ( 
.A(n_4209),
.Y(n_5471)
);

CKINVDCx20_ASAP7_75t_R g5472 ( 
.A(n_4724),
.Y(n_5472)
);

INVx1_ASAP7_75t_L g5473 ( 
.A(n_4381),
.Y(n_5473)
);

AOI21xp5_ASAP7_75t_L g5474 ( 
.A1(n_4691),
.A2(n_3436),
.B(n_3450),
.Y(n_5474)
);

OAI22xp5_ASAP7_75t_L g5475 ( 
.A1(n_4477),
.A2(n_3572),
.B1(n_3323),
.B2(n_3700),
.Y(n_5475)
);

OR2x2_ASAP7_75t_L g5476 ( 
.A(n_4714),
.B(n_4036),
.Y(n_5476)
);

HB1xp67_ASAP7_75t_L g5477 ( 
.A(n_4156),
.Y(n_5477)
);

INVx1_ASAP7_75t_L g5478 ( 
.A(n_4381),
.Y(n_5478)
);

HB1xp67_ASAP7_75t_L g5479 ( 
.A(n_4181),
.Y(n_5479)
);

INVx2_ASAP7_75t_L g5480 ( 
.A(n_4209),
.Y(n_5480)
);

AOI22xp33_ASAP7_75t_L g5481 ( 
.A1(n_4431),
.A2(n_4089),
.B1(n_4070),
.B2(n_4036),
.Y(n_5481)
);

NAND2xp5_ASAP7_75t_L g5482 ( 
.A(n_4778),
.B(n_3430),
.Y(n_5482)
);

INVx1_ASAP7_75t_L g5483 ( 
.A(n_4386),
.Y(n_5483)
);

NOR2x1_ASAP7_75t_L g5484 ( 
.A(n_4862),
.B(n_4778),
.Y(n_5484)
);

INVx1_ASAP7_75t_L g5485 ( 
.A(n_4386),
.Y(n_5485)
);

INVx1_ASAP7_75t_L g5486 ( 
.A(n_4386),
.Y(n_5486)
);

INVx2_ASAP7_75t_L g5487 ( 
.A(n_4209),
.Y(n_5487)
);

INVx3_ASAP7_75t_L g5488 ( 
.A(n_4578),
.Y(n_5488)
);

O2A1O1Ixp33_ASAP7_75t_L g5489 ( 
.A1(n_4516),
.A2(n_3539),
.B(n_3158),
.C(n_3700),
.Y(n_5489)
);

HB1xp67_ASAP7_75t_L g5490 ( 
.A(n_4181),
.Y(n_5490)
);

A2O1A1Ixp33_ASAP7_75t_L g5491 ( 
.A1(n_4891),
.A2(n_3444),
.B(n_3434),
.C(n_3450),
.Y(n_5491)
);

AOI22xp33_ASAP7_75t_L g5492 ( 
.A1(n_4825),
.A2(n_4379),
.B1(n_4852),
.B2(n_4831),
.Y(n_5492)
);

INVx4_ASAP7_75t_L g5493 ( 
.A(n_5102),
.Y(n_5493)
);

INVx2_ASAP7_75t_L g5494 ( 
.A(n_4209),
.Y(n_5494)
);

OAI21xp33_ASAP7_75t_L g5495 ( 
.A1(n_4831),
.A2(n_3620),
.B(n_3475),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_4394),
.Y(n_5496)
);

AOI222xp33_ASAP7_75t_L g5497 ( 
.A1(n_5033),
.A2(n_4409),
.B1(n_4779),
.B2(n_4227),
.C1(n_4852),
.C2(n_4379),
.Y(n_5497)
);

BUFx2_ASAP7_75t_L g5498 ( 
.A(n_4886),
.Y(n_5498)
);

AND2x2_ASAP7_75t_L g5499 ( 
.A(n_4731),
.B(n_4038),
.Y(n_5499)
);

AO32x2_ASAP7_75t_L g5500 ( 
.A1(n_5069),
.A2(n_4591),
.A3(n_4679),
.B1(n_4516),
.B2(n_4202),
.Y(n_5500)
);

INVx3_ASAP7_75t_L g5501 ( 
.A(n_4578),
.Y(n_5501)
);

AOI21xp5_ASAP7_75t_L g5502 ( 
.A1(n_4329),
.A2(n_3445),
.B(n_3448),
.Y(n_5502)
);

AOI21xp5_ASAP7_75t_L g5503 ( 
.A1(n_4329),
.A2(n_3434),
.B(n_3445),
.Y(n_5503)
);

A2O1A1Ixp33_ASAP7_75t_L g5504 ( 
.A1(n_4892),
.A2(n_3435),
.B(n_3431),
.C(n_3443),
.Y(n_5504)
);

OAI22xp5_ASAP7_75t_SL g5505 ( 
.A1(n_4525),
.A2(n_3853),
.B1(n_3810),
.B2(n_3313),
.Y(n_5505)
);

INVx1_ASAP7_75t_L g5506 ( 
.A(n_4394),
.Y(n_5506)
);

AOI22xp33_ASAP7_75t_SL g5507 ( 
.A1(n_4892),
.A2(n_3460),
.B1(n_3491),
.B2(n_4068),
.Y(n_5507)
);

AOI21xp5_ASAP7_75t_L g5508 ( 
.A1(n_4275),
.A2(n_3435),
.B(n_3431),
.Y(n_5508)
);

INVxp67_ASAP7_75t_SL g5509 ( 
.A(n_5007),
.Y(n_5509)
);

A2O1A1Ixp33_ASAP7_75t_L g5510 ( 
.A1(n_4865),
.A2(n_3474),
.B(n_3309),
.C(n_3327),
.Y(n_5510)
);

INVx1_ASAP7_75t_L g5511 ( 
.A(n_4394),
.Y(n_5511)
);

AOI22xp5_ASAP7_75t_L g5512 ( 
.A1(n_4536),
.A2(n_4066),
.B1(n_4038),
.B2(n_4042),
.Y(n_5512)
);

HB1xp67_ASAP7_75t_L g5513 ( 
.A(n_4186),
.Y(n_5513)
);

CKINVDCx5p33_ASAP7_75t_R g5514 ( 
.A(n_4153),
.Y(n_5514)
);

A2O1A1Ixp33_ASAP7_75t_L g5515 ( 
.A1(n_4865),
.A2(n_3474),
.B(n_3326),
.C(n_3318),
.Y(n_5515)
);

AOI21xp5_ASAP7_75t_L g5516 ( 
.A1(n_4326),
.A2(n_3634),
.B(n_3313),
.Y(n_5516)
);

NOR2xp33_ASAP7_75t_L g5517 ( 
.A(n_4692),
.B(n_3620),
.Y(n_5517)
);

AOI21xp5_ASAP7_75t_L g5518 ( 
.A1(n_4326),
.A2(n_3634),
.B(n_3978),
.Y(n_5518)
);

HB1xp67_ASAP7_75t_L g5519 ( 
.A(n_4186),
.Y(n_5519)
);

NAND2xp5_ASAP7_75t_SL g5520 ( 
.A(n_4577),
.B(n_3643),
.Y(n_5520)
);

INVx2_ASAP7_75t_L g5521 ( 
.A(n_4214),
.Y(n_5521)
);

INVx2_ASAP7_75t_L g5522 ( 
.A(n_4214),
.Y(n_5522)
);

AOI22xp5_ASAP7_75t_L g5523 ( 
.A1(n_4536),
.A2(n_4066),
.B1(n_4038),
.B2(n_4042),
.Y(n_5523)
);

AOI21xp5_ASAP7_75t_L g5524 ( 
.A1(n_4362),
.A2(n_3978),
.B(n_3681),
.Y(n_5524)
);

INVx2_ASAP7_75t_L g5525 ( 
.A(n_4214),
.Y(n_5525)
);

BUFx2_ASAP7_75t_L g5526 ( 
.A(n_4888),
.Y(n_5526)
);

INVx1_ASAP7_75t_SL g5527 ( 
.A(n_4793),
.Y(n_5527)
);

INVx3_ASAP7_75t_SL g5528 ( 
.A(n_4692),
.Y(n_5528)
);

INVx1_ASAP7_75t_L g5529 ( 
.A(n_4396),
.Y(n_5529)
);

NOR2xp33_ASAP7_75t_SL g5530 ( 
.A(n_4340),
.B(n_3853),
.Y(n_5530)
);

BUFx12f_ASAP7_75t_L g5531 ( 
.A(n_4896),
.Y(n_5531)
);

AOI21xp5_ASAP7_75t_L g5532 ( 
.A1(n_4362),
.A2(n_3669),
.B(n_3681),
.Y(n_5532)
);

BUFx2_ASAP7_75t_L g5533 ( 
.A(n_4888),
.Y(n_5533)
);

A2O1A1Ixp33_ASAP7_75t_L g5534 ( 
.A1(n_4606),
.A2(n_3324),
.B(n_3318),
.C(n_3475),
.Y(n_5534)
);

AOI22xp5_ASAP7_75t_L g5535 ( 
.A1(n_4227),
.A2(n_4065),
.B1(n_4042),
.B2(n_4044),
.Y(n_5535)
);

INVx1_ASAP7_75t_L g5536 ( 
.A(n_4396),
.Y(n_5536)
);

AOI22xp5_ASAP7_75t_L g5537 ( 
.A1(n_4605),
.A2(n_4065),
.B1(n_4044),
.B2(n_4046),
.Y(n_5537)
);

O2A1O1Ixp33_ASAP7_75t_L g5538 ( 
.A1(n_4572),
.A2(n_4580),
.B(n_4547),
.C(n_4591),
.Y(n_5538)
);

AOI21xp5_ASAP7_75t_L g5539 ( 
.A1(n_4389),
.A2(n_3643),
.B(n_3437),
.Y(n_5539)
);

AOI22xp33_ASAP7_75t_L g5540 ( 
.A1(n_4825),
.A2(n_4065),
.B1(n_4064),
.B2(n_4061),
.Y(n_5540)
);

A2O1A1Ixp33_ASAP7_75t_L g5541 ( 
.A1(n_4606),
.A2(n_3669),
.B(n_3437),
.C(n_3438),
.Y(n_5541)
);

CKINVDCx8_ASAP7_75t_R g5542 ( 
.A(n_4292),
.Y(n_5542)
);

NAND2xp5_ASAP7_75t_L g5543 ( 
.A(n_4142),
.B(n_4064),
.Y(n_5543)
);

NOR2xp33_ASAP7_75t_L g5544 ( 
.A(n_4696),
.B(n_3451),
.Y(n_5544)
);

AOI21xp5_ASAP7_75t_L g5545 ( 
.A1(n_4389),
.A2(n_3784),
.B(n_3810),
.Y(n_5545)
);

INVx3_ASAP7_75t_L g5546 ( 
.A(n_4587),
.Y(n_5546)
);

BUFx2_ASAP7_75t_L g5547 ( 
.A(n_4897),
.Y(n_5547)
);

NAND2xp5_ASAP7_75t_L g5548 ( 
.A(n_4142),
.B(n_4064),
.Y(n_5548)
);

BUFx2_ASAP7_75t_L g5549 ( 
.A(n_4897),
.Y(n_5549)
);

INVx1_ASAP7_75t_L g5550 ( 
.A(n_4396),
.Y(n_5550)
);

NAND2xp5_ASAP7_75t_L g5551 ( 
.A(n_4146),
.B(n_4061),
.Y(n_5551)
);

INVx2_ASAP7_75t_L g5552 ( 
.A(n_4214),
.Y(n_5552)
);

INVx2_ASAP7_75t_L g5553 ( 
.A(n_4221),
.Y(n_5553)
);

OAI22xp5_ASAP7_75t_L g5554 ( 
.A1(n_4341),
.A2(n_3784),
.B1(n_3853),
.B2(n_4061),
.Y(n_5554)
);

INVx1_ASAP7_75t_L g5555 ( 
.A(n_4398),
.Y(n_5555)
);

AOI22xp5_ASAP7_75t_L g5556 ( 
.A1(n_4716),
.A2(n_4046),
.B1(n_4044),
.B2(n_3460),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_4398),
.Y(n_5557)
);

INVx1_ASAP7_75t_L g5558 ( 
.A(n_4398),
.Y(n_5558)
);

HB1xp67_ASAP7_75t_L g5559 ( 
.A(n_4294),
.Y(n_5559)
);

O2A1O1Ixp33_ASAP7_75t_L g5560 ( 
.A1(n_4572),
.A2(n_3492),
.B(n_3505),
.C(n_3514),
.Y(n_5560)
);

AOI21xp5_ASAP7_75t_L g5561 ( 
.A1(n_4407),
.A2(n_3490),
.B(n_3513),
.Y(n_5561)
);

HB1xp67_ASAP7_75t_L g5562 ( 
.A(n_4294),
.Y(n_5562)
);

AND2x2_ASAP7_75t_L g5563 ( 
.A(n_4731),
.B(n_4046),
.Y(n_5563)
);

O2A1O1Ixp33_ASAP7_75t_L g5564 ( 
.A1(n_4580),
.A2(n_3492),
.B(n_3498),
.C(n_3514),
.Y(n_5564)
);

INVx3_ASAP7_75t_L g5565 ( 
.A(n_5031),
.Y(n_5565)
);

AOI22xp33_ASAP7_75t_L g5566 ( 
.A1(n_4409),
.A2(n_3491),
.B1(n_3462),
.B2(n_3493),
.Y(n_5566)
);

INVx2_ASAP7_75t_L g5567 ( 
.A(n_4221),
.Y(n_5567)
);

OAI21xp5_ASAP7_75t_L g5568 ( 
.A1(n_4341),
.A2(n_3464),
.B(n_3099),
.Y(n_5568)
);

AOI21xp5_ASAP7_75t_L g5569 ( 
.A1(n_4407),
.A2(n_3487),
.B(n_3513),
.Y(n_5569)
);

OAI22xp5_ASAP7_75t_L g5570 ( 
.A1(n_4215),
.A2(n_3480),
.B1(n_3462),
.B2(n_3488),
.Y(n_5570)
);

AND2x4_ASAP7_75t_L g5571 ( 
.A(n_5091),
.B(n_3099),
.Y(n_5571)
);

NOR2xp33_ASAP7_75t_L g5572 ( 
.A(n_4696),
.B(n_3099),
.Y(n_5572)
);

INVx2_ASAP7_75t_L g5573 ( 
.A(n_4221),
.Y(n_5573)
);

AOI21xp5_ASAP7_75t_L g5574 ( 
.A1(n_4411),
.A2(n_3495),
.B(n_3490),
.Y(n_5574)
);

CKINVDCx8_ASAP7_75t_R g5575 ( 
.A(n_5074),
.Y(n_5575)
);

OR2x6_ASAP7_75t_L g5576 ( 
.A(n_4246),
.B(n_3487),
.Y(n_5576)
);

O2A1O1Ixp33_ASAP7_75t_L g5577 ( 
.A1(n_4547),
.A2(n_3483),
.B(n_3510),
.C(n_3471),
.Y(n_5577)
);

HB1xp67_ASAP7_75t_L g5578 ( 
.A(n_4370),
.Y(n_5578)
);

INVx2_ASAP7_75t_L g5579 ( 
.A(n_4221),
.Y(n_5579)
);

HB1xp67_ASAP7_75t_L g5580 ( 
.A(n_4370),
.Y(n_5580)
);

OAI21xp33_ASAP7_75t_L g5581 ( 
.A1(n_4620),
.A2(n_3488),
.B(n_3493),
.Y(n_5581)
);

INVx2_ASAP7_75t_L g5582 ( 
.A(n_4223),
.Y(n_5582)
);

INVx2_ASAP7_75t_L g5583 ( 
.A(n_4223),
.Y(n_5583)
);

NAND2xp5_ASAP7_75t_L g5584 ( 
.A(n_4146),
.B(n_3518),
.Y(n_5584)
);

AOI21xp5_ASAP7_75t_L g5585 ( 
.A1(n_4411),
.A2(n_3485),
.B(n_3495),
.Y(n_5585)
);

NAND3xp33_ASAP7_75t_L g5586 ( 
.A(n_4215),
.B(n_3480),
.C(n_3473),
.Y(n_5586)
);

AND2x2_ASAP7_75t_L g5587 ( 
.A(n_4150),
.B(n_3518),
.Y(n_5587)
);

OR2x6_ASAP7_75t_L g5588 ( 
.A(n_4246),
.B(n_4351),
.Y(n_5588)
);

O2A1O1Ixp33_ASAP7_75t_L g5589 ( 
.A1(n_4548),
.A2(n_3486),
.B(n_3505),
.C(n_3471),
.Y(n_5589)
);

AOI21xp5_ASAP7_75t_L g5590 ( 
.A1(n_4463),
.A2(n_3485),
.B(n_3509),
.Y(n_5590)
);

BUFx8_ASAP7_75t_SL g5591 ( 
.A(n_4761),
.Y(n_5591)
);

NOR2xp33_ASAP7_75t_L g5592 ( 
.A(n_4705),
.B(n_3464),
.Y(n_5592)
);

OAI22xp5_ASAP7_75t_L g5593 ( 
.A1(n_4548),
.A2(n_3473),
.B1(n_3472),
.B2(n_3486),
.Y(n_5593)
);

O2A1O1Ixp33_ASAP7_75t_L g5594 ( 
.A1(n_4574),
.A2(n_4620),
.B(n_4861),
.C(n_4969),
.Y(n_5594)
);

O2A1O1Ixp5_ASAP7_75t_L g5595 ( 
.A1(n_4963),
.A2(n_3476),
.B(n_3477),
.C(n_3469),
.Y(n_5595)
);

O2A1O1Ixp5_ASAP7_75t_L g5596 ( 
.A1(n_4963),
.A2(n_3476),
.B(n_3469),
.C(n_3499),
.Y(n_5596)
);

AOI22xp5_ASAP7_75t_L g5597 ( 
.A1(n_4716),
.A2(n_3472),
.B1(n_3496),
.B2(n_3499),
.Y(n_5597)
);

CKINVDCx5p33_ASAP7_75t_R g5598 ( 
.A(n_4896),
.Y(n_5598)
);

AOI21xp5_ASAP7_75t_L g5599 ( 
.A1(n_4463),
.A2(n_4500),
.B(n_4471),
.Y(n_5599)
);

INVx1_ASAP7_75t_SL g5600 ( 
.A(n_4916),
.Y(n_5600)
);

OAI21x1_ASAP7_75t_L g5601 ( 
.A1(n_4421),
.A2(n_3483),
.B(n_3489),
.Y(n_5601)
);

INVxp67_ASAP7_75t_L g5602 ( 
.A(n_4689),
.Y(n_5602)
);

AOI21xp5_ASAP7_75t_L g5603 ( 
.A1(n_4471),
.A2(n_3489),
.B(n_3498),
.Y(n_5603)
);

INVx2_ASAP7_75t_L g5604 ( 
.A(n_4223),
.Y(n_5604)
);

AOI22xp5_ASAP7_75t_L g5605 ( 
.A1(n_4577),
.A2(n_3496),
.B1(n_3499),
.B2(n_3510),
.Y(n_5605)
);

NOR2xp33_ASAP7_75t_L g5606 ( 
.A(n_4705),
.B(n_3496),
.Y(n_5606)
);

OAI22xp5_ASAP7_75t_L g5607 ( 
.A1(n_4574),
.A2(n_4496),
.B1(n_4664),
.B2(n_4657),
.Y(n_5607)
);

BUFx4f_ASAP7_75t_SL g5608 ( 
.A(n_4480),
.Y(n_5608)
);

INVx2_ASAP7_75t_L g5609 ( 
.A(n_4223),
.Y(n_5609)
);

AOI21xp5_ASAP7_75t_L g5610 ( 
.A1(n_4500),
.A2(n_4514),
.B(n_4506),
.Y(n_5610)
);

BUFx2_ASAP7_75t_L g5611 ( 
.A(n_4916),
.Y(n_5611)
);

HB1xp67_ASAP7_75t_L g5612 ( 
.A(n_4189),
.Y(n_5612)
);

NAND2xp5_ASAP7_75t_L g5613 ( 
.A(n_4783),
.B(n_4147),
.Y(n_5613)
);

NAND2xp5_ASAP7_75t_L g5614 ( 
.A(n_4783),
.B(n_4147),
.Y(n_5614)
);

INVx3_ASAP7_75t_L g5615 ( 
.A(n_4587),
.Y(n_5615)
);

A2O1A1Ixp33_ASAP7_75t_L g5616 ( 
.A1(n_5033),
.A2(n_4618),
.B(n_4820),
.C(n_4992),
.Y(n_5616)
);

AND2x2_ASAP7_75t_L g5617 ( 
.A(n_4150),
.B(n_4180),
.Y(n_5617)
);

NAND2xp5_ASAP7_75t_L g5618 ( 
.A(n_4161),
.B(n_4579),
.Y(n_5618)
);

AOI22xp33_ASAP7_75t_L g5619 ( 
.A1(n_4861),
.A2(n_4820),
.B1(n_4855),
.B2(n_4992),
.Y(n_5619)
);

NAND2xp5_ASAP7_75t_L g5620 ( 
.A(n_4161),
.B(n_4579),
.Y(n_5620)
);

AOI21xp5_ASAP7_75t_L g5621 ( 
.A1(n_4506),
.A2(n_4542),
.B(n_4514),
.Y(n_5621)
);

AOI21xp5_ASAP7_75t_L g5622 ( 
.A1(n_4542),
.A2(n_4546),
.B(n_4764),
.Y(n_5622)
);

NOR2x1_ASAP7_75t_L g5623 ( 
.A(n_4725),
.B(n_4863),
.Y(n_5623)
);

CKINVDCx5p33_ASAP7_75t_R g5624 ( 
.A(n_4975),
.Y(n_5624)
);

AOI21xp5_ASAP7_75t_L g5625 ( 
.A1(n_4546),
.A2(n_4764),
.B(n_4556),
.Y(n_5625)
);

AOI22xp5_ASAP7_75t_L g5626 ( 
.A1(n_4664),
.A2(n_4414),
.B1(n_5015),
.B2(n_4496),
.Y(n_5626)
);

OAI22xp5_ASAP7_75t_L g5627 ( 
.A1(n_4652),
.A2(n_4657),
.B1(n_4669),
.B2(n_4668),
.Y(n_5627)
);

CKINVDCx20_ASAP7_75t_R g5628 ( 
.A(n_4761),
.Y(n_5628)
);

AOI21xp5_ASAP7_75t_L g5629 ( 
.A1(n_4556),
.A2(n_5007),
.B(n_4384),
.Y(n_5629)
);

AND3x1_ASAP7_75t_SL g5630 ( 
.A(n_4414),
.B(n_4816),
.C(n_4863),
.Y(n_5630)
);

CKINVDCx8_ASAP7_75t_R g5631 ( 
.A(n_5074),
.Y(n_5631)
);

AOI21xp5_ASAP7_75t_L g5632 ( 
.A1(n_4384),
.A2(n_4421),
.B(n_4187),
.Y(n_5632)
);

AOI21xp5_ASAP7_75t_L g5633 ( 
.A1(n_4421),
.A2(n_4187),
.B(n_4172),
.Y(n_5633)
);

NAND2xp5_ASAP7_75t_L g5634 ( 
.A(n_4610),
.B(n_4168),
.Y(n_5634)
);

AO32x2_ASAP7_75t_L g5635 ( 
.A1(n_4679),
.A2(n_4143),
.A3(n_4204),
.B1(n_4202),
.B2(n_4170),
.Y(n_5635)
);

AOI21xp5_ASAP7_75t_L g5636 ( 
.A1(n_4421),
.A2(n_4188),
.B(n_4172),
.Y(n_5636)
);

BUFx2_ASAP7_75t_L g5637 ( 
.A(n_4916),
.Y(n_5637)
);

AOI21xp5_ASAP7_75t_L g5638 ( 
.A1(n_4188),
.A2(n_4194),
.B(n_4193),
.Y(n_5638)
);

AOI22xp33_ASAP7_75t_SL g5639 ( 
.A1(n_4560),
.A2(n_4618),
.B1(n_4453),
.B2(n_4946),
.Y(n_5639)
);

AOI22xp33_ASAP7_75t_L g5640 ( 
.A1(n_4855),
.A2(n_5015),
.B1(n_4969),
.B2(n_4652),
.Y(n_5640)
);

OAI22xp5_ASAP7_75t_L g5641 ( 
.A1(n_4668),
.A2(n_4669),
.B1(n_4796),
.B2(n_4792),
.Y(n_5641)
);

INVx3_ASAP7_75t_SL g5642 ( 
.A(n_4725),
.Y(n_5642)
);

BUFx12f_ASAP7_75t_L g5643 ( 
.A(n_4253),
.Y(n_5643)
);

A2O1A1Ixp33_ASAP7_75t_L g5644 ( 
.A1(n_4751),
.A2(n_4690),
.B(n_4898),
.C(n_4648),
.Y(n_5644)
);

OAI22xp5_ASAP7_75t_L g5645 ( 
.A1(n_4796),
.A2(n_4786),
.B1(n_4792),
.B2(n_4690),
.Y(n_5645)
);

A2O1A1Ixp33_ASAP7_75t_L g5646 ( 
.A1(n_4898),
.A2(n_4648),
.B(n_5005),
.C(n_4697),
.Y(n_5646)
);

AOI21xp5_ASAP7_75t_L g5647 ( 
.A1(n_4193),
.A2(n_4197),
.B(n_4194),
.Y(n_5647)
);

AO31x2_ASAP7_75t_L g5648 ( 
.A1(n_4182),
.A2(n_4183),
.A3(n_4207),
.B(n_4177),
.Y(n_5648)
);

BUFx2_ASAP7_75t_L g5649 ( 
.A(n_4932),
.Y(n_5649)
);

HB1xp67_ASAP7_75t_L g5650 ( 
.A(n_4189),
.Y(n_5650)
);

O2A1O1Ixp33_ASAP7_75t_L g5651 ( 
.A1(n_4727),
.A2(n_4941),
.B(n_4972),
.C(n_4639),
.Y(n_5651)
);

O2A1O1Ixp5_ASAP7_75t_SL g5652 ( 
.A1(n_4177),
.A2(n_4183),
.B(n_4207),
.C(n_4182),
.Y(n_5652)
);

BUFx2_ASAP7_75t_L g5653 ( 
.A(n_4932),
.Y(n_5653)
);

AND2x2_ASAP7_75t_L g5654 ( 
.A(n_4150),
.B(n_4180),
.Y(n_5654)
);

OAI22xp5_ASAP7_75t_L g5655 ( 
.A1(n_4786),
.A2(n_4972),
.B1(n_4823),
.B2(n_5098),
.Y(n_5655)
);

INVx3_ASAP7_75t_L g5656 ( 
.A(n_4587),
.Y(n_5656)
);

AOI21xp5_ASAP7_75t_L g5657 ( 
.A1(n_4197),
.A2(n_4218),
.B(n_4212),
.Y(n_5657)
);

NAND2xp5_ASAP7_75t_SL g5658 ( 
.A(n_4300),
.B(n_5008),
.Y(n_5658)
);

NAND2xp5_ASAP7_75t_L g5659 ( 
.A(n_4610),
.B(n_4168),
.Y(n_5659)
);

O2A1O1Ixp33_ASAP7_75t_L g5660 ( 
.A1(n_4727),
.A2(n_4941),
.B(n_4639),
.C(n_4651),
.Y(n_5660)
);

INVx8_ASAP7_75t_L g5661 ( 
.A(n_4537),
.Y(n_5661)
);

NAND2xp5_ASAP7_75t_L g5662 ( 
.A(n_4169),
.B(n_4746),
.Y(n_5662)
);

INVx1_ASAP7_75t_L g5663 ( 
.A(n_4433),
.Y(n_5663)
);

NAND2x1p5_ASAP7_75t_L g5664 ( 
.A(n_4416),
.B(n_4490),
.Y(n_5664)
);

NAND2xp5_ASAP7_75t_SL g5665 ( 
.A(n_4300),
.B(n_5008),
.Y(n_5665)
);

NAND2x1p5_ASAP7_75t_L g5666 ( 
.A(n_4416),
.B(n_4490),
.Y(n_5666)
);

INVx1_ASAP7_75t_L g5667 ( 
.A(n_4433),
.Y(n_5667)
);

NOR2xp33_ASAP7_75t_L g5668 ( 
.A(n_4300),
.B(n_4738),
.Y(n_5668)
);

INVx2_ASAP7_75t_L g5669 ( 
.A(n_4234),
.Y(n_5669)
);

AND2x4_ASAP7_75t_L g5670 ( 
.A(n_4195),
.B(n_4416),
.Y(n_5670)
);

INVx5_ASAP7_75t_L g5671 ( 
.A(n_4195),
.Y(n_5671)
);

AND2x6_ASAP7_75t_L g5672 ( 
.A(n_4785),
.B(n_4839),
.Y(n_5672)
);

AND2x4_ASAP7_75t_L g5673 ( 
.A(n_4195),
.B(n_4416),
.Y(n_5673)
);

AOI21xp5_ASAP7_75t_L g5674 ( 
.A1(n_4212),
.A2(n_4224),
.B(n_4218),
.Y(n_5674)
);

OAI22xp5_ASAP7_75t_L g5675 ( 
.A1(n_4823),
.A2(n_5098),
.B1(n_4770),
.B2(n_4743),
.Y(n_5675)
);

INVx1_ASAP7_75t_L g5676 ( 
.A(n_4434),
.Y(n_5676)
);

BUFx2_ASAP7_75t_L g5677 ( 
.A(n_4934),
.Y(n_5677)
);

OR2x6_ASAP7_75t_L g5678 ( 
.A(n_4246),
.B(n_4351),
.Y(n_5678)
);

NOR2xp33_ASAP7_75t_L g5679 ( 
.A(n_4300),
.B(n_4738),
.Y(n_5679)
);

HB1xp67_ASAP7_75t_L g5680 ( 
.A(n_4189),
.Y(n_5680)
);

NAND2xp5_ASAP7_75t_L g5681 ( 
.A(n_4169),
.B(n_4746),
.Y(n_5681)
);

CKINVDCx6p67_ASAP7_75t_R g5682 ( 
.A(n_4480),
.Y(n_5682)
);

AOI22xp5_ASAP7_75t_L g5683 ( 
.A1(n_4811),
.A2(n_4560),
.B1(n_5005),
.B2(n_4925),
.Y(n_5683)
);

INVx3_ASAP7_75t_L g5684 ( 
.A(n_4587),
.Y(n_5684)
);

NAND2xp5_ASAP7_75t_L g5685 ( 
.A(n_4781),
.B(n_4827),
.Y(n_5685)
);

INVx2_ASAP7_75t_L g5686 ( 
.A(n_4234),
.Y(n_5686)
);

AND2x2_ASAP7_75t_L g5687 ( 
.A(n_4180),
.B(n_4650),
.Y(n_5687)
);

HB1xp67_ASAP7_75t_L g5688 ( 
.A(n_4206),
.Y(n_5688)
);

A2O1A1Ixp33_ASAP7_75t_L g5689 ( 
.A1(n_4697),
.A2(n_4952),
.B(n_4811),
.C(n_5065),
.Y(n_5689)
);

INVx3_ASAP7_75t_L g5690 ( 
.A(n_4587),
.Y(n_5690)
);

OA22x2_ASAP7_75t_L g5691 ( 
.A1(n_4931),
.A2(n_5004),
.B1(n_5099),
.B2(n_5041),
.Y(n_5691)
);

INVx2_ASAP7_75t_L g5692 ( 
.A(n_4234),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_4434),
.Y(n_5693)
);

CKINVDCx14_ASAP7_75t_R g5694 ( 
.A(n_4844),
.Y(n_5694)
);

INVx1_ASAP7_75t_L g5695 ( 
.A(n_4434),
.Y(n_5695)
);

NAND2xp5_ASAP7_75t_L g5696 ( 
.A(n_4781),
.B(n_4827),
.Y(n_5696)
);

AOI21xp5_ASAP7_75t_L g5697 ( 
.A1(n_4224),
.A2(n_4231),
.B(n_4228),
.Y(n_5697)
);

AOI21xp5_ASAP7_75t_L g5698 ( 
.A1(n_4228),
.A2(n_4233),
.B(n_4231),
.Y(n_5698)
);

OAI21xp33_ASAP7_75t_L g5699 ( 
.A1(n_4233),
.A2(n_4239),
.B(n_4238),
.Y(n_5699)
);

INVx1_ASAP7_75t_SL g5700 ( 
.A(n_4948),
.Y(n_5700)
);

INVx1_ASAP7_75t_L g5701 ( 
.A(n_4435),
.Y(n_5701)
);

BUFx2_ASAP7_75t_L g5702 ( 
.A(n_4962),
.Y(n_5702)
);

AND2x2_ASAP7_75t_L g5703 ( 
.A(n_4650),
.B(n_4654),
.Y(n_5703)
);

OAI21xp5_ASAP7_75t_L g5704 ( 
.A1(n_4631),
.A2(n_4651),
.B(n_5065),
.Y(n_5704)
);

INVx3_ASAP7_75t_L g5705 ( 
.A(n_4587),
.Y(n_5705)
);

INVx2_ASAP7_75t_L g5706 ( 
.A(n_4244),
.Y(n_5706)
);

OR2x2_ASAP7_75t_L g5707 ( 
.A(n_4728),
.B(n_4782),
.Y(n_5707)
);

NOR2xp33_ASAP7_75t_L g5708 ( 
.A(n_4300),
.B(n_4743),
.Y(n_5708)
);

AOI21xp5_ASAP7_75t_L g5709 ( 
.A1(n_4238),
.A2(n_4240),
.B(n_4239),
.Y(n_5709)
);

AOI21xp5_ASAP7_75t_L g5710 ( 
.A1(n_4240),
.A2(n_4263),
.B(n_4252),
.Y(n_5710)
);

INVx1_ASAP7_75t_L g5711 ( 
.A(n_4435),
.Y(n_5711)
);

AOI22xp33_ASAP7_75t_L g5712 ( 
.A1(n_4890),
.A2(n_4560),
.B1(n_4952),
.B2(n_4797),
.Y(n_5712)
);

O2A1O1Ixp33_ASAP7_75t_L g5713 ( 
.A1(n_4631),
.A2(n_5025),
.B(n_4933),
.C(n_4640),
.Y(n_5713)
);

OR2x6_ASAP7_75t_SL g5714 ( 
.A(n_4688),
.B(n_4252),
.Y(n_5714)
);

AND2x2_ASAP7_75t_L g5715 ( 
.A(n_4650),
.B(n_4654),
.Y(n_5715)
);

INVx1_ASAP7_75t_L g5716 ( 
.A(n_4435),
.Y(n_5716)
);

O2A1O1Ixp33_ASAP7_75t_L g5717 ( 
.A1(n_5025),
.A2(n_4933),
.B(n_4640),
.C(n_4643),
.Y(n_5717)
);

AOI22xp5_ASAP7_75t_L g5718 ( 
.A1(n_4560),
.A2(n_4921),
.B1(n_4938),
.B2(n_4925),
.Y(n_5718)
);

AOI22xp33_ASAP7_75t_L g5719 ( 
.A1(n_4890),
.A2(n_4560),
.B1(n_4797),
.B2(n_4859),
.Y(n_5719)
);

AOI21xp5_ASAP7_75t_L g5720 ( 
.A1(n_4263),
.A2(n_4267),
.B(n_4264),
.Y(n_5720)
);

NAND2xp5_ASAP7_75t_L g5721 ( 
.A(n_4832),
.B(n_4846),
.Y(n_5721)
);

OA22x2_ASAP7_75t_L g5722 ( 
.A1(n_5101),
.A2(n_4931),
.B1(n_5041),
.B2(n_5004),
.Y(n_5722)
);

CKINVDCx5p33_ASAP7_75t_R g5723 ( 
.A(n_4975),
.Y(n_5723)
);

CKINVDCx20_ASAP7_75t_R g5724 ( 
.A(n_4844),
.Y(n_5724)
);

INVx2_ASAP7_75t_L g5725 ( 
.A(n_4249),
.Y(n_5725)
);

HB1xp67_ASAP7_75t_L g5726 ( 
.A(n_4206),
.Y(n_5726)
);

CKINVDCx5p33_ASAP7_75t_R g5727 ( 
.A(n_4237),
.Y(n_5727)
);

INVx1_ASAP7_75t_L g5728 ( 
.A(n_4444),
.Y(n_5728)
);

OAI22xp33_ASAP7_75t_L g5729 ( 
.A1(n_4757),
.A2(n_4688),
.B1(n_4453),
.B2(n_5099),
.Y(n_5729)
);

NAND2xp5_ASAP7_75t_L g5730 ( 
.A(n_4832),
.B(n_4846),
.Y(n_5730)
);

NAND2xp5_ASAP7_75t_L g5731 ( 
.A(n_4851),
.B(n_4857),
.Y(n_5731)
);

INVx4_ASAP7_75t_L g5732 ( 
.A(n_4416),
.Y(n_5732)
);

NAND2xp5_ASAP7_75t_L g5733 ( 
.A(n_4851),
.B(n_4857),
.Y(n_5733)
);

BUFx2_ASAP7_75t_L g5734 ( 
.A(n_5000),
.Y(n_5734)
);

INVx3_ASAP7_75t_L g5735 ( 
.A(n_4694),
.Y(n_5735)
);

AOI22xp33_ASAP7_75t_L g5736 ( 
.A1(n_4560),
.A2(n_4859),
.B1(n_4300),
.B2(n_4921),
.Y(n_5736)
);

BUFx2_ASAP7_75t_L g5737 ( 
.A(n_5000),
.Y(n_5737)
);

INVx3_ASAP7_75t_SL g5738 ( 
.A(n_4517),
.Y(n_5738)
);

NAND2xp5_ASAP7_75t_SL g5739 ( 
.A(n_4748),
.B(n_4767),
.Y(n_5739)
);

AOI22xp33_ASAP7_75t_L g5740 ( 
.A1(n_4560),
.A2(n_4938),
.B1(n_4979),
.B2(n_4944),
.Y(n_5740)
);

AOI21xp5_ASAP7_75t_L g5741 ( 
.A1(n_4264),
.A2(n_4282),
.B(n_4267),
.Y(n_5741)
);

INVx1_ASAP7_75t_L g5742 ( 
.A(n_4444),
.Y(n_5742)
);

INVx1_ASAP7_75t_L g5743 ( 
.A(n_4444),
.Y(n_5743)
);

AOI222xp33_ASAP7_75t_L g5744 ( 
.A1(n_4944),
.A2(n_4979),
.B1(n_4560),
.B2(n_4910),
.C1(n_4807),
.C2(n_4804),
.Y(n_5744)
);

NAND2xp5_ASAP7_75t_SL g5745 ( 
.A(n_4748),
.B(n_4767),
.Y(n_5745)
);

CKINVDCx20_ASAP7_75t_R g5746 ( 
.A(n_5011),
.Y(n_5746)
);

A2O1A1Ixp33_ASAP7_75t_L g5747 ( 
.A1(n_4884),
.A2(n_4854),
.B(n_4929),
.C(n_5049),
.Y(n_5747)
);

NOR2xp33_ASAP7_75t_L g5748 ( 
.A(n_4768),
.B(n_4770),
.Y(n_5748)
);

CKINVDCx20_ASAP7_75t_R g5749 ( 
.A(n_5011),
.Y(n_5749)
);

CKINVDCx5p33_ASAP7_75t_R g5750 ( 
.A(n_4237),
.Y(n_5750)
);

HB1xp67_ASAP7_75t_L g5751 ( 
.A(n_4206),
.Y(n_5751)
);

AND2x2_ASAP7_75t_L g5752 ( 
.A(n_4654),
.B(n_4728),
.Y(n_5752)
);

A2O1A1Ixp33_ASAP7_75t_L g5753 ( 
.A1(n_4884),
.A2(n_4854),
.B(n_4929),
.C(n_5049),
.Y(n_5753)
);

INVx1_ASAP7_75t_L g5754 ( 
.A(n_4448),
.Y(n_5754)
);

CKINVDCx11_ASAP7_75t_R g5755 ( 
.A(n_4422),
.Y(n_5755)
);

INVx2_ASAP7_75t_L g5756 ( 
.A(n_4249),
.Y(n_5756)
);

BUFx4f_ASAP7_75t_L g5757 ( 
.A(n_4537),
.Y(n_5757)
);

A2O1A1Ixp33_ASAP7_75t_L g5758 ( 
.A1(n_4905),
.A2(n_4910),
.B(n_4768),
.C(n_4726),
.Y(n_5758)
);

INVx3_ASAP7_75t_L g5759 ( 
.A(n_4694),
.Y(n_5759)
);

OR2x6_ASAP7_75t_L g5760 ( 
.A(n_4246),
.B(n_4351),
.Y(n_5760)
);

INVx2_ASAP7_75t_L g5761 ( 
.A(n_4249),
.Y(n_5761)
);

INVx4_ASAP7_75t_L g5762 ( 
.A(n_4416),
.Y(n_5762)
);

INVx2_ASAP7_75t_L g5763 ( 
.A(n_4249),
.Y(n_5763)
);

INVx1_ASAP7_75t_L g5764 ( 
.A(n_4448),
.Y(n_5764)
);

AND2x4_ASAP7_75t_L g5765 ( 
.A(n_4416),
.B(n_4490),
.Y(n_5765)
);

NAND2xp5_ASAP7_75t_L g5766 ( 
.A(n_4866),
.B(n_4895),
.Y(n_5766)
);

OAI22xp5_ASAP7_75t_L g5767 ( 
.A1(n_4636),
.A2(n_4647),
.B1(n_4653),
.B2(n_4643),
.Y(n_5767)
);

INVx1_ASAP7_75t_L g5768 ( 
.A(n_4448),
.Y(n_5768)
);

A2O1A1Ixp33_ASAP7_75t_L g5769 ( 
.A1(n_4905),
.A2(n_4726),
.B(n_5029),
.C(n_4872),
.Y(n_5769)
);

AND2x4_ASAP7_75t_L g5770 ( 
.A(n_4416),
.B(n_4490),
.Y(n_5770)
);

NOR2xp33_ASAP7_75t_R g5771 ( 
.A(n_4480),
.B(n_4517),
.Y(n_5771)
);

NAND3xp33_ASAP7_75t_L g5772 ( 
.A(n_4798),
.B(n_4946),
.C(n_4290),
.Y(n_5772)
);

AND2x4_ASAP7_75t_L g5773 ( 
.A(n_4416),
.B(n_4490),
.Y(n_5773)
);

INVx2_ASAP7_75t_L g5774 ( 
.A(n_4295),
.Y(n_5774)
);

NAND2xp5_ASAP7_75t_L g5775 ( 
.A(n_4866),
.B(n_4895),
.Y(n_5775)
);

OAI22xp5_ASAP7_75t_L g5776 ( 
.A1(n_4647),
.A2(n_4655),
.B1(n_4658),
.B2(n_4653),
.Y(n_5776)
);

AOI21xp33_ASAP7_75t_L g5777 ( 
.A1(n_4282),
.A2(n_4301),
.B(n_4290),
.Y(n_5777)
);

INVx1_ASAP7_75t_L g5778 ( 
.A(n_4456),
.Y(n_5778)
);

INVx1_ASAP7_75t_L g5779 ( 
.A(n_4456),
.Y(n_5779)
);

AOI22xp5_ASAP7_75t_L g5780 ( 
.A1(n_4560),
.A2(n_4557),
.B1(n_5101),
.B2(n_4757),
.Y(n_5780)
);

CKINVDCx6p67_ASAP7_75t_R g5781 ( 
.A(n_4817),
.Y(n_5781)
);

NAND2xp5_ASAP7_75t_L g5782 ( 
.A(n_4900),
.B(n_4908),
.Y(n_5782)
);

AOI21xp5_ASAP7_75t_L g5783 ( 
.A1(n_4301),
.A2(n_4310),
.B(n_4304),
.Y(n_5783)
);

INVx1_ASAP7_75t_L g5784 ( 
.A(n_4456),
.Y(n_5784)
);

OAI22x1_ASAP7_75t_L g5785 ( 
.A1(n_4182),
.A2(n_4207),
.B1(n_4183),
.B2(n_4782),
.Y(n_5785)
);

OR2x2_ASAP7_75t_L g5786 ( 
.A(n_4782),
.B(n_4876),
.Y(n_5786)
);

AND2x2_ASAP7_75t_L g5787 ( 
.A(n_4754),
.B(n_4756),
.Y(n_5787)
);

INVx1_ASAP7_75t_L g5788 ( 
.A(n_4457),
.Y(n_5788)
);

AOI22xp33_ASAP7_75t_L g5789 ( 
.A1(n_4560),
.A2(n_4798),
.B1(n_4946),
.B2(n_4537),
.Y(n_5789)
);

NAND2xp5_ASAP7_75t_L g5790 ( 
.A(n_4900),
.B(n_4908),
.Y(n_5790)
);

NOR2xp33_ASAP7_75t_L g5791 ( 
.A(n_4655),
.B(n_4658),
.Y(n_5791)
);

INVx1_ASAP7_75t_L g5792 ( 
.A(n_4457),
.Y(n_5792)
);

NAND2xp5_ASAP7_75t_L g5793 ( 
.A(n_4920),
.B(n_4958),
.Y(n_5793)
);

AND2x4_ASAP7_75t_L g5794 ( 
.A(n_4490),
.B(n_4520),
.Y(n_5794)
);

INVx4_ASAP7_75t_L g5795 ( 
.A(n_4490),
.Y(n_5795)
);

A2O1A1Ixp33_ASAP7_75t_L g5796 ( 
.A1(n_5029),
.A2(n_4872),
.B(n_4803),
.C(n_5079),
.Y(n_5796)
);

AND2x2_ASAP7_75t_L g5797 ( 
.A(n_4754),
.B(n_4756),
.Y(n_5797)
);

INVx1_ASAP7_75t_L g5798 ( 
.A(n_4457),
.Y(n_5798)
);

AOI21xp5_ASAP7_75t_L g5799 ( 
.A1(n_4304),
.A2(n_4312),
.B(n_4310),
.Y(n_5799)
);

OAI22xp5_ASAP7_75t_L g5800 ( 
.A1(n_4667),
.A2(n_4672),
.B1(n_4677),
.B2(n_4671),
.Y(n_5800)
);

O2A1O1Ixp33_ASAP7_75t_L g5801 ( 
.A1(n_4667),
.A2(n_4672),
.B(n_4677),
.C(n_4671),
.Y(n_5801)
);

OR2x2_ASAP7_75t_L g5802 ( 
.A(n_4876),
.B(n_4688),
.Y(n_5802)
);

NAND2xp5_ASAP7_75t_L g5803 ( 
.A(n_4920),
.B(n_4958),
.Y(n_5803)
);

INVxp67_ASAP7_75t_L g5804 ( 
.A(n_4399),
.Y(n_5804)
);

A2O1A1Ixp33_ASAP7_75t_L g5805 ( 
.A1(n_4803),
.A2(n_5079),
.B(n_4428),
.C(n_4328),
.Y(n_5805)
);

BUFx2_ASAP7_75t_L g5806 ( 
.A(n_5016),
.Y(n_5806)
);

INVx8_ASAP7_75t_L g5807 ( 
.A(n_4537),
.Y(n_5807)
);

INVx1_ASAP7_75t_SL g5808 ( 
.A(n_5021),
.Y(n_5808)
);

AND2x2_ASAP7_75t_L g5809 ( 
.A(n_4754),
.B(n_4756),
.Y(n_5809)
);

AOI22xp33_ASAP7_75t_L g5810 ( 
.A1(n_4560),
.A2(n_4798),
.B1(n_4537),
.B2(n_4858),
.Y(n_5810)
);

INVx4_ASAP7_75t_L g5811 ( 
.A(n_4490),
.Y(n_5811)
);

AOI21xp5_ASAP7_75t_L g5812 ( 
.A1(n_4312),
.A2(n_4319),
.B(n_4314),
.Y(n_5812)
);

INVx4_ASAP7_75t_L g5813 ( 
.A(n_4490),
.Y(n_5813)
);

INVx2_ASAP7_75t_L g5814 ( 
.A(n_4295),
.Y(n_5814)
);

INVxp67_ASAP7_75t_L g5815 ( 
.A(n_4399),
.Y(n_5815)
);

INVx2_ASAP7_75t_L g5816 ( 
.A(n_4309),
.Y(n_5816)
);

CKINVDCx11_ASAP7_75t_R g5817 ( 
.A(n_4422),
.Y(n_5817)
);

INVx4_ASAP7_75t_L g5818 ( 
.A(n_4490),
.Y(n_5818)
);

OAI22x1_ASAP7_75t_L g5819 ( 
.A1(n_4288),
.A2(n_4143),
.B1(n_4202),
.B2(n_4170),
.Y(n_5819)
);

INVxp67_ASAP7_75t_L g5820 ( 
.A(n_4400),
.Y(n_5820)
);

NAND2xp5_ASAP7_75t_L g5821 ( 
.A(n_4974),
.B(n_4986),
.Y(n_5821)
);

OR2x6_ASAP7_75t_L g5822 ( 
.A(n_4246),
.B(n_4351),
.Y(n_5822)
);

AND2x4_ASAP7_75t_L g5823 ( 
.A(n_4520),
.B(n_4523),
.Y(n_5823)
);

OAI22xp5_ASAP7_75t_L g5824 ( 
.A1(n_4822),
.A2(n_4833),
.B1(n_4835),
.B2(n_4828),
.Y(n_5824)
);

AOI21xp5_ASAP7_75t_L g5825 ( 
.A1(n_4314),
.A2(n_4325),
.B(n_4319),
.Y(n_5825)
);

AND2x4_ASAP7_75t_L g5826 ( 
.A(n_4520),
.B(n_4523),
.Y(n_5826)
);

NAND2xp5_ASAP7_75t_L g5827 ( 
.A(n_4974),
.B(n_4986),
.Y(n_5827)
);

NAND2xp5_ASAP7_75t_SL g5828 ( 
.A(n_4805),
.B(n_4683),
.Y(n_5828)
);

OAI22xp5_ASAP7_75t_L g5829 ( 
.A1(n_4822),
.A2(n_4833),
.B1(n_4835),
.B2(n_4828),
.Y(n_5829)
);

BUFx8_ASAP7_75t_L g5830 ( 
.A(n_4537),
.Y(n_5830)
);

OR2x2_ASAP7_75t_L g5831 ( 
.A(n_4876),
.B(n_4873),
.Y(n_5831)
);

OAI22xp5_ASAP7_75t_L g5832 ( 
.A1(n_4325),
.A2(n_4334),
.B1(n_4337),
.B2(n_4335),
.Y(n_5832)
);

BUFx6f_ASAP7_75t_SL g5833 ( 
.A(n_4537),
.Y(n_5833)
);

INVx2_ASAP7_75t_L g5834 ( 
.A(n_4309),
.Y(n_5834)
);

NAND2xp5_ASAP7_75t_L g5835 ( 
.A(n_4987),
.B(n_4997),
.Y(n_5835)
);

A2O1A1Ixp33_ASAP7_75t_SL g5836 ( 
.A1(n_4334),
.A2(n_4337),
.B(n_4342),
.C(n_4335),
.Y(n_5836)
);

OR2x2_ASAP7_75t_L g5837 ( 
.A(n_4873),
.B(n_4875),
.Y(n_5837)
);

NAND2xp5_ASAP7_75t_SL g5838 ( 
.A(n_4805),
.B(n_4683),
.Y(n_5838)
);

AOI22xp5_ASAP7_75t_L g5839 ( 
.A1(n_4560),
.A2(n_4557),
.B1(n_4453),
.B2(n_5104),
.Y(n_5839)
);

AOI22xp5_ASAP7_75t_L g5840 ( 
.A1(n_5104),
.A2(n_5078),
.B1(n_4807),
.B2(n_4804),
.Y(n_5840)
);

NAND2xp5_ASAP7_75t_L g5841 ( 
.A(n_4987),
.B(n_4997),
.Y(n_5841)
);

BUFx2_ASAP7_75t_L g5842 ( 
.A(n_5021),
.Y(n_5842)
);

O2A1O1Ixp33_ASAP7_75t_L g5843 ( 
.A1(n_4342),
.A2(n_4345),
.B(n_4348),
.C(n_4344),
.Y(n_5843)
);

HB1xp67_ASAP7_75t_L g5844 ( 
.A(n_5014),
.Y(n_5844)
);

INVx2_ASAP7_75t_L g5845 ( 
.A(n_4309),
.Y(n_5845)
);

INVxp67_ASAP7_75t_L g5846 ( 
.A(n_4400),
.Y(n_5846)
);

INVx2_ASAP7_75t_L g5847 ( 
.A(n_4313),
.Y(n_5847)
);

INVxp67_ASAP7_75t_L g5848 ( 
.A(n_4404),
.Y(n_5848)
);

NAND2xp5_ASAP7_75t_L g5849 ( 
.A(n_5014),
.B(n_5058),
.Y(n_5849)
);

INVx2_ASAP7_75t_L g5850 ( 
.A(n_4313),
.Y(n_5850)
);

CKINVDCx20_ASAP7_75t_R g5851 ( 
.A(n_4190),
.Y(n_5851)
);

O2A1O1Ixp5_ASAP7_75t_L g5852 ( 
.A1(n_4344),
.A2(n_4348),
.B(n_4355),
.C(n_4345),
.Y(n_5852)
);

NAND2xp5_ASAP7_75t_L g5853 ( 
.A(n_5058),
.B(n_5066),
.Y(n_5853)
);

AND2x4_ASAP7_75t_L g5854 ( 
.A(n_4520),
.B(n_4523),
.Y(n_5854)
);

AND2x4_ASAP7_75t_SL g5855 ( 
.A(n_4246),
.B(n_4417),
.Y(n_5855)
);

CKINVDCx16_ASAP7_75t_R g5856 ( 
.A(n_4982),
.Y(n_5856)
);

BUFx8_ASAP7_75t_L g5857 ( 
.A(n_4537),
.Y(n_5857)
);

O2A1O1Ixp5_ASAP7_75t_SL g5858 ( 
.A1(n_4154),
.A2(n_4167),
.B(n_4173),
.C(n_4157),
.Y(n_5858)
);

NAND2xp5_ASAP7_75t_L g5859 ( 
.A(n_5066),
.B(n_5071),
.Y(n_5859)
);

NOR3xp33_ASAP7_75t_L g5860 ( 
.A(n_4355),
.B(n_4358),
.C(n_4356),
.Y(n_5860)
);

INVx3_ASAP7_75t_L g5861 ( 
.A(n_4694),
.Y(n_5861)
);

CKINVDCx5p33_ASAP7_75t_R g5862 ( 
.A(n_4242),
.Y(n_5862)
);

HB1xp67_ASAP7_75t_L g5863 ( 
.A(n_5071),
.Y(n_5863)
);

AND2x2_ASAP7_75t_L g5864 ( 
.A(n_4776),
.B(n_4802),
.Y(n_5864)
);

BUFx12f_ASAP7_75t_L g5865 ( 
.A(n_4253),
.Y(n_5865)
);

AO22x1_ASAP7_75t_L g5866 ( 
.A1(n_4537),
.A2(n_4288),
.B1(n_4924),
.B2(n_4864),
.Y(n_5866)
);

A2O1A1Ixp33_ASAP7_75t_L g5867 ( 
.A1(n_4803),
.A2(n_4328),
.B(n_4428),
.C(n_4698),
.Y(n_5867)
);

AND2x2_ASAP7_75t_L g5868 ( 
.A(n_4776),
.B(n_4802),
.Y(n_5868)
);

NAND2x1p5_ASAP7_75t_L g5869 ( 
.A(n_4520),
.B(n_4523),
.Y(n_5869)
);

NAND2xp5_ASAP7_75t_SL g5870 ( 
.A(n_4635),
.B(n_4608),
.Y(n_5870)
);

NAND2xp5_ASAP7_75t_SL g5871 ( 
.A(n_4635),
.B(n_4608),
.Y(n_5871)
);

CKINVDCx14_ASAP7_75t_R g5872 ( 
.A(n_4978),
.Y(n_5872)
);

HB1xp67_ASAP7_75t_L g5873 ( 
.A(n_4638),
.Y(n_5873)
);

OR2x6_ASAP7_75t_L g5874 ( 
.A(n_4246),
.B(n_4351),
.Y(n_5874)
);

O2A1O1Ixp5_ASAP7_75t_L g5875 ( 
.A1(n_4356),
.A2(n_4359),
.B(n_4366),
.C(n_4358),
.Y(n_5875)
);

AOI22xp33_ASAP7_75t_L g5876 ( 
.A1(n_4537),
.A2(n_4858),
.B1(n_4922),
.B2(n_4909),
.Y(n_5876)
);

NAND2xp5_ASAP7_75t_SL g5877 ( 
.A(n_4570),
.B(n_5062),
.Y(n_5877)
);

AND2x6_ASAP7_75t_SL g5878 ( 
.A(n_4983),
.B(n_4996),
.Y(n_5878)
);

AOI22xp5_ASAP7_75t_L g5879 ( 
.A1(n_5078),
.A2(n_4909),
.B1(n_4968),
.B2(n_4922),
.Y(n_5879)
);

AND2x4_ASAP7_75t_L g5880 ( 
.A(n_4520),
.B(n_4523),
.Y(n_5880)
);

AOI22xp33_ASAP7_75t_L g5881 ( 
.A1(n_4968),
.A2(n_5050),
.B1(n_5063),
.B2(n_4999),
.Y(n_5881)
);

OR2x6_ASAP7_75t_L g5882 ( 
.A(n_4246),
.B(n_4351),
.Y(n_5882)
);

INVxp67_ASAP7_75t_L g5883 ( 
.A(n_4404),
.Y(n_5883)
);

A2O1A1Ixp33_ASAP7_75t_L g5884 ( 
.A1(n_4803),
.A2(n_4698),
.B(n_4766),
.C(n_4359),
.Y(n_5884)
);

INVx4_ASAP7_75t_L g5885 ( 
.A(n_4520),
.Y(n_5885)
);

OAI22xp33_ASAP7_75t_L g5886 ( 
.A1(n_4982),
.A2(n_4575),
.B1(n_4940),
.B2(n_4928),
.Y(n_5886)
);

AOI22xp5_ASAP7_75t_L g5887 ( 
.A1(n_4999),
.A2(n_5050),
.B1(n_5076),
.B2(n_5063),
.Y(n_5887)
);

AND2x2_ASAP7_75t_L g5888 ( 
.A(n_4776),
.B(n_4802),
.Y(n_5888)
);

BUFx2_ASAP7_75t_L g5889 ( 
.A(n_5022),
.Y(n_5889)
);

OAI22xp5_ASAP7_75t_L g5890 ( 
.A1(n_4366),
.A2(n_4390),
.B1(n_4397),
.B2(n_4378),
.Y(n_5890)
);

INVx3_ASAP7_75t_L g5891 ( 
.A(n_4694),
.Y(n_5891)
);

AND2x2_ASAP7_75t_SL g5892 ( 
.A(n_4899),
.B(n_4912),
.Y(n_5892)
);

INVx1_ASAP7_75t_SL g5893 ( 
.A(n_5022),
.Y(n_5893)
);

NAND2xp5_ASAP7_75t_L g5894 ( 
.A(n_4749),
.B(n_4774),
.Y(n_5894)
);

AOI21xp5_ASAP7_75t_L g5895 ( 
.A1(n_4378),
.A2(n_4397),
.B(n_4390),
.Y(n_5895)
);

HAxp5_ASAP7_75t_L g5896 ( 
.A(n_4816),
.B(n_4403),
.CON(n_5896),
.SN(n_5896)
);

BUFx4f_ASAP7_75t_SL g5897 ( 
.A(n_4817),
.Y(n_5897)
);

A2O1A1Ixp33_ASAP7_75t_L g5898 ( 
.A1(n_4803),
.A2(n_4766),
.B(n_4403),
.C(n_4415),
.Y(n_5898)
);

AOI22xp5_ASAP7_75t_L g5899 ( 
.A1(n_5076),
.A2(n_5085),
.B1(n_5064),
.B2(n_4575),
.Y(n_5899)
);

AND2x2_ASAP7_75t_L g5900 ( 
.A(n_4830),
.B(n_4269),
.Y(n_5900)
);

AND2x2_ASAP7_75t_L g5901 ( 
.A(n_4830),
.B(n_4269),
.Y(n_5901)
);

NOR2xp33_ASAP7_75t_SL g5902 ( 
.A(n_4340),
.B(n_4417),
.Y(n_5902)
);

OAI22x1_ASAP7_75t_L g5903 ( 
.A1(n_4288),
.A2(n_4143),
.B1(n_4202),
.B2(n_4170),
.Y(n_5903)
);

AOI22xp5_ASAP7_75t_L g5904 ( 
.A1(n_5085),
.A2(n_5064),
.B1(n_4810),
.B2(n_4834),
.Y(n_5904)
);

NAND2x1p5_ASAP7_75t_L g5905 ( 
.A(n_4520),
.B(n_4523),
.Y(n_5905)
);

O2A1O1Ixp33_ASAP7_75t_L g5906 ( 
.A1(n_4413),
.A2(n_4418),
.B(n_4439),
.C(n_4415),
.Y(n_5906)
);

NAND2xp5_ASAP7_75t_L g5907 ( 
.A(n_4749),
.B(n_4774),
.Y(n_5907)
);

CKINVDCx20_ASAP7_75t_R g5908 ( 
.A(n_4190),
.Y(n_5908)
);

NAND2xp5_ASAP7_75t_L g5909 ( 
.A(n_4413),
.B(n_4418),
.Y(n_5909)
);

OAI21xp33_ASAP7_75t_L g5910 ( 
.A1(n_4439),
.A2(n_4447),
.B(n_4441),
.Y(n_5910)
);

AOI21xp5_ASAP7_75t_L g5911 ( 
.A1(n_4441),
.A2(n_4452),
.B(n_4447),
.Y(n_5911)
);

OAI22xp5_ASAP7_75t_L g5912 ( 
.A1(n_4452),
.A2(n_4458),
.B1(n_4459),
.B2(n_4454),
.Y(n_5912)
);

NAND2xp5_ASAP7_75t_SL g5913 ( 
.A(n_4570),
.B(n_5062),
.Y(n_5913)
);

AOI22xp33_ASAP7_75t_SL g5914 ( 
.A1(n_4985),
.A2(n_4408),
.B1(n_4450),
.B2(n_4405),
.Y(n_5914)
);

NAND2xp5_ASAP7_75t_SL g5915 ( 
.A(n_5062),
.B(n_4451),
.Y(n_5915)
);

NAND2x1p5_ASAP7_75t_L g5916 ( 
.A(n_4523),
.B(n_4417),
.Y(n_5916)
);

AND2x4_ASAP7_75t_L g5917 ( 
.A(n_4523),
.B(n_4361),
.Y(n_5917)
);

HB1xp67_ASAP7_75t_L g5918 ( 
.A(n_4638),
.Y(n_5918)
);

NAND2xp5_ASAP7_75t_L g5919 ( 
.A(n_4454),
.B(n_4458),
.Y(n_5919)
);

BUFx2_ASAP7_75t_L g5920 ( 
.A(n_5037),
.Y(n_5920)
);

A2O1A1Ixp33_ASAP7_75t_SL g5921 ( 
.A1(n_4459),
.A2(n_4474),
.B(n_4478),
.C(n_4470),
.Y(n_5921)
);

NOR2xp33_ASAP7_75t_L g5922 ( 
.A(n_5097),
.B(n_4983),
.Y(n_5922)
);

HB1xp67_ASAP7_75t_L g5923 ( 
.A(n_4405),
.Y(n_5923)
);

NAND2xp5_ASAP7_75t_SL g5924 ( 
.A(n_5062),
.B(n_4451),
.Y(n_5924)
);

NAND2xp5_ASAP7_75t_L g5925 ( 
.A(n_4470),
.B(n_4474),
.Y(n_5925)
);

INVx1_ASAP7_75t_SL g5926 ( 
.A(n_5037),
.Y(n_5926)
);

AND2x4_ASAP7_75t_L g5927 ( 
.A(n_4523),
.B(n_4361),
.Y(n_5927)
);

O2A1O1Ixp33_ASAP7_75t_L g5928 ( 
.A1(n_4478),
.A2(n_4482),
.B(n_4489),
.C(n_4481),
.Y(n_5928)
);

NAND2xp5_ASAP7_75t_L g5929 ( 
.A(n_4481),
.B(n_4482),
.Y(n_5929)
);

NOR2xp33_ASAP7_75t_L g5930 ( 
.A(n_4996),
.B(n_5030),
.Y(n_5930)
);

NOR2xp33_ASAP7_75t_L g5931 ( 
.A(n_5030),
.B(n_5097),
.Y(n_5931)
);

O2A1O1Ixp5_ASAP7_75t_L g5932 ( 
.A1(n_4489),
.A2(n_4494),
.B(n_4495),
.C(n_4492),
.Y(n_5932)
);

A2O1A1Ixp33_ASAP7_75t_L g5933 ( 
.A1(n_4492),
.A2(n_4494),
.B(n_4498),
.C(n_4495),
.Y(n_5933)
);

AND2x2_ASAP7_75t_L g5934 ( 
.A(n_4830),
.B(n_4269),
.Y(n_5934)
);

OAI22xp5_ASAP7_75t_L g5935 ( 
.A1(n_4498),
.A2(n_4508),
.B1(n_4509),
.B2(n_4499),
.Y(n_5935)
);

AOI22xp33_ASAP7_75t_L g5936 ( 
.A1(n_4928),
.A2(n_4940),
.B1(n_4989),
.B2(n_4950),
.Y(n_5936)
);

OAI21xp5_ASAP7_75t_L g5937 ( 
.A1(n_4499),
.A2(n_4509),
.B(n_4508),
.Y(n_5937)
);

OAI21x1_ASAP7_75t_L g5938 ( 
.A1(n_4281),
.A2(n_4771),
.B(n_4596),
.Y(n_5938)
);

INVx1_ASAP7_75t_SL g5939 ( 
.A(n_5054),
.Y(n_5939)
);

O2A1O1Ixp5_ASAP7_75t_L g5940 ( 
.A1(n_4510),
.A2(n_4524),
.B(n_4534),
.C(n_4512),
.Y(n_5940)
);

BUFx8_ASAP7_75t_SL g5941 ( 
.A(n_4297),
.Y(n_5941)
);

NAND2xp5_ASAP7_75t_L g5942 ( 
.A(n_4510),
.B(n_4512),
.Y(n_5942)
);

NAND2xp5_ASAP7_75t_L g5943 ( 
.A(n_4524),
.B(n_4534),
.Y(n_5943)
);

BUFx8_ASAP7_75t_L g5944 ( 
.A(n_4817),
.Y(n_5944)
);

A2O1A1Ixp33_ASAP7_75t_L g5945 ( 
.A1(n_4539),
.A2(n_4540),
.B(n_4549),
.C(n_4541),
.Y(n_5945)
);

NAND2xp5_ASAP7_75t_L g5946 ( 
.A(n_4539),
.B(n_4540),
.Y(n_5946)
);

NAND2xp5_ASAP7_75t_L g5947 ( 
.A(n_4541),
.B(n_4549),
.Y(n_5947)
);

HB1xp67_ASAP7_75t_L g5948 ( 
.A(n_4408),
.Y(n_5948)
);

CKINVDCx5p33_ASAP7_75t_R g5949 ( 
.A(n_4242),
.Y(n_5949)
);

AND2x2_ASAP7_75t_L g5950 ( 
.A(n_4330),
.B(n_4333),
.Y(n_5950)
);

NOR2xp33_ASAP7_75t_L g5951 ( 
.A(n_4819),
.B(n_4821),
.Y(n_5951)
);

INVx8_ASAP7_75t_L g5952 ( 
.A(n_5077),
.Y(n_5952)
);

A2O1A1Ixp33_ASAP7_75t_L g5953 ( 
.A1(n_4550),
.A2(n_4268),
.B(n_4596),
.C(n_4585),
.Y(n_5953)
);

A2O1A1Ixp33_ASAP7_75t_L g5954 ( 
.A1(n_4550),
.A2(n_4268),
.B(n_4599),
.C(n_4585),
.Y(n_5954)
);

NAND2xp5_ASAP7_75t_L g5955 ( 
.A(n_4450),
.B(n_4465),
.Y(n_5955)
);

AOI22xp33_ASAP7_75t_L g5956 ( 
.A1(n_4928),
.A2(n_4950),
.B1(n_4989),
.B2(n_4940),
.Y(n_5956)
);

O2A1O1Ixp33_ASAP7_75t_L g5957 ( 
.A1(n_4599),
.A2(n_4607),
.B(n_4602),
.C(n_4465),
.Y(n_5957)
);

INVx4_ASAP7_75t_L g5958 ( 
.A(n_4623),
.Y(n_5958)
);

CKINVDCx20_ASAP7_75t_R g5959 ( 
.A(n_4260),
.Y(n_5959)
);

BUFx2_ASAP7_75t_L g5960 ( 
.A(n_5056),
.Y(n_5960)
);

CKINVDCx5p33_ASAP7_75t_R g5961 ( 
.A(n_4297),
.Y(n_5961)
);

AOI22xp33_ASAP7_75t_L g5962 ( 
.A1(n_4950),
.A2(n_4991),
.B1(n_5053),
.B2(n_4989),
.Y(n_5962)
);

INVx1_ASAP7_75t_SL g5963 ( 
.A(n_5056),
.Y(n_5963)
);

AND3x2_ASAP7_75t_L g5964 ( 
.A(n_4864),
.B(n_4924),
.C(n_4476),
.Y(n_5964)
);

AOI21xp5_ASAP7_75t_L g5965 ( 
.A1(n_4602),
.A2(n_4607),
.B(n_4287),
.Y(n_5965)
);

OAI22x1_ASAP7_75t_L g5966 ( 
.A1(n_4288),
.A2(n_4143),
.B1(n_4204),
.B2(n_4170),
.Y(n_5966)
);

INVxp67_ASAP7_75t_SL g5967 ( 
.A(n_4192),
.Y(n_5967)
);

AOI21xp5_ASAP7_75t_L g5968 ( 
.A1(n_4287),
.A2(n_5062),
.B(n_4752),
.Y(n_5968)
);

A2O1A1Ixp33_ASAP7_75t_SL g5969 ( 
.A1(n_4145),
.A2(n_4213),
.B(n_4259),
.C(n_4178),
.Y(n_5969)
);

BUFx12f_ASAP7_75t_L g5970 ( 
.A(n_4364),
.Y(n_5970)
);

OAI22xp5_ASAP7_75t_L g5971 ( 
.A1(n_4982),
.A2(n_4991),
.B1(n_5083),
.B2(n_5053),
.Y(n_5971)
);

NAND2xp5_ASAP7_75t_L g5972 ( 
.A(n_4491),
.B(n_4497),
.Y(n_5972)
);

NAND2xp5_ASAP7_75t_L g5973 ( 
.A(n_4491),
.B(n_4497),
.Y(n_5973)
);

OAI22x1_ASAP7_75t_L g5974 ( 
.A1(n_4204),
.A2(n_4302),
.B1(n_4446),
.B2(n_4332),
.Y(n_5974)
);

NAND2xp5_ASAP7_75t_L g5975 ( 
.A(n_4504),
.B(n_4513),
.Y(n_5975)
);

NAND2xp5_ASAP7_75t_L g5976 ( 
.A(n_4504),
.B(n_4513),
.Y(n_5976)
);

NAND2xp5_ASAP7_75t_SL g5977 ( 
.A(n_4451),
.B(n_4461),
.Y(n_5977)
);

A2O1A1Ixp33_ASAP7_75t_L g5978 ( 
.A1(n_4902),
.A2(n_4526),
.B(n_4930),
.C(n_4912),
.Y(n_5978)
);

NAND2xp5_ASAP7_75t_SL g5979 ( 
.A(n_4451),
.B(n_4461),
.Y(n_5979)
);

AND2x2_ASAP7_75t_L g5980 ( 
.A(n_4330),
.B(n_4333),
.Y(n_5980)
);

INVx3_ASAP7_75t_L g5981 ( 
.A(n_4708),
.Y(n_5981)
);

AND2x6_ASAP7_75t_L g5982 ( 
.A(n_4785),
.B(n_4839),
.Y(n_5982)
);

AOI22xp5_ASAP7_75t_L g5983 ( 
.A1(n_4799),
.A2(n_4814),
.B1(n_4849),
.B2(n_4834),
.Y(n_5983)
);

INVxp67_ASAP7_75t_L g5984 ( 
.A(n_4526),
.Y(n_5984)
);

OAI21x1_ASAP7_75t_SL g5985 ( 
.A1(n_4985),
.A2(n_4559),
.B(n_4462),
.Y(n_5985)
);

NOR2xp33_ASAP7_75t_SL g5986 ( 
.A(n_4340),
.B(n_4417),
.Y(n_5986)
);

HB1xp67_ASAP7_75t_L g5987 ( 
.A(n_4154),
.Y(n_5987)
);

AOI22xp5_ASAP7_75t_L g5988 ( 
.A1(n_4799),
.A2(n_4814),
.B1(n_4810),
.B2(n_4849),
.Y(n_5988)
);

INVx4_ASAP7_75t_L g5989 ( 
.A(n_4623),
.Y(n_5989)
);

BUFx12f_ASAP7_75t_L g5990 ( 
.A(n_4364),
.Y(n_5990)
);

AOI21xp5_ASAP7_75t_L g5991 ( 
.A1(n_4287),
.A2(n_4752),
.B(n_4745),
.Y(n_5991)
);

AND2x4_ASAP7_75t_L g5992 ( 
.A(n_4361),
.B(n_4382),
.Y(n_5992)
);

OAI22xp5_ASAP7_75t_L g5993 ( 
.A1(n_4991),
.A2(n_5083),
.B1(n_5053),
.B2(n_5040),
.Y(n_5993)
);

NOR2xp33_ASAP7_75t_L g5994 ( 
.A(n_4819),
.B(n_4821),
.Y(n_5994)
);

AO21x2_ASAP7_75t_L g5995 ( 
.A1(n_4737),
.A2(n_4740),
.B(n_4739),
.Y(n_5995)
);

AOI21xp5_ASAP7_75t_L g5996 ( 
.A1(n_4745),
.A2(n_4760),
.B(n_4752),
.Y(n_5996)
);

AOI21xp5_ASAP7_75t_L g5997 ( 
.A1(n_4745),
.A2(n_4763),
.B(n_4760),
.Y(n_5997)
);

BUFx2_ASAP7_75t_SL g5998 ( 
.A(n_4340),
.Y(n_5998)
);

A2O1A1Ixp33_ASAP7_75t_L g5999 ( 
.A1(n_4902),
.A2(n_4930),
.B(n_4912),
.C(n_4203),
.Y(n_5999)
);

AOI21xp5_ASAP7_75t_L g6000 ( 
.A1(n_4760),
.A2(n_4765),
.B(n_4763),
.Y(n_6000)
);

O2A1O1Ixp33_ASAP7_75t_L g6001 ( 
.A1(n_4808),
.A2(n_4818),
.B(n_4531),
.C(n_4565),
.Y(n_6001)
);

BUFx8_ASAP7_75t_L g6002 ( 
.A(n_4817),
.Y(n_6002)
);

OAI22xp5_ASAP7_75t_L g6003 ( 
.A1(n_5083),
.A2(n_5040),
.B1(n_4985),
.B2(n_4843),
.Y(n_6003)
);

A2O1A1Ixp33_ASAP7_75t_L g6004 ( 
.A1(n_4912),
.A2(n_4930),
.B(n_4203),
.C(n_4208),
.Y(n_6004)
);

NOR2xp33_ASAP7_75t_L g6005 ( 
.A(n_4887),
.B(n_4889),
.Y(n_6005)
);

BUFx3_ASAP7_75t_L g6006 ( 
.A(n_4483),
.Y(n_6006)
);

AND2x4_ASAP7_75t_L g6007 ( 
.A(n_4361),
.B(n_4382),
.Y(n_6007)
);

CKINVDCx14_ASAP7_75t_R g6008 ( 
.A(n_4978),
.Y(n_6008)
);

AND2x2_ASAP7_75t_L g6009 ( 
.A(n_4372),
.B(n_4388),
.Y(n_6009)
);

HB1xp67_ASAP7_75t_L g6010 ( 
.A(n_4154),
.Y(n_6010)
);

AOI21xp5_ASAP7_75t_L g6011 ( 
.A1(n_4763),
.A2(n_4769),
.B(n_4765),
.Y(n_6011)
);

NAND2xp5_ASAP7_75t_L g6012 ( 
.A(n_4808),
.B(n_4818),
.Y(n_6012)
);

INVx3_ASAP7_75t_L g6013 ( 
.A(n_4708),
.Y(n_6013)
);

A2O1A1Ixp33_ASAP7_75t_L g6014 ( 
.A1(n_4912),
.A2(n_4930),
.B(n_4203),
.C(n_4208),
.Y(n_6014)
);

O2A1O1Ixp33_ASAP7_75t_SL g6015 ( 
.A1(n_4586),
.A2(n_4260),
.B(n_4371),
.C(n_4265),
.Y(n_6015)
);

INVx3_ASAP7_75t_L g6016 ( 
.A(n_4755),
.Y(n_6016)
);

A2O1A1Ixp33_ASAP7_75t_L g6017 ( 
.A1(n_4930),
.A2(n_4203),
.B(n_4208),
.C(n_4199),
.Y(n_6017)
);

AND2x4_ASAP7_75t_L g6018 ( 
.A(n_4361),
.B(n_4382),
.Y(n_6018)
);

NAND2xp5_ASAP7_75t_L g6019 ( 
.A(n_4787),
.B(n_4791),
.Y(n_6019)
);

CKINVDCx5p33_ASAP7_75t_R g6020 ( 
.A(n_4376),
.Y(n_6020)
);

AOI222xp33_ASAP7_75t_L g6021 ( 
.A1(n_4887),
.A2(n_4889),
.B1(n_4903),
.B2(n_4906),
.C1(n_4904),
.C2(n_4893),
.Y(n_6021)
);

NAND2xp5_ASAP7_75t_SL g6022 ( 
.A(n_4451),
.B(n_4461),
.Y(n_6022)
);

AND2x4_ASAP7_75t_L g6023 ( 
.A(n_4361),
.B(n_4382),
.Y(n_6023)
);

NAND2xp5_ASAP7_75t_L g6024 ( 
.A(n_4787),
.B(n_4791),
.Y(n_6024)
);

INVx2_ASAP7_75t_SL g6025 ( 
.A(n_4623),
.Y(n_6025)
);

NAND2xp5_ASAP7_75t_SL g6026 ( 
.A(n_4461),
.B(n_4584),
.Y(n_6026)
);

INVx3_ASAP7_75t_L g6027 ( 
.A(n_4755),
.Y(n_6027)
);

AND2x2_ASAP7_75t_L g6028 ( 
.A(n_4372),
.B(n_4388),
.Y(n_6028)
);

INVx4_ASAP7_75t_L g6029 ( 
.A(n_4623),
.Y(n_6029)
);

A2O1A1Ixp33_ASAP7_75t_L g6030 ( 
.A1(n_4199),
.A2(n_4208),
.B(n_4211),
.C(n_4203),
.Y(n_6030)
);

AND2x4_ASAP7_75t_L g6031 ( 
.A(n_4382),
.B(n_4383),
.Y(n_6031)
);

NOR2x1_ASAP7_75t_L g6032 ( 
.A(n_4945),
.B(n_5009),
.Y(n_6032)
);

NAND2xp5_ASAP7_75t_L g6033 ( 
.A(n_4788),
.B(n_4789),
.Y(n_6033)
);

A2O1A1Ixp33_ASAP7_75t_SL g6034 ( 
.A1(n_4145),
.A2(n_4213),
.B(n_4259),
.C(n_4178),
.Y(n_6034)
);

INVxp67_ASAP7_75t_L g6035 ( 
.A(n_4192),
.Y(n_6035)
);

INVx1_ASAP7_75t_SL g6036 ( 
.A(n_5061),
.Y(n_6036)
);

AOI22xp33_ASAP7_75t_L g6037 ( 
.A1(n_4918),
.A2(n_4956),
.B1(n_4960),
.B2(n_4919),
.Y(n_6037)
);

AND2x4_ASAP7_75t_L g6038 ( 
.A(n_4382),
.B(n_4383),
.Y(n_6038)
);

AND2x2_ASAP7_75t_L g6039 ( 
.A(n_4372),
.B(n_4388),
.Y(n_6039)
);

NAND2xp5_ASAP7_75t_L g6040 ( 
.A(n_4788),
.B(n_4789),
.Y(n_6040)
);

INVx4_ASAP7_75t_L g6041 ( 
.A(n_4623),
.Y(n_6041)
);

A2O1A1Ixp33_ASAP7_75t_L g6042 ( 
.A1(n_4199),
.A2(n_4203),
.B(n_4211),
.C(n_4208),
.Y(n_6042)
);

INVxp67_ASAP7_75t_SL g6043 ( 
.A(n_4765),
.Y(n_6043)
);

NOR2xp67_ASAP7_75t_L g6044 ( 
.A(n_4737),
.B(n_4739),
.Y(n_6044)
);

AOI21xp5_ASAP7_75t_L g6045 ( 
.A1(n_4769),
.A2(n_4777),
.B(n_4775),
.Y(n_6045)
);

INVx3_ASAP7_75t_SL g6046 ( 
.A(n_4543),
.Y(n_6046)
);

CKINVDCx20_ASAP7_75t_R g6047 ( 
.A(n_4265),
.Y(n_6047)
);

A2O1A1Ixp33_ASAP7_75t_L g6048 ( 
.A1(n_4199),
.A2(n_4203),
.B(n_4211),
.C(n_4208),
.Y(n_6048)
);

O2A1O1Ixp5_ASAP7_75t_L g6049 ( 
.A1(n_4281),
.A2(n_4815),
.B(n_4755),
.C(n_5038),
.Y(n_6049)
);

BUFx2_ASAP7_75t_L g6050 ( 
.A(n_4402),
.Y(n_6050)
);

AOI22xp33_ASAP7_75t_L g6051 ( 
.A1(n_4913),
.A2(n_4980),
.B1(n_4990),
.B2(n_4973),
.Y(n_6051)
);

AOI21xp5_ASAP7_75t_L g6052 ( 
.A1(n_4769),
.A2(n_4777),
.B(n_4775),
.Y(n_6052)
);

AOI222xp33_ASAP7_75t_L g6053 ( 
.A1(n_4893),
.A2(n_4903),
.B1(n_4906),
.B2(n_4918),
.C1(n_4913),
.C2(n_4904),
.Y(n_6053)
);

INVxp67_ASAP7_75t_SL g6054 ( 
.A(n_4775),
.Y(n_6054)
);

AOI21xp5_ASAP7_75t_L g6055 ( 
.A1(n_4777),
.A2(n_4784),
.B(n_4780),
.Y(n_6055)
);

AOI22xp5_ASAP7_75t_L g6056 ( 
.A1(n_4919),
.A2(n_4926),
.B1(n_4927),
.B2(n_4923),
.Y(n_6056)
);

AND2x4_ASAP7_75t_L g6057 ( 
.A(n_4383),
.B(n_4385),
.Y(n_6057)
);

BUFx2_ASAP7_75t_L g6058 ( 
.A(n_4402),
.Y(n_6058)
);

OAI22xp5_ASAP7_75t_L g6059 ( 
.A1(n_4841),
.A2(n_4843),
.B1(n_4926),
.B2(n_4923),
.Y(n_6059)
);

INVx2_ASAP7_75t_SL g6060 ( 
.A(n_4623),
.Y(n_6060)
);

OAI22xp5_ASAP7_75t_SL g6061 ( 
.A1(n_4371),
.A2(n_4742),
.B1(n_4614),
.B2(n_4837),
.Y(n_6061)
);

NAND2xp5_ASAP7_75t_SL g6062 ( 
.A(n_4461),
.B(n_4584),
.Y(n_6062)
);

INVx2_ASAP7_75t_SL g6063 ( 
.A(n_4623),
.Y(n_6063)
);

OAI22xp5_ASAP7_75t_SL g6064 ( 
.A1(n_4614),
.A2(n_4742),
.B1(n_4874),
.B2(n_4837),
.Y(n_6064)
);

HB1xp67_ASAP7_75t_L g6065 ( 
.A(n_4157),
.Y(n_6065)
);

INVx8_ASAP7_75t_L g6066 ( 
.A(n_5077),
.Y(n_6066)
);

BUFx3_ASAP7_75t_L g6067 ( 
.A(n_4483),
.Y(n_6067)
);

INVx1_ASAP7_75t_SL g6068 ( 
.A(n_5061),
.Y(n_6068)
);

INVx3_ASAP7_75t_L g6069 ( 
.A(n_4755),
.Y(n_6069)
);

AND2x2_ASAP7_75t_L g6070 ( 
.A(n_4410),
.B(n_4445),
.Y(n_6070)
);

OAI22xp5_ASAP7_75t_L g6071 ( 
.A1(n_4841),
.A2(n_4943),
.B1(n_4949),
.B2(n_4927),
.Y(n_6071)
);

NOR2xp33_ASAP7_75t_R g6072 ( 
.A(n_4543),
.B(n_4632),
.Y(n_6072)
);

NOR2xp33_ASAP7_75t_L g6073 ( 
.A(n_4943),
.B(n_4949),
.Y(n_6073)
);

AOI21xp5_ASAP7_75t_L g6074 ( 
.A1(n_4780),
.A2(n_4790),
.B(n_4784),
.Y(n_6074)
);

AND2x4_ASAP7_75t_L g6075 ( 
.A(n_4383),
.B(n_4385),
.Y(n_6075)
);

OAI22xp5_ASAP7_75t_L g6076 ( 
.A1(n_4951),
.A2(n_4956),
.B1(n_4957),
.B2(n_4953),
.Y(n_6076)
);

BUFx2_ASAP7_75t_L g6077 ( 
.A(n_4438),
.Y(n_6077)
);

AOI22xp5_ASAP7_75t_L g6078 ( 
.A1(n_4951),
.A2(n_4957),
.B1(n_4960),
.B2(n_4953),
.Y(n_6078)
);

OAI22xp5_ASAP7_75t_L g6079 ( 
.A1(n_4966),
.A2(n_4970),
.B1(n_4971),
.B2(n_4967),
.Y(n_6079)
);

BUFx8_ASAP7_75t_L g6080 ( 
.A(n_4907),
.Y(n_6080)
);

OAI22xp5_ASAP7_75t_L g6081 ( 
.A1(n_4966),
.A2(n_4970),
.B1(n_4971),
.B2(n_4967),
.Y(n_6081)
);

AND2x4_ASAP7_75t_L g6082 ( 
.A(n_4383),
.B(n_4385),
.Y(n_6082)
);

INVx1_ASAP7_75t_SL g6083 ( 
.A(n_5068),
.Y(n_6083)
);

AOI22xp33_ASAP7_75t_L g6084 ( 
.A1(n_5032),
.A2(n_5057),
.B1(n_5075),
.B2(n_5034),
.Y(n_6084)
);

HB1xp67_ASAP7_75t_L g6085 ( 
.A(n_4157),
.Y(n_6085)
);

O2A1O1Ixp33_ASAP7_75t_L g6086 ( 
.A1(n_4531),
.A2(n_4565),
.B(n_4571),
.C(n_4554),
.Y(n_6086)
);

INVx1_ASAP7_75t_L g6087 ( 
.A(n_4511),
.Y(n_6087)
);

AOI21xp5_ASAP7_75t_L g6088 ( 
.A1(n_4780),
.A2(n_4790),
.B(n_4784),
.Y(n_6088)
);

BUFx3_ASAP7_75t_L g6089 ( 
.A(n_4483),
.Y(n_6089)
);

INVx2_ASAP7_75t_L g6090 ( 
.A(n_4365),
.Y(n_6090)
);

OAI22xp5_ASAP7_75t_L g6091 ( 
.A1(n_4973),
.A2(n_4977),
.B1(n_4980),
.B2(n_4976),
.Y(n_6091)
);

HB1xp67_ASAP7_75t_L g6092 ( 
.A(n_4167),
.Y(n_6092)
);

OAI21xp5_ASAP7_75t_L g6093 ( 
.A1(n_4554),
.A2(n_4571),
.B(n_4790),
.Y(n_6093)
);

O2A1O1Ixp33_ASAP7_75t_L g6094 ( 
.A1(n_4794),
.A2(n_4977),
.B(n_4984),
.C(n_4976),
.Y(n_6094)
);

AO32x2_ASAP7_75t_L g6095 ( 
.A1(n_4204),
.A2(n_4446),
.A3(n_4598),
.B1(n_4332),
.B2(n_4302),
.Y(n_6095)
);

CKINVDCx5p33_ASAP7_75t_R g6096 ( 
.A(n_4376),
.Y(n_6096)
);

INVx6_ASAP7_75t_L g6097 ( 
.A(n_4772),
.Y(n_6097)
);

CKINVDCx11_ASAP7_75t_R g6098 ( 
.A(n_4907),
.Y(n_6098)
);

INVx1_ASAP7_75t_L g6099 ( 
.A(n_4511),
.Y(n_6099)
);

CKINVDCx20_ASAP7_75t_R g6100 ( 
.A(n_4406),
.Y(n_6100)
);

O2A1O1Ixp33_ASAP7_75t_L g6101 ( 
.A1(n_4794),
.A2(n_4990),
.B(n_4998),
.C(n_4984),
.Y(n_6101)
);

INVx3_ASAP7_75t_L g6102 ( 
.A(n_4755),
.Y(n_6102)
);

CKINVDCx20_ASAP7_75t_R g6103 ( 
.A(n_4406),
.Y(n_6103)
);

AOI221xp5_ASAP7_75t_L g6104 ( 
.A1(n_4994),
.A2(n_5012),
.B1(n_5013),
.B2(n_5001),
.C(n_4998),
.Y(n_6104)
);

INVx2_ASAP7_75t_L g6105 ( 
.A(n_4367),
.Y(n_6105)
);

AOI22xp33_ASAP7_75t_L g6106 ( 
.A1(n_5019),
.A2(n_5089),
.B1(n_5072),
.B2(n_5001),
.Y(n_6106)
);

INVx1_ASAP7_75t_L g6107 ( 
.A(n_4518),
.Y(n_6107)
);

BUFx3_ASAP7_75t_L g6108 ( 
.A(n_4601),
.Y(n_6108)
);

AND2x2_ASAP7_75t_L g6109 ( 
.A(n_4410),
.B(n_4445),
.Y(n_6109)
);

INVx2_ASAP7_75t_L g6110 ( 
.A(n_4367),
.Y(n_6110)
);

INVx3_ASAP7_75t_L g6111 ( 
.A(n_4755),
.Y(n_6111)
);

INVx1_ASAP7_75t_SL g6112 ( 
.A(n_5068),
.Y(n_6112)
);

INVx2_ASAP7_75t_L g6113 ( 
.A(n_4367),
.Y(n_6113)
);

AOI22xp33_ASAP7_75t_L g6114 ( 
.A1(n_5013),
.A2(n_5039),
.B1(n_5075),
.B2(n_5032),
.Y(n_6114)
);

INVx2_ASAP7_75t_L g6115 ( 
.A(n_4367),
.Y(n_6115)
);

INVx3_ASAP7_75t_L g6116 ( 
.A(n_4815),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_4518),
.Y(n_6117)
);

NOR2xp33_ASAP7_75t_L g6118 ( 
.A(n_4994),
.B(n_5012),
.Y(n_6118)
);

CKINVDCx5p33_ASAP7_75t_R g6119 ( 
.A(n_4423),
.Y(n_6119)
);

INVx2_ASAP7_75t_L g6120 ( 
.A(n_4369),
.Y(n_6120)
);

NAND2xp5_ASAP7_75t_L g6121 ( 
.A(n_4656),
.B(n_4662),
.Y(n_6121)
);

NAND2xp5_ASAP7_75t_L g6122 ( 
.A(n_4656),
.B(n_4662),
.Y(n_6122)
);

AOI21x1_ASAP7_75t_L g6123 ( 
.A1(n_4167),
.A2(n_4174),
.B(n_4173),
.Y(n_6123)
);

O2A1O1Ixp5_ASAP7_75t_SL g6124 ( 
.A1(n_4173),
.A2(n_4174),
.B(n_4247),
.C(n_4232),
.Y(n_6124)
);

OAI22xp5_ASAP7_75t_L g6125 ( 
.A1(n_5017),
.A2(n_5019),
.B1(n_5027),
.B2(n_5018),
.Y(n_6125)
);

BUFx3_ASAP7_75t_L g6126 ( 
.A(n_4601),
.Y(n_6126)
);

NAND2xp5_ASAP7_75t_L g6127 ( 
.A(n_4656),
.B(n_4662),
.Y(n_6127)
);

AND2x4_ASAP7_75t_L g6128 ( 
.A(n_5174),
.B(n_5670),
.Y(n_6128)
);

OAI22xp5_ASAP7_75t_L g6129 ( 
.A1(n_5197),
.A2(n_5103),
.B1(n_5100),
.B2(n_5018),
.Y(n_6129)
);

INVx1_ASAP7_75t_L g6130 ( 
.A(n_5113),
.Y(n_6130)
);

AND2x2_ASAP7_75t_L g6131 ( 
.A(n_5687),
.B(n_4410),
.Y(n_6131)
);

BUFx3_ASAP7_75t_L g6132 ( 
.A(n_5672),
.Y(n_6132)
);

HB1xp67_ASAP7_75t_L g6133 ( 
.A(n_5109),
.Y(n_6133)
);

AND2x4_ASAP7_75t_SL g6134 ( 
.A(n_5571),
.B(n_4144),
.Y(n_6134)
);

INVx8_ASAP7_75t_L g6135 ( 
.A(n_5198),
.Y(n_6135)
);

INVx2_ASAP7_75t_L g6136 ( 
.A(n_5114),
.Y(n_6136)
);

BUFx6f_ASAP7_75t_L g6137 ( 
.A(n_5115),
.Y(n_6137)
);

INVx2_ASAP7_75t_L g6138 ( 
.A(n_5114),
.Y(n_6138)
);

INVx1_ASAP7_75t_L g6139 ( 
.A(n_5113),
.Y(n_6139)
);

INVx3_ASAP7_75t_L g6140 ( 
.A(n_5115),
.Y(n_6140)
);

NAND2x1p5_ASAP7_75t_L g6141 ( 
.A(n_5118),
.B(n_5757),
.Y(n_6141)
);

BUFx2_ASAP7_75t_SL g6142 ( 
.A(n_5438),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_5119),
.Y(n_6143)
);

INVx2_ASAP7_75t_L g6144 ( 
.A(n_5114),
.Y(n_6144)
);

BUFx2_ASAP7_75t_L g6145 ( 
.A(n_6095),
.Y(n_6145)
);

OAI22xp5_ASAP7_75t_L g6146 ( 
.A1(n_5197),
.A2(n_5607),
.B1(n_5626),
.B2(n_5270),
.Y(n_6146)
);

INVx3_ASAP7_75t_L g6147 ( 
.A(n_5115),
.Y(n_6147)
);

AOI21xp5_ASAP7_75t_L g6148 ( 
.A1(n_5965),
.A2(n_4794),
.B(n_4476),
.Y(n_6148)
);

BUFx6f_ASAP7_75t_L g6149 ( 
.A(n_5115),
.Y(n_6149)
);

INVx2_ASAP7_75t_L g6150 ( 
.A(n_5121),
.Y(n_6150)
);

NAND2xp5_ASAP7_75t_L g6151 ( 
.A(n_5791),
.B(n_4663),
.Y(n_6151)
);

INVx1_ASAP7_75t_SL g6152 ( 
.A(n_5528),
.Y(n_6152)
);

INVx2_ASAP7_75t_SL g6153 ( 
.A(n_5974),
.Y(n_6153)
);

CKINVDCx5p33_ASAP7_75t_R g6154 ( 
.A(n_5300),
.Y(n_6154)
);

AND2x2_ASAP7_75t_L g6155 ( 
.A(n_5687),
.B(n_4445),
.Y(n_6155)
);

INVx2_ASAP7_75t_SL g6156 ( 
.A(n_5974),
.Y(n_6156)
);

INVx1_ASAP7_75t_SL g6157 ( 
.A(n_5528),
.Y(n_6157)
);

AOI21xp5_ASAP7_75t_L g6158 ( 
.A1(n_5965),
.A2(n_5038),
.B(n_4584),
.Y(n_6158)
);

INVx3_ASAP7_75t_L g6159 ( 
.A(n_5115),
.Y(n_6159)
);

AOI22xp33_ASAP7_75t_L g6160 ( 
.A1(n_5607),
.A2(n_5027),
.B1(n_5028),
.B2(n_5017),
.Y(n_6160)
);

INVx3_ASAP7_75t_L g6161 ( 
.A(n_5115),
.Y(n_6161)
);

NAND2xp5_ASAP7_75t_L g6162 ( 
.A(n_5791),
.B(n_4663),
.Y(n_6162)
);

INVx2_ASAP7_75t_L g6163 ( 
.A(n_5121),
.Y(n_6163)
);

CKINVDCx5p33_ASAP7_75t_R g6164 ( 
.A(n_5300),
.Y(n_6164)
);

NOR2xp33_ASAP7_75t_L g6165 ( 
.A(n_5170),
.B(n_5042),
.Y(n_6165)
);

NOR2xp33_ASAP7_75t_L g6166 ( 
.A(n_5170),
.B(n_5042),
.Y(n_6166)
);

CKINVDCx20_ASAP7_75t_R g6167 ( 
.A(n_5229),
.Y(n_6167)
);

INVx1_ASAP7_75t_L g6168 ( 
.A(n_5119),
.Y(n_6168)
);

AOI22xp5_ASAP7_75t_L g6169 ( 
.A1(n_5645),
.A2(n_4847),
.B1(n_5034),
.B2(n_5028),
.Y(n_6169)
);

AND2x2_ASAP7_75t_SL g6170 ( 
.A(n_5118),
.B(n_4383),
.Y(n_6170)
);

AND2x2_ASAP7_75t_L g6171 ( 
.A(n_5687),
.B(n_4464),
.Y(n_6171)
);

NAND2xp5_ASAP7_75t_L g6172 ( 
.A(n_5860),
.B(n_4663),
.Y(n_6172)
);

AOI21xp5_ASAP7_75t_L g6173 ( 
.A1(n_5352),
.A2(n_5038),
.B(n_4584),
.Y(n_6173)
);

INVx1_ASAP7_75t_L g6174 ( 
.A(n_5126),
.Y(n_6174)
);

AOI21xp5_ASAP7_75t_L g6175 ( 
.A1(n_5352),
.A2(n_5038),
.B(n_4584),
.Y(n_6175)
);

HB1xp67_ASAP7_75t_L g6176 ( 
.A(n_5109),
.Y(n_6176)
);

BUFx6f_ASAP7_75t_L g6177 ( 
.A(n_5129),
.Y(n_6177)
);

AND2x2_ASAP7_75t_L g6178 ( 
.A(n_5436),
.B(n_4464),
.Y(n_6178)
);

BUFx6f_ASAP7_75t_L g6179 ( 
.A(n_5129),
.Y(n_6179)
);

BUFx2_ASAP7_75t_L g6180 ( 
.A(n_6095),
.Y(n_6180)
);

INVx1_ASAP7_75t_SL g6181 ( 
.A(n_5528),
.Y(n_6181)
);

CKINVDCx6p67_ASAP7_75t_R g6182 ( 
.A(n_5361),
.Y(n_6182)
);

OAI22xp5_ASAP7_75t_L g6183 ( 
.A1(n_5626),
.A2(n_5100),
.B1(n_5103),
.B2(n_5094),
.Y(n_6183)
);

AND2x2_ASAP7_75t_L g6184 ( 
.A(n_5436),
.B(n_4464),
.Y(n_6184)
);

CKINVDCx6p67_ASAP7_75t_R g6185 ( 
.A(n_5361),
.Y(n_6185)
);

INVx1_ASAP7_75t_L g6186 ( 
.A(n_5126),
.Y(n_6186)
);

INVx2_ASAP7_75t_L g6187 ( 
.A(n_5121),
.Y(n_6187)
);

CKINVDCx5p33_ASAP7_75t_R g6188 ( 
.A(n_5362),
.Y(n_6188)
);

AND2x2_ASAP7_75t_L g6189 ( 
.A(n_5436),
.B(n_4469),
.Y(n_6189)
);

OAI22xp5_ASAP7_75t_L g6190 ( 
.A1(n_5492),
.A2(n_5094),
.B1(n_5036),
.B2(n_5039),
.Y(n_6190)
);

AOI21xp5_ASAP7_75t_L g6191 ( 
.A1(n_5163),
.A2(n_5038),
.B(n_4771),
.Y(n_6191)
);

BUFx6f_ASAP7_75t_L g6192 ( 
.A(n_5129),
.Y(n_6192)
);

AND2x2_ASAP7_75t_L g6193 ( 
.A(n_5617),
.B(n_4469),
.Y(n_6193)
);

NAND2xp5_ASAP7_75t_L g6194 ( 
.A(n_5860),
.B(n_4665),
.Y(n_6194)
);

INVx4_ASAP7_75t_L g6195 ( 
.A(n_5964),
.Y(n_6195)
);

BUFx3_ASAP7_75t_L g6196 ( 
.A(n_5672),
.Y(n_6196)
);

CKINVDCx8_ASAP7_75t_R g6197 ( 
.A(n_5998),
.Y(n_6197)
);

INVx1_ASAP7_75t_L g6198 ( 
.A(n_5130),
.Y(n_6198)
);

AOI21xp5_ASAP7_75t_L g6199 ( 
.A1(n_5163),
.A2(n_4771),
.B(n_4203),
.Y(n_6199)
);

INVx3_ASAP7_75t_L g6200 ( 
.A(n_5129),
.Y(n_6200)
);

BUFx2_ASAP7_75t_L g6201 ( 
.A(n_6095),
.Y(n_6201)
);

NAND2xp5_ASAP7_75t_L g6202 ( 
.A(n_5634),
.B(n_4665),
.Y(n_6202)
);

AOI22xp33_ASAP7_75t_L g6203 ( 
.A1(n_5645),
.A2(n_5497),
.B1(n_5492),
.B2(n_5641),
.Y(n_6203)
);

INVx1_ASAP7_75t_L g6204 ( 
.A(n_5130),
.Y(n_6204)
);

NAND2xp5_ASAP7_75t_L g6205 ( 
.A(n_5634),
.B(n_5659),
.Y(n_6205)
);

AOI21xp5_ASAP7_75t_L g6206 ( 
.A1(n_5341),
.A2(n_4771),
.B(n_4203),
.Y(n_6206)
);

AOI21xp5_ASAP7_75t_L g6207 ( 
.A1(n_5341),
.A2(n_4208),
.B(n_4199),
.Y(n_6207)
);

INVx3_ASAP7_75t_L g6208 ( 
.A(n_5129),
.Y(n_6208)
);

OAI21x1_ASAP7_75t_SL g6209 ( 
.A1(n_5247),
.A2(n_4559),
.B(n_4945),
.Y(n_6209)
);

AND2x4_ASAP7_75t_L g6210 ( 
.A(n_5174),
.B(n_5670),
.Y(n_6210)
);

BUFx2_ASAP7_75t_L g6211 ( 
.A(n_6095),
.Y(n_6211)
);

INVx2_ASAP7_75t_L g6212 ( 
.A(n_5154),
.Y(n_6212)
);

BUFx6f_ASAP7_75t_L g6213 ( 
.A(n_5129),
.Y(n_6213)
);

INVx2_ASAP7_75t_L g6214 ( 
.A(n_5154),
.Y(n_6214)
);

BUFx6f_ASAP7_75t_L g6215 ( 
.A(n_5129),
.Y(n_6215)
);

AND2x4_ASAP7_75t_L g6216 ( 
.A(n_5670),
.B(n_4144),
.Y(n_6216)
);

AND2x2_ASAP7_75t_L g6217 ( 
.A(n_5617),
.B(n_4469),
.Y(n_6217)
);

BUFx3_ASAP7_75t_L g6218 ( 
.A(n_5672),
.Y(n_6218)
);

AND2x4_ASAP7_75t_L g6219 ( 
.A(n_5670),
.B(n_4144),
.Y(n_6219)
);

BUFx2_ASAP7_75t_L g6220 ( 
.A(n_6095),
.Y(n_6220)
);

NAND2xp5_ASAP7_75t_SL g6221 ( 
.A(n_5856),
.B(n_5370),
.Y(n_6221)
);

OR2x6_ASAP7_75t_L g6222 ( 
.A(n_5198),
.B(n_4351),
.Y(n_6222)
);

CKINVDCx5p33_ASAP7_75t_R g6223 ( 
.A(n_5362),
.Y(n_6223)
);

INVx1_ASAP7_75t_L g6224 ( 
.A(n_5136),
.Y(n_6224)
);

OAI22xp5_ASAP7_75t_L g6225 ( 
.A1(n_5640),
.A2(n_5036),
.B1(n_5043),
.B2(n_5035),
.Y(n_6225)
);

INVx1_ASAP7_75t_L g6226 ( 
.A(n_5136),
.Y(n_6226)
);

INVx3_ASAP7_75t_L g6227 ( 
.A(n_5135),
.Y(n_6227)
);

NAND2xp5_ASAP7_75t_L g6228 ( 
.A(n_5659),
.B(n_4665),
.Y(n_6228)
);

AOI22xp5_ASAP7_75t_L g6229 ( 
.A1(n_5497),
.A2(n_4847),
.B1(n_5043),
.B2(n_5035),
.Y(n_6229)
);

INVx2_ASAP7_75t_SL g6230 ( 
.A(n_5974),
.Y(n_6230)
);

HB1xp67_ASAP7_75t_L g6231 ( 
.A(n_5251),
.Y(n_6231)
);

INVx2_ASAP7_75t_L g6232 ( 
.A(n_5154),
.Y(n_6232)
);

AOI21xp5_ASAP7_75t_L g6233 ( 
.A1(n_5509),
.A2(n_4208),
.B(n_4199),
.Y(n_6233)
);

AND2x2_ASAP7_75t_L g6234 ( 
.A(n_5617),
.B(n_4488),
.Y(n_6234)
);

INVx3_ASAP7_75t_L g6235 ( 
.A(n_5135),
.Y(n_6235)
);

INVx5_ASAP7_75t_L g6236 ( 
.A(n_5264),
.Y(n_6236)
);

BUFx12f_ASAP7_75t_L g6237 ( 
.A(n_5361),
.Y(n_6237)
);

A2O1A1Ixp33_ASAP7_75t_L g6238 ( 
.A1(n_5538),
.A2(n_4199),
.B(n_4211),
.C(n_4208),
.Y(n_6238)
);

HB1xp67_ASAP7_75t_L g6239 ( 
.A(n_5251),
.Y(n_6239)
);

INVxp67_ASAP7_75t_SL g6240 ( 
.A(n_5432),
.Y(n_6240)
);

BUFx3_ASAP7_75t_L g6241 ( 
.A(n_5672),
.Y(n_6241)
);

INVx1_ASAP7_75t_L g6242 ( 
.A(n_5146),
.Y(n_6242)
);

AOI21xp5_ASAP7_75t_L g6243 ( 
.A1(n_5509),
.A2(n_4211),
.B(n_4199),
.Y(n_6243)
);

INVx2_ASAP7_75t_L g6244 ( 
.A(n_5191),
.Y(n_6244)
);

INVx2_ASAP7_75t_SL g6245 ( 
.A(n_5964),
.Y(n_6245)
);

INVx1_ASAP7_75t_L g6246 ( 
.A(n_5146),
.Y(n_6246)
);

INVx2_ASAP7_75t_L g6247 ( 
.A(n_5191),
.Y(n_6247)
);

INVx6_ASAP7_75t_L g6248 ( 
.A(n_5830),
.Y(n_6248)
);

A2O1A1Ixp33_ASAP7_75t_L g6249 ( 
.A1(n_5538),
.A2(n_5594),
.B(n_5247),
.C(n_5616),
.Y(n_6249)
);

BUFx6f_ASAP7_75t_L g6250 ( 
.A(n_5135),
.Y(n_6250)
);

INVx2_ASAP7_75t_L g6251 ( 
.A(n_5191),
.Y(n_6251)
);

AND2x4_ASAP7_75t_L g6252 ( 
.A(n_5670),
.B(n_4225),
.Y(n_6252)
);

AOI22xp5_ASAP7_75t_L g6253 ( 
.A1(n_5641),
.A2(n_4847),
.B1(n_5051),
.B2(n_5046),
.Y(n_6253)
);

INVx3_ASAP7_75t_L g6254 ( 
.A(n_5135),
.Y(n_6254)
);

NAND2x1p5_ASAP7_75t_L g6255 ( 
.A(n_5118),
.B(n_4225),
.Y(n_6255)
);

AND2x2_ASAP7_75t_L g6256 ( 
.A(n_5654),
.B(n_4488),
.Y(n_6256)
);

AND2x2_ASAP7_75t_L g6257 ( 
.A(n_5654),
.B(n_4488),
.Y(n_6257)
);

AOI21xp5_ASAP7_75t_L g6258 ( 
.A1(n_5116),
.A2(n_4211),
.B(n_4199),
.Y(n_6258)
);

CKINVDCx5p33_ASAP7_75t_R g6259 ( 
.A(n_5591),
.Y(n_6259)
);

INVx1_ASAP7_75t_SL g6260 ( 
.A(n_5642),
.Y(n_6260)
);

AOI22xp5_ASAP7_75t_L g6261 ( 
.A1(n_5627),
.A2(n_5051),
.B1(n_5057),
.B2(n_5046),
.Y(n_6261)
);

OAI22xp5_ASAP7_75t_L g6262 ( 
.A1(n_5640),
.A2(n_5619),
.B1(n_5740),
.B2(n_5627),
.Y(n_6262)
);

NOR2xp33_ASAP7_75t_L g6263 ( 
.A(n_5120),
.B(n_5048),
.Y(n_6263)
);

OAI22xp5_ASAP7_75t_L g6264 ( 
.A1(n_5619),
.A2(n_5740),
.B1(n_5655),
.B2(n_5718),
.Y(n_6264)
);

INVx3_ASAP7_75t_L g6265 ( 
.A(n_5135),
.Y(n_6265)
);

OR2x6_ASAP7_75t_SL g6266 ( 
.A(n_5971),
.B(n_4874),
.Y(n_6266)
);

BUFx6f_ASAP7_75t_L g6267 ( 
.A(n_5135),
.Y(n_6267)
);

INVx2_ASAP7_75t_L g6268 ( 
.A(n_5195),
.Y(n_6268)
);

BUFx3_ASAP7_75t_L g6269 ( 
.A(n_5672),
.Y(n_6269)
);

INVx1_ASAP7_75t_L g6270 ( 
.A(n_5156),
.Y(n_6270)
);

INVx2_ASAP7_75t_R g6271 ( 
.A(n_5370),
.Y(n_6271)
);

CKINVDCx5p33_ASAP7_75t_R g6272 ( 
.A(n_5222),
.Y(n_6272)
);

INVx3_ASAP7_75t_SL g6273 ( 
.A(n_5370),
.Y(n_6273)
);

INVx1_ASAP7_75t_L g6274 ( 
.A(n_5156),
.Y(n_6274)
);

INVx1_ASAP7_75t_L g6275 ( 
.A(n_5179),
.Y(n_6275)
);

INVx3_ASAP7_75t_L g6276 ( 
.A(n_5135),
.Y(n_6276)
);

CKINVDCx20_ASAP7_75t_R g6277 ( 
.A(n_5357),
.Y(n_6277)
);

AOI21xp5_ASAP7_75t_L g6278 ( 
.A1(n_5116),
.A2(n_5594),
.B(n_5632),
.Y(n_6278)
);

HB1xp67_ASAP7_75t_L g6279 ( 
.A(n_5293),
.Y(n_6279)
);

NAND2xp5_ASAP7_75t_L g6280 ( 
.A(n_5618),
.B(n_4674),
.Y(n_6280)
);

O2A1O1Ixp5_ASAP7_75t_L g6281 ( 
.A1(n_5457),
.A2(n_4178),
.B(n_4213),
.C(n_4145),
.Y(n_6281)
);

AOI21xp5_ASAP7_75t_L g6282 ( 
.A1(n_5632),
.A2(n_4230),
.B(n_4211),
.Y(n_6282)
);

OAI22xp5_ASAP7_75t_L g6283 ( 
.A1(n_5655),
.A2(n_5072),
.B1(n_5080),
.B2(n_5070),
.Y(n_6283)
);

NAND2xp5_ASAP7_75t_L g6284 ( 
.A(n_5618),
.B(n_4674),
.Y(n_6284)
);

BUFx5_ASAP7_75t_L g6285 ( 
.A(n_5765),
.Y(n_6285)
);

INVx2_ASAP7_75t_L g6286 ( 
.A(n_5195),
.Y(n_6286)
);

NAND2xp5_ASAP7_75t_L g6287 ( 
.A(n_5620),
.B(n_4674),
.Y(n_6287)
);

INVx2_ASAP7_75t_L g6288 ( 
.A(n_5195),
.Y(n_6288)
);

OAI22xp5_ASAP7_75t_L g6289 ( 
.A1(n_5718),
.A2(n_5683),
.B1(n_5839),
.B2(n_5736),
.Y(n_6289)
);

AOI21xp5_ASAP7_75t_L g6290 ( 
.A1(n_5123),
.A2(n_4230),
.B(n_4211),
.Y(n_6290)
);

INVx1_ASAP7_75t_L g6291 ( 
.A(n_5179),
.Y(n_6291)
);

INVx1_ASAP7_75t_SL g6292 ( 
.A(n_5642),
.Y(n_6292)
);

AOI221xp5_ASAP7_75t_L g6293 ( 
.A1(n_5237),
.A2(n_5081),
.B1(n_5082),
.B2(n_5080),
.C(n_5070),
.Y(n_6293)
);

AOI21xp5_ASAP7_75t_L g6294 ( 
.A1(n_5123),
.A2(n_5629),
.B(n_5991),
.Y(n_6294)
);

HB1xp67_ASAP7_75t_L g6295 ( 
.A(n_5293),
.Y(n_6295)
);

AOI21xp5_ASAP7_75t_L g6296 ( 
.A1(n_5629),
.A2(n_4230),
.B(n_4211),
.Y(n_6296)
);

BUFx6f_ASAP7_75t_L g6297 ( 
.A(n_5140),
.Y(n_6297)
);

INVx1_ASAP7_75t_L g6298 ( 
.A(n_5189),
.Y(n_6298)
);

BUFx2_ASAP7_75t_L g6299 ( 
.A(n_6095),
.Y(n_6299)
);

INVx1_ASAP7_75t_L g6300 ( 
.A(n_5189),
.Y(n_6300)
);

INVx2_ASAP7_75t_L g6301 ( 
.A(n_5210),
.Y(n_6301)
);

O2A1O1Ixp33_ASAP7_75t_L g6302 ( 
.A1(n_5367),
.A2(n_4737),
.B(n_4740),
.C(n_4739),
.Y(n_6302)
);

AOI22xp5_ASAP7_75t_L g6303 ( 
.A1(n_5691),
.A2(n_5082),
.B1(n_5087),
.B2(n_5081),
.Y(n_6303)
);

AND2x4_ASAP7_75t_L g6304 ( 
.A(n_5673),
.B(n_4225),
.Y(n_6304)
);

AOI22xp33_ASAP7_75t_L g6305 ( 
.A1(n_5691),
.A2(n_5088),
.B1(n_5089),
.B2(n_5087),
.Y(n_6305)
);

AOI222xp33_ASAP7_75t_L g6306 ( 
.A1(n_5186),
.A2(n_4586),
.B1(n_5088),
.B2(n_5092),
.C1(n_5090),
.C2(n_4885),
.Y(n_6306)
);

BUFx2_ASAP7_75t_L g6307 ( 
.A(n_6095),
.Y(n_6307)
);

INVx1_ASAP7_75t_L g6308 ( 
.A(n_5190),
.Y(n_6308)
);

INVx5_ASAP7_75t_L g6309 ( 
.A(n_5264),
.Y(n_6309)
);

BUFx3_ASAP7_75t_L g6310 ( 
.A(n_5672),
.Y(n_6310)
);

OAI21x1_ASAP7_75t_L g6311 ( 
.A1(n_5938),
.A2(n_4744),
.B(n_4740),
.Y(n_6311)
);

INVx1_ASAP7_75t_L g6312 ( 
.A(n_5190),
.Y(n_6312)
);

AND2x4_ASAP7_75t_L g6313 ( 
.A(n_5673),
.B(n_4225),
.Y(n_6313)
);

INVxp67_ASAP7_75t_L g6314 ( 
.A(n_5714),
.Y(n_6314)
);

BUFx3_ASAP7_75t_L g6315 ( 
.A(n_5672),
.Y(n_6315)
);

INVx1_ASAP7_75t_L g6316 ( 
.A(n_5194),
.Y(n_6316)
);

NAND2xp5_ASAP7_75t_SL g6317 ( 
.A(n_5856),
.B(n_4302),
.Y(n_6317)
);

INVx2_ASAP7_75t_L g6318 ( 
.A(n_5210),
.Y(n_6318)
);

BUFx2_ASAP7_75t_SL g6319 ( 
.A(n_5438),
.Y(n_6319)
);

AOI21xp5_ASAP7_75t_L g6320 ( 
.A1(n_5991),
.A2(n_4235),
.B(n_4230),
.Y(n_6320)
);

INVx2_ASAP7_75t_L g6321 ( 
.A(n_5210),
.Y(n_6321)
);

NAND2xp5_ASAP7_75t_L g6322 ( 
.A(n_5620),
.B(n_4675),
.Y(n_6322)
);

INVx1_ASAP7_75t_L g6323 ( 
.A(n_5194),
.Y(n_6323)
);

INVx2_ASAP7_75t_L g6324 ( 
.A(n_5218),
.Y(n_6324)
);

INVx3_ASAP7_75t_L g6325 ( 
.A(n_5149),
.Y(n_6325)
);

O2A1O1Ixp33_ASAP7_75t_L g6326 ( 
.A1(n_5237),
.A2(n_4744),
.B(n_5092),
.C(n_5090),
.Y(n_6326)
);

AND2x2_ASAP7_75t_L g6327 ( 
.A(n_5654),
.B(n_4502),
.Y(n_6327)
);

AOI21xp5_ASAP7_75t_L g6328 ( 
.A1(n_5633),
.A2(n_4235),
.B(n_4230),
.Y(n_6328)
);

INVx3_ASAP7_75t_L g6329 ( 
.A(n_5149),
.Y(n_6329)
);

INVx1_ASAP7_75t_L g6330 ( 
.A(n_5204),
.Y(n_6330)
);

NAND2xp5_ASAP7_75t_L g6331 ( 
.A(n_5933),
.B(n_5945),
.Y(n_6331)
);

INVx1_ASAP7_75t_L g6332 ( 
.A(n_5204),
.Y(n_6332)
);

NAND2xp5_ASAP7_75t_L g6333 ( 
.A(n_5613),
.B(n_5614),
.Y(n_6333)
);

AND2x2_ASAP7_75t_SL g6334 ( 
.A(n_5118),
.B(n_4385),
.Y(n_6334)
);

INVx2_ASAP7_75t_SL g6335 ( 
.A(n_5992),
.Y(n_6335)
);

INVx1_ASAP7_75t_L g6336 ( 
.A(n_5214),
.Y(n_6336)
);

INVx2_ASAP7_75t_L g6337 ( 
.A(n_5218),
.Y(n_6337)
);

AOI21xp5_ASAP7_75t_L g6338 ( 
.A1(n_5633),
.A2(n_5636),
.B(n_5651),
.Y(n_6338)
);

BUFx12f_ASAP7_75t_L g6339 ( 
.A(n_5463),
.Y(n_6339)
);

BUFx2_ASAP7_75t_L g6340 ( 
.A(n_5635),
.Y(n_6340)
);

INVx2_ASAP7_75t_L g6341 ( 
.A(n_5218),
.Y(n_6341)
);

INVx1_ASAP7_75t_L g6342 ( 
.A(n_5214),
.Y(n_6342)
);

NOR2xp33_ASAP7_75t_L g6343 ( 
.A(n_5120),
.B(n_5048),
.Y(n_6343)
);

HB1xp67_ASAP7_75t_L g6344 ( 
.A(n_5303),
.Y(n_6344)
);

INVx3_ASAP7_75t_L g6345 ( 
.A(n_5149),
.Y(n_6345)
);

CKINVDCx20_ASAP7_75t_R g6346 ( 
.A(n_5746),
.Y(n_6346)
);

NAND2x1p5_ASAP7_75t_L g6347 ( 
.A(n_5757),
.B(n_4225),
.Y(n_6347)
);

AND2x2_ASAP7_75t_L g6348 ( 
.A(n_5787),
.B(n_4502),
.Y(n_6348)
);

INVx1_ASAP7_75t_L g6349 ( 
.A(n_5230),
.Y(n_6349)
);

AND2x2_ASAP7_75t_L g6350 ( 
.A(n_5787),
.B(n_4502),
.Y(n_6350)
);

AOI22xp33_ASAP7_75t_L g6351 ( 
.A1(n_5691),
.A2(n_4885),
.B1(n_4883),
.B2(n_4877),
.Y(n_6351)
);

NAND2x1p5_ASAP7_75t_L g6352 ( 
.A(n_5757),
.B(n_4229),
.Y(n_6352)
);

CKINVDCx5p33_ASAP7_75t_R g6353 ( 
.A(n_5222),
.Y(n_6353)
);

AOI22xp33_ASAP7_75t_L g6354 ( 
.A1(n_5691),
.A2(n_4883),
.B1(n_4877),
.B2(n_4880),
.Y(n_6354)
);

NOR2x1_ASAP7_75t_SL g6355 ( 
.A(n_5457),
.B(n_5074),
.Y(n_6355)
);

BUFx3_ASAP7_75t_L g6356 ( 
.A(n_5672),
.Y(n_6356)
);

INVx2_ASAP7_75t_L g6357 ( 
.A(n_5228),
.Y(n_6357)
);

BUFx3_ASAP7_75t_L g6358 ( 
.A(n_5672),
.Y(n_6358)
);

INVx4_ASAP7_75t_L g6359 ( 
.A(n_5757),
.Y(n_6359)
);

CKINVDCx12_ASAP7_75t_R g6360 ( 
.A(n_6061),
.Y(n_6360)
);

INVx3_ASAP7_75t_L g6361 ( 
.A(n_5149),
.Y(n_6361)
);

AOI22xp33_ASAP7_75t_L g6362 ( 
.A1(n_5722),
.A2(n_5133),
.B1(n_5382),
.B2(n_5186),
.Y(n_6362)
);

NAND2xp5_ASAP7_75t_L g6363 ( 
.A(n_5613),
.B(n_4675),
.Y(n_6363)
);

OR2x2_ASAP7_75t_L g6364 ( 
.A(n_5802),
.B(n_5707),
.Y(n_6364)
);

INVx1_ASAP7_75t_L g6365 ( 
.A(n_5230),
.Y(n_6365)
);

AOI22xp5_ASAP7_75t_L g6366 ( 
.A1(n_5722),
.A2(n_4880),
.B1(n_4878),
.B2(n_4627),
.Y(n_6366)
);

INVx3_ASAP7_75t_L g6367 ( 
.A(n_5153),
.Y(n_6367)
);

INVx1_ASAP7_75t_L g6368 ( 
.A(n_5242),
.Y(n_6368)
);

INVx2_ASAP7_75t_L g6369 ( 
.A(n_5228),
.Y(n_6369)
);

BUFx2_ASAP7_75t_L g6370 ( 
.A(n_5635),
.Y(n_6370)
);

AOI21xp5_ASAP7_75t_L g6371 ( 
.A1(n_5636),
.A2(n_4235),
.B(n_4230),
.Y(n_6371)
);

NAND2xp5_ASAP7_75t_L g6372 ( 
.A(n_5614),
.B(n_4675),
.Y(n_6372)
);

INVx2_ASAP7_75t_L g6373 ( 
.A(n_5228),
.Y(n_6373)
);

BUFx2_ASAP7_75t_L g6374 ( 
.A(n_5635),
.Y(n_6374)
);

INVx2_ASAP7_75t_L g6375 ( 
.A(n_5240),
.Y(n_6375)
);

INVx1_ASAP7_75t_L g6376 ( 
.A(n_5242),
.Y(n_6376)
);

AOI22xp33_ASAP7_75t_SL g6377 ( 
.A1(n_5722),
.A2(n_4235),
.B1(n_4241),
.B2(n_4230),
.Y(n_6377)
);

BUFx3_ASAP7_75t_L g6378 ( 
.A(n_5982),
.Y(n_6378)
);

AOI22xp5_ASAP7_75t_L g6379 ( 
.A1(n_5722),
.A2(n_4878),
.B1(n_4627),
.B2(n_4634),
.Y(n_6379)
);

CKINVDCx5p33_ASAP7_75t_R g6380 ( 
.A(n_5463),
.Y(n_6380)
);

INVx1_ASAP7_75t_L g6381 ( 
.A(n_5252),
.Y(n_6381)
);

BUFx2_ASAP7_75t_L g6382 ( 
.A(n_5635),
.Y(n_6382)
);

BUFx12f_ASAP7_75t_L g6383 ( 
.A(n_5463),
.Y(n_6383)
);

BUFx2_ASAP7_75t_L g6384 ( 
.A(n_5635),
.Y(n_6384)
);

INVx1_ASAP7_75t_SL g6385 ( 
.A(n_5642),
.Y(n_6385)
);

BUFx3_ASAP7_75t_L g6386 ( 
.A(n_5982),
.Y(n_6386)
);

BUFx2_ASAP7_75t_L g6387 ( 
.A(n_5635),
.Y(n_6387)
);

AOI21xp5_ASAP7_75t_L g6388 ( 
.A1(n_5651),
.A2(n_4235),
.B(n_4230),
.Y(n_6388)
);

BUFx3_ASAP7_75t_L g6389 ( 
.A(n_5982),
.Y(n_6389)
);

INVx1_ASAP7_75t_L g6390 ( 
.A(n_5252),
.Y(n_6390)
);

OAI22xp5_ASAP7_75t_L g6391 ( 
.A1(n_5683),
.A2(n_4875),
.B1(n_4601),
.B2(n_4332),
.Y(n_6391)
);

INVx2_ASAP7_75t_L g6392 ( 
.A(n_5240),
.Y(n_6392)
);

NOR2xp33_ASAP7_75t_L g6393 ( 
.A(n_5748),
.B(n_5451),
.Y(n_6393)
);

CKINVDCx5p33_ASAP7_75t_R g6394 ( 
.A(n_5531),
.Y(n_6394)
);

INVx2_ASAP7_75t_SL g6395 ( 
.A(n_5992),
.Y(n_6395)
);

OAI22xp5_ASAP7_75t_L g6396 ( 
.A1(n_5839),
.A2(n_4332),
.B1(n_4446),
.B2(n_4302),
.Y(n_6396)
);

INVx1_ASAP7_75t_L g6397 ( 
.A(n_5254),
.Y(n_6397)
);

AOI22xp5_ASAP7_75t_L g6398 ( 
.A1(n_5133),
.A2(n_4613),
.B1(n_4634),
.B2(n_4576),
.Y(n_6398)
);

CKINVDCx5p33_ASAP7_75t_R g6399 ( 
.A(n_5531),
.Y(n_6399)
);

INVx3_ASAP7_75t_L g6400 ( 
.A(n_5153),
.Y(n_6400)
);

NAND2xp5_ASAP7_75t_L g6401 ( 
.A(n_5699),
.B(n_4680),
.Y(n_6401)
);

OR2x6_ASAP7_75t_L g6402 ( 
.A(n_5198),
.B(n_4351),
.Y(n_6402)
);

AOI22xp33_ASAP7_75t_L g6403 ( 
.A1(n_5382),
.A2(n_5111),
.B1(n_5311),
.B2(n_5744),
.Y(n_6403)
);

INVx1_ASAP7_75t_L g6404 ( 
.A(n_5254),
.Y(n_6404)
);

BUFx3_ASAP7_75t_L g6405 ( 
.A(n_5982),
.Y(n_6405)
);

NAND2xp5_ASAP7_75t_L g6406 ( 
.A(n_5699),
.B(n_5910),
.Y(n_6406)
);

AOI22xp33_ASAP7_75t_SL g6407 ( 
.A1(n_5221),
.A2(n_4235),
.B1(n_4241),
.B2(n_4230),
.Y(n_6407)
);

HB1xp67_ASAP7_75t_L g6408 ( 
.A(n_5303),
.Y(n_6408)
);

AOI22xp5_ASAP7_75t_L g6409 ( 
.A1(n_5744),
.A2(n_4613),
.B1(n_4576),
.B2(n_4611),
.Y(n_6409)
);

AOI21xp5_ASAP7_75t_L g6410 ( 
.A1(n_5772),
.A2(n_5789),
.B(n_5443),
.Y(n_6410)
);

NAND2xp5_ASAP7_75t_L g6411 ( 
.A(n_5910),
.B(n_4680),
.Y(n_6411)
);

AND2x2_ASAP7_75t_SL g6412 ( 
.A(n_5892),
.B(n_4424),
.Y(n_6412)
);

INVx1_ASAP7_75t_SL g6413 ( 
.A(n_5152),
.Y(n_6413)
);

NAND2xp5_ASAP7_75t_L g6414 ( 
.A(n_5767),
.B(n_4680),
.Y(n_6414)
);

INVx1_ASAP7_75t_L g6415 ( 
.A(n_5256),
.Y(n_6415)
);

INVx1_ASAP7_75t_L g6416 ( 
.A(n_5256),
.Y(n_6416)
);

BUFx6f_ASAP7_75t_SL g6417 ( 
.A(n_5892),
.Y(n_6417)
);

INVx1_ASAP7_75t_SL g6418 ( 
.A(n_5152),
.Y(n_6418)
);

AND2x2_ASAP7_75t_L g6419 ( 
.A(n_5787),
.B(n_4503),
.Y(n_6419)
);

INVx1_ASAP7_75t_L g6420 ( 
.A(n_5258),
.Y(n_6420)
);

INVx1_ASAP7_75t_L g6421 ( 
.A(n_5258),
.Y(n_6421)
);

BUFx10_ASAP7_75t_L g6422 ( 
.A(n_5187),
.Y(n_6422)
);

AND2x2_ASAP7_75t_L g6423 ( 
.A(n_5797),
.B(n_4503),
.Y(n_6423)
);

OR2x2_ASAP7_75t_L g6424 ( 
.A(n_5802),
.B(n_4545),
.Y(n_6424)
);

INVx2_ASAP7_75t_SL g6425 ( 
.A(n_5992),
.Y(n_6425)
);

HB1xp67_ASAP7_75t_L g6426 ( 
.A(n_5321),
.Y(n_6426)
);

CKINVDCx5p33_ASAP7_75t_R g6427 ( 
.A(n_5531),
.Y(n_6427)
);

BUFx12f_ASAP7_75t_L g6428 ( 
.A(n_5598),
.Y(n_6428)
);

HB1xp67_ASAP7_75t_L g6429 ( 
.A(n_5321),
.Y(n_6429)
);

INVx4_ASAP7_75t_L g6430 ( 
.A(n_5982),
.Y(n_6430)
);

AOI22xp33_ASAP7_75t_L g6431 ( 
.A1(n_5111),
.A2(n_5311),
.B1(n_5297),
.B2(n_5348),
.Y(n_6431)
);

AOI21xp5_ASAP7_75t_L g6432 ( 
.A1(n_5772),
.A2(n_4241),
.B(n_4235),
.Y(n_6432)
);

AOI22xp33_ASAP7_75t_L g6433 ( 
.A1(n_5297),
.A2(n_4907),
.B1(n_4993),
.B2(n_4744),
.Y(n_6433)
);

BUFx12f_ASAP7_75t_L g6434 ( 
.A(n_5643),
.Y(n_6434)
);

NAND2xp5_ASAP7_75t_L g6435 ( 
.A(n_5767),
.B(n_5776),
.Y(n_6435)
);

INVx3_ASAP7_75t_L g6436 ( 
.A(n_5153),
.Y(n_6436)
);

NAND2xp5_ASAP7_75t_L g6437 ( 
.A(n_5776),
.B(n_4681),
.Y(n_6437)
);

AND2x4_ASAP7_75t_L g6438 ( 
.A(n_5320),
.B(n_5328),
.Y(n_6438)
);

INVx2_ASAP7_75t_L g6439 ( 
.A(n_5240),
.Y(n_6439)
);

INVx2_ASAP7_75t_SL g6440 ( 
.A(n_5992),
.Y(n_6440)
);

INVx2_ASAP7_75t_L g6441 ( 
.A(n_5241),
.Y(n_6441)
);

NAND2xp5_ASAP7_75t_L g6442 ( 
.A(n_5800),
.B(n_4681),
.Y(n_6442)
);

INVx3_ASAP7_75t_L g6443 ( 
.A(n_5155),
.Y(n_6443)
);

INVx2_ASAP7_75t_L g6444 ( 
.A(n_5241),
.Y(n_6444)
);

INVx3_ASAP7_75t_L g6445 ( 
.A(n_5155),
.Y(n_6445)
);

OR2x2_ASAP7_75t_L g6446 ( 
.A(n_5802),
.B(n_4545),
.Y(n_6446)
);

INVx1_ASAP7_75t_L g6447 ( 
.A(n_5261),
.Y(n_6447)
);

NAND2xp5_ASAP7_75t_L g6448 ( 
.A(n_5800),
.B(n_4681),
.Y(n_6448)
);

INVx2_ASAP7_75t_L g6449 ( 
.A(n_5241),
.Y(n_6449)
);

NAND2x1p5_ASAP7_75t_L g6450 ( 
.A(n_5892),
.B(n_4229),
.Y(n_6450)
);

NOR2xp67_ASAP7_75t_L g6451 ( 
.A(n_5819),
.B(n_4232),
.Y(n_6451)
);

AOI22xp5_ASAP7_75t_L g6452 ( 
.A1(n_5223),
.A2(n_4611),
.B1(n_4993),
.B2(n_4907),
.Y(n_6452)
);

AOI22xp33_ASAP7_75t_SL g6453 ( 
.A1(n_5221),
.A2(n_4235),
.B1(n_4250),
.B2(n_4241),
.Y(n_6453)
);

OAI22xp33_ASAP7_75t_L g6454 ( 
.A1(n_5780),
.A2(n_4462),
.B1(n_4417),
.B2(n_4642),
.Y(n_6454)
);

NAND2xp5_ASAP7_75t_L g6455 ( 
.A(n_5909),
.B(n_4695),
.Y(n_6455)
);

INVx1_ASAP7_75t_L g6456 ( 
.A(n_5261),
.Y(n_6456)
);

INVx3_ASAP7_75t_L g6457 ( 
.A(n_5155),
.Y(n_6457)
);

AOI21xp5_ASAP7_75t_L g6458 ( 
.A1(n_5789),
.A2(n_4241),
.B(n_4235),
.Y(n_6458)
);

INVx2_ASAP7_75t_SL g6459 ( 
.A(n_5992),
.Y(n_6459)
);

INVx1_ASAP7_75t_L g6460 ( 
.A(n_5263),
.Y(n_6460)
);

INVxp67_ASAP7_75t_SL g6461 ( 
.A(n_5432),
.Y(n_6461)
);

BUFx4f_ASAP7_75t_L g6462 ( 
.A(n_5388),
.Y(n_6462)
);

OA21x2_ASAP7_75t_L g6463 ( 
.A1(n_5938),
.A2(n_4247),
.B(n_4232),
.Y(n_6463)
);

NAND2xp5_ASAP7_75t_L g6464 ( 
.A(n_5909),
.B(n_4695),
.Y(n_6464)
);

NOR3xp33_ASAP7_75t_L g6465 ( 
.A(n_5660),
.B(n_4493),
.C(n_4438),
.Y(n_6465)
);

AOI22xp33_ASAP7_75t_L g6466 ( 
.A1(n_5348),
.A2(n_4993),
.B1(n_4462),
.B2(n_4250),
.Y(n_6466)
);

INVx1_ASAP7_75t_L g6467 ( 
.A(n_5263),
.Y(n_6467)
);

BUFx2_ASAP7_75t_L g6468 ( 
.A(n_5635),
.Y(n_6468)
);

INVx3_ASAP7_75t_L g6469 ( 
.A(n_5155),
.Y(n_6469)
);

INVx1_ASAP7_75t_SL g6470 ( 
.A(n_5161),
.Y(n_6470)
);

INVx1_ASAP7_75t_L g6471 ( 
.A(n_5268),
.Y(n_6471)
);

INVx1_ASAP7_75t_L g6472 ( 
.A(n_5268),
.Y(n_6472)
);

AOI21xp5_ASAP7_75t_SL g6473 ( 
.A1(n_5644),
.A2(n_4462),
.B(n_4959),
.Y(n_6473)
);

INVx1_ASAP7_75t_L g6474 ( 
.A(n_5289),
.Y(n_6474)
);

NAND2xp5_ASAP7_75t_L g6475 ( 
.A(n_5919),
.B(n_4695),
.Y(n_6475)
);

HB1xp67_ASAP7_75t_L g6476 ( 
.A(n_5329),
.Y(n_6476)
);

INVx1_ASAP7_75t_L g6477 ( 
.A(n_5289),
.Y(n_6477)
);

AND2x2_ASAP7_75t_L g6478 ( 
.A(n_5797),
.B(n_5809),
.Y(n_6478)
);

BUFx3_ASAP7_75t_L g6479 ( 
.A(n_5982),
.Y(n_6479)
);

AND2x2_ASAP7_75t_L g6480 ( 
.A(n_5797),
.B(n_4503),
.Y(n_6480)
);

INVx2_ASAP7_75t_SL g6481 ( 
.A(n_6007),
.Y(n_6481)
);

INVx1_ASAP7_75t_L g6482 ( 
.A(n_5295),
.Y(n_6482)
);

AOI22xp33_ASAP7_75t_SL g6483 ( 
.A1(n_5971),
.A2(n_4250),
.B1(n_4258),
.B2(n_4241),
.Y(n_6483)
);

AOI21x1_ASAP7_75t_L g6484 ( 
.A1(n_5287),
.A2(n_4171),
.B(n_4174),
.Y(n_6484)
);

BUFx4_ASAP7_75t_SL g6485 ( 
.A(n_6100),
.Y(n_6485)
);

NAND2xp5_ASAP7_75t_L g6486 ( 
.A(n_5919),
.B(n_4699),
.Y(n_6486)
);

NAND2xp5_ASAP7_75t_SL g6487 ( 
.A(n_5639),
.B(n_4446),
.Y(n_6487)
);

AOI21xp5_ASAP7_75t_L g6488 ( 
.A1(n_5443),
.A2(n_4250),
.B(n_4241),
.Y(n_6488)
);

INVxp67_ASAP7_75t_L g6489 ( 
.A(n_5714),
.Y(n_6489)
);

AOI22xp33_ASAP7_75t_L g6490 ( 
.A1(n_5124),
.A2(n_5314),
.B1(n_5712),
.B2(n_5675),
.Y(n_6490)
);

INVx3_ASAP7_75t_L g6491 ( 
.A(n_5169),
.Y(n_6491)
);

BUFx2_ASAP7_75t_L g6492 ( 
.A(n_5982),
.Y(n_6492)
);

AOI22xp33_ASAP7_75t_L g6493 ( 
.A1(n_5124),
.A2(n_4993),
.B1(n_4462),
.B2(n_4241),
.Y(n_6493)
);

AOI22xp33_ASAP7_75t_L g6494 ( 
.A1(n_5314),
.A2(n_5712),
.B1(n_5675),
.B2(n_5755),
.Y(n_6494)
);

BUFx3_ASAP7_75t_L g6495 ( 
.A(n_5982),
.Y(n_6495)
);

BUFx2_ASAP7_75t_SL g6496 ( 
.A(n_5438),
.Y(n_6496)
);

OAI22xp5_ASAP7_75t_L g6497 ( 
.A1(n_5736),
.A2(n_4609),
.B1(n_4713),
.B2(n_4598),
.Y(n_6497)
);

INVx1_ASAP7_75t_L g6498 ( 
.A(n_5295),
.Y(n_6498)
);

CKINVDCx5p33_ASAP7_75t_R g6499 ( 
.A(n_5643),
.Y(n_6499)
);

NAND3xp33_ASAP7_75t_L g6500 ( 
.A(n_5660),
.B(n_5704),
.C(n_5689),
.Y(n_6500)
);

BUFx2_ASAP7_75t_L g6501 ( 
.A(n_5982),
.Y(n_6501)
);

INVx3_ASAP7_75t_L g6502 ( 
.A(n_5169),
.Y(n_6502)
);

A2O1A1Ixp33_ASAP7_75t_L g6503 ( 
.A1(n_5796),
.A2(n_4250),
.B(n_4258),
.C(n_4241),
.Y(n_6503)
);

AND2x2_ASAP7_75t_L g6504 ( 
.A(n_5809),
.B(n_4532),
.Y(n_6504)
);

AOI21xp5_ASAP7_75t_L g6505 ( 
.A1(n_6043),
.A2(n_4258),
.B(n_4250),
.Y(n_6505)
);

BUFx2_ASAP7_75t_L g6506 ( 
.A(n_5714),
.Y(n_6506)
);

CKINVDCx20_ASAP7_75t_R g6507 ( 
.A(n_5749),
.Y(n_6507)
);

AOI21xp5_ASAP7_75t_L g6508 ( 
.A1(n_6043),
.A2(n_6054),
.B(n_5302),
.Y(n_6508)
);

NAND2xp5_ASAP7_75t_L g6509 ( 
.A(n_5925),
.B(n_4699),
.Y(n_6509)
);

INVx1_ASAP7_75t_L g6510 ( 
.A(n_5296),
.Y(n_6510)
);

INVx1_ASAP7_75t_L g6511 ( 
.A(n_5296),
.Y(n_6511)
);

INVx1_ASAP7_75t_L g6512 ( 
.A(n_5304),
.Y(n_6512)
);

AOI21xp5_ASAP7_75t_L g6513 ( 
.A1(n_6054),
.A2(n_4258),
.B(n_4250),
.Y(n_6513)
);

O2A1O1Ixp33_ASAP7_75t_L g6514 ( 
.A1(n_5704),
.A2(n_4553),
.B(n_4842),
.C(n_4493),
.Y(n_6514)
);

BUFx2_ASAP7_75t_SL g6515 ( 
.A(n_5542),
.Y(n_6515)
);

INVx8_ASAP7_75t_L g6516 ( 
.A(n_5198),
.Y(n_6516)
);

OAI21x1_ASAP7_75t_L g6517 ( 
.A1(n_5938),
.A2(n_4262),
.B(n_4247),
.Y(n_6517)
);

NOR2xp33_ASAP7_75t_L g6518 ( 
.A(n_5748),
.B(n_5059),
.Y(n_6518)
);

INVx2_ASAP7_75t_SL g6519 ( 
.A(n_6007),
.Y(n_6519)
);

INVx2_ASAP7_75t_SL g6520 ( 
.A(n_6007),
.Y(n_6520)
);

INVx1_ASAP7_75t_L g6521 ( 
.A(n_5304),
.Y(n_6521)
);

AND2x4_ASAP7_75t_L g6522 ( 
.A(n_5320),
.B(n_5328),
.Y(n_6522)
);

NAND2xp5_ASAP7_75t_L g6523 ( 
.A(n_5925),
.B(n_4699),
.Y(n_6523)
);

INVx1_ASAP7_75t_L g6524 ( 
.A(n_5309),
.Y(n_6524)
);

INVx2_ASAP7_75t_SL g6525 ( 
.A(n_6007),
.Y(n_6525)
);

CKINVDCx20_ASAP7_75t_R g6526 ( 
.A(n_5450),
.Y(n_6526)
);

OAI21xp33_ASAP7_75t_L g6527 ( 
.A1(n_5623),
.A2(n_4710),
.B(n_4709),
.Y(n_6527)
);

NAND2xp5_ASAP7_75t_SL g6528 ( 
.A(n_5639),
.B(n_4598),
.Y(n_6528)
);

INVx1_ASAP7_75t_L g6529 ( 
.A(n_5309),
.Y(n_6529)
);

INVx1_ASAP7_75t_SL g6530 ( 
.A(n_5161),
.Y(n_6530)
);

OAI21x1_ASAP7_75t_L g6531 ( 
.A1(n_5287),
.A2(n_4262),
.B(n_4256),
.Y(n_6531)
);

INVx3_ASAP7_75t_L g6532 ( 
.A(n_5169),
.Y(n_6532)
);

O2A1O1Ixp33_ASAP7_75t_L g6533 ( 
.A1(n_5122),
.A2(n_4553),
.B(n_4882),
.C(n_4842),
.Y(n_6533)
);

HB1xp67_ASAP7_75t_L g6534 ( 
.A(n_5329),
.Y(n_6534)
);

AOI21xp5_ASAP7_75t_L g6535 ( 
.A1(n_5302),
.A2(n_4258),
.B(n_4250),
.Y(n_6535)
);

INVx3_ASAP7_75t_L g6536 ( 
.A(n_5173),
.Y(n_6536)
);

OR2x2_ASAP7_75t_L g6537 ( 
.A(n_5707),
.B(n_4545),
.Y(n_6537)
);

AOI221xp5_ASAP7_75t_L g6538 ( 
.A1(n_5122),
.A2(n_4710),
.B1(n_4721),
.B2(n_4718),
.C(n_4709),
.Y(n_6538)
);

AOI22xp5_ASAP7_75t_L g6539 ( 
.A1(n_5223),
.A2(n_4899),
.B1(n_4443),
.B2(n_4505),
.Y(n_6539)
);

AND2x2_ASAP7_75t_L g6540 ( 
.A(n_5809),
.B(n_4532),
.Y(n_6540)
);

OAI21xp5_ASAP7_75t_L g6541 ( 
.A1(n_5623),
.A2(n_5086),
.B(n_4995),
.Y(n_6541)
);

CKINVDCx5p33_ASAP7_75t_R g6542 ( 
.A(n_5643),
.Y(n_6542)
);

NOR2x1_ASAP7_75t_L g6543 ( 
.A(n_5484),
.B(n_4945),
.Y(n_6543)
);

INVx3_ASAP7_75t_L g6544 ( 
.A(n_5173),
.Y(n_6544)
);

AOI21xp5_ASAP7_75t_L g6545 ( 
.A1(n_5638),
.A2(n_4258),
.B(n_4250),
.Y(n_6545)
);

AND2x2_ASAP7_75t_L g6546 ( 
.A(n_5864),
.B(n_4532),
.Y(n_6546)
);

INVx3_ASAP7_75t_SL g6547 ( 
.A(n_5682),
.Y(n_6547)
);

INVx1_ASAP7_75t_L g6548 ( 
.A(n_5317),
.Y(n_6548)
);

BUFx2_ASAP7_75t_L g6549 ( 
.A(n_5117),
.Y(n_6549)
);

NAND2xp5_ASAP7_75t_L g6550 ( 
.A(n_5929),
.B(n_4709),
.Y(n_6550)
);

INVx1_ASAP7_75t_L g6551 ( 
.A(n_5317),
.Y(n_6551)
);

AOI21xp5_ASAP7_75t_L g6552 ( 
.A1(n_5638),
.A2(n_5657),
.B(n_5647),
.Y(n_6552)
);

INVx1_ASAP7_75t_L g6553 ( 
.A(n_5322),
.Y(n_6553)
);

AND3x1_ASAP7_75t_SL g6554 ( 
.A(n_5630),
.B(n_4649),
.C(n_4632),
.Y(n_6554)
);

AOI21xp5_ASAP7_75t_L g6555 ( 
.A1(n_5647),
.A2(n_4321),
.B(n_4258),
.Y(n_6555)
);

INVx2_ASAP7_75t_SL g6556 ( 
.A(n_6007),
.Y(n_6556)
);

BUFx2_ASAP7_75t_L g6557 ( 
.A(n_5117),
.Y(n_6557)
);

AOI22xp5_ASAP7_75t_L g6558 ( 
.A1(n_5145),
.A2(n_4899),
.B1(n_4430),
.B2(n_4505),
.Y(n_6558)
);

AOI21xp5_ASAP7_75t_L g6559 ( 
.A1(n_5657),
.A2(n_4321),
.B(n_4258),
.Y(n_6559)
);

NOR2xp33_ASAP7_75t_L g6560 ( 
.A(n_5451),
.B(n_5059),
.Y(n_6560)
);

CKINVDCx5p33_ASAP7_75t_R g6561 ( 
.A(n_5865),
.Y(n_6561)
);

INVx3_ASAP7_75t_L g6562 ( 
.A(n_5206),
.Y(n_6562)
);

CKINVDCx20_ASAP7_75t_R g6563 ( 
.A(n_5472),
.Y(n_6563)
);

AND2x2_ASAP7_75t_L g6564 ( 
.A(n_5864),
.B(n_4561),
.Y(n_6564)
);

OAI22xp5_ASAP7_75t_L g6565 ( 
.A1(n_5780),
.A2(n_4598),
.B1(n_4713),
.B2(n_4609),
.Y(n_6565)
);

INVx3_ASAP7_75t_L g6566 ( 
.A(n_5206),
.Y(n_6566)
);

BUFx12f_ASAP7_75t_L g6567 ( 
.A(n_5865),
.Y(n_6567)
);

OR2x2_ASAP7_75t_L g6568 ( 
.A(n_5707),
.B(n_4552),
.Y(n_6568)
);

BUFx3_ASAP7_75t_L g6569 ( 
.A(n_5298),
.Y(n_6569)
);

BUFx10_ASAP7_75t_L g6570 ( 
.A(n_5187),
.Y(n_6570)
);

INVx1_ASAP7_75t_L g6571 ( 
.A(n_5322),
.Y(n_6571)
);

OR2x2_ASAP7_75t_SL g6572 ( 
.A(n_5500),
.B(n_5398),
.Y(n_6572)
);

INVx1_ASAP7_75t_L g6573 ( 
.A(n_5327),
.Y(n_6573)
);

INVxp67_ASAP7_75t_SL g6574 ( 
.A(n_5484),
.Y(n_6574)
);

OR2x2_ASAP7_75t_L g6575 ( 
.A(n_5786),
.B(n_4552),
.Y(n_6575)
);

AOI21xp5_ASAP7_75t_L g6576 ( 
.A1(n_5674),
.A2(n_4321),
.B(n_4258),
.Y(n_6576)
);

AOI21xp5_ASAP7_75t_L g6577 ( 
.A1(n_5674),
.A2(n_4349),
.B(n_4321),
.Y(n_6577)
);

BUFx3_ASAP7_75t_L g6578 ( 
.A(n_5298),
.Y(n_6578)
);

BUFx12f_ASAP7_75t_L g6579 ( 
.A(n_5865),
.Y(n_6579)
);

AOI22xp5_ASAP7_75t_L g6580 ( 
.A1(n_5145),
.A2(n_4899),
.B1(n_4443),
.B2(n_4430),
.Y(n_6580)
);

AOI21xp5_ASAP7_75t_L g6581 ( 
.A1(n_5697),
.A2(n_4349),
.B(n_4321),
.Y(n_6581)
);

AOI22xp5_ASAP7_75t_L g6582 ( 
.A1(n_5719),
.A2(n_5084),
.B1(n_5023),
.B2(n_4642),
.Y(n_6582)
);

BUFx2_ASAP7_75t_R g6583 ( 
.A(n_5157),
.Y(n_6583)
);

OAI22xp5_ASAP7_75t_L g6584 ( 
.A1(n_5719),
.A2(n_4609),
.B1(n_4713),
.B2(n_4710),
.Y(n_6584)
);

BUFx3_ASAP7_75t_L g6585 ( 
.A(n_5298),
.Y(n_6585)
);

NOR2xp33_ASAP7_75t_L g6586 ( 
.A(n_5739),
.B(n_5060),
.Y(n_6586)
);

INVx1_ASAP7_75t_L g6587 ( 
.A(n_5327),
.Y(n_6587)
);

INVx1_ASAP7_75t_L g6588 ( 
.A(n_5330),
.Y(n_6588)
);

NAND2x1p5_ASAP7_75t_L g6589 ( 
.A(n_5138),
.B(n_4276),
.Y(n_6589)
);

AND2x2_ASAP7_75t_L g6590 ( 
.A(n_5864),
.B(n_5868),
.Y(n_6590)
);

OAI21x1_ASAP7_75t_L g6591 ( 
.A1(n_5291),
.A2(n_4262),
.B(n_4256),
.Y(n_6591)
);

NOR2xp33_ASAP7_75t_L g6592 ( 
.A(n_5745),
.B(n_5060),
.Y(n_6592)
);

INVx1_ASAP7_75t_L g6593 ( 
.A(n_5330),
.Y(n_6593)
);

HB1xp67_ASAP7_75t_L g6594 ( 
.A(n_5368),
.Y(n_6594)
);

INVx5_ASAP7_75t_L g6595 ( 
.A(n_5264),
.Y(n_6595)
);

INVx3_ASAP7_75t_L g6596 ( 
.A(n_5206),
.Y(n_6596)
);

AOI22xp33_ASAP7_75t_L g6597 ( 
.A1(n_5817),
.A2(n_4321),
.B1(n_4352),
.B2(n_4349),
.Y(n_6597)
);

BUFx3_ASAP7_75t_L g6598 ( 
.A(n_5298),
.Y(n_6598)
);

BUFx3_ASAP7_75t_L g6599 ( 
.A(n_5298),
.Y(n_6599)
);

INVx6_ASAP7_75t_L g6600 ( 
.A(n_5830),
.Y(n_6600)
);

CKINVDCx11_ASAP7_75t_R g6601 ( 
.A(n_6103),
.Y(n_6601)
);

NAND2xp5_ASAP7_75t_L g6602 ( 
.A(n_5929),
.B(n_4718),
.Y(n_6602)
);

INVx1_ASAP7_75t_L g6603 ( 
.A(n_5340),
.Y(n_6603)
);

INVx1_ASAP7_75t_L g6604 ( 
.A(n_5340),
.Y(n_6604)
);

AOI22xp33_ASAP7_75t_L g6605 ( 
.A1(n_5132),
.A2(n_4321),
.B1(n_4352),
.B2(n_4349),
.Y(n_6605)
);

BUFx2_ASAP7_75t_L g6606 ( 
.A(n_5117),
.Y(n_6606)
);

BUFx2_ASAP7_75t_L g6607 ( 
.A(n_5117),
.Y(n_6607)
);

CKINVDCx20_ASAP7_75t_R g6608 ( 
.A(n_5628),
.Y(n_6608)
);

INVx1_ASAP7_75t_L g6609 ( 
.A(n_5351),
.Y(n_6609)
);

AND2x2_ASAP7_75t_L g6610 ( 
.A(n_5868),
.B(n_4561),
.Y(n_6610)
);

INVx2_ASAP7_75t_SL g6611 ( 
.A(n_6018),
.Y(n_6611)
);

INVx1_ASAP7_75t_L g6612 ( 
.A(n_5351),
.Y(n_6612)
);

NAND2xp5_ASAP7_75t_L g6613 ( 
.A(n_5942),
.B(n_4718),
.Y(n_6613)
);

BUFx12f_ASAP7_75t_L g6614 ( 
.A(n_5970),
.Y(n_6614)
);

NAND2xp33_ASAP7_75t_SL g6615 ( 
.A(n_6072),
.B(n_4649),
.Y(n_6615)
);

NAND2xp5_ASAP7_75t_L g6616 ( 
.A(n_5942),
.B(n_4721),
.Y(n_6616)
);

BUFx2_ASAP7_75t_L g6617 ( 
.A(n_5117),
.Y(n_6617)
);

INVx1_ASAP7_75t_L g6618 ( 
.A(n_5354),
.Y(n_6618)
);

OAI22xp33_ASAP7_75t_L g6619 ( 
.A1(n_5141),
.A2(n_4642),
.B1(n_4981),
.B2(n_4713),
.Y(n_6619)
);

OAI22xp5_ASAP7_75t_L g6620 ( 
.A1(n_5810),
.A2(n_4609),
.B1(n_4723),
.B2(n_4721),
.Y(n_6620)
);

INVx1_ASAP7_75t_L g6621 ( 
.A(n_5354),
.Y(n_6621)
);

INVx1_ASAP7_75t_L g6622 ( 
.A(n_5355),
.Y(n_6622)
);

INVxp67_ASAP7_75t_SL g6623 ( 
.A(n_5662),
.Y(n_6623)
);

AND2x2_ASAP7_75t_L g6624 ( 
.A(n_5868),
.B(n_4561),
.Y(n_6624)
);

INVxp67_ASAP7_75t_SL g6625 ( 
.A(n_5662),
.Y(n_6625)
);

INVx1_ASAP7_75t_L g6626 ( 
.A(n_5355),
.Y(n_6626)
);

NAND2xp5_ASAP7_75t_L g6627 ( 
.A(n_5943),
.B(n_4723),
.Y(n_6627)
);

INVx1_ASAP7_75t_L g6628 ( 
.A(n_5372),
.Y(n_6628)
);

BUFx12f_ASAP7_75t_L g6629 ( 
.A(n_5970),
.Y(n_6629)
);

OA21x2_ASAP7_75t_L g6630 ( 
.A1(n_6030),
.A2(n_4171),
.B(n_4935),
.Y(n_6630)
);

NAND2xp33_ASAP7_75t_L g6631 ( 
.A(n_6072),
.B(n_4936),
.Y(n_6631)
);

INVx1_ASAP7_75t_L g6632 ( 
.A(n_5372),
.Y(n_6632)
);

AOI21xp33_ASAP7_75t_L g6633 ( 
.A1(n_5713),
.A2(n_4349),
.B(n_4321),
.Y(n_6633)
);

OAI22xp5_ASAP7_75t_L g6634 ( 
.A1(n_5810),
.A2(n_4736),
.B1(n_4723),
.B2(n_4945),
.Y(n_6634)
);

AND2x4_ASAP7_75t_L g6635 ( 
.A(n_5462),
.B(n_5917),
.Y(n_6635)
);

OR2x2_ASAP7_75t_SL g6636 ( 
.A(n_5500),
.B(n_4321),
.Y(n_6636)
);

BUFx12f_ASAP7_75t_L g6637 ( 
.A(n_5970),
.Y(n_6637)
);

NAND2xp5_ASAP7_75t_L g6638 ( 
.A(n_5943),
.B(n_4736),
.Y(n_6638)
);

HB1xp67_ASAP7_75t_L g6639 ( 
.A(n_5368),
.Y(n_6639)
);

INVx8_ASAP7_75t_L g6640 ( 
.A(n_5661),
.Y(n_6640)
);

AOI222xp33_ASAP7_75t_L g6641 ( 
.A1(n_5108),
.A2(n_4838),
.B1(n_4826),
.B2(n_4845),
.C1(n_4829),
.C2(n_4824),
.Y(n_6641)
);

INVx1_ASAP7_75t_L g6642 ( 
.A(n_5375),
.Y(n_6642)
);

CKINVDCx20_ASAP7_75t_R g6643 ( 
.A(n_5724),
.Y(n_6643)
);

INVx1_ASAP7_75t_L g6644 ( 
.A(n_5375),
.Y(n_6644)
);

NOR2xp33_ASAP7_75t_SL g6645 ( 
.A(n_5530),
.B(n_4981),
.Y(n_6645)
);

BUFx2_ASAP7_75t_L g6646 ( 
.A(n_5137),
.Y(n_6646)
);

BUFx12f_ASAP7_75t_L g6647 ( 
.A(n_5990),
.Y(n_6647)
);

OR2x2_ASAP7_75t_L g6648 ( 
.A(n_5786),
.B(n_4552),
.Y(n_6648)
);

BUFx12f_ASAP7_75t_L g6649 ( 
.A(n_5990),
.Y(n_6649)
);

AOI21x1_ASAP7_75t_L g6650 ( 
.A1(n_5291),
.A2(n_4171),
.B(n_5086),
.Y(n_6650)
);

INVx2_ASAP7_75t_SL g6651 ( 
.A(n_6018),
.Y(n_6651)
);

OAI22xp5_ASAP7_75t_L g6652 ( 
.A1(n_5881),
.A2(n_4736),
.B1(n_5009),
.B2(n_4945),
.Y(n_6652)
);

INVx1_ASAP7_75t_L g6653 ( 
.A(n_5378),
.Y(n_6653)
);

AO22x1_ASAP7_75t_L g6654 ( 
.A1(n_6006),
.A2(n_4666),
.B1(n_4380),
.B2(n_4642),
.Y(n_6654)
);

AND2x2_ASAP7_75t_L g6655 ( 
.A(n_5888),
.B(n_5703),
.Y(n_6655)
);

BUFx3_ASAP7_75t_L g6656 ( 
.A(n_5298),
.Y(n_6656)
);

AOI21x1_ASAP7_75t_L g6657 ( 
.A1(n_6123),
.A2(n_4171),
.B(n_4935),
.Y(n_6657)
);

HB1xp67_ASAP7_75t_L g6658 ( 
.A(n_5383),
.Y(n_6658)
);

INVx1_ASAP7_75t_L g6659 ( 
.A(n_5378),
.Y(n_6659)
);

NAND2xp5_ASAP7_75t_L g6660 ( 
.A(n_5946),
.B(n_5947),
.Y(n_6660)
);

INVx1_ASAP7_75t_L g6661 ( 
.A(n_5379),
.Y(n_6661)
);

AOI21xp5_ASAP7_75t_L g6662 ( 
.A1(n_5697),
.A2(n_4352),
.B(n_4349),
.Y(n_6662)
);

NAND2xp5_ASAP7_75t_L g6663 ( 
.A(n_5946),
.B(n_4573),
.Y(n_6663)
);

AOI21xp5_ASAP7_75t_L g6664 ( 
.A1(n_5698),
.A2(n_5710),
.B(n_5709),
.Y(n_6664)
);

OAI22xp5_ASAP7_75t_L g6665 ( 
.A1(n_5881),
.A2(n_5009),
.B1(n_4945),
.B2(n_4628),
.Y(n_6665)
);

CKINVDCx6p67_ASAP7_75t_R g6666 ( 
.A(n_5738),
.Y(n_6666)
);

BUFx2_ASAP7_75t_L g6667 ( 
.A(n_5137),
.Y(n_6667)
);

OR2x2_ASAP7_75t_L g6668 ( 
.A(n_5786),
.B(n_4628),
.Y(n_6668)
);

NAND2xp5_ASAP7_75t_L g6669 ( 
.A(n_5947),
.B(n_4573),
.Y(n_6669)
);

AOI22xp33_ASAP7_75t_L g6670 ( 
.A1(n_5323),
.A2(n_4349),
.B1(n_4360),
.B2(n_4352),
.Y(n_6670)
);

AOI21xp5_ASAP7_75t_L g6671 ( 
.A1(n_5698),
.A2(n_4352),
.B(n_4349),
.Y(n_6671)
);

INVx1_ASAP7_75t_L g6672 ( 
.A(n_5379),
.Y(n_6672)
);

AND2x2_ASAP7_75t_L g6673 ( 
.A(n_5888),
.B(n_4573),
.Y(n_6673)
);

BUFx3_ASAP7_75t_L g6674 ( 
.A(n_5298),
.Y(n_6674)
);

AND2x2_ASAP7_75t_L g6675 ( 
.A(n_5888),
.B(n_4582),
.Y(n_6675)
);

HB1xp67_ASAP7_75t_L g6676 ( 
.A(n_5383),
.Y(n_6676)
);

INVxp67_ASAP7_75t_L g6677 ( 
.A(n_5409),
.Y(n_6677)
);

AO22x1_ASAP7_75t_L g6678 ( 
.A1(n_6006),
.A2(n_4666),
.B1(n_4380),
.B2(n_4981),
.Y(n_6678)
);

AND2x2_ASAP7_75t_SL g6679 ( 
.A(n_5388),
.B(n_4432),
.Y(n_6679)
);

INVx1_ASAP7_75t_L g6680 ( 
.A(n_5387),
.Y(n_6680)
);

OAI21x1_ASAP7_75t_SL g6681 ( 
.A1(n_5713),
.A2(n_4559),
.B(n_5009),
.Y(n_6681)
);

AOI22xp5_ASAP7_75t_L g6682 ( 
.A1(n_5141),
.A2(n_5084),
.B1(n_5023),
.B2(n_4839),
.Y(n_6682)
);

BUFx2_ASAP7_75t_L g6683 ( 
.A(n_5137),
.Y(n_6683)
);

INVx1_ASAP7_75t_L g6684 ( 
.A(n_5387),
.Y(n_6684)
);

AOI21xp5_ASAP7_75t_L g6685 ( 
.A1(n_5709),
.A2(n_4352),
.B(n_4349),
.Y(n_6685)
);

OR2x6_ASAP7_75t_L g6686 ( 
.A(n_5661),
.B(n_5807),
.Y(n_6686)
);

INVx3_ASAP7_75t_SL g6687 ( 
.A(n_5682),
.Y(n_6687)
);

INVx1_ASAP7_75t_L g6688 ( 
.A(n_5396),
.Y(n_6688)
);

AOI21xp5_ASAP7_75t_L g6689 ( 
.A1(n_5710),
.A2(n_4360),
.B(n_4352),
.Y(n_6689)
);

INVx1_ASAP7_75t_L g6690 ( 
.A(n_5396),
.Y(n_6690)
);

BUFx4f_ASAP7_75t_L g6691 ( 
.A(n_5388),
.Y(n_6691)
);

INVx1_ASAP7_75t_L g6692 ( 
.A(n_5402),
.Y(n_6692)
);

OAI22xp33_ASAP7_75t_L g6693 ( 
.A1(n_5887),
.A2(n_5879),
.B1(n_5899),
.B2(n_5398),
.Y(n_6693)
);

INVx1_ASAP7_75t_SL g6694 ( 
.A(n_5217),
.Y(n_6694)
);

AND2x4_ASAP7_75t_L g6695 ( 
.A(n_5917),
.B(n_4472),
.Y(n_6695)
);

AND2x4_ASAP7_75t_L g6696 ( 
.A(n_5917),
.B(n_5927),
.Y(n_6696)
);

BUFx2_ASAP7_75t_L g6697 ( 
.A(n_5137),
.Y(n_6697)
);

NAND2xp5_ASAP7_75t_SL g6698 ( 
.A(n_5886),
.B(n_4472),
.Y(n_6698)
);

AOI21x1_ASAP7_75t_L g6699 ( 
.A1(n_6123),
.A2(n_5610),
.B(n_5599),
.Y(n_6699)
);

BUFx3_ASAP7_75t_L g6700 ( 
.A(n_5298),
.Y(n_6700)
);

OR2x2_ASAP7_75t_L g6701 ( 
.A(n_5612),
.B(n_5650),
.Y(n_6701)
);

BUFx3_ASAP7_75t_L g6702 ( 
.A(n_5298),
.Y(n_6702)
);

INVx3_ASAP7_75t_SL g6703 ( 
.A(n_5682),
.Y(n_6703)
);

HB1xp67_ASAP7_75t_L g6704 ( 
.A(n_5409),
.Y(n_6704)
);

OR2x2_ASAP7_75t_SL g6705 ( 
.A(n_5500),
.B(n_4352),
.Y(n_6705)
);

BUFx3_ASAP7_75t_L g6706 ( 
.A(n_5830),
.Y(n_6706)
);

AND2x2_ASAP7_75t_L g6707 ( 
.A(n_5703),
.B(n_4582),
.Y(n_6707)
);

INVxp67_ASAP7_75t_SL g6708 ( 
.A(n_5681),
.Y(n_6708)
);

BUFx3_ASAP7_75t_L g6709 ( 
.A(n_5830),
.Y(n_6709)
);

INVx1_ASAP7_75t_L g6710 ( 
.A(n_5402),
.Y(n_6710)
);

AOI21xp33_ASAP7_75t_L g6711 ( 
.A1(n_5717),
.A2(n_4360),
.B(n_4352),
.Y(n_6711)
);

INVx1_ASAP7_75t_L g6712 ( 
.A(n_5404),
.Y(n_6712)
);

INVx3_ASAP7_75t_L g6713 ( 
.A(n_5215),
.Y(n_6713)
);

INVx4_ASAP7_75t_L g6714 ( 
.A(n_5661),
.Y(n_6714)
);

AOI22xp5_ASAP7_75t_L g6715 ( 
.A1(n_5630),
.A2(n_5084),
.B1(n_5023),
.B2(n_4839),
.Y(n_6715)
);

INVx1_ASAP7_75t_L g6716 ( 
.A(n_5404),
.Y(n_6716)
);

INVx1_ASAP7_75t_L g6717 ( 
.A(n_5421),
.Y(n_6717)
);

OR2x2_ASAP7_75t_L g6718 ( 
.A(n_5612),
.B(n_4628),
.Y(n_6718)
);

OAI22xp5_ASAP7_75t_L g6719 ( 
.A1(n_5887),
.A2(n_5009),
.B1(n_5096),
.B2(n_4882),
.Y(n_6719)
);

AOI22xp33_ASAP7_75t_L g6720 ( 
.A1(n_5323),
.A2(n_4363),
.B1(n_4392),
.B2(n_4360),
.Y(n_6720)
);

OR2x2_ASAP7_75t_L g6721 ( 
.A(n_5650),
.B(n_5680),
.Y(n_6721)
);

OAI22xp5_ASAP7_75t_L g6722 ( 
.A1(n_5876),
.A2(n_5009),
.B1(n_5096),
.B2(n_4995),
.Y(n_6722)
);

BUFx2_ASAP7_75t_L g6723 ( 
.A(n_5137),
.Y(n_6723)
);

NOR2xp33_ASAP7_75t_SL g6724 ( 
.A(n_5530),
.B(n_5444),
.Y(n_6724)
);

NAND2x1p5_ASAP7_75t_L g6725 ( 
.A(n_5138),
.B(n_5150),
.Y(n_6725)
);

HB1xp67_ASAP7_75t_L g6726 ( 
.A(n_5446),
.Y(n_6726)
);

INVx1_ASAP7_75t_SL g6727 ( 
.A(n_5217),
.Y(n_6727)
);

INVx1_ASAP7_75t_L g6728 ( 
.A(n_5421),
.Y(n_6728)
);

AND2x2_ASAP7_75t_L g6729 ( 
.A(n_5703),
.B(n_4582),
.Y(n_6729)
);

AND2x2_ASAP7_75t_L g6730 ( 
.A(n_5715),
.B(n_4612),
.Y(n_6730)
);

HB1xp67_ASAP7_75t_L g6731 ( 
.A(n_5446),
.Y(n_6731)
);

INVx1_ASAP7_75t_L g6732 ( 
.A(n_5430),
.Y(n_6732)
);

AOI222xp33_ASAP7_75t_L g6733 ( 
.A1(n_5108),
.A2(n_4838),
.B1(n_4826),
.B2(n_4845),
.C1(n_4829),
.C2(n_4824),
.Y(n_6733)
);

INVx1_ASAP7_75t_L g6734 ( 
.A(n_5430),
.Y(n_6734)
);

BUFx3_ASAP7_75t_L g6735 ( 
.A(n_5830),
.Y(n_6735)
);

INVx3_ASAP7_75t_L g6736 ( 
.A(n_5215),
.Y(n_6736)
);

INVx2_ASAP7_75t_SL g6737 ( 
.A(n_6018),
.Y(n_6737)
);

OAI22xp5_ASAP7_75t_L g6738 ( 
.A1(n_5876),
.A2(n_5096),
.B1(n_5002),
.B2(n_5006),
.Y(n_6738)
);

NAND2xp5_ASAP7_75t_SL g6739 ( 
.A(n_5886),
.B(n_4485),
.Y(n_6739)
);

OAI22xp5_ASAP7_75t_L g6740 ( 
.A1(n_5168),
.A2(n_5096),
.B1(n_5002),
.B2(n_5006),
.Y(n_6740)
);

HB1xp67_ASAP7_75t_L g6741 ( 
.A(n_5455),
.Y(n_6741)
);

INVx1_ASAP7_75t_L g6742 ( 
.A(n_5435),
.Y(n_6742)
);

AND2x2_ASAP7_75t_SL g6743 ( 
.A(n_5444),
.B(n_6018),
.Y(n_6743)
);

OR2x2_ASAP7_75t_L g6744 ( 
.A(n_5680),
.B(n_4521),
.Y(n_6744)
);

AOI21xp5_ASAP7_75t_L g6745 ( 
.A1(n_5720),
.A2(n_4363),
.B(n_4360),
.Y(n_6745)
);

INVx2_ASAP7_75t_SL g6746 ( 
.A(n_6018),
.Y(n_6746)
);

INVx1_ASAP7_75t_L g6747 ( 
.A(n_5435),
.Y(n_6747)
);

NAND2xp5_ASAP7_75t_SL g6748 ( 
.A(n_5769),
.B(n_4485),
.Y(n_6748)
);

NOR2xp33_ASAP7_75t_L g6749 ( 
.A(n_5878),
.B(n_5067),
.Y(n_6749)
);

INVx1_ASAP7_75t_L g6750 ( 
.A(n_5441),
.Y(n_6750)
);

O2A1O1Ixp33_ASAP7_75t_L g6751 ( 
.A1(n_5164),
.A2(n_5003),
.B(n_5020),
.C(n_4947),
.Y(n_6751)
);

AOI22xp33_ASAP7_75t_L g6752 ( 
.A1(n_5151),
.A2(n_4363),
.B1(n_4392),
.B2(n_4360),
.Y(n_6752)
);

BUFx6f_ASAP7_75t_SL g6753 ( 
.A(n_5444),
.Y(n_6753)
);

OAI22xp5_ASAP7_75t_L g6754 ( 
.A1(n_5208),
.A2(n_5003),
.B1(n_5067),
.B2(n_4559),
.Y(n_6754)
);

OAI22xp5_ASAP7_75t_L g6755 ( 
.A1(n_5208),
.A2(n_4559),
.B1(n_4485),
.B2(n_4487),
.Y(n_6755)
);

NAND2xp5_ASAP7_75t_L g6756 ( 
.A(n_5720),
.B(n_4616),
.Y(n_6756)
);

BUFx3_ASAP7_75t_L g6757 ( 
.A(n_5857),
.Y(n_6757)
);

AOI22xp5_ASAP7_75t_L g6758 ( 
.A1(n_5294),
.A2(n_5084),
.B1(n_5023),
.B2(n_4839),
.Y(n_6758)
);

BUFx2_ASAP7_75t_L g6759 ( 
.A(n_5211),
.Y(n_6759)
);

AOI22xp5_ASAP7_75t_L g6760 ( 
.A1(n_5294),
.A2(n_5084),
.B1(n_5023),
.B2(n_4839),
.Y(n_6760)
);

AOI22xp33_ASAP7_75t_L g6761 ( 
.A1(n_5151),
.A2(n_4363),
.B1(n_4392),
.B2(n_4360),
.Y(n_6761)
);

INVx6_ASAP7_75t_L g6762 ( 
.A(n_5857),
.Y(n_6762)
);

BUFx2_ASAP7_75t_L g6763 ( 
.A(n_5211),
.Y(n_6763)
);

OR2x2_ASAP7_75t_L g6764 ( 
.A(n_5688),
.B(n_4521),
.Y(n_6764)
);

INVx3_ASAP7_75t_L g6765 ( 
.A(n_5259),
.Y(n_6765)
);

AND2x4_ASAP7_75t_SL g6766 ( 
.A(n_5927),
.B(n_4485),
.Y(n_6766)
);

BUFx2_ASAP7_75t_L g6767 ( 
.A(n_5211),
.Y(n_6767)
);

NAND2xp5_ASAP7_75t_L g6768 ( 
.A(n_5741),
.B(n_4616),
.Y(n_6768)
);

O2A1O1Ixp5_ASAP7_75t_SL g6769 ( 
.A1(n_5777),
.A2(n_4806),
.B(n_4813),
.C(n_4800),
.Y(n_6769)
);

INVx3_ASAP7_75t_L g6770 ( 
.A(n_5259),
.Y(n_6770)
);

CKINVDCx5p33_ASAP7_75t_R g6771 ( 
.A(n_5990),
.Y(n_6771)
);

OAI22xp5_ASAP7_75t_L g6772 ( 
.A1(n_5248),
.A2(n_4559),
.B1(n_4486),
.B2(n_4507),
.Y(n_6772)
);

INVx2_ASAP7_75t_SL g6773 ( 
.A(n_6023),
.Y(n_6773)
);

CKINVDCx20_ASAP7_75t_R g6774 ( 
.A(n_5941),
.Y(n_6774)
);

NOR2xp33_ASAP7_75t_SL g6775 ( 
.A(n_5833),
.B(n_4981),
.Y(n_6775)
);

INVx1_ASAP7_75t_SL g6776 ( 
.A(n_5243),
.Y(n_6776)
);

INVx1_ASAP7_75t_L g6777 ( 
.A(n_5441),
.Y(n_6777)
);

AND2x2_ASAP7_75t_L g6778 ( 
.A(n_5900),
.B(n_5901),
.Y(n_6778)
);

CKINVDCx5p33_ASAP7_75t_R g6779 ( 
.A(n_5262),
.Y(n_6779)
);

AOI22xp33_ASAP7_75t_L g6780 ( 
.A1(n_5316),
.A2(n_4363),
.B1(n_4392),
.B2(n_4360),
.Y(n_6780)
);

INVx1_ASAP7_75t_L g6781 ( 
.A(n_5442),
.Y(n_6781)
);

CKINVDCx9p33_ASAP7_75t_R g6782 ( 
.A(n_5165),
.Y(n_6782)
);

INVx6_ASAP7_75t_L g6783 ( 
.A(n_5857),
.Y(n_6783)
);

INVx1_ASAP7_75t_L g6784 ( 
.A(n_5442),
.Y(n_6784)
);

BUFx12f_ASAP7_75t_L g6785 ( 
.A(n_6098),
.Y(n_6785)
);

INVx5_ASAP7_75t_L g6786 ( 
.A(n_5264),
.Y(n_6786)
);

HB1xp67_ASAP7_75t_L g6787 ( 
.A(n_5455),
.Y(n_6787)
);

HB1xp67_ASAP7_75t_L g6788 ( 
.A(n_5477),
.Y(n_6788)
);

OAI21xp33_ASAP7_75t_L g6789 ( 
.A1(n_5646),
.A2(n_4626),
.B(n_4616),
.Y(n_6789)
);

INVx1_ASAP7_75t_SL g6790 ( 
.A(n_5243),
.Y(n_6790)
);

NAND2xp5_ASAP7_75t_L g6791 ( 
.A(n_5741),
.B(n_4626),
.Y(n_6791)
);

OA22x2_ASAP7_75t_L g6792 ( 
.A1(n_5879),
.A2(n_4486),
.B1(n_4507),
.B2(n_4487),
.Y(n_6792)
);

INVx1_ASAP7_75t_L g6793 ( 
.A(n_5454),
.Y(n_6793)
);

NOR2x1_ASAP7_75t_SL g6794 ( 
.A(n_5998),
.B(n_5264),
.Y(n_6794)
);

AOI22xp33_ASAP7_75t_L g6795 ( 
.A1(n_5316),
.A2(n_4363),
.B1(n_4392),
.B2(n_4360),
.Y(n_6795)
);

A2O1A1Ixp33_ASAP7_75t_L g6796 ( 
.A1(n_5747),
.A2(n_4363),
.B(n_4440),
.C(n_4392),
.Y(n_6796)
);

INVx1_ASAP7_75t_SL g6797 ( 
.A(n_5299),
.Y(n_6797)
);

AOI21xp5_ASAP7_75t_L g6798 ( 
.A1(n_5783),
.A2(n_4392),
.B(n_4363),
.Y(n_6798)
);

INVx2_ASAP7_75t_SL g6799 ( 
.A(n_6023),
.Y(n_6799)
);

AOI22xp5_ASAP7_75t_L g6800 ( 
.A1(n_5729),
.A2(n_5110),
.B1(n_5391),
.B2(n_5257),
.Y(n_6800)
);

AOI21xp33_ASAP7_75t_L g6801 ( 
.A1(n_5717),
.A2(n_4392),
.B(n_4363),
.Y(n_6801)
);

AOI21xp5_ASAP7_75t_L g6802 ( 
.A1(n_5783),
.A2(n_4440),
.B(n_4392),
.Y(n_6802)
);

INVx6_ASAP7_75t_SL g6803 ( 
.A(n_5264),
.Y(n_6803)
);

AOI21xp5_ASAP7_75t_L g6804 ( 
.A1(n_5799),
.A2(n_4479),
.B(n_4440),
.Y(n_6804)
);

BUFx2_ASAP7_75t_L g6805 ( 
.A(n_5211),
.Y(n_6805)
);

AOI22xp33_ASAP7_75t_L g6806 ( 
.A1(n_5540),
.A2(n_4440),
.B1(n_4515),
.B2(n_4479),
.Y(n_6806)
);

NAND2xp5_ASAP7_75t_L g6807 ( 
.A(n_5799),
.B(n_4626),
.Y(n_6807)
);

INVx1_ASAP7_75t_L g6808 ( 
.A(n_5454),
.Y(n_6808)
);

NOR2xp33_ASAP7_75t_SL g6809 ( 
.A(n_5833),
.B(n_4437),
.Y(n_6809)
);

NAND2xp5_ASAP7_75t_L g6810 ( 
.A(n_5812),
.B(n_4633),
.Y(n_6810)
);

INVx1_ASAP7_75t_L g6811 ( 
.A(n_5459),
.Y(n_6811)
);

INVx1_ASAP7_75t_L g6812 ( 
.A(n_5459),
.Y(n_6812)
);

BUFx2_ASAP7_75t_L g6813 ( 
.A(n_5211),
.Y(n_6813)
);

INVx2_ASAP7_75t_SL g6814 ( 
.A(n_6023),
.Y(n_6814)
);

CKINVDCx20_ASAP7_75t_R g6815 ( 
.A(n_5694),
.Y(n_6815)
);

HB1xp67_ASAP7_75t_L g6816 ( 
.A(n_5477),
.Y(n_6816)
);

AOI22xp33_ASAP7_75t_L g6817 ( 
.A1(n_5540),
.A2(n_4440),
.B1(n_4515),
.B2(n_4479),
.Y(n_6817)
);

AOI22xp33_ASAP7_75t_L g6818 ( 
.A1(n_5729),
.A2(n_4440),
.B1(n_4515),
.B2(n_4479),
.Y(n_6818)
);

AND2x2_ASAP7_75t_L g6819 ( 
.A(n_5900),
.B(n_4633),
.Y(n_6819)
);

BUFx2_ASAP7_75t_L g6820 ( 
.A(n_5219),
.Y(n_6820)
);

INVx1_ASAP7_75t_SL g6821 ( 
.A(n_5299),
.Y(n_6821)
);

BUFx3_ASAP7_75t_L g6822 ( 
.A(n_5857),
.Y(n_6822)
);

INVx5_ASAP7_75t_L g6823 ( 
.A(n_5301),
.Y(n_6823)
);

BUFx2_ASAP7_75t_L g6824 ( 
.A(n_5219),
.Y(n_6824)
);

INVxp67_ASAP7_75t_L g6825 ( 
.A(n_5479),
.Y(n_6825)
);

OR2x2_ASAP7_75t_L g6826 ( 
.A(n_5688),
.B(n_4522),
.Y(n_6826)
);

AOI21xp5_ASAP7_75t_L g6827 ( 
.A1(n_5812),
.A2(n_4479),
.B(n_4440),
.Y(n_6827)
);

INVx1_ASAP7_75t_SL g6828 ( 
.A(n_5326),
.Y(n_6828)
);

AND3x1_ASAP7_75t_SL g6829 ( 
.A(n_5896),
.B(n_6008),
.C(n_5872),
.Y(n_6829)
);

INVx1_ASAP7_75t_L g6830 ( 
.A(n_5460),
.Y(n_6830)
);

AOI22xp33_ASAP7_75t_L g6831 ( 
.A1(n_5220),
.A2(n_4440),
.B1(n_4515),
.B2(n_4479),
.Y(n_6831)
);

INVx1_ASAP7_75t_L g6832 ( 
.A(n_5460),
.Y(n_6832)
);

INVx1_ASAP7_75t_L g6833 ( 
.A(n_5469),
.Y(n_6833)
);

NAND2xp5_ASAP7_75t_SL g6834 ( 
.A(n_6006),
.B(n_6067),
.Y(n_6834)
);

AOI22xp33_ASAP7_75t_SL g6835 ( 
.A1(n_5568),
.A2(n_4479),
.B1(n_4515),
.B2(n_4440),
.Y(n_6835)
);

INVx1_ASAP7_75t_L g6836 ( 
.A(n_5469),
.Y(n_6836)
);

OAI22xp5_ASAP7_75t_L g6837 ( 
.A1(n_5248),
.A2(n_4507),
.B1(n_4659),
.B2(n_4487),
.Y(n_6837)
);

INVx4_ASAP7_75t_L g6838 ( 
.A(n_5807),
.Y(n_6838)
);

BUFx2_ASAP7_75t_L g6839 ( 
.A(n_5219),
.Y(n_6839)
);

CKINVDCx20_ASAP7_75t_R g6840 ( 
.A(n_5851),
.Y(n_6840)
);

AOI22xp33_ASAP7_75t_L g6841 ( 
.A1(n_5257),
.A2(n_4479),
.B1(n_4530),
.B2(n_4515),
.Y(n_6841)
);

AOI21xp5_ASAP7_75t_L g6842 ( 
.A1(n_5825),
.A2(n_4515),
.B(n_4479),
.Y(n_6842)
);

INVx1_ASAP7_75t_L g6843 ( 
.A(n_5473),
.Y(n_6843)
);

NAND2xp5_ASAP7_75t_L g6844 ( 
.A(n_5825),
.B(n_5895),
.Y(n_6844)
);

AOI22xp5_ASAP7_75t_L g6845 ( 
.A1(n_5110),
.A2(n_5084),
.B1(n_5023),
.B2(n_4881),
.Y(n_6845)
);

HB1xp67_ASAP7_75t_L g6846 ( 
.A(n_5479),
.Y(n_6846)
);

HB1xp67_ASAP7_75t_L g6847 ( 
.A(n_5490),
.Y(n_6847)
);

OR2x2_ASAP7_75t_L g6848 ( 
.A(n_5726),
.B(n_4522),
.Y(n_6848)
);

OAI21xp5_ASAP7_75t_L g6849 ( 
.A1(n_5753),
.A2(n_4449),
.B(n_4427),
.Y(n_6849)
);

INVxp67_ASAP7_75t_L g6850 ( 
.A(n_5490),
.Y(n_6850)
);

INVx1_ASAP7_75t_L g6851 ( 
.A(n_5473),
.Y(n_6851)
);

BUFx2_ASAP7_75t_L g6852 ( 
.A(n_5219),
.Y(n_6852)
);

BUFx3_ASAP7_75t_L g6853 ( 
.A(n_5857),
.Y(n_6853)
);

NAND2xp5_ASAP7_75t_L g6854 ( 
.A(n_5895),
.B(n_4644),
.Y(n_6854)
);

OAI22xp5_ASAP7_75t_L g6855 ( 
.A1(n_5165),
.A2(n_5143),
.B1(n_5899),
.B2(n_5249),
.Y(n_6855)
);

AOI22xp33_ASAP7_75t_L g6856 ( 
.A1(n_5391),
.A2(n_4515),
.B1(n_4535),
.B2(n_4530),
.Y(n_6856)
);

OR2x2_ASAP7_75t_L g6857 ( 
.A(n_5726),
.B(n_4522),
.Y(n_6857)
);

HB1xp67_ASAP7_75t_L g6858 ( 
.A(n_5873),
.Y(n_6858)
);

INVx4_ASAP7_75t_L g6859 ( 
.A(n_5807),
.Y(n_6859)
);

INVx4_ASAP7_75t_L g6860 ( 
.A(n_5807),
.Y(n_6860)
);

INVx1_ASAP7_75t_L g6861 ( 
.A(n_5478),
.Y(n_6861)
);

BUFx2_ASAP7_75t_L g6862 ( 
.A(n_5219),
.Y(n_6862)
);

INVx1_ASAP7_75t_L g6863 ( 
.A(n_5478),
.Y(n_6863)
);

INVx1_ASAP7_75t_L g6864 ( 
.A(n_5483),
.Y(n_6864)
);

NOR2xp33_ASAP7_75t_L g6865 ( 
.A(n_5878),
.B(n_4936),
.Y(n_6865)
);

INVx4_ASAP7_75t_L g6866 ( 
.A(n_5833),
.Y(n_6866)
);

BUFx12f_ASAP7_75t_L g6867 ( 
.A(n_5514),
.Y(n_6867)
);

NAND2xp5_ASAP7_75t_L g6868 ( 
.A(n_5911),
.B(n_4646),
.Y(n_6868)
);

NAND2xp5_ASAP7_75t_L g6869 ( 
.A(n_5911),
.B(n_4646),
.Y(n_6869)
);

AOI22xp5_ASAP7_75t_L g6870 ( 
.A1(n_5143),
.A2(n_4881),
.B1(n_4785),
.B2(n_4959),
.Y(n_6870)
);

BUFx3_ASAP7_75t_L g6871 ( 
.A(n_5819),
.Y(n_6871)
);

HB1xp67_ASAP7_75t_L g6872 ( 
.A(n_5873),
.Y(n_6872)
);

OAI22xp5_ASAP7_75t_L g6873 ( 
.A1(n_5249),
.A2(n_4507),
.B1(n_4659),
.B2(n_4487),
.Y(n_6873)
);

AND2x2_ASAP7_75t_SL g6874 ( 
.A(n_6023),
.B(n_6031),
.Y(n_6874)
);

NOR2xp33_ASAP7_75t_SL g6875 ( 
.A(n_5833),
.B(n_4437),
.Y(n_6875)
);

NOR2xp33_ASAP7_75t_L g6876 ( 
.A(n_5212),
.B(n_4937),
.Y(n_6876)
);

AND2x2_ASAP7_75t_L g6877 ( 
.A(n_5934),
.B(n_5385),
.Y(n_6877)
);

INVx1_ASAP7_75t_L g6878 ( 
.A(n_5483),
.Y(n_6878)
);

O2A1O1Ixp5_ASAP7_75t_L g6879 ( 
.A1(n_5658),
.A2(n_4178),
.B(n_4213),
.C(n_4145),
.Y(n_6879)
);

OR2x2_ASAP7_75t_L g6880 ( 
.A(n_5751),
.B(n_4527),
.Y(n_6880)
);

NAND2xp5_ASAP7_75t_L g6881 ( 
.A(n_5937),
.B(n_4527),
.Y(n_6881)
);

BUFx3_ASAP7_75t_L g6882 ( 
.A(n_5819),
.Y(n_6882)
);

NAND2xp5_ASAP7_75t_L g6883 ( 
.A(n_5937),
.B(n_4527),
.Y(n_6883)
);

HB1xp67_ASAP7_75t_L g6884 ( 
.A(n_5918),
.Y(n_6884)
);

INVx1_ASAP7_75t_L g6885 ( 
.A(n_5485),
.Y(n_6885)
);

AOI21xp5_ASAP7_75t_L g6886 ( 
.A1(n_5599),
.A2(n_5621),
.B(n_5610),
.Y(n_6886)
);

INVx1_ASAP7_75t_L g6887 ( 
.A(n_5485),
.Y(n_6887)
);

HB1xp67_ASAP7_75t_L g6888 ( 
.A(n_5918),
.Y(n_6888)
);

INVx1_ASAP7_75t_L g6889 ( 
.A(n_5486),
.Y(n_6889)
);

INVx1_ASAP7_75t_L g6890 ( 
.A(n_5486),
.Y(n_6890)
);

BUFx2_ASAP7_75t_L g6891 ( 
.A(n_5225),
.Y(n_6891)
);

AOI21xp5_ASAP7_75t_L g6892 ( 
.A1(n_5621),
.A2(n_4530),
.B(n_4515),
.Y(n_6892)
);

CKINVDCx20_ASAP7_75t_R g6893 ( 
.A(n_5908),
.Y(n_6893)
);

NOR2xp33_ASAP7_75t_R g6894 ( 
.A(n_5961),
.B(n_4670),
.Y(n_6894)
);

NAND2xp5_ASAP7_75t_L g6895 ( 
.A(n_5836),
.B(n_4538),
.Y(n_6895)
);

NOR2xp33_ASAP7_75t_L g6896 ( 
.A(n_5212),
.B(n_4937),
.Y(n_6896)
);

NAND2xp5_ASAP7_75t_L g6897 ( 
.A(n_5921),
.B(n_4538),
.Y(n_6897)
);

CKINVDCx11_ASAP7_75t_R g6898 ( 
.A(n_5959),
.Y(n_6898)
);

CKINVDCx5p33_ASAP7_75t_R g6899 ( 
.A(n_5624),
.Y(n_6899)
);

AOI21xp5_ASAP7_75t_L g6900 ( 
.A1(n_5502),
.A2(n_4535),
.B(n_4530),
.Y(n_6900)
);

INVx1_ASAP7_75t_L g6901 ( 
.A(n_5496),
.Y(n_6901)
);

AND2x2_ASAP7_75t_L g6902 ( 
.A(n_5385),
.B(n_4427),
.Y(n_6902)
);

BUFx3_ASAP7_75t_L g6903 ( 
.A(n_5903),
.Y(n_6903)
);

NAND2xp5_ASAP7_75t_L g6904 ( 
.A(n_5238),
.B(n_4538),
.Y(n_6904)
);

CKINVDCx5p33_ASAP7_75t_R g6905 ( 
.A(n_5723),
.Y(n_6905)
);

AOI22xp33_ASAP7_75t_L g6906 ( 
.A1(n_5172),
.A2(n_4530),
.B1(n_4535),
.B2(n_4380),
.Y(n_6906)
);

NAND2xp5_ASAP7_75t_L g6907 ( 
.A(n_5238),
.B(n_5434),
.Y(n_6907)
);

INVx1_ASAP7_75t_L g6908 ( 
.A(n_5496),
.Y(n_6908)
);

INVx1_ASAP7_75t_L g6909 ( 
.A(n_5506),
.Y(n_6909)
);

AND2x2_ASAP7_75t_L g6910 ( 
.A(n_5385),
.B(n_4449),
.Y(n_6910)
);

CKINVDCx20_ASAP7_75t_R g6911 ( 
.A(n_6047),
.Y(n_6911)
);

AND2x2_ASAP7_75t_L g6912 ( 
.A(n_5356),
.B(n_4449),
.Y(n_6912)
);

OA21x2_ASAP7_75t_L g6913 ( 
.A1(n_6042),
.A2(n_4939),
.B(n_4935),
.Y(n_6913)
);

HB1xp67_ASAP7_75t_L g6914 ( 
.A(n_5923),
.Y(n_6914)
);

AOI21xp5_ASAP7_75t_L g6915 ( 
.A1(n_5502),
.A2(n_4535),
.B(n_4530),
.Y(n_6915)
);

NAND2xp5_ASAP7_75t_L g6916 ( 
.A(n_5434),
.B(n_4544),
.Y(n_6916)
);

INVx1_ASAP7_75t_L g6917 ( 
.A(n_5506),
.Y(n_6917)
);

AOI21xp5_ASAP7_75t_L g6918 ( 
.A1(n_5503),
.A2(n_4535),
.B(n_4530),
.Y(n_6918)
);

AOI22xp33_ASAP7_75t_L g6919 ( 
.A1(n_5172),
.A2(n_4530),
.B1(n_4535),
.B2(n_4380),
.Y(n_6919)
);

OR2x6_ASAP7_75t_L g6920 ( 
.A(n_5866),
.B(n_4437),
.Y(n_6920)
);

OR2x2_ASAP7_75t_L g6921 ( 
.A(n_5751),
.B(n_4544),
.Y(n_6921)
);

AOI21xp5_ASAP7_75t_L g6922 ( 
.A1(n_5503),
.A2(n_4535),
.B(n_4530),
.Y(n_6922)
);

BUFx8_ASAP7_75t_L g6923 ( 
.A(n_5500),
.Y(n_6923)
);

HB1xp67_ASAP7_75t_L g6924 ( 
.A(n_5923),
.Y(n_6924)
);

INVx1_ASAP7_75t_L g6925 ( 
.A(n_5511),
.Y(n_6925)
);

AOI22xp33_ASAP7_75t_L g6926 ( 
.A1(n_5586),
.A2(n_4535),
.B1(n_4666),
.B2(n_4380),
.Y(n_6926)
);

INVx4_ASAP7_75t_L g6927 ( 
.A(n_5187),
.Y(n_6927)
);

INVx1_ASAP7_75t_L g6928 ( 
.A(n_5511),
.Y(n_6928)
);

INVx1_ASAP7_75t_L g6929 ( 
.A(n_5529),
.Y(n_6929)
);

AND2x2_ASAP7_75t_L g6930 ( 
.A(n_5356),
.B(n_4455),
.Y(n_6930)
);

OR2x2_ASAP7_75t_L g6931 ( 
.A(n_5955),
.B(n_4544),
.Y(n_6931)
);

BUFx2_ASAP7_75t_L g6932 ( 
.A(n_5225),
.Y(n_6932)
);

INVx1_ASAP7_75t_SL g6933 ( 
.A(n_5326),
.Y(n_6933)
);

NAND2xp5_ASAP7_75t_L g6934 ( 
.A(n_5832),
.B(n_4551),
.Y(n_6934)
);

INVx8_ASAP7_75t_L g6935 ( 
.A(n_5952),
.Y(n_6935)
);

OAI22xp5_ASAP7_75t_L g6936 ( 
.A1(n_5226),
.A2(n_4676),
.B1(n_4686),
.B2(n_4659),
.Y(n_6936)
);

AOI22xp33_ASAP7_75t_L g6937 ( 
.A1(n_5586),
.A2(n_4535),
.B1(n_4666),
.B2(n_4380),
.Y(n_6937)
);

BUFx3_ASAP7_75t_L g6938 ( 
.A(n_5903),
.Y(n_6938)
);

BUFx12f_ASAP7_75t_L g6939 ( 
.A(n_5944),
.Y(n_6939)
);

AND2x2_ASAP7_75t_L g6940 ( 
.A(n_5356),
.B(n_4455),
.Y(n_6940)
);

CKINVDCx5p33_ASAP7_75t_R g6941 ( 
.A(n_5727),
.Y(n_6941)
);

OAI22xp33_ASAP7_75t_L g6942 ( 
.A1(n_5904),
.A2(n_4795),
.B1(n_4809),
.B2(n_4747),
.Y(n_6942)
);

OR2x6_ASAP7_75t_L g6943 ( 
.A(n_5866),
.B(n_4473),
.Y(n_6943)
);

BUFx3_ASAP7_75t_L g6944 ( 
.A(n_5903),
.Y(n_6944)
);

NAND2xp5_ASAP7_75t_L g6945 ( 
.A(n_5832),
.B(n_4551),
.Y(n_6945)
);

AOI22xp5_ASAP7_75t_L g6946 ( 
.A1(n_5134),
.A2(n_4881),
.B1(n_4785),
.B2(n_4959),
.Y(n_6946)
);

NAND2xp5_ASAP7_75t_SL g6947 ( 
.A(n_6067),
.B(n_4676),
.Y(n_6947)
);

NAND2xp5_ASAP7_75t_L g6948 ( 
.A(n_5890),
.B(n_4551),
.Y(n_6948)
);

INVx5_ASAP7_75t_L g6949 ( 
.A(n_5301),
.Y(n_6949)
);

AOI221xp5_ASAP7_75t_L g6950 ( 
.A1(n_5785),
.A2(n_4562),
.B1(n_4568),
.B2(n_4566),
.C(n_4558),
.Y(n_6950)
);

BUFx2_ASAP7_75t_L g6951 ( 
.A(n_5225),
.Y(n_6951)
);

INVx2_ASAP7_75t_SL g6952 ( 
.A(n_6023),
.Y(n_6952)
);

NAND2xp5_ASAP7_75t_L g6953 ( 
.A(n_5890),
.B(n_5912),
.Y(n_6953)
);

AOI21xp5_ASAP7_75t_L g6954 ( 
.A1(n_5867),
.A2(n_4460),
.B(n_4455),
.Y(n_6954)
);

INVx1_ASAP7_75t_L g6955 ( 
.A(n_5529),
.Y(n_6955)
);

AND2x2_ASAP7_75t_L g6956 ( 
.A(n_5369),
.B(n_4460),
.Y(n_6956)
);

HB1xp67_ASAP7_75t_L g6957 ( 
.A(n_5948),
.Y(n_6957)
);

INVx1_ASAP7_75t_L g6958 ( 
.A(n_5536),
.Y(n_6958)
);

INVxp67_ASAP7_75t_SL g6959 ( 
.A(n_5681),
.Y(n_6959)
);

CKINVDCx5p33_ASAP7_75t_R g6960 ( 
.A(n_5750),
.Y(n_6960)
);

BUFx2_ASAP7_75t_L g6961 ( 
.A(n_5225),
.Y(n_6961)
);

BUFx2_ASAP7_75t_L g6962 ( 
.A(n_5225),
.Y(n_6962)
);

INVx1_ASAP7_75t_L g6963 ( 
.A(n_5536),
.Y(n_6963)
);

BUFx12f_ASAP7_75t_L g6964 ( 
.A(n_5944),
.Y(n_6964)
);

CKINVDCx20_ASAP7_75t_R g6965 ( 
.A(n_6020),
.Y(n_6965)
);

INVx5_ASAP7_75t_L g6966 ( 
.A(n_5301),
.Y(n_6966)
);

OR2x2_ASAP7_75t_L g6967 ( 
.A(n_5955),
.B(n_4558),
.Y(n_6967)
);

INVx1_ASAP7_75t_L g6968 ( 
.A(n_5550),
.Y(n_6968)
);

INVx1_ASAP7_75t_L g6969 ( 
.A(n_5550),
.Y(n_6969)
);

O2A1O1Ixp33_ASAP7_75t_SL g6970 ( 
.A1(n_5665),
.A2(n_5093),
.B(n_5044),
.C(n_4558),
.Y(n_6970)
);

CKINVDCx5p33_ASAP7_75t_R g6971 ( 
.A(n_5862),
.Y(n_6971)
);

NAND2xp5_ASAP7_75t_L g6972 ( 
.A(n_5912),
.B(n_4562),
.Y(n_6972)
);

INVx1_ASAP7_75t_L g6973 ( 
.A(n_5555),
.Y(n_6973)
);

INVx1_ASAP7_75t_L g6974 ( 
.A(n_5555),
.Y(n_6974)
);

NOR3xp33_ASAP7_75t_L g6975 ( 
.A(n_5428),
.B(n_5269),
.C(n_5226),
.Y(n_6975)
);

NAND2x1_ASAP7_75t_L g6976 ( 
.A(n_5985),
.B(n_4815),
.Y(n_6976)
);

INVx1_ASAP7_75t_L g6977 ( 
.A(n_5557),
.Y(n_6977)
);

BUFx2_ASAP7_75t_L g6978 ( 
.A(n_5232),
.Y(n_6978)
);

OAI22xp5_ASAP7_75t_L g6979 ( 
.A1(n_5339),
.A2(n_4686),
.B1(n_4733),
.B2(n_4676),
.Y(n_6979)
);

BUFx2_ASAP7_75t_SL g6980 ( 
.A(n_5542),
.Y(n_6980)
);

AO22x1_ASAP7_75t_L g6981 ( 
.A1(n_6067),
.A2(n_6089),
.B1(n_6126),
.B2(n_6108),
.Y(n_6981)
);

AOI222xp33_ASAP7_75t_L g6982 ( 
.A1(n_5785),
.A2(n_4838),
.B1(n_4826),
.B2(n_4845),
.C1(n_4829),
.C2(n_4824),
.Y(n_6982)
);

INVx8_ASAP7_75t_L g6983 ( 
.A(n_5952),
.Y(n_6983)
);

NAND2xp5_ASAP7_75t_L g6984 ( 
.A(n_5935),
.B(n_4562),
.Y(n_6984)
);

AOI22xp33_ASAP7_75t_L g6985 ( 
.A1(n_5785),
.A2(n_4666),
.B1(n_5095),
.B2(n_4529),
.Y(n_6985)
);

HB1xp67_ASAP7_75t_L g6986 ( 
.A(n_5948),
.Y(n_6986)
);

BUFx2_ASAP7_75t_SL g6987 ( 
.A(n_5542),
.Y(n_6987)
);

CKINVDCx8_ASAP7_75t_R g6988 ( 
.A(n_5415),
.Y(n_6988)
);

OR2x2_ASAP7_75t_L g6989 ( 
.A(n_5972),
.B(n_4566),
.Y(n_6989)
);

INVx4_ASAP7_75t_L g6990 ( 
.A(n_5187),
.Y(n_6990)
);

INVx1_ASAP7_75t_L g6991 ( 
.A(n_5557),
.Y(n_6991)
);

INVx3_ASAP7_75t_SL g6992 ( 
.A(n_5781),
.Y(n_6992)
);

OAI22xp5_ASAP7_75t_L g6993 ( 
.A1(n_5180),
.A2(n_4733),
.B1(n_4686),
.B2(n_4964),
.Y(n_6993)
);

INVx1_ASAP7_75t_L g6994 ( 
.A(n_5558),
.Y(n_6994)
);

OAI21xp5_ASAP7_75t_L g6995 ( 
.A1(n_5381),
.A2(n_5622),
.B(n_5147),
.Y(n_6995)
);

AOI21xp33_ASAP7_75t_L g6996 ( 
.A1(n_5957),
.A2(n_4860),
.B(n_4853),
.Y(n_6996)
);

AOI22xp33_ASAP7_75t_SL g6997 ( 
.A1(n_5568),
.A2(n_5500),
.B1(n_6108),
.B2(n_6089),
.Y(n_6997)
);

OR2x2_ASAP7_75t_L g6998 ( 
.A(n_5972),
.B(n_4566),
.Y(n_6998)
);

INVx4_ASAP7_75t_L g6999 ( 
.A(n_5187),
.Y(n_6999)
);

NAND2xp5_ASAP7_75t_SL g7000 ( 
.A(n_6089),
.B(n_4686),
.Y(n_7000)
);

CKINVDCx16_ASAP7_75t_R g7001 ( 
.A(n_5902),
.Y(n_7001)
);

HB1xp67_ASAP7_75t_L g7002 ( 
.A(n_5844),
.Y(n_7002)
);

NAND2xp5_ASAP7_75t_L g7003 ( 
.A(n_5935),
.B(n_4568),
.Y(n_7003)
);

CKINVDCx5p33_ASAP7_75t_R g7004 ( 
.A(n_5949),
.Y(n_7004)
);

NAND2xp5_ASAP7_75t_L g7005 ( 
.A(n_6012),
.B(n_4568),
.Y(n_7005)
);

A2O1A1Ixp33_ASAP7_75t_L g7006 ( 
.A1(n_5207),
.A2(n_4733),
.B(n_4686),
.C(n_4785),
.Y(n_7006)
);

NOR3xp33_ASAP7_75t_L g7007 ( 
.A(n_5269),
.B(n_5026),
.C(n_4423),
.Y(n_7007)
);

BUFx3_ASAP7_75t_L g7008 ( 
.A(n_5966),
.Y(n_7008)
);

AOI22xp33_ASAP7_75t_L g7009 ( 
.A1(n_5512),
.A2(n_5523),
.B1(n_5180),
.B2(n_5581),
.Y(n_7009)
);

AOI22xp33_ASAP7_75t_L g7010 ( 
.A1(n_5512),
.A2(n_4666),
.B1(n_5095),
.B2(n_4529),
.Y(n_7010)
);

OR2x6_ASAP7_75t_L g7011 ( 
.A(n_5588),
.B(n_4473),
.Y(n_7011)
);

BUFx3_ASAP7_75t_L g7012 ( 
.A(n_5966),
.Y(n_7012)
);

NAND2xp5_ASAP7_75t_L g7013 ( 
.A(n_6012),
.B(n_4569),
.Y(n_7013)
);

AOI22xp33_ASAP7_75t_L g7014 ( 
.A1(n_5523),
.A2(n_5095),
.B1(n_4529),
.B2(n_4583),
.Y(n_7014)
);

AOI21xp5_ASAP7_75t_L g7015 ( 
.A1(n_5306),
.A2(n_4533),
.B(n_4468),
.Y(n_7015)
);

AOI21xp5_ASAP7_75t_L g7016 ( 
.A1(n_5306),
.A2(n_4533),
.B(n_4468),
.Y(n_7016)
);

AOI222xp33_ASAP7_75t_L g7017 ( 
.A1(n_5581),
.A2(n_4870),
.B1(n_4860),
.B2(n_4871),
.C1(n_4867),
.C2(n_4853),
.Y(n_7017)
);

OR2x2_ASAP7_75t_SL g7018 ( 
.A(n_5500),
.B(n_4274),
.Y(n_7018)
);

NAND2xp5_ASAP7_75t_L g7019 ( 
.A(n_6094),
.B(n_4569),
.Y(n_7019)
);

INVx2_ASAP7_75t_SL g7020 ( 
.A(n_6031),
.Y(n_7020)
);

AOI21xp5_ASAP7_75t_L g7021 ( 
.A1(n_5957),
.A2(n_4533),
.B(n_4468),
.Y(n_7021)
);

NAND2xp5_ASAP7_75t_L g7022 ( 
.A(n_6094),
.B(n_4569),
.Y(n_7022)
);

BUFx12f_ASAP7_75t_L g7023 ( 
.A(n_5944),
.Y(n_7023)
);

INVxp67_ASAP7_75t_L g7024 ( 
.A(n_5973),
.Y(n_7024)
);

INVxp67_ASAP7_75t_SL g7025 ( 
.A(n_6001),
.Y(n_7025)
);

INVx8_ASAP7_75t_L g7026 ( 
.A(n_5952),
.Y(n_7026)
);

INVx1_ASAP7_75t_SL g7027 ( 
.A(n_5332),
.Y(n_7027)
);

INVx1_ASAP7_75t_SL g7028 ( 
.A(n_5332),
.Y(n_7028)
);

A2O1A1Ixp33_ASAP7_75t_L g7029 ( 
.A1(n_5207),
.A2(n_4733),
.B(n_4686),
.C(n_4785),
.Y(n_7029)
);

INVx4_ASAP7_75t_L g7030 ( 
.A(n_6097),
.Y(n_7030)
);

AOI22xp5_ASAP7_75t_L g7031 ( 
.A1(n_5392),
.A2(n_4881),
.B1(n_5093),
.B2(n_4529),
.Y(n_7031)
);

CKINVDCx6p67_ASAP7_75t_R g7032 ( 
.A(n_5738),
.Y(n_7032)
);

CKINVDCx5p33_ASAP7_75t_R g7033 ( 
.A(n_5342),
.Y(n_7033)
);

AOI21xp5_ASAP7_75t_L g7034 ( 
.A1(n_5625),
.A2(n_4593),
.B(n_4564),
.Y(n_7034)
);

NAND2xp5_ASAP7_75t_L g7035 ( 
.A(n_6101),
.B(n_5801),
.Y(n_7035)
);

HB1xp67_ASAP7_75t_L g7036 ( 
.A(n_5844),
.Y(n_7036)
);

AOI21xp5_ASAP7_75t_L g7037 ( 
.A1(n_5625),
.A2(n_4593),
.B(n_4564),
.Y(n_7037)
);

AND2x2_ASAP7_75t_L g7038 ( 
.A(n_5950),
.B(n_5980),
.Y(n_7038)
);

BUFx12f_ASAP7_75t_L g7039 ( 
.A(n_5944),
.Y(n_7039)
);

AOI22xp5_ASAP7_75t_L g7040 ( 
.A1(n_5392),
.A2(n_4881),
.B1(n_4529),
.B2(n_4583),
.Y(n_7040)
);

AOI22xp33_ASAP7_75t_L g7041 ( 
.A1(n_5202),
.A2(n_5095),
.B1(n_4529),
.B2(n_4583),
.Y(n_7041)
);

NAND2xp5_ASAP7_75t_L g7042 ( 
.A(n_6101),
.B(n_5801),
.Y(n_7042)
);

CKINVDCx6p67_ASAP7_75t_R g7043 ( 
.A(n_5738),
.Y(n_7043)
);

AOI221xp5_ASAP7_75t_L g7044 ( 
.A1(n_5777),
.A2(n_4600),
.B1(n_4603),
.B2(n_4597),
.C(n_4592),
.Y(n_7044)
);

INVx1_ASAP7_75t_SL g7045 ( 
.A(n_5338),
.Y(n_7045)
);

OAI21x1_ASAP7_75t_L g7046 ( 
.A1(n_6049),
.A2(n_5652),
.B(n_5996),
.Y(n_7046)
);

HB1xp67_ASAP7_75t_L g7047 ( 
.A(n_5863),
.Y(n_7047)
);

INVx4_ASAP7_75t_L g7048 ( 
.A(n_6097),
.Y(n_7048)
);

NOR2xp33_ASAP7_75t_L g7049 ( 
.A(n_5828),
.B(n_4964),
.Y(n_7049)
);

INVxp67_ASAP7_75t_L g7050 ( 
.A(n_5973),
.Y(n_7050)
);

INVx4_ASAP7_75t_L g7051 ( 
.A(n_6097),
.Y(n_7051)
);

CKINVDCx8_ASAP7_75t_R g7052 ( 
.A(n_5415),
.Y(n_7052)
);

INVx2_ASAP7_75t_SL g7053 ( 
.A(n_6031),
.Y(n_7053)
);

NOR2xp67_ASAP7_75t_L g7054 ( 
.A(n_5966),
.B(n_4747),
.Y(n_7054)
);

AOI21xp5_ASAP7_75t_L g7055 ( 
.A1(n_5622),
.A2(n_4617),
.B(n_4593),
.Y(n_7055)
);

BUFx8_ASAP7_75t_SL g7056 ( 
.A(n_6096),
.Y(n_7056)
);

AOI21xp5_ASAP7_75t_L g7057 ( 
.A1(n_5843),
.A2(n_5928),
.B(n_5906),
.Y(n_7057)
);

INVxp67_ASAP7_75t_L g7058 ( 
.A(n_5975),
.Y(n_7058)
);

OR2x6_ASAP7_75t_L g7059 ( 
.A(n_5588),
.B(n_4473),
.Y(n_7059)
);

AND3x1_ASAP7_75t_SL g7060 ( 
.A(n_5896),
.B(n_4682),
.C(n_4670),
.Y(n_7060)
);

INVxp67_ASAP7_75t_SL g7061 ( 
.A(n_6001),
.Y(n_7061)
);

INVx2_ASAP7_75t_SL g7062 ( 
.A(n_6031),
.Y(n_7062)
);

NAND2xp5_ASAP7_75t_SL g7063 ( 
.A(n_6108),
.B(n_4747),
.Y(n_7063)
);

NOR2x1_ASAP7_75t_L g7064 ( 
.A(n_5315),
.B(n_4815),
.Y(n_7064)
);

O2A1O1Ixp5_ASAP7_75t_L g7065 ( 
.A1(n_6003),
.A2(n_4178),
.B(n_4213),
.C(n_4145),
.Y(n_7065)
);

OR2x2_ASAP7_75t_L g7066 ( 
.A(n_5975),
.B(n_4592),
.Y(n_7066)
);

HB1xp67_ASAP7_75t_L g7067 ( 
.A(n_5863),
.Y(n_7067)
);

AOI21xp5_ASAP7_75t_L g7068 ( 
.A1(n_5843),
.A2(n_4660),
.B(n_4617),
.Y(n_7068)
);

NAND2xp5_ASAP7_75t_L g7069 ( 
.A(n_5906),
.B(n_4592),
.Y(n_7069)
);

OR2x6_ASAP7_75t_L g7070 ( 
.A(n_5588),
.B(n_4473),
.Y(n_7070)
);

INVx4_ASAP7_75t_L g7071 ( 
.A(n_6097),
.Y(n_7071)
);

NAND2xp5_ASAP7_75t_L g7072 ( 
.A(n_5928),
.B(n_4597),
.Y(n_7072)
);

INVx2_ASAP7_75t_SL g7073 ( 
.A(n_6031),
.Y(n_7073)
);

CKINVDCx5p33_ASAP7_75t_R g7074 ( 
.A(n_5347),
.Y(n_7074)
);

NAND2xp5_ASAP7_75t_L g7075 ( 
.A(n_5840),
.B(n_5976),
.Y(n_7075)
);

NAND2xp5_ASAP7_75t_L g7076 ( 
.A(n_5840),
.B(n_4597),
.Y(n_7076)
);

CKINVDCx5p33_ASAP7_75t_R g7077 ( 
.A(n_6119),
.Y(n_7077)
);

OAI22xp5_ASAP7_75t_L g7078 ( 
.A1(n_5904),
.A2(n_5914),
.B1(n_5930),
.B2(n_5922),
.Y(n_7078)
);

AOI21xp33_ASAP7_75t_L g7079 ( 
.A1(n_5397),
.A2(n_4860),
.B(n_4853),
.Y(n_7079)
);

CKINVDCx5p33_ASAP7_75t_R g7080 ( 
.A(n_6064),
.Y(n_7080)
);

BUFx12f_ASAP7_75t_L g7081 ( 
.A(n_5944),
.Y(n_7081)
);

NOR2xp33_ASAP7_75t_L g7082 ( 
.A(n_5838),
.B(n_4673),
.Y(n_7082)
);

INVx5_ASAP7_75t_L g7083 ( 
.A(n_5301),
.Y(n_7083)
);

INVxp67_ASAP7_75t_L g7084 ( 
.A(n_5976),
.Y(n_7084)
);

OAI22xp5_ASAP7_75t_L g7085 ( 
.A1(n_5914),
.A2(n_4603),
.B1(n_4604),
.B2(n_4600),
.Y(n_7085)
);

NOR2xp33_ASAP7_75t_L g7086 ( 
.A(n_5922),
.B(n_5930),
.Y(n_7086)
);

INVx5_ASAP7_75t_L g7087 ( 
.A(n_5301),
.Y(n_7087)
);

CKINVDCx5p33_ASAP7_75t_R g7088 ( 
.A(n_6064),
.Y(n_7088)
);

INVx4_ASAP7_75t_SL g7089 ( 
.A(n_5588),
.Y(n_7089)
);

NOR2xp33_ASAP7_75t_L g7090 ( 
.A(n_5931),
.B(n_4687),
.Y(n_7090)
);

AND2x2_ASAP7_75t_L g7091 ( 
.A(n_6009),
.B(n_6028),
.Y(n_7091)
);

AOI22xp5_ASAP7_75t_L g7092 ( 
.A1(n_5278),
.A2(n_4881),
.B1(n_4529),
.B2(n_4583),
.Y(n_7092)
);

HB1xp67_ASAP7_75t_L g7093 ( 
.A(n_5513),
.Y(n_7093)
);

NAND2xp5_ASAP7_75t_L g7094 ( 
.A(n_6021),
.B(n_4600),
.Y(n_7094)
);

AOI21xp5_ASAP7_75t_L g7095 ( 
.A1(n_5968),
.A2(n_4704),
.B(n_4693),
.Y(n_7095)
);

INVx2_ASAP7_75t_SL g7096 ( 
.A(n_6038),
.Y(n_7096)
);

INVxp67_ASAP7_75t_L g7097 ( 
.A(n_5513),
.Y(n_7097)
);

BUFx3_ASAP7_75t_L g7098 ( 
.A(n_5106),
.Y(n_7098)
);

NAND2xp5_ASAP7_75t_L g7099 ( 
.A(n_6021),
.B(n_4603),
.Y(n_7099)
);

AOI21xp5_ASAP7_75t_L g7100 ( 
.A1(n_5968),
.A2(n_4704),
.B(n_4693),
.Y(n_7100)
);

HB1xp67_ASAP7_75t_L g7101 ( 
.A(n_5519),
.Y(n_7101)
);

BUFx3_ASAP7_75t_L g7102 ( 
.A(n_5106),
.Y(n_7102)
);

OR2x6_ASAP7_75t_L g7103 ( 
.A(n_5588),
.B(n_4473),
.Y(n_7103)
);

OAI21xp33_ASAP7_75t_L g7104 ( 
.A1(n_5758),
.A2(n_4615),
.B(n_4604),
.Y(n_7104)
);

NAND2xp5_ASAP7_75t_SL g7105 ( 
.A(n_6126),
.B(n_4747),
.Y(n_7105)
);

OAI22xp33_ASAP7_75t_L g7106 ( 
.A1(n_6126),
.A2(n_4795),
.B1(n_4809),
.B2(n_4747),
.Y(n_7106)
);

AOI21xp5_ASAP7_75t_L g7107 ( 
.A1(n_5805),
.A2(n_4704),
.B(n_4693),
.Y(n_7107)
);

INVx2_ASAP7_75t_SL g7108 ( 
.A(n_6038),
.Y(n_7108)
);

BUFx3_ASAP7_75t_L g7109 ( 
.A(n_5106),
.Y(n_7109)
);

BUFx3_ASAP7_75t_L g7110 ( 
.A(n_5106),
.Y(n_7110)
);

BUFx6f_ASAP7_75t_SL g7111 ( 
.A(n_5765),
.Y(n_7111)
);

AND2x4_ASAP7_75t_SL g7112 ( 
.A(n_6038),
.B(n_4501),
.Y(n_7112)
);

OR2x2_ASAP7_75t_L g7113 ( 
.A(n_5213),
.B(n_4604),
.Y(n_7113)
);

NAND2xp5_ASAP7_75t_L g7114 ( 
.A(n_6053),
.B(n_4615),
.Y(n_7114)
);

NAND2xp5_ASAP7_75t_L g7115 ( 
.A(n_6053),
.B(n_4615),
.Y(n_7115)
);

NAND2x1_ASAP7_75t_L g7116 ( 
.A(n_5985),
.B(n_4815),
.Y(n_7116)
);

AOI22xp33_ASAP7_75t_L g7117 ( 
.A1(n_5202),
.A2(n_5095),
.B1(n_4529),
.B2(n_4583),
.Y(n_7117)
);

CKINVDCx20_ASAP7_75t_R g7118 ( 
.A(n_6061),
.Y(n_7118)
);

AOI22xp33_ASAP7_75t_L g7119 ( 
.A1(n_5570),
.A2(n_5095),
.B1(n_4583),
.B2(n_4595),
.Y(n_7119)
);

BUFx3_ASAP7_75t_L g7120 ( 
.A(n_5106),
.Y(n_7120)
);

A2O1A1Ixp33_ASAP7_75t_L g7121 ( 
.A1(n_5260),
.A2(n_4965),
.B(n_4961),
.C(n_4420),
.Y(n_7121)
);

HB1xp67_ASAP7_75t_L g7122 ( 
.A(n_5519),
.Y(n_7122)
);

HB1xp67_ASAP7_75t_L g7123 ( 
.A(n_5559),
.Y(n_7123)
);

OR2x2_ASAP7_75t_L g7124 ( 
.A(n_5213),
.B(n_4619),
.Y(n_7124)
);

NAND2xp5_ASAP7_75t_L g7125 ( 
.A(n_5804),
.B(n_4619),
.Y(n_7125)
);

OAI22xp5_ASAP7_75t_L g7126 ( 
.A1(n_5931),
.A2(n_4619),
.B1(n_4625),
.B2(n_4622),
.Y(n_7126)
);

OAI22xp5_ASAP7_75t_L g7127 ( 
.A1(n_5898),
.A2(n_4622),
.B1(n_4630),
.B2(n_4625),
.Y(n_7127)
);

BUFx6f_ASAP7_75t_L g7128 ( 
.A(n_5333),
.Y(n_7128)
);

BUFx6f_ASAP7_75t_L g7129 ( 
.A(n_5333),
.Y(n_7129)
);

HB1xp67_ASAP7_75t_L g7130 ( 
.A(n_5559),
.Y(n_7130)
);

HB1xp67_ASAP7_75t_L g7131 ( 
.A(n_5562),
.Y(n_7131)
);

INVx3_ASAP7_75t_SL g7132 ( 
.A(n_5781),
.Y(n_7132)
);

NOR2xp67_ASAP7_75t_L g7133 ( 
.A(n_5138),
.B(n_4795),
.Y(n_7133)
);

INVx3_ASAP7_75t_L g7134 ( 
.A(n_5250),
.Y(n_7134)
);

NOR2xp33_ASAP7_75t_L g7135 ( 
.A(n_5668),
.B(n_5679),
.Y(n_7135)
);

BUFx6f_ASAP7_75t_L g7136 ( 
.A(n_5333),
.Y(n_7136)
);

INVx8_ASAP7_75t_L g7137 ( 
.A(n_5952),
.Y(n_7137)
);

INVx2_ASAP7_75t_SL g7138 ( 
.A(n_6038),
.Y(n_7138)
);

NAND2xp5_ASAP7_75t_L g7139 ( 
.A(n_5804),
.B(n_4622),
.Y(n_7139)
);

OR2x2_ASAP7_75t_L g7140 ( 
.A(n_5213),
.B(n_4625),
.Y(n_7140)
);

AOI21xp5_ASAP7_75t_L g7141 ( 
.A1(n_5474),
.A2(n_4732),
.B(n_4717),
.Y(n_7141)
);

CKINVDCx5p33_ASAP7_75t_R g7142 ( 
.A(n_6046),
.Y(n_7142)
);

NOR2xp33_ASAP7_75t_SL g7143 ( 
.A(n_5902),
.B(n_4795),
.Y(n_7143)
);

BUFx2_ASAP7_75t_L g7144 ( 
.A(n_5250),
.Y(n_7144)
);

AOI22xp33_ASAP7_75t_L g7145 ( 
.A1(n_5570),
.A2(n_4583),
.B1(n_4595),
.B2(n_4501),
.Y(n_7145)
);

BUFx2_ASAP7_75t_L g7146 ( 
.A(n_5250),
.Y(n_7146)
);

NAND2xp5_ASAP7_75t_L g7147 ( 
.A(n_5815),
.B(n_5820),
.Y(n_7147)
);

NOR2xp33_ASAP7_75t_SL g7148 ( 
.A(n_5986),
.B(n_4795),
.Y(n_7148)
);

O2A1O1Ixp33_ASAP7_75t_L g7149 ( 
.A1(n_5896),
.A2(n_5020),
.B(n_5045),
.C(n_4947),
.Y(n_7149)
);

NAND2xp5_ASAP7_75t_L g7150 ( 
.A(n_5815),
.B(n_5820),
.Y(n_7150)
);

INVx6_ASAP7_75t_L g7151 ( 
.A(n_5127),
.Y(n_7151)
);

HB1xp67_ASAP7_75t_L g7152 ( 
.A(n_5562),
.Y(n_7152)
);

INVx3_ASAP7_75t_L g7153 ( 
.A(n_5250),
.Y(n_7153)
);

BUFx6f_ASAP7_75t_L g7154 ( 
.A(n_5333),
.Y(n_7154)
);

BUFx2_ASAP7_75t_SL g7155 ( 
.A(n_5575),
.Y(n_7155)
);

INVx1_ASAP7_75t_L g7156 ( 
.A(n_6130),
.Y(n_7156)
);

AOI222xp33_ASAP7_75t_L g7157 ( 
.A1(n_6203),
.A2(n_5203),
.B1(n_5381),
.B2(n_5255),
.C1(n_5593),
.C2(n_5216),
.Y(n_7157)
);

INVx4_ASAP7_75t_L g7158 ( 
.A(n_6237),
.Y(n_7158)
);

INVx3_ASAP7_75t_SL g7159 ( 
.A(n_6182),
.Y(n_7159)
);

OAI22x1_ASAP7_75t_L g7160 ( 
.A1(n_6379),
.A2(n_5397),
.B1(n_5602),
.B2(n_5535),
.Y(n_7160)
);

INVx3_ASAP7_75t_L g7161 ( 
.A(n_6132),
.Y(n_7161)
);

OAI21x1_ASAP7_75t_L g7162 ( 
.A1(n_6320),
.A2(n_6049),
.B(n_5439),
.Y(n_7162)
);

INVx1_ASAP7_75t_L g7163 ( 
.A(n_6130),
.Y(n_7163)
);

NAND2x1p5_ASAP7_75t_L g7164 ( 
.A(n_6462),
.B(n_5138),
.Y(n_7164)
);

AOI22x1_ASAP7_75t_L g7165 ( 
.A1(n_6995),
.A2(n_6278),
.B1(n_6886),
.B2(n_7057),
.Y(n_7165)
);

NOR2xp33_ASAP7_75t_L g7166 ( 
.A(n_6500),
.B(n_6059),
.Y(n_7166)
);

OAI21x1_ASAP7_75t_L g7167 ( 
.A1(n_6320),
.A2(n_5439),
.B(n_5652),
.Y(n_7167)
);

OA21x2_ASAP7_75t_L g7168 ( 
.A1(n_6294),
.A2(n_6048),
.B(n_5875),
.Y(n_7168)
);

AO32x2_ASAP7_75t_L g7169 ( 
.A1(n_7126),
.A2(n_6059),
.A3(n_6071),
.B1(n_5829),
.B2(n_5824),
.Y(n_7169)
);

AOI21xp5_ASAP7_75t_L g7170 ( 
.A1(n_6508),
.A2(n_6294),
.B(n_6278),
.Y(n_7170)
);

AND2x4_ASAP7_75t_L g7171 ( 
.A(n_6132),
.B(n_6038),
.Y(n_7171)
);

AOI221x1_ASAP7_75t_L g7172 ( 
.A1(n_6146),
.A2(n_6003),
.B1(n_5308),
.B2(n_5592),
.C(n_5349),
.Y(n_7172)
);

BUFx6f_ASAP7_75t_L g7173 ( 
.A(n_6137),
.Y(n_7173)
);

AND2x4_ASAP7_75t_L g7174 ( 
.A(n_6132),
.B(n_6196),
.Y(n_7174)
);

OAI21x1_ASAP7_75t_L g7175 ( 
.A1(n_6488),
.A2(n_5997),
.B(n_5996),
.Y(n_7175)
);

HB1xp67_ASAP7_75t_L g7176 ( 
.A(n_6914),
.Y(n_7176)
);

OAI21x1_ASAP7_75t_L g7177 ( 
.A1(n_6488),
.A2(n_6000),
.B(n_5997),
.Y(n_7177)
);

AND2x4_ASAP7_75t_L g7178 ( 
.A(n_6132),
.B(n_6057),
.Y(n_7178)
);

AO31x2_ASAP7_75t_L g7179 ( 
.A1(n_7085),
.A2(n_5954),
.A3(n_5953),
.B(n_5884),
.Y(n_7179)
);

AND2x2_ASAP7_75t_L g7180 ( 
.A(n_6145),
.B(n_5752),
.Y(n_7180)
);

OA21x2_ASAP7_75t_L g7181 ( 
.A1(n_7046),
.A2(n_5875),
.B(n_5852),
.Y(n_7181)
);

AO31x2_ASAP7_75t_L g7182 ( 
.A1(n_7085),
.A2(n_6338),
.A3(n_7127),
.B(n_6238),
.Y(n_7182)
);

INVx2_ASAP7_75t_L g7183 ( 
.A(n_6657),
.Y(n_7183)
);

INVx1_ASAP7_75t_SL g7184 ( 
.A(n_6152),
.Y(n_7184)
);

AOI21xp5_ASAP7_75t_L g7185 ( 
.A1(n_6508),
.A2(n_5470),
.B(n_5508),
.Y(n_7185)
);

OAI21x1_ASAP7_75t_L g7186 ( 
.A1(n_6328),
.A2(n_6011),
.B(n_6000),
.Y(n_7186)
);

BUFx6f_ASAP7_75t_L g7187 ( 
.A(n_6137),
.Y(n_7187)
);

OAI21x1_ASAP7_75t_L g7188 ( 
.A1(n_6328),
.A2(n_6045),
.B(n_6011),
.Y(n_7188)
);

INVx1_ASAP7_75t_L g7189 ( 
.A(n_6130),
.Y(n_7189)
);

BUFx3_ASAP7_75t_L g7190 ( 
.A(n_6636),
.Y(n_7190)
);

OR2x6_ASAP7_75t_L g7191 ( 
.A(n_6222),
.B(n_5588),
.Y(n_7191)
);

INVx1_ASAP7_75t_L g7192 ( 
.A(n_6139),
.Y(n_7192)
);

AOI221xp5_ASAP7_75t_L g7193 ( 
.A1(n_6693),
.A2(n_5602),
.B1(n_5940),
.B2(n_5932),
.C(n_5852),
.Y(n_7193)
);

NAND2xp5_ASAP7_75t_L g7194 ( 
.A(n_7035),
.B(n_7042),
.Y(n_7194)
);

BUFx2_ASAP7_75t_SL g7195 ( 
.A(n_7054),
.Y(n_7195)
);

OAI21x1_ASAP7_75t_L g7196 ( 
.A1(n_6371),
.A2(n_6915),
.B(n_6900),
.Y(n_7196)
);

CKINVDCx5p33_ASAP7_75t_R g7197 ( 
.A(n_6601),
.Y(n_7197)
);

OAI21x1_ASAP7_75t_L g7198 ( 
.A1(n_6371),
.A2(n_6052),
.B(n_6045),
.Y(n_7198)
);

NAND2xp5_ASAP7_75t_L g7199 ( 
.A(n_7035),
.B(n_5846),
.Y(n_7199)
);

NAND2x1p5_ASAP7_75t_L g7200 ( 
.A(n_6462),
.B(n_5150),
.Y(n_7200)
);

AO31x2_ASAP7_75t_L g7201 ( 
.A1(n_6338),
.A2(n_5592),
.A3(n_5504),
.B(n_5593),
.Y(n_7201)
);

HB1xp67_ASAP7_75t_L g7202 ( 
.A(n_6914),
.Y(n_7202)
);

AND2x2_ASAP7_75t_L g7203 ( 
.A(n_6145),
.B(n_5752),
.Y(n_7203)
);

INVx1_ASAP7_75t_L g7204 ( 
.A(n_6139),
.Y(n_7204)
);

OAI21x1_ASAP7_75t_L g7205 ( 
.A1(n_6900),
.A2(n_6055),
.B(n_6052),
.Y(n_7205)
);

BUFx6f_ASAP7_75t_L g7206 ( 
.A(n_6137),
.Y(n_7206)
);

AND2x4_ASAP7_75t_L g7207 ( 
.A(n_6196),
.B(n_6057),
.Y(n_7207)
);

INVx1_ASAP7_75t_L g7208 ( 
.A(n_6139),
.Y(n_7208)
);

INVx2_ASAP7_75t_L g7209 ( 
.A(n_6657),
.Y(n_7209)
);

INVx2_ASAP7_75t_L g7210 ( 
.A(n_6657),
.Y(n_7210)
);

OAI21x1_ASAP7_75t_L g7211 ( 
.A1(n_6915),
.A2(n_6074),
.B(n_6055),
.Y(n_7211)
);

NOR3xp33_ASAP7_75t_SL g7212 ( 
.A(n_6500),
.B(n_4706),
.C(n_4682),
.Y(n_7212)
);

OAI21x1_ASAP7_75t_L g7213 ( 
.A1(n_6918),
.A2(n_6088),
.B(n_6074),
.Y(n_7213)
);

INVx1_ASAP7_75t_L g7214 ( 
.A(n_6143),
.Y(n_7214)
);

AO21x2_ASAP7_75t_L g7215 ( 
.A1(n_6918),
.A2(n_5508),
.B(n_5470),
.Y(n_7215)
);

INVx1_ASAP7_75t_L g7216 ( 
.A(n_6143),
.Y(n_7216)
);

INVx1_ASAP7_75t_L g7217 ( 
.A(n_6143),
.Y(n_7217)
);

OAI21x1_ASAP7_75t_L g7218 ( 
.A1(n_6922),
.A2(n_6088),
.B(n_5596),
.Y(n_7218)
);

INVxp67_ASAP7_75t_L g7219 ( 
.A(n_6172),
.Y(n_7219)
);

OA21x2_ASAP7_75t_L g7220 ( 
.A1(n_7046),
.A2(n_5940),
.B(n_5932),
.Y(n_7220)
);

OR2x6_ASAP7_75t_L g7221 ( 
.A(n_6222),
.B(n_5678),
.Y(n_7221)
);

O2A1O1Ixp33_ASAP7_75t_SL g7222 ( 
.A1(n_6249),
.A2(n_5244),
.B(n_5331),
.C(n_5668),
.Y(n_7222)
);

INVx1_ASAP7_75t_L g7223 ( 
.A(n_6168),
.Y(n_7223)
);

OAI21x1_ASAP7_75t_L g7224 ( 
.A1(n_6922),
.A2(n_5596),
.B(n_6124),
.Y(n_7224)
);

OR2x2_ASAP7_75t_L g7225 ( 
.A(n_6340),
.B(n_5236),
.Y(n_7225)
);

INVx2_ASAP7_75t_L g7226 ( 
.A(n_6136),
.Y(n_7226)
);

A2O1A1Ixp33_ASAP7_75t_L g7227 ( 
.A1(n_6249),
.A2(n_5260),
.B(n_5184),
.C(n_5177),
.Y(n_7227)
);

INVx1_ASAP7_75t_L g7228 ( 
.A(n_6168),
.Y(n_7228)
);

CKINVDCx5p33_ASAP7_75t_R g7229 ( 
.A(n_6601),
.Y(n_7229)
);

O2A1O1Ixp33_ASAP7_75t_SL g7230 ( 
.A1(n_6146),
.A2(n_5679),
.B(n_5708),
.C(n_5870),
.Y(n_7230)
);

BUFx3_ASAP7_75t_L g7231 ( 
.A(n_6636),
.Y(n_7231)
);

OAI21x1_ASAP7_75t_L g7232 ( 
.A1(n_6281),
.A2(n_6513),
.B(n_6505),
.Y(n_7232)
);

AND2x4_ASAP7_75t_L g7233 ( 
.A(n_6196),
.B(n_6057),
.Y(n_7233)
);

AO21x2_ASAP7_75t_L g7234 ( 
.A1(n_6388),
.A2(n_5535),
.B(n_6044),
.Y(n_7234)
);

OAI21x1_ASAP7_75t_L g7235 ( 
.A1(n_6281),
.A2(n_6124),
.B(n_6086),
.Y(n_7235)
);

INVx1_ASAP7_75t_L g7236 ( 
.A(n_6168),
.Y(n_7236)
);

INVx1_ASAP7_75t_L g7237 ( 
.A(n_6174),
.Y(n_7237)
);

OAI21x1_ASAP7_75t_L g7238 ( 
.A1(n_6505),
.A2(n_6086),
.B(n_5595),
.Y(n_7238)
);

INVx2_ASAP7_75t_L g7239 ( 
.A(n_6136),
.Y(n_7239)
);

OAI21x1_ASAP7_75t_L g7240 ( 
.A1(n_6513),
.A2(n_5595),
.B(n_5277),
.Y(n_7240)
);

OAI21x1_ASAP7_75t_L g7241 ( 
.A1(n_6545),
.A2(n_5277),
.B(n_5265),
.Y(n_7241)
);

CKINVDCx6p67_ASAP7_75t_R g7242 ( 
.A(n_6237),
.Y(n_7242)
);

INVxp67_ASAP7_75t_L g7243 ( 
.A(n_6172),
.Y(n_7243)
);

NAND2xp5_ASAP7_75t_L g7244 ( 
.A(n_7042),
.B(n_6435),
.Y(n_7244)
);

CKINVDCx11_ASAP7_75t_R g7245 ( 
.A(n_6774),
.Y(n_7245)
);

BUFx3_ASAP7_75t_L g7246 ( 
.A(n_6636),
.Y(n_7246)
);

OA21x2_ASAP7_75t_L g7247 ( 
.A1(n_7046),
.A2(n_6093),
.B(n_5193),
.Y(n_7247)
);

OAI21x1_ASAP7_75t_L g7248 ( 
.A1(n_6545),
.A2(n_5265),
.B(n_5561),
.Y(n_7248)
);

OAI21x1_ASAP7_75t_L g7249 ( 
.A1(n_6555),
.A2(n_5569),
.B(n_5561),
.Y(n_7249)
);

INVx1_ASAP7_75t_L g7250 ( 
.A(n_6174),
.Y(n_7250)
);

INVx1_ASAP7_75t_SL g7251 ( 
.A(n_6152),
.Y(n_7251)
);

INVx1_ASAP7_75t_L g7252 ( 
.A(n_6174),
.Y(n_7252)
);

INVx1_ASAP7_75t_L g7253 ( 
.A(n_6186),
.Y(n_7253)
);

OAI21x1_ASAP7_75t_L g7254 ( 
.A1(n_6555),
.A2(n_5574),
.B(n_5569),
.Y(n_7254)
);

OAI21x1_ASAP7_75t_L g7255 ( 
.A1(n_6559),
.A2(n_5585),
.B(n_5574),
.Y(n_7255)
);

AOI22xp5_ASAP7_75t_L g7256 ( 
.A1(n_6203),
.A2(n_5453),
.B1(n_5371),
.B2(n_5554),
.Y(n_7256)
);

OR2x4_ASAP7_75t_L g7257 ( 
.A(n_6393),
.B(n_6865),
.Y(n_7257)
);

INVx1_ASAP7_75t_L g7258 ( 
.A(n_6186),
.Y(n_7258)
);

OAI21xp5_ASAP7_75t_L g7259 ( 
.A1(n_7078),
.A2(n_5271),
.B(n_5184),
.Y(n_7259)
);

INVx1_ASAP7_75t_L g7260 ( 
.A(n_6186),
.Y(n_7260)
);

OAI21x1_ASAP7_75t_L g7261 ( 
.A1(n_6559),
.A2(n_5590),
.B(n_5585),
.Y(n_7261)
);

CKINVDCx5p33_ASAP7_75t_R g7262 ( 
.A(n_6485),
.Y(n_7262)
);

INVx2_ASAP7_75t_L g7263 ( 
.A(n_6136),
.Y(n_7263)
);

BUFx3_ASAP7_75t_L g7264 ( 
.A(n_6705),
.Y(n_7264)
);

INVx8_ASAP7_75t_L g7265 ( 
.A(n_6237),
.Y(n_7265)
);

AOI21x1_ASAP7_75t_L g7266 ( 
.A1(n_6484),
.A2(n_6044),
.B(n_6010),
.Y(n_7266)
);

INVx2_ASAP7_75t_L g7267 ( 
.A(n_6136),
.Y(n_7267)
);

OAI31xp33_ASAP7_75t_L g7268 ( 
.A1(n_6693),
.A2(n_5414),
.A3(n_5554),
.B(n_5337),
.Y(n_7268)
);

AOI21xp5_ASAP7_75t_L g7269 ( 
.A1(n_6552),
.A2(n_6034),
.B(n_5969),
.Y(n_7269)
);

OAI21x1_ASAP7_75t_SL g7270 ( 
.A1(n_6995),
.A2(n_5177),
.B(n_5993),
.Y(n_7270)
);

AND2x6_ASAP7_75t_L g7271 ( 
.A(n_6706),
.B(n_4942),
.Y(n_7271)
);

OAI21x1_ASAP7_75t_L g7272 ( 
.A1(n_6576),
.A2(n_5590),
.B(n_5474),
.Y(n_7272)
);

OAI22xp5_ASAP7_75t_L g7273 ( 
.A1(n_6572),
.A2(n_5708),
.B1(n_5253),
.B2(n_5290),
.Y(n_7273)
);

INVx1_ASAP7_75t_L g7274 ( 
.A(n_6198),
.Y(n_7274)
);

OAI21x1_ASAP7_75t_L g7275 ( 
.A1(n_6576),
.A2(n_5162),
.B(n_6093),
.Y(n_7275)
);

INVx4_ASAP7_75t_L g7276 ( 
.A(n_6237),
.Y(n_7276)
);

BUFx2_ASAP7_75t_L g7277 ( 
.A(n_6492),
.Y(n_7277)
);

INVx1_ASAP7_75t_L g7278 ( 
.A(n_6198),
.Y(n_7278)
);

OA21x2_ASAP7_75t_L g7279 ( 
.A1(n_7046),
.A2(n_5193),
.B(n_5176),
.Y(n_7279)
);

NAND2xp5_ASAP7_75t_L g7280 ( 
.A(n_6435),
.B(n_5846),
.Y(n_7280)
);

NAND2x1p5_ASAP7_75t_L g7281 ( 
.A(n_6462),
.B(n_5150),
.Y(n_7281)
);

AOI22xp33_ASAP7_75t_L g7282 ( 
.A1(n_6362),
.A2(n_5337),
.B1(n_5440),
.B2(n_5433),
.Y(n_7282)
);

BUFx12f_ASAP7_75t_L g7283 ( 
.A(n_6339),
.Y(n_7283)
);

AND2x4_ASAP7_75t_L g7284 ( 
.A(n_6196),
.B(n_6218),
.Y(n_7284)
);

AOI22xp33_ASAP7_75t_L g7285 ( 
.A1(n_6362),
.A2(n_5433),
.B1(n_5440),
.B2(n_5537),
.Y(n_7285)
);

OAI21xp5_ASAP7_75t_L g7286 ( 
.A1(n_7078),
.A2(n_5271),
.B(n_5534),
.Y(n_7286)
);

AOI22xp33_ASAP7_75t_L g7287 ( 
.A1(n_6262),
.A2(n_5537),
.B1(n_5556),
.B2(n_5566),
.Y(n_7287)
);

AOI21xp5_ASAP7_75t_L g7288 ( 
.A1(n_6552),
.A2(n_6017),
.B(n_5390),
.Y(n_7288)
);

OAI21x1_ASAP7_75t_L g7289 ( 
.A1(n_6577),
.A2(n_6662),
.B(n_6581),
.Y(n_7289)
);

INVx1_ASAP7_75t_L g7290 ( 
.A(n_6198),
.Y(n_7290)
);

AND2x2_ASAP7_75t_L g7291 ( 
.A(n_6145),
.B(n_5752),
.Y(n_7291)
);

AOI221xp5_ASAP7_75t_L g7292 ( 
.A1(n_6262),
.A2(n_6076),
.B1(n_6091),
.B2(n_6081),
.C(n_6079),
.Y(n_7292)
);

OAI21x1_ASAP7_75t_L g7293 ( 
.A1(n_6577),
.A2(n_6662),
.B(n_6581),
.Y(n_7293)
);

OAI21x1_ASAP7_75t_L g7294 ( 
.A1(n_6671),
.A2(n_5162),
.B(n_5416),
.Y(n_7294)
);

INVx1_ASAP7_75t_L g7295 ( 
.A(n_6204),
.Y(n_7295)
);

OAI21x1_ASAP7_75t_L g7296 ( 
.A1(n_6671),
.A2(n_5416),
.B(n_5284),
.Y(n_7296)
);

NOR2xp33_ASAP7_75t_L g7297 ( 
.A(n_6393),
.B(n_5253),
.Y(n_7297)
);

BUFx2_ASAP7_75t_L g7298 ( 
.A(n_6492),
.Y(n_7298)
);

INVx2_ASAP7_75t_SL g7299 ( 
.A(n_6874),
.Y(n_7299)
);

OAI21xp5_ASAP7_75t_L g7300 ( 
.A1(n_6975),
.A2(n_5489),
.B(n_5871),
.Y(n_7300)
);

AOI22xp33_ASAP7_75t_L g7301 ( 
.A1(n_6431),
.A2(n_5556),
.B1(n_5566),
.B2(n_5481),
.Y(n_7301)
);

OAI22xp33_ASAP7_75t_L g7302 ( 
.A1(n_6800),
.A2(n_5453),
.B1(n_5158),
.B2(n_5500),
.Y(n_7302)
);

OAI21x1_ASAP7_75t_L g7303 ( 
.A1(n_6685),
.A2(n_5284),
.B(n_5250),
.Y(n_7303)
);

INVx1_ASAP7_75t_L g7304 ( 
.A(n_6204),
.Y(n_7304)
);

OAI21x1_ASAP7_75t_L g7305 ( 
.A1(n_6685),
.A2(n_5284),
.B(n_5431),
.Y(n_7305)
);

INVx1_ASAP7_75t_L g7306 ( 
.A(n_6204),
.Y(n_7306)
);

INVx1_ASAP7_75t_SL g7307 ( 
.A(n_6157),
.Y(n_7307)
);

OR2x2_ASAP7_75t_L g7308 ( 
.A(n_6340),
.B(n_6370),
.Y(n_7308)
);

AO21x2_ASAP7_75t_L g7309 ( 
.A1(n_6388),
.A2(n_6801),
.B(n_6711),
.Y(n_7309)
);

NAND2xp5_ASAP7_75t_L g7310 ( 
.A(n_7025),
.B(n_5848),
.Y(n_7310)
);

OAI21x1_ASAP7_75t_L g7311 ( 
.A1(n_6689),
.A2(n_5284),
.B(n_5431),
.Y(n_7311)
);

OA21x2_ASAP7_75t_L g7312 ( 
.A1(n_6664),
.A2(n_5390),
.B(n_5176),
.Y(n_7312)
);

AND2x4_ASAP7_75t_L g7313 ( 
.A(n_6218),
.B(n_6057),
.Y(n_7313)
);

CKINVDCx20_ASAP7_75t_R g7314 ( 
.A(n_6774),
.Y(n_7314)
);

NAND2xp5_ASAP7_75t_L g7315 ( 
.A(n_7025),
.B(n_5848),
.Y(n_7315)
);

INVx2_ASAP7_75t_SL g7316 ( 
.A(n_6874),
.Y(n_7316)
);

BUFx2_ASAP7_75t_L g7317 ( 
.A(n_6492),
.Y(n_7317)
);

INVx2_ASAP7_75t_L g7318 ( 
.A(n_6138),
.Y(n_7318)
);

OAI21x1_ASAP7_75t_L g7319 ( 
.A1(n_6689),
.A2(n_6798),
.B(n_6745),
.Y(n_7319)
);

OAI21xp5_ASAP7_75t_L g7320 ( 
.A1(n_6975),
.A2(n_5489),
.B(n_5308),
.Y(n_7320)
);

OAI21x1_ASAP7_75t_L g7321 ( 
.A1(n_6745),
.A2(n_5284),
.B(n_5858),
.Y(n_7321)
);

HB1xp67_ASAP7_75t_L g7322 ( 
.A(n_6924),
.Y(n_7322)
);

CKINVDCx5p33_ASAP7_75t_R g7323 ( 
.A(n_6485),
.Y(n_7323)
);

HB1xp67_ASAP7_75t_L g7324 ( 
.A(n_6924),
.Y(n_7324)
);

AOI21xp5_ASAP7_75t_L g7325 ( 
.A1(n_6664),
.A2(n_5319),
.B(n_5301),
.Y(n_7325)
);

INVx2_ASAP7_75t_L g7326 ( 
.A(n_6138),
.Y(n_7326)
);

INVx1_ASAP7_75t_L g7327 ( 
.A(n_6224),
.Y(n_7327)
);

CKINVDCx6p67_ASAP7_75t_R g7328 ( 
.A(n_6339),
.Y(n_7328)
);

INVx2_ASAP7_75t_L g7329 ( 
.A(n_6138),
.Y(n_7329)
);

OAI21xp5_ASAP7_75t_L g7330 ( 
.A1(n_6264),
.A2(n_5491),
.B(n_5452),
.Y(n_7330)
);

INVx2_ASAP7_75t_SL g7331 ( 
.A(n_6874),
.Y(n_7331)
);

A2O1A1Ixp33_ASAP7_75t_L g7332 ( 
.A1(n_6379),
.A2(n_5408),
.B(n_5449),
.C(n_5605),
.Y(n_7332)
);

OAI21x1_ASAP7_75t_L g7333 ( 
.A1(n_6798),
.A2(n_6804),
.B(n_6802),
.Y(n_7333)
);

INVx3_ASAP7_75t_L g7334 ( 
.A(n_6218),
.Y(n_7334)
);

AND2x2_ASAP7_75t_L g7335 ( 
.A(n_6180),
.B(n_6039),
.Y(n_7335)
);

INVx1_ASAP7_75t_L g7336 ( 
.A(n_6224),
.Y(n_7336)
);

AOI21xp5_ASAP7_75t_L g7337 ( 
.A1(n_6410),
.A2(n_5319),
.B(n_5273),
.Y(n_7337)
);

AO21x2_ASAP7_75t_L g7338 ( 
.A1(n_6711),
.A2(n_5995),
.B(n_5597),
.Y(n_7338)
);

BUFx12f_ASAP7_75t_L g7339 ( 
.A(n_6339),
.Y(n_7339)
);

INVx2_ASAP7_75t_L g7340 ( 
.A(n_6138),
.Y(n_7340)
);

NAND2xp33_ASAP7_75t_L g7341 ( 
.A(n_7007),
.B(n_6894),
.Y(n_7341)
);

OA21x2_ASAP7_75t_L g7342 ( 
.A1(n_6282),
.A2(n_6035),
.B(n_5364),
.Y(n_7342)
);

OAI21x1_ASAP7_75t_L g7343 ( 
.A1(n_6802),
.A2(n_5858),
.B(n_5411),
.Y(n_7343)
);

OAI21xp5_ASAP7_75t_L g7344 ( 
.A1(n_6264),
.A2(n_5452),
.B(n_5510),
.Y(n_7344)
);

BUFx2_ASAP7_75t_L g7345 ( 
.A(n_6501),
.Y(n_7345)
);

BUFx2_ASAP7_75t_SL g7346 ( 
.A(n_7054),
.Y(n_7346)
);

BUFx2_ASAP7_75t_L g7347 ( 
.A(n_6501),
.Y(n_7347)
);

INVx1_ASAP7_75t_L g7348 ( 
.A(n_6224),
.Y(n_7348)
);

NAND2xp5_ASAP7_75t_L g7349 ( 
.A(n_7061),
.B(n_5883),
.Y(n_7349)
);

BUFx2_ASAP7_75t_L g7350 ( 
.A(n_6501),
.Y(n_7350)
);

HB1xp67_ASAP7_75t_L g7351 ( 
.A(n_6957),
.Y(n_7351)
);

OAI21xp5_ASAP7_75t_L g7352 ( 
.A1(n_6303),
.A2(n_5515),
.B(n_5883),
.Y(n_7352)
);

OA21x2_ASAP7_75t_L g7353 ( 
.A1(n_6282),
.A2(n_6035),
.B(n_5364),
.Y(n_7353)
);

OAI21x1_ASAP7_75t_L g7354 ( 
.A1(n_6804),
.A2(n_5411),
.B(n_5373),
.Y(n_7354)
);

AO21x2_ASAP7_75t_L g7355 ( 
.A1(n_6801),
.A2(n_5995),
.B(n_5597),
.Y(n_7355)
);

INVx1_ASAP7_75t_L g7356 ( 
.A(n_6226),
.Y(n_7356)
);

INVx1_ASAP7_75t_L g7357 ( 
.A(n_6226),
.Y(n_7357)
);

OA21x2_ASAP7_75t_L g7358 ( 
.A1(n_6827),
.A2(n_5373),
.B(n_5334),
.Y(n_7358)
);

OA21x2_ASAP7_75t_L g7359 ( 
.A1(n_6827),
.A2(n_5374),
.B(n_5334),
.Y(n_7359)
);

NAND2xp5_ASAP7_75t_L g7360 ( 
.A(n_7061),
.B(n_5984),
.Y(n_7360)
);

INVx1_ASAP7_75t_L g7361 ( 
.A(n_6226),
.Y(n_7361)
);

INVx3_ASAP7_75t_L g7362 ( 
.A(n_6218),
.Y(n_7362)
);

CKINVDCx5p33_ASAP7_75t_R g7363 ( 
.A(n_6898),
.Y(n_7363)
);

INVx1_ASAP7_75t_L g7364 ( 
.A(n_6242),
.Y(n_7364)
);

BUFx6f_ASAP7_75t_L g7365 ( 
.A(n_6137),
.Y(n_7365)
);

NAND2xp5_ASAP7_75t_SL g7366 ( 
.A(n_6923),
.B(n_5993),
.Y(n_7366)
);

HB1xp67_ASAP7_75t_L g7367 ( 
.A(n_6957),
.Y(n_7367)
);

INVx1_ASAP7_75t_SL g7368 ( 
.A(n_6157),
.Y(n_7368)
);

BUFx6f_ASAP7_75t_L g7369 ( 
.A(n_6137),
.Y(n_7369)
);

OAI21xp33_ASAP7_75t_SL g7370 ( 
.A1(n_6874),
.A2(n_6109),
.B(n_6070),
.Y(n_7370)
);

AND2x2_ASAP7_75t_L g7371 ( 
.A(n_6180),
.B(n_6070),
.Y(n_7371)
);

INVx2_ASAP7_75t_L g7372 ( 
.A(n_6144),
.Y(n_7372)
);

INVx2_ASAP7_75t_L g7373 ( 
.A(n_6144),
.Y(n_7373)
);

AND2x2_ASAP7_75t_L g7374 ( 
.A(n_6180),
.B(n_6070),
.Y(n_7374)
);

CKINVDCx20_ASAP7_75t_R g7375 ( 
.A(n_6167),
.Y(n_7375)
);

AOI21xp5_ASAP7_75t_L g7376 ( 
.A1(n_6410),
.A2(n_5319),
.B(n_5273),
.Y(n_7376)
);

AO21x2_ASAP7_75t_L g7377 ( 
.A1(n_6633),
.A2(n_5995),
.B(n_5605),
.Y(n_7377)
);

BUFx2_ASAP7_75t_R g7378 ( 
.A(n_6259),
.Y(n_7378)
);

HB1xp67_ASAP7_75t_L g7379 ( 
.A(n_6986),
.Y(n_7379)
);

AOI22xp33_ASAP7_75t_L g7380 ( 
.A1(n_6431),
.A2(n_5481),
.B1(n_5414),
.B2(n_5445),
.Y(n_7380)
);

BUFx3_ASAP7_75t_L g7381 ( 
.A(n_6705),
.Y(n_7381)
);

AND2x2_ASAP7_75t_L g7382 ( 
.A(n_6201),
.B(n_6109),
.Y(n_7382)
);

BUFx3_ASAP7_75t_L g7383 ( 
.A(n_6705),
.Y(n_7383)
);

OAI21x1_ASAP7_75t_L g7384 ( 
.A1(n_6842),
.A2(n_5395),
.B(n_5374),
.Y(n_7384)
);

NAND2x1p5_ASAP7_75t_L g7385 ( 
.A(n_6462),
.B(n_5150),
.Y(n_7385)
);

INVx2_ASAP7_75t_L g7386 ( 
.A(n_6144),
.Y(n_7386)
);

BUFx3_ASAP7_75t_L g7387 ( 
.A(n_6339),
.Y(n_7387)
);

OAI21x1_ASAP7_75t_L g7388 ( 
.A1(n_6842),
.A2(n_5407),
.B(n_5395),
.Y(n_7388)
);

INVx1_ASAP7_75t_L g7389 ( 
.A(n_6242),
.Y(n_7389)
);

INVx2_ASAP7_75t_L g7390 ( 
.A(n_6144),
.Y(n_7390)
);

OAI21x1_ASAP7_75t_L g7391 ( 
.A1(n_6432),
.A2(n_5410),
.B(n_5407),
.Y(n_7391)
);

AOI21xp5_ASAP7_75t_L g7392 ( 
.A1(n_6886),
.A2(n_5319),
.B(n_5280),
.Y(n_7392)
);

OR2x2_ASAP7_75t_L g7393 ( 
.A(n_6340),
.B(n_5236),
.Y(n_7393)
);

OAI21xp5_ASAP7_75t_L g7394 ( 
.A1(n_6303),
.A2(n_6366),
.B(n_6800),
.Y(n_7394)
);

A2O1A1Ixp33_ASAP7_75t_L g7395 ( 
.A1(n_6997),
.A2(n_5449),
.B(n_5495),
.C(n_5359),
.Y(n_7395)
);

INVx2_ASAP7_75t_L g7396 ( 
.A(n_6150),
.Y(n_7396)
);

OAI21x1_ASAP7_75t_L g7397 ( 
.A1(n_6432),
.A2(n_6535),
.B(n_6258),
.Y(n_7397)
);

AOI22xp33_ASAP7_75t_SL g7398 ( 
.A1(n_6923),
.A2(n_5158),
.B1(n_5313),
.B2(n_5150),
.Y(n_7398)
);

O2A1O1Ixp5_ASAP7_75t_L g7399 ( 
.A1(n_6855),
.A2(n_5175),
.B(n_5406),
.C(n_5376),
.Y(n_7399)
);

HB1xp67_ASAP7_75t_L g7400 ( 
.A(n_6986),
.Y(n_7400)
);

AOI22xp33_ASAP7_75t_L g7401 ( 
.A1(n_6403),
.A2(n_5445),
.B1(n_5312),
.B2(n_5995),
.Y(n_7401)
);

NAND2x1p5_ASAP7_75t_L g7402 ( 
.A(n_6462),
.B(n_5150),
.Y(n_7402)
);

OAI22xp5_ASAP7_75t_L g7403 ( 
.A1(n_6572),
.A2(n_5275),
.B1(n_5290),
.B2(n_5158),
.Y(n_7403)
);

BUFx3_ASAP7_75t_L g7404 ( 
.A(n_6383),
.Y(n_7404)
);

NAND2xp5_ASAP7_75t_L g7405 ( 
.A(n_6623),
.B(n_5984),
.Y(n_7405)
);

OAI221xp5_ASAP7_75t_L g7406 ( 
.A1(n_6997),
.A2(n_5393),
.B1(n_5507),
.B2(n_5495),
.C(n_5359),
.Y(n_7406)
);

AO32x2_ASAP7_75t_L g7407 ( 
.A1(n_7126),
.A2(n_6071),
.A3(n_5829),
.B1(n_5824),
.B2(n_6076),
.Y(n_7407)
);

BUFx2_ASAP7_75t_L g7408 ( 
.A(n_6241),
.Y(n_7408)
);

OAI21x1_ASAP7_75t_L g7409 ( 
.A1(n_6535),
.A2(n_6258),
.B(n_6206),
.Y(n_7409)
);

AOI22xp33_ASAP7_75t_SL g7410 ( 
.A1(n_6923),
.A2(n_6370),
.B1(n_6382),
.B2(n_6374),
.Y(n_7410)
);

NAND2x1p5_ASAP7_75t_L g7411 ( 
.A(n_6691),
.B(n_5150),
.Y(n_7411)
);

OA21x2_ASAP7_75t_L g7412 ( 
.A1(n_6199),
.A2(n_5437),
.B(n_5410),
.Y(n_7412)
);

AND2x2_ASAP7_75t_L g7413 ( 
.A(n_6201),
.B(n_6109),
.Y(n_7413)
);

NAND2xp5_ASAP7_75t_L g7414 ( 
.A(n_6623),
.B(n_6079),
.Y(n_7414)
);

INVxp67_ASAP7_75t_SL g7415 ( 
.A(n_6331),
.Y(n_7415)
);

INVx1_ASAP7_75t_L g7416 ( 
.A(n_6242),
.Y(n_7416)
);

AO21x2_ASAP7_75t_L g7417 ( 
.A1(n_6633),
.A2(n_5967),
.B(n_5467),
.Y(n_7417)
);

OAI21x1_ASAP7_75t_L g7418 ( 
.A1(n_6199),
.A2(n_5467),
.B(n_5437),
.Y(n_7418)
);

OAI21x1_ASAP7_75t_L g7419 ( 
.A1(n_6206),
.A2(n_5482),
.B(n_5664),
.Y(n_7419)
);

CKINVDCx5p33_ASAP7_75t_R g7420 ( 
.A(n_6898),
.Y(n_7420)
);

INVx1_ASAP7_75t_L g7421 ( 
.A(n_6246),
.Y(n_7421)
);

INVx4_ASAP7_75t_L g7422 ( 
.A(n_6383),
.Y(n_7422)
);

OAI21x1_ASAP7_75t_L g7423 ( 
.A1(n_6207),
.A2(n_5482),
.B(n_5664),
.Y(n_7423)
);

OAI21x1_ASAP7_75t_L g7424 ( 
.A1(n_6207),
.A2(n_5666),
.B(n_5664),
.Y(n_7424)
);

OAI21x1_ASAP7_75t_L g7425 ( 
.A1(n_6233),
.A2(n_5666),
.B(n_5664),
.Y(n_7425)
);

INVx2_ASAP7_75t_L g7426 ( 
.A(n_6150),
.Y(n_7426)
);

INVx1_ASAP7_75t_L g7427 ( 
.A(n_6246),
.Y(n_7427)
);

OAI21x1_ASAP7_75t_L g7428 ( 
.A1(n_6233),
.A2(n_5869),
.B(n_5666),
.Y(n_7428)
);

INVx3_ASAP7_75t_L g7429 ( 
.A(n_6241),
.Y(n_7429)
);

A2O1A1Ixp33_ASAP7_75t_L g7430 ( 
.A1(n_6366),
.A2(n_5577),
.B(n_5572),
.C(n_6004),
.Y(n_7430)
);

INVx1_ASAP7_75t_SL g7431 ( 
.A(n_6181),
.Y(n_7431)
);

INVx2_ASAP7_75t_L g7432 ( 
.A(n_6150),
.Y(n_7432)
);

BUFx3_ASAP7_75t_L g7433 ( 
.A(n_6383),
.Y(n_7433)
);

INVx1_ASAP7_75t_L g7434 ( 
.A(n_6246),
.Y(n_7434)
);

HB1xp67_ASAP7_75t_L g7435 ( 
.A(n_6858),
.Y(n_7435)
);

OAI21x1_ASAP7_75t_SL g7436 ( 
.A1(n_6355),
.A2(n_6849),
.B(n_6794),
.Y(n_7436)
);

OAI22xp5_ASAP7_75t_L g7437 ( 
.A1(n_6572),
.A2(n_5275),
.B1(n_5956),
.B2(n_5936),
.Y(n_7437)
);

NOR2xp67_ASAP7_75t_L g7438 ( 
.A(n_6195),
.B(n_5150),
.Y(n_7438)
);

NOR2xp67_ASAP7_75t_L g7439 ( 
.A(n_6195),
.B(n_5313),
.Y(n_7439)
);

O2A1O1Ixp33_ASAP7_75t_L g7440 ( 
.A1(n_6331),
.A2(n_5406),
.B(n_5376),
.C(n_5475),
.Y(n_7440)
);

OAI21x1_ASAP7_75t_SL g7441 ( 
.A1(n_6355),
.A2(n_5429),
.B(n_5353),
.Y(n_7441)
);

NOR2xp67_ASAP7_75t_L g7442 ( 
.A(n_6195),
.B(n_5313),
.Y(n_7442)
);

OA21x2_ASAP7_75t_L g7443 ( 
.A1(n_6296),
.A2(n_5967),
.B(n_5280),
.Y(n_7443)
);

AOI21xp5_ASAP7_75t_L g7444 ( 
.A1(n_6953),
.A2(n_5319),
.B(n_5310),
.Y(n_7444)
);

AND2x4_ASAP7_75t_L g7445 ( 
.A(n_6241),
.B(n_6057),
.Y(n_7445)
);

INVx1_ASAP7_75t_L g7446 ( 
.A(n_6270),
.Y(n_7446)
);

INVx2_ASAP7_75t_L g7447 ( 
.A(n_6150),
.Y(n_7447)
);

OAI21x1_ASAP7_75t_L g7448 ( 
.A1(n_6243),
.A2(n_5869),
.B(n_5666),
.Y(n_7448)
);

INVx1_ASAP7_75t_L g7449 ( 
.A(n_6270),
.Y(n_7449)
);

NAND2xp33_ASAP7_75t_L g7450 ( 
.A(n_7007),
.B(n_5771),
.Y(n_7450)
);

A2O1A1Ixp33_ASAP7_75t_L g7451 ( 
.A1(n_6326),
.A2(n_5577),
.B(n_5572),
.C(n_6014),
.Y(n_7451)
);

BUFx2_ASAP7_75t_L g7452 ( 
.A(n_6241),
.Y(n_7452)
);

CKINVDCx20_ASAP7_75t_R g7453 ( 
.A(n_6167),
.Y(n_7453)
);

AND2x4_ASAP7_75t_L g7454 ( 
.A(n_6269),
.B(n_6075),
.Y(n_7454)
);

INVx1_ASAP7_75t_L g7455 ( 
.A(n_6270),
.Y(n_7455)
);

OAI21x1_ASAP7_75t_L g7456 ( 
.A1(n_6243),
.A2(n_5905),
.B(n_5869),
.Y(n_7456)
);

OAI21x1_ASAP7_75t_L g7457 ( 
.A1(n_6650),
.A2(n_6290),
.B(n_6296),
.Y(n_7457)
);

AO21x2_ASAP7_75t_L g7458 ( 
.A1(n_6290),
.A2(n_5603),
.B(n_5564),
.Y(n_7458)
);

OAI21xp5_ASAP7_75t_L g7459 ( 
.A1(n_7057),
.A2(n_5475),
.B(n_5458),
.Y(n_7459)
);

OA21x2_ASAP7_75t_L g7460 ( 
.A1(n_7065),
.A2(n_5310),
.B(n_5272),
.Y(n_7460)
);

AOI21xp5_ASAP7_75t_L g7461 ( 
.A1(n_6953),
.A2(n_5319),
.B(n_5272),
.Y(n_7461)
);

OAI21x1_ASAP7_75t_L g7462 ( 
.A1(n_6650),
.A2(n_5905),
.B(n_5869),
.Y(n_7462)
);

NOR2xp33_ASAP7_75t_L g7463 ( 
.A(n_7086),
.B(n_6560),
.Y(n_7463)
);

OAI21x1_ASAP7_75t_SL g7464 ( 
.A1(n_6355),
.A2(n_5429),
.B(n_5353),
.Y(n_7464)
);

OAI21x1_ASAP7_75t_L g7465 ( 
.A1(n_6650),
.A2(n_5905),
.B(n_5315),
.Y(n_7465)
);

BUFx2_ASAP7_75t_L g7466 ( 
.A(n_6269),
.Y(n_7466)
);

OAI21x1_ASAP7_75t_L g7467 ( 
.A1(n_6892),
.A2(n_5905),
.B(n_5601),
.Y(n_7467)
);

INVx1_ASAP7_75t_L g7468 ( 
.A(n_6274),
.Y(n_7468)
);

BUFx2_ASAP7_75t_L g7469 ( 
.A(n_6269),
.Y(n_7469)
);

AO21x2_ASAP7_75t_L g7470 ( 
.A1(n_6892),
.A2(n_5603),
.B(n_5564),
.Y(n_7470)
);

NOR2xp33_ASAP7_75t_L g7471 ( 
.A(n_7086),
.B(n_6560),
.Y(n_7471)
);

OAI21x1_ASAP7_75t_L g7472 ( 
.A1(n_6458),
.A2(n_6311),
.B(n_6591),
.Y(n_7472)
);

OAI21x1_ASAP7_75t_L g7473 ( 
.A1(n_6458),
.A2(n_5601),
.B(n_5283),
.Y(n_7473)
);

OAI21x1_ASAP7_75t_L g7474 ( 
.A1(n_6311),
.A2(n_5601),
.B(n_5283),
.Y(n_7474)
);

INVx2_ASAP7_75t_L g7475 ( 
.A(n_6163),
.Y(n_7475)
);

CKINVDCx12_ASAP7_75t_R g7476 ( 
.A(n_6277),
.Y(n_7476)
);

NAND2xp5_ASAP7_75t_SL g7477 ( 
.A(n_6923),
.B(n_5575),
.Y(n_7477)
);

BUFx6f_ASAP7_75t_L g7478 ( 
.A(n_6137),
.Y(n_7478)
);

NOR2xp33_ASAP7_75t_L g7479 ( 
.A(n_6263),
.B(n_5951),
.Y(n_7479)
);

OAI21xp5_ASAP7_75t_L g7480 ( 
.A1(n_6855),
.A2(n_5458),
.B(n_5560),
.Y(n_7480)
);

INVx1_ASAP7_75t_L g7481 ( 
.A(n_6274),
.Y(n_7481)
);

INVx1_ASAP7_75t_L g7482 ( 
.A(n_6274),
.Y(n_7482)
);

OAI21x1_ASAP7_75t_L g7483 ( 
.A1(n_6311),
.A2(n_5405),
.B(n_5377),
.Y(n_7483)
);

OAI21x1_ASAP7_75t_L g7484 ( 
.A1(n_6311),
.A2(n_5405),
.B(n_5377),
.Y(n_7484)
);

OAI21x1_ASAP7_75t_L g7485 ( 
.A1(n_6591),
.A2(n_5324),
.B(n_5545),
.Y(n_7485)
);

NOR2xp33_ASAP7_75t_L g7486 ( 
.A(n_6263),
.B(n_5951),
.Y(n_7486)
);

OAI21x1_ASAP7_75t_L g7487 ( 
.A1(n_6591),
.A2(n_5324),
.B(n_5545),
.Y(n_7487)
);

INVx2_ASAP7_75t_L g7488 ( 
.A(n_6163),
.Y(n_7488)
);

BUFx3_ASAP7_75t_L g7489 ( 
.A(n_6383),
.Y(n_7489)
);

INVx1_ASAP7_75t_L g7490 ( 
.A(n_6275),
.Y(n_7490)
);

AND2x2_ASAP7_75t_L g7491 ( 
.A(n_6201),
.B(n_6211),
.Y(n_7491)
);

BUFx2_ASAP7_75t_L g7492 ( 
.A(n_6269),
.Y(n_7492)
);

BUFx6f_ASAP7_75t_L g7493 ( 
.A(n_6137),
.Y(n_7493)
);

NAND2xp5_ASAP7_75t_L g7494 ( 
.A(n_6625),
.B(n_6081),
.Y(n_7494)
);

OAI21x1_ASAP7_75t_L g7495 ( 
.A1(n_6591),
.A2(n_5916),
.B(n_5560),
.Y(n_7495)
);

INVx2_ASAP7_75t_L g7496 ( 
.A(n_6163),
.Y(n_7496)
);

OAI21xp5_ASAP7_75t_L g7497 ( 
.A1(n_6305),
.A2(n_5520),
.B(n_5371),
.Y(n_7497)
);

NOR2xp67_ASAP7_75t_L g7498 ( 
.A(n_6195),
.B(n_5313),
.Y(n_7498)
);

INVx1_ASAP7_75t_L g7499 ( 
.A(n_6275),
.Y(n_7499)
);

AOI22xp33_ASAP7_75t_L g7500 ( 
.A1(n_6403),
.A2(n_5312),
.B1(n_5466),
.B2(n_5235),
.Y(n_7500)
);

INVx2_ASAP7_75t_L g7501 ( 
.A(n_6163),
.Y(n_7501)
);

AO31x2_ASAP7_75t_L g7502 ( 
.A1(n_7127),
.A2(n_5606),
.A3(n_6091),
.B(n_6125),
.Y(n_7502)
);

OAI21x1_ASAP7_75t_L g7503 ( 
.A1(n_6699),
.A2(n_5916),
.B(n_5589),
.Y(n_7503)
);

AOI21xp5_ASAP7_75t_L g7504 ( 
.A1(n_6148),
.A2(n_5986),
.B(n_5175),
.Y(n_7504)
);

AO31x2_ASAP7_75t_L g7505 ( 
.A1(n_6238),
.A2(n_5606),
.A3(n_6125),
.B(n_5178),
.Y(n_7505)
);

INVx2_ASAP7_75t_L g7506 ( 
.A(n_6187),
.Y(n_7506)
);

INVx2_ASAP7_75t_L g7507 ( 
.A(n_6187),
.Y(n_7507)
);

AOI21xp5_ASAP7_75t_L g7508 ( 
.A1(n_6148),
.A2(n_5216),
.B(n_5403),
.Y(n_7508)
);

OAI21x1_ASAP7_75t_SL g7509 ( 
.A1(n_6849),
.A2(n_6032),
.B(n_5350),
.Y(n_7509)
);

NAND2x1p5_ASAP7_75t_L g7510 ( 
.A(n_6691),
.B(n_5313),
.Y(n_7510)
);

NAND2xp5_ASAP7_75t_L g7511 ( 
.A(n_6625),
.B(n_6005),
.Y(n_7511)
);

NAND2x1p5_ASAP7_75t_L g7512 ( 
.A(n_6691),
.B(n_5313),
.Y(n_7512)
);

NAND2x1p5_ASAP7_75t_L g7513 ( 
.A(n_6691),
.B(n_5313),
.Y(n_7513)
);

OAI21x1_ASAP7_75t_L g7514 ( 
.A1(n_6699),
.A2(n_5916),
.B(n_5589),
.Y(n_7514)
);

NAND3xp33_ASAP7_75t_L g7515 ( 
.A(n_6306),
.B(n_6104),
.C(n_5422),
.Y(n_7515)
);

OA21x2_ASAP7_75t_L g7516 ( 
.A1(n_7065),
.A2(n_5541),
.B(n_5518),
.Y(n_7516)
);

INVx1_ASAP7_75t_SL g7517 ( 
.A(n_6181),
.Y(n_7517)
);

INVx1_ASAP7_75t_SL g7518 ( 
.A(n_6260),
.Y(n_7518)
);

AND2x4_ASAP7_75t_L g7519 ( 
.A(n_6310),
.B(n_6075),
.Y(n_7519)
);

OAI21x1_ASAP7_75t_L g7520 ( 
.A1(n_6699),
.A2(n_5916),
.B(n_5418),
.Y(n_7520)
);

CKINVDCx5p33_ASAP7_75t_R g7521 ( 
.A(n_7056),
.Y(n_7521)
);

BUFx2_ASAP7_75t_L g7522 ( 
.A(n_6310),
.Y(n_7522)
);

HB1xp67_ASAP7_75t_L g7523 ( 
.A(n_6858),
.Y(n_7523)
);

INVx1_ASAP7_75t_L g7524 ( 
.A(n_6275),
.Y(n_7524)
);

AOI22xp33_ASAP7_75t_L g7525 ( 
.A1(n_6923),
.A2(n_5466),
.B1(n_5235),
.B2(n_5234),
.Y(n_7525)
);

OAI21x1_ASAP7_75t_L g7526 ( 
.A1(n_6531),
.A2(n_5418),
.B(n_5366),
.Y(n_7526)
);

INVx1_ASAP7_75t_L g7527 ( 
.A(n_6291),
.Y(n_7527)
);

INVx1_ASAP7_75t_L g7528 ( 
.A(n_6291),
.Y(n_7528)
);

OA21x2_ASAP7_75t_L g7529 ( 
.A1(n_6844),
.A2(n_6796),
.B(n_6531),
.Y(n_7529)
);

OAI21x1_ASAP7_75t_L g7530 ( 
.A1(n_6531),
.A2(n_5418),
.B(n_5366),
.Y(n_7530)
);

INVx2_ASAP7_75t_SL g7531 ( 
.A(n_6310),
.Y(n_7531)
);

OAI21x1_ASAP7_75t_L g7532 ( 
.A1(n_6484),
.A2(n_5418),
.B(n_5366),
.Y(n_7532)
);

AND2x4_ASAP7_75t_L g7533 ( 
.A(n_6310),
.B(n_6075),
.Y(n_7533)
);

INVx2_ASAP7_75t_L g7534 ( 
.A(n_6187),
.Y(n_7534)
);

AND2x2_ASAP7_75t_L g7535 ( 
.A(n_6211),
.B(n_6220),
.Y(n_7535)
);

AND2x2_ASAP7_75t_L g7536 ( 
.A(n_6211),
.B(n_5285),
.Y(n_7536)
);

INVx1_ASAP7_75t_L g7537 ( 
.A(n_6291),
.Y(n_7537)
);

AOI22xp33_ASAP7_75t_SL g7538 ( 
.A1(n_6923),
.A2(n_5344),
.B1(n_5384),
.B2(n_5313),
.Y(n_7538)
);

OAI21x1_ASAP7_75t_L g7539 ( 
.A1(n_6484),
.A2(n_5448),
.B(n_5366),
.Y(n_7539)
);

AND2x2_ASAP7_75t_L g7540 ( 
.A(n_6220),
.B(n_5285),
.Y(n_7540)
);

BUFx6f_ASAP7_75t_L g7541 ( 
.A(n_6137),
.Y(n_7541)
);

INVx2_ASAP7_75t_L g7542 ( 
.A(n_6187),
.Y(n_7542)
);

BUFx6f_ASAP7_75t_L g7543 ( 
.A(n_6137),
.Y(n_7543)
);

AO21x2_ASAP7_75t_L g7544 ( 
.A1(n_6796),
.A2(n_4939),
.B(n_5516),
.Y(n_7544)
);

AOI22xp33_ASAP7_75t_SL g7545 ( 
.A1(n_6370),
.A2(n_5384),
.B1(n_5671),
.B2(n_5344),
.Y(n_7545)
);

AOI21xp5_ASAP7_75t_L g7546 ( 
.A1(n_6844),
.A2(n_5403),
.B(n_5978),
.Y(n_7546)
);

AND2x2_ASAP7_75t_L g7547 ( 
.A(n_6220),
.B(n_5285),
.Y(n_7547)
);

AND2x4_ASAP7_75t_L g7548 ( 
.A(n_6315),
.B(n_6075),
.Y(n_7548)
);

OA21x2_ASAP7_75t_L g7549 ( 
.A1(n_6517),
.A2(n_5518),
.B(n_5516),
.Y(n_7549)
);

INVx2_ASAP7_75t_L g7550 ( 
.A(n_6212),
.Y(n_7550)
);

HB1xp67_ASAP7_75t_L g7551 ( 
.A(n_6872),
.Y(n_7551)
);

OR2x6_ASAP7_75t_L g7552 ( 
.A(n_6222),
.B(n_5678),
.Y(n_7552)
);

INVx2_ASAP7_75t_L g7553 ( 
.A(n_6212),
.Y(n_7553)
);

OR2x2_ASAP7_75t_L g7554 ( 
.A(n_6374),
.B(n_5236),
.Y(n_7554)
);

BUFx6f_ASAP7_75t_L g7555 ( 
.A(n_6149),
.Y(n_7555)
);

INVx1_ASAP7_75t_L g7556 ( 
.A(n_6298),
.Y(n_7556)
);

INVx2_ASAP7_75t_L g7557 ( 
.A(n_6212),
.Y(n_7557)
);

INVx1_ASAP7_75t_L g7558 ( 
.A(n_6298),
.Y(n_7558)
);

NAND2xp5_ASAP7_75t_L g7559 ( 
.A(n_6708),
.B(n_6005),
.Y(n_7559)
);

AO21x2_ASAP7_75t_L g7560 ( 
.A1(n_6503),
.A2(n_4939),
.B(n_5524),
.Y(n_7560)
);

NAND3xp33_ASAP7_75t_L g7561 ( 
.A(n_6306),
.B(n_6104),
.C(n_5422),
.Y(n_7561)
);

INVxp67_ASAP7_75t_SL g7562 ( 
.A(n_7069),
.Y(n_7562)
);

OAI21x1_ASAP7_75t_SL g7563 ( 
.A1(n_6794),
.A2(n_6032),
.B(n_5350),
.Y(n_7563)
);

AND2x4_ASAP7_75t_L g7564 ( 
.A(n_6356),
.B(n_6075),
.Y(n_7564)
);

INVxp67_ASAP7_75t_L g7565 ( 
.A(n_6194),
.Y(n_7565)
);

INVx2_ASAP7_75t_L g7566 ( 
.A(n_6212),
.Y(n_7566)
);

O2A1O1Ixp33_ASAP7_75t_SL g7567 ( 
.A1(n_6749),
.A2(n_5386),
.B(n_6015),
.C(n_5426),
.Y(n_7567)
);

AND2x4_ASAP7_75t_L g7568 ( 
.A(n_6315),
.B(n_6082),
.Y(n_7568)
);

INVx1_ASAP7_75t_L g7569 ( 
.A(n_6298),
.Y(n_7569)
);

HB1xp67_ASAP7_75t_L g7570 ( 
.A(n_6872),
.Y(n_7570)
);

OAI21x1_ASAP7_75t_L g7571 ( 
.A1(n_6191),
.A2(n_5464),
.B(n_5448),
.Y(n_7571)
);

OAI21x1_ASAP7_75t_L g7572 ( 
.A1(n_6191),
.A2(n_5488),
.B(n_5464),
.Y(n_7572)
);

OAI221xp5_ASAP7_75t_L g7573 ( 
.A1(n_6305),
.A2(n_5393),
.B1(n_5507),
.B2(n_5234),
.C(n_5426),
.Y(n_7573)
);

INVx1_ASAP7_75t_L g7574 ( 
.A(n_6300),
.Y(n_7574)
);

OAI21x1_ASAP7_75t_L g7575 ( 
.A1(n_6976),
.A2(n_5501),
.B(n_5488),
.Y(n_7575)
);

OAI21x1_ASAP7_75t_L g7576 ( 
.A1(n_6976),
.A2(n_7116),
.B(n_6769),
.Y(n_7576)
);

OAI21xp5_ASAP7_75t_L g7577 ( 
.A1(n_7104),
.A2(n_5349),
.B(n_5425),
.Y(n_7577)
);

INVx1_ASAP7_75t_L g7578 ( 
.A(n_6300),
.Y(n_7578)
);

OR2x2_ASAP7_75t_L g7579 ( 
.A(n_6374),
.B(n_6382),
.Y(n_7579)
);

OAI21xp33_ASAP7_75t_SL g7580 ( 
.A1(n_6792),
.A2(n_5360),
.B(n_5958),
.Y(n_7580)
);

BUFx3_ASAP7_75t_L g7581 ( 
.A(n_6315),
.Y(n_7581)
);

BUFx3_ASAP7_75t_L g7582 ( 
.A(n_6315),
.Y(n_7582)
);

INVxp67_ASAP7_75t_L g7583 ( 
.A(n_6194),
.Y(n_7583)
);

OAI21xp5_ASAP7_75t_L g7584 ( 
.A1(n_7104),
.A2(n_5425),
.B(n_5427),
.Y(n_7584)
);

OAI21x1_ASAP7_75t_L g7585 ( 
.A1(n_6769),
.A2(n_5546),
.B(n_5501),
.Y(n_7585)
);

OAI21x1_ASAP7_75t_SL g7586 ( 
.A1(n_6794),
.A2(n_6063),
.B(n_6060),
.Y(n_7586)
);

INVx2_ASAP7_75t_L g7587 ( 
.A(n_6214),
.Y(n_7587)
);

AO21x2_ASAP7_75t_L g7588 ( 
.A1(n_6503),
.A2(n_5532),
.B(n_5524),
.Y(n_7588)
);

BUFx6f_ASAP7_75t_L g7589 ( 
.A(n_6149),
.Y(n_7589)
);

NAND2xp5_ASAP7_75t_L g7590 ( 
.A(n_6708),
.B(n_6073),
.Y(n_7590)
);

OAI21xp5_ASAP7_75t_L g7591 ( 
.A1(n_6326),
.A2(n_5427),
.B(n_5178),
.Y(n_7591)
);

AND2x4_ASAP7_75t_L g7592 ( 
.A(n_6356),
.B(n_6082),
.Y(n_7592)
);

OA21x2_ASAP7_75t_L g7593 ( 
.A1(n_6299),
.A2(n_6307),
.B(n_6382),
.Y(n_7593)
);

AOI21xp5_ASAP7_75t_L g7594 ( 
.A1(n_6527),
.A2(n_5403),
.B(n_5384),
.Y(n_7594)
);

AOI22xp33_ASAP7_75t_L g7595 ( 
.A1(n_6490),
.A2(n_5461),
.B1(n_5346),
.B2(n_5384),
.Y(n_7595)
);

INVx3_ASAP7_75t_L g7596 ( 
.A(n_6356),
.Y(n_7596)
);

OAI21xp5_ASAP7_75t_L g7597 ( 
.A1(n_6302),
.A2(n_5181),
.B(n_5167),
.Y(n_7597)
);

OAI22xp5_ASAP7_75t_L g7598 ( 
.A1(n_6490),
.A2(n_5936),
.B1(n_5962),
.B2(n_5956),
.Y(n_7598)
);

OAI22xp5_ASAP7_75t_L g7599 ( 
.A1(n_7018),
.A2(n_5962),
.B1(n_6051),
.B2(n_6037),
.Y(n_7599)
);

CKINVDCx11_ASAP7_75t_R g7600 ( 
.A(n_6277),
.Y(n_7600)
);

OA21x2_ASAP7_75t_L g7601 ( 
.A1(n_6299),
.A2(n_6307),
.B(n_6384),
.Y(n_7601)
);

OAI21x1_ASAP7_75t_L g7602 ( 
.A1(n_6769),
.A2(n_5615),
.B(n_5546),
.Y(n_7602)
);

AOI22xp33_ASAP7_75t_L g7603 ( 
.A1(n_6494),
.A2(n_5461),
.B1(n_5346),
.B2(n_5384),
.Y(n_7603)
);

O2A1O1Ixp33_ASAP7_75t_L g7604 ( 
.A1(n_6970),
.A2(n_6527),
.B(n_6283),
.C(n_6289),
.Y(n_7604)
);

OR2x2_ASAP7_75t_L g7605 ( 
.A(n_6384),
.B(n_5831),
.Y(n_7605)
);

OAI21x1_ASAP7_75t_L g7606 ( 
.A1(n_7141),
.A2(n_5615),
.B(n_5546),
.Y(n_7606)
);

INVx2_ASAP7_75t_L g7607 ( 
.A(n_6214),
.Y(n_7607)
);

OAI21x1_ASAP7_75t_L g7608 ( 
.A1(n_7141),
.A2(n_5615),
.B(n_5546),
.Y(n_7608)
);

OAI22xp5_ASAP7_75t_L g7609 ( 
.A1(n_7018),
.A2(n_6051),
.B1(n_6084),
.B2(n_6037),
.Y(n_7609)
);

INVx1_ASAP7_75t_SL g7610 ( 
.A(n_6260),
.Y(n_7610)
);

AND2x2_ASAP7_75t_L g7611 ( 
.A(n_6299),
.B(n_5285),
.Y(n_7611)
);

NOR2xp33_ASAP7_75t_L g7612 ( 
.A(n_6343),
.B(n_5994),
.Y(n_7612)
);

OAI21x1_ASAP7_75t_L g7613 ( 
.A1(n_7021),
.A2(n_6879),
.B(n_6725),
.Y(n_7613)
);

INVx1_ASAP7_75t_L g7614 ( 
.A(n_6300),
.Y(n_7614)
);

OAI21x1_ASAP7_75t_L g7615 ( 
.A1(n_7021),
.A2(n_5615),
.B(n_5546),
.Y(n_7615)
);

AOI22xp33_ASAP7_75t_L g7616 ( 
.A1(n_6494),
.A2(n_5344),
.B1(n_5671),
.B2(n_5384),
.Y(n_7616)
);

INVx1_ASAP7_75t_L g7617 ( 
.A(n_6308),
.Y(n_7617)
);

OAI21x1_ASAP7_75t_SL g7618 ( 
.A1(n_6751),
.A2(n_6060),
.B(n_6025),
.Y(n_7618)
);

A2O1A1Ixp33_ASAP7_75t_L g7619 ( 
.A1(n_7092),
.A2(n_6229),
.B(n_6377),
.C(n_6487),
.Y(n_7619)
);

INVx2_ASAP7_75t_L g7620 ( 
.A(n_6214),
.Y(n_7620)
);

OAI21x1_ASAP7_75t_L g7621 ( 
.A1(n_6879),
.A2(n_5656),
.B(n_5615),
.Y(n_7621)
);

OAI21x1_ASAP7_75t_L g7622 ( 
.A1(n_6725),
.A2(n_5684),
.B(n_5656),
.Y(n_7622)
);

OAI21x1_ASAP7_75t_L g7623 ( 
.A1(n_6725),
.A2(n_5684),
.B(n_5656),
.Y(n_7623)
);

OAI21x1_ASAP7_75t_L g7624 ( 
.A1(n_6725),
.A2(n_5684),
.B(n_5656),
.Y(n_7624)
);

HB1xp67_ASAP7_75t_L g7625 ( 
.A(n_6884),
.Y(n_7625)
);

AOI21xp5_ASAP7_75t_L g7626 ( 
.A1(n_6406),
.A2(n_5403),
.B(n_5384),
.Y(n_7626)
);

OAI21x1_ASAP7_75t_L g7627 ( 
.A1(n_6725),
.A2(n_5684),
.B(n_5656),
.Y(n_7627)
);

NAND2xp5_ASAP7_75t_L g7628 ( 
.A(n_6959),
.B(n_6073),
.Y(n_7628)
);

OAI21xp33_ASAP7_75t_L g7629 ( 
.A1(n_6406),
.A2(n_6789),
.B(n_6489),
.Y(n_7629)
);

AOI22xp33_ASAP7_75t_L g7630 ( 
.A1(n_6229),
.A2(n_5344),
.B1(n_5671),
.B2(n_5384),
.Y(n_7630)
);

INVx1_ASAP7_75t_L g7631 ( 
.A(n_6308),
.Y(n_7631)
);

OA21x2_ASAP7_75t_L g7632 ( 
.A1(n_6307),
.A2(n_5539),
.B(n_5532),
.Y(n_7632)
);

OAI21xp5_ASAP7_75t_L g7633 ( 
.A1(n_6302),
.A2(n_5181),
.B(n_5167),
.Y(n_7633)
);

OAI21x1_ASAP7_75t_L g7634 ( 
.A1(n_7068),
.A2(n_5690),
.B(n_5684),
.Y(n_7634)
);

NAND2x1p5_ASAP7_75t_L g7635 ( 
.A(n_6691),
.B(n_5344),
.Y(n_7635)
);

OR2x6_ASAP7_75t_L g7636 ( 
.A(n_6222),
.B(n_5678),
.Y(n_7636)
);

OAI21x1_ASAP7_75t_L g7637 ( 
.A1(n_7068),
.A2(n_5705),
.B(n_5690),
.Y(n_7637)
);

OA21x2_ASAP7_75t_L g7638 ( 
.A1(n_6384),
.A2(n_5539),
.B(n_5201),
.Y(n_7638)
);

CKINVDCx11_ASAP7_75t_R g7639 ( 
.A(n_6428),
.Y(n_7639)
);

OAI21x1_ASAP7_75t_L g7640 ( 
.A1(n_7149),
.A2(n_7100),
.B(n_7095),
.Y(n_7640)
);

OAI21x1_ASAP7_75t_L g7641 ( 
.A1(n_7149),
.A2(n_5705),
.B(n_5690),
.Y(n_7641)
);

INVx1_ASAP7_75t_SL g7642 ( 
.A(n_6292),
.Y(n_7642)
);

OAI211xp5_ASAP7_75t_L g7643 ( 
.A1(n_6506),
.A2(n_5771),
.B(n_5125),
.C(n_5183),
.Y(n_7643)
);

OAI21x1_ASAP7_75t_L g7644 ( 
.A1(n_7095),
.A2(n_5705),
.B(n_5690),
.Y(n_7644)
);

NAND2xp5_ASAP7_75t_SL g7645 ( 
.A(n_6743),
.B(n_5575),
.Y(n_7645)
);

AND2x4_ASAP7_75t_L g7646 ( 
.A(n_6356),
.B(n_6082),
.Y(n_7646)
);

INVx1_ASAP7_75t_L g7647 ( 
.A(n_6308),
.Y(n_7647)
);

BUFx12f_ASAP7_75t_L g7648 ( 
.A(n_6380),
.Y(n_7648)
);

OAI21x1_ASAP7_75t_L g7649 ( 
.A1(n_7100),
.A2(n_5705),
.B(n_5690),
.Y(n_7649)
);

INVxp67_ASAP7_75t_SL g7650 ( 
.A(n_7069),
.Y(n_7650)
);

INVx1_ASAP7_75t_L g7651 ( 
.A(n_6312),
.Y(n_7651)
);

AO21x1_ASAP7_75t_L g7652 ( 
.A1(n_7094),
.A2(n_5139),
.B(n_5131),
.Y(n_7652)
);

INVxp33_ASAP7_75t_L g7653 ( 
.A(n_6894),
.Y(n_7653)
);

O2A1O1Ixp33_ASAP7_75t_SL g7654 ( 
.A1(n_6749),
.A2(n_5578),
.B(n_5580),
.C(n_5205),
.Y(n_7654)
);

INVx3_ASAP7_75t_L g7655 ( 
.A(n_6358),
.Y(n_7655)
);

INVx2_ASAP7_75t_L g7656 ( 
.A(n_6214),
.Y(n_7656)
);

OAI21x1_ASAP7_75t_L g7657 ( 
.A1(n_7015),
.A2(n_5735),
.B(n_5705),
.Y(n_7657)
);

OAI21x1_ASAP7_75t_L g7658 ( 
.A1(n_7015),
.A2(n_5759),
.B(n_5735),
.Y(n_7658)
);

INVx2_ASAP7_75t_L g7659 ( 
.A(n_6232),
.Y(n_7659)
);

OA21x2_ASAP7_75t_L g7660 ( 
.A1(n_6387),
.A2(n_5201),
.B(n_5192),
.Y(n_7660)
);

AND2x2_ASAP7_75t_SL g7661 ( 
.A(n_6743),
.B(n_6082),
.Y(n_7661)
);

OA21x2_ASAP7_75t_L g7662 ( 
.A1(n_6387),
.A2(n_5224),
.B(n_5192),
.Y(n_7662)
);

INVx1_ASAP7_75t_L g7663 ( 
.A(n_6312),
.Y(n_7663)
);

INVx1_ASAP7_75t_L g7664 ( 
.A(n_6312),
.Y(n_7664)
);

NAND2x1p5_ASAP7_75t_L g7665 ( 
.A(n_6743),
.B(n_6679),
.Y(n_7665)
);

INVx3_ASAP7_75t_L g7666 ( 
.A(n_6358),
.Y(n_7666)
);

OAI21x1_ASAP7_75t_L g7667 ( 
.A1(n_7016),
.A2(n_5759),
.B(n_5735),
.Y(n_7667)
);

INVx2_ASAP7_75t_L g7668 ( 
.A(n_6232),
.Y(n_7668)
);

OR2x2_ASAP7_75t_L g7669 ( 
.A(n_6387),
.B(n_6468),
.Y(n_7669)
);

INVx2_ASAP7_75t_L g7670 ( 
.A(n_6232),
.Y(n_7670)
);

AND2x4_ASAP7_75t_L g7671 ( 
.A(n_6358),
.B(n_6082),
.Y(n_7671)
);

INVx1_ASAP7_75t_L g7672 ( 
.A(n_6316),
.Y(n_7672)
);

INVx1_ASAP7_75t_L g7673 ( 
.A(n_6316),
.Y(n_7673)
);

AO31x2_ASAP7_75t_L g7674 ( 
.A1(n_6468),
.A2(n_5231),
.A3(n_5233),
.B(n_5224),
.Y(n_7674)
);

OAI21x1_ASAP7_75t_L g7675 ( 
.A1(n_7016),
.A2(n_5759),
.B(n_5735),
.Y(n_7675)
);

INVx1_ASAP7_75t_SL g7676 ( 
.A(n_6292),
.Y(n_7676)
);

NAND2x1p5_ASAP7_75t_L g7677 ( 
.A(n_6743),
.B(n_5344),
.Y(n_7677)
);

INVx2_ASAP7_75t_L g7678 ( 
.A(n_6232),
.Y(n_7678)
);

NAND2xp5_ASAP7_75t_L g7679 ( 
.A(n_6959),
.B(n_6118),
.Y(n_7679)
);

AOI21xp5_ASAP7_75t_L g7680 ( 
.A1(n_6970),
.A2(n_5403),
.B(n_5344),
.Y(n_7680)
);

INVx2_ASAP7_75t_R g7681 ( 
.A(n_6236),
.Y(n_7681)
);

NOR2xp33_ASAP7_75t_SL g7682 ( 
.A(n_6988),
.B(n_5631),
.Y(n_7682)
);

AO31x2_ASAP7_75t_L g7683 ( 
.A1(n_6468),
.A2(n_5233),
.A3(n_5239),
.B(n_5231),
.Y(n_7683)
);

INVx1_ASAP7_75t_L g7684 ( 
.A(n_6316),
.Y(n_7684)
);

INVx2_ASAP7_75t_L g7685 ( 
.A(n_6244),
.Y(n_7685)
);

NAND2x1p5_ASAP7_75t_L g7686 ( 
.A(n_6679),
.B(n_5344),
.Y(n_7686)
);

OAI21x1_ASAP7_75t_L g7687 ( 
.A1(n_7034),
.A2(n_5759),
.B(n_5735),
.Y(n_7687)
);

OA21x2_ASAP7_75t_L g7688 ( 
.A1(n_6954),
.A2(n_5267),
.B(n_5239),
.Y(n_7688)
);

BUFx3_ASAP7_75t_L g7689 ( 
.A(n_6386),
.Y(n_7689)
);

INVx2_ASAP7_75t_L g7690 ( 
.A(n_6244),
.Y(n_7690)
);

OAI21xp5_ASAP7_75t_L g7691 ( 
.A1(n_6354),
.A2(n_5267),
.B(n_5360),
.Y(n_7691)
);

OAI21x1_ASAP7_75t_L g7692 ( 
.A1(n_7034),
.A2(n_5861),
.B(n_5759),
.Y(n_7692)
);

OAI21x1_ASAP7_75t_L g7693 ( 
.A1(n_7037),
.A2(n_5891),
.B(n_5861),
.Y(n_7693)
);

INVx4_ASAP7_75t_L g7694 ( 
.A(n_6785),
.Y(n_7694)
);

OAI21x1_ASAP7_75t_L g7695 ( 
.A1(n_7037),
.A2(n_5891),
.B(n_5861),
.Y(n_7695)
);

INVx1_ASAP7_75t_SL g7696 ( 
.A(n_6385),
.Y(n_7696)
);

INVx2_ASAP7_75t_L g7697 ( 
.A(n_6244),
.Y(n_7697)
);

AO21x2_ASAP7_75t_L g7698 ( 
.A1(n_6895),
.A2(n_6010),
.B(n_5987),
.Y(n_7698)
);

OAI22xp33_ASAP7_75t_L g7699 ( 
.A1(n_6398),
.A2(n_5424),
.B1(n_6078),
.B2(n_6056),
.Y(n_7699)
);

AND2x4_ASAP7_75t_L g7700 ( 
.A(n_6358),
.B(n_5671),
.Y(n_7700)
);

NOR2x1_ASAP7_75t_SL g7701 ( 
.A(n_6195),
.B(n_5403),
.Y(n_7701)
);

OAI221xp5_ASAP7_75t_L g7702 ( 
.A1(n_6354),
.A2(n_5424),
.B1(n_6106),
.B2(n_6114),
.C(n_6084),
.Y(n_7702)
);

INVx1_ASAP7_75t_L g7703 ( 
.A(n_6323),
.Y(n_7703)
);

OR2x2_ASAP7_75t_L g7704 ( 
.A(n_7018),
.B(n_5831),
.Y(n_7704)
);

AND2x4_ASAP7_75t_L g7705 ( 
.A(n_6378),
.B(n_5671),
.Y(n_7705)
);

AOI22xp33_ASAP7_75t_L g7706 ( 
.A1(n_6351),
.A2(n_5671),
.B1(n_5576),
.B2(n_5401),
.Y(n_7706)
);

AOI221xp5_ASAP7_75t_L g7707 ( 
.A1(n_6283),
.A2(n_5139),
.B1(n_5131),
.B2(n_6118),
.C(n_5159),
.Y(n_7707)
);

NAND2xp5_ASAP7_75t_L g7708 ( 
.A(n_6414),
.B(n_6056),
.Y(n_7708)
);

AND2x4_ASAP7_75t_L g7709 ( 
.A(n_6378),
.B(n_5671),
.Y(n_7709)
);

INVx2_ASAP7_75t_L g7710 ( 
.A(n_6244),
.Y(n_7710)
);

INVx2_ASAP7_75t_L g7711 ( 
.A(n_6247),
.Y(n_7711)
);

AND2x2_ASAP7_75t_L g7712 ( 
.A(n_6655),
.B(n_6478),
.Y(n_7712)
);

AOI21xp5_ASAP7_75t_L g7713 ( 
.A1(n_7006),
.A2(n_5671),
.B(n_5505),
.Y(n_7713)
);

INVx1_ASAP7_75t_L g7714 ( 
.A(n_6323),
.Y(n_7714)
);

AOI222xp33_ASAP7_75t_SL g7715 ( 
.A1(n_6506),
.A2(n_5199),
.B1(n_5166),
.B2(n_5209),
.C1(n_5183),
.C2(n_5125),
.Y(n_7715)
);

OAI22xp33_ASAP7_75t_L g7716 ( 
.A1(n_6398),
.A2(n_6078),
.B1(n_5983),
.B2(n_5988),
.Y(n_7716)
);

OAI21xp5_ASAP7_75t_L g7717 ( 
.A1(n_6351),
.A2(n_5343),
.B(n_5338),
.Y(n_7717)
);

AO31x2_ASAP7_75t_L g7718 ( 
.A1(n_6289),
.A2(n_5667),
.A3(n_5676),
.B(n_5663),
.Y(n_7718)
);

INVx2_ASAP7_75t_L g7719 ( 
.A(n_6247),
.Y(n_7719)
);

AO21x2_ASAP7_75t_L g7720 ( 
.A1(n_6895),
.A2(n_6065),
.B(n_5987),
.Y(n_7720)
);

BUFx2_ASAP7_75t_L g7721 ( 
.A(n_6378),
.Y(n_7721)
);

OAI22xp5_ASAP7_75t_L g7722 ( 
.A1(n_6539),
.A2(n_6114),
.B1(n_6106),
.B2(n_5994),
.Y(n_7722)
);

INVx2_ASAP7_75t_L g7723 ( 
.A(n_6247),
.Y(n_7723)
);

AO21x2_ASAP7_75t_L g7724 ( 
.A1(n_6897),
.A2(n_6085),
.B(n_6065),
.Y(n_7724)
);

INVx2_ASAP7_75t_L g7725 ( 
.A(n_6247),
.Y(n_7725)
);

INVx4_ASAP7_75t_L g7726 ( 
.A(n_6785),
.Y(n_7726)
);

INVx1_ASAP7_75t_SL g7727 ( 
.A(n_6385),
.Y(n_7727)
);

AND2x2_ASAP7_75t_L g7728 ( 
.A(n_6655),
.B(n_5285),
.Y(n_7728)
);

INVx1_ASAP7_75t_L g7729 ( 
.A(n_6323),
.Y(n_7729)
);

INVx2_ASAP7_75t_SL g7730 ( 
.A(n_6378),
.Y(n_7730)
);

AOI21xp33_ASAP7_75t_SL g7731 ( 
.A1(n_6154),
.A2(n_6164),
.B(n_6343),
.Y(n_7731)
);

AND2x2_ASAP7_75t_L g7732 ( 
.A(n_6655),
.B(n_6478),
.Y(n_7732)
);

OA21x2_ASAP7_75t_L g7733 ( 
.A1(n_6954),
.A2(n_5480),
.B(n_5471),
.Y(n_7733)
);

INVx2_ASAP7_75t_L g7734 ( 
.A(n_6251),
.Y(n_7734)
);

AOI21xp5_ASAP7_75t_L g7735 ( 
.A1(n_7006),
.A2(n_5505),
.B(n_5999),
.Y(n_7735)
);

OAI22xp33_ASAP7_75t_L g7736 ( 
.A1(n_6409),
.A2(n_5983),
.B1(n_5988),
.B2(n_5831),
.Y(n_7736)
);

NOR2xp33_ASAP7_75t_L g7737 ( 
.A(n_6165),
.B(n_5343),
.Y(n_7737)
);

INVx2_ASAP7_75t_L g7738 ( 
.A(n_6251),
.Y(n_7738)
);

INVx1_ASAP7_75t_L g7739 ( 
.A(n_6330),
.Y(n_7739)
);

OAI222xp33_ASAP7_75t_L g7740 ( 
.A1(n_6988),
.A2(n_5822),
.B1(n_5678),
.B2(n_5882),
.C1(n_5874),
.C2(n_5760),
.Y(n_7740)
);

OA21x2_ASAP7_75t_L g7741 ( 
.A1(n_7029),
.A2(n_5480),
.B(n_5471),
.Y(n_7741)
);

INVx1_ASAP7_75t_SL g7742 ( 
.A(n_6413),
.Y(n_7742)
);

CKINVDCx5p33_ASAP7_75t_R g7743 ( 
.A(n_7056),
.Y(n_7743)
);

INVx2_ASAP7_75t_L g7744 ( 
.A(n_6251),
.Y(n_7744)
);

INVx1_ASAP7_75t_L g7745 ( 
.A(n_6330),
.Y(n_7745)
);

INVx2_ASAP7_75t_L g7746 ( 
.A(n_6251),
.Y(n_7746)
);

NOR2xp67_ASAP7_75t_L g7747 ( 
.A(n_6195),
.B(n_5345),
.Y(n_7747)
);

INVx1_ASAP7_75t_L g7748 ( 
.A(n_6330),
.Y(n_7748)
);

O2A1O1Ixp33_ASAP7_75t_L g7749 ( 
.A1(n_6190),
.A2(n_5417),
.B(n_5527),
.C(n_5400),
.Y(n_7749)
);

AOI221xp5_ASAP7_75t_L g7750 ( 
.A1(n_6225),
.A2(n_5159),
.B1(n_5142),
.B2(n_6024),
.C(n_6019),
.Y(n_7750)
);

AO21x2_ASAP7_75t_L g7751 ( 
.A1(n_6897),
.A2(n_6092),
.B(n_6085),
.Y(n_7751)
);

A2O1A1Ixp33_ASAP7_75t_L g7752 ( 
.A1(n_7092),
.A2(n_5285),
.B(n_5855),
.C(n_5281),
.Y(n_7752)
);

OA21x2_ASAP7_75t_L g7753 ( 
.A1(n_7029),
.A2(n_5487),
.B(n_5480),
.Y(n_7753)
);

INVx4_ASAP7_75t_SL g7754 ( 
.A(n_6753),
.Y(n_7754)
);

INVx2_ASAP7_75t_SL g7755 ( 
.A(n_6386),
.Y(n_7755)
);

AND2x2_ASAP7_75t_L g7756 ( 
.A(n_6478),
.B(n_6590),
.Y(n_7756)
);

OAI22xp33_ASAP7_75t_L g7757 ( 
.A1(n_6409),
.A2(n_5837),
.B1(n_5678),
.B2(n_5822),
.Y(n_7757)
);

INVx1_ASAP7_75t_L g7758 ( 
.A(n_6332),
.Y(n_7758)
);

OAI21x1_ASAP7_75t_SL g7759 ( 
.A1(n_6751),
.A2(n_6060),
.B(n_6025),
.Y(n_7759)
);

OA21x2_ASAP7_75t_L g7760 ( 
.A1(n_7055),
.A2(n_5494),
.B(n_5487),
.Y(n_7760)
);

AND2x2_ASAP7_75t_L g7761 ( 
.A(n_6590),
.B(n_5285),
.Y(n_7761)
);

INVx1_ASAP7_75t_L g7762 ( 
.A(n_6332),
.Y(n_7762)
);

OAI21xp5_ASAP7_75t_L g7763 ( 
.A1(n_6377),
.A2(n_5417),
.B(n_5400),
.Y(n_7763)
);

AO31x2_ASAP7_75t_L g7764 ( 
.A1(n_6620),
.A2(n_5667),
.A3(n_5693),
.B(n_5676),
.Y(n_7764)
);

INVx5_ASAP7_75t_L g7765 ( 
.A(n_6920),
.Y(n_7765)
);

AND2x2_ASAP7_75t_L g7766 ( 
.A(n_6590),
.B(n_5171),
.Y(n_7766)
);

HB1xp67_ASAP7_75t_L g7767 ( 
.A(n_6884),
.Y(n_7767)
);

NOR2xp67_ASAP7_75t_L g7768 ( 
.A(n_6430),
.B(n_5345),
.Y(n_7768)
);

A2O1A1Ixp33_ASAP7_75t_L g7769 ( 
.A1(n_6487),
.A2(n_5855),
.B(n_5281),
.C(n_5282),
.Y(n_7769)
);

INVx1_ASAP7_75t_L g7770 ( 
.A(n_6332),
.Y(n_7770)
);

INVx1_ASAP7_75t_L g7771 ( 
.A(n_6336),
.Y(n_7771)
);

AOI22xp33_ASAP7_75t_SL g7772 ( 
.A1(n_6506),
.A2(n_5281),
.B1(n_5855),
.B2(n_5576),
.Y(n_7772)
);

INVx2_ASAP7_75t_L g7773 ( 
.A(n_6268),
.Y(n_7773)
);

INVx1_ASAP7_75t_L g7774 ( 
.A(n_6336),
.Y(n_7774)
);

INVx2_ASAP7_75t_L g7775 ( 
.A(n_6268),
.Y(n_7775)
);

OR2x6_ASAP7_75t_L g7776 ( 
.A(n_6222),
.B(n_5678),
.Y(n_7776)
);

AND2x4_ASAP7_75t_L g7777 ( 
.A(n_6389),
.B(n_5365),
.Y(n_7777)
);

INVx1_ASAP7_75t_L g7778 ( 
.A(n_6336),
.Y(n_7778)
);

AOI21xp33_ASAP7_75t_L g7779 ( 
.A1(n_6533),
.A2(n_5527),
.B(n_6092),
.Y(n_7779)
);

INVx1_ASAP7_75t_L g7780 ( 
.A(n_6342),
.Y(n_7780)
);

BUFx2_ASAP7_75t_L g7781 ( 
.A(n_6386),
.Y(n_7781)
);

BUFx2_ASAP7_75t_L g7782 ( 
.A(n_6386),
.Y(n_7782)
);

NAND2xp5_ASAP7_75t_L g7783 ( 
.A(n_6414),
.B(n_5685),
.Y(n_7783)
);

INVx6_ASAP7_75t_SL g7784 ( 
.A(n_6686),
.Y(n_7784)
);

AND2x4_ASAP7_75t_L g7785 ( 
.A(n_6389),
.B(n_5365),
.Y(n_7785)
);

AOI21xp5_ASAP7_75t_L g7786 ( 
.A1(n_6528),
.A2(n_5696),
.B(n_5685),
.Y(n_7786)
);

CKINVDCx6p67_ASAP7_75t_R g7787 ( 
.A(n_6182),
.Y(n_7787)
);

OAI21x1_ASAP7_75t_L g7788 ( 
.A1(n_6158),
.A2(n_6027),
.B(n_6013),
.Y(n_7788)
);

OAI21x1_ASAP7_75t_L g7789 ( 
.A1(n_6158),
.A2(n_6027),
.B(n_6013),
.Y(n_7789)
);

CKINVDCx5p33_ASAP7_75t_R g7790 ( 
.A(n_6840),
.Y(n_7790)
);

INVx1_ASAP7_75t_L g7791 ( 
.A(n_6342),
.Y(n_7791)
);

AOI22xp33_ASAP7_75t_L g7792 ( 
.A1(n_6190),
.A2(n_5576),
.B1(n_5401),
.B2(n_4583),
.Y(n_7792)
);

HB1xp67_ASAP7_75t_L g7793 ( 
.A(n_6888),
.Y(n_7793)
);

INVx2_ASAP7_75t_L g7794 ( 
.A(n_6268),
.Y(n_7794)
);

AOI22x1_ASAP7_75t_L g7795 ( 
.A1(n_6188),
.A2(n_4706),
.B1(n_6046),
.B2(n_4735),
.Y(n_7795)
);

HB1xp67_ASAP7_75t_L g7796 ( 
.A(n_6888),
.Y(n_7796)
);

O2A1O1Ixp5_ASAP7_75t_L g7797 ( 
.A1(n_6528),
.A2(n_5721),
.B(n_5730),
.C(n_5696),
.Y(n_7797)
);

OA21x2_ASAP7_75t_L g7798 ( 
.A1(n_7055),
.A2(n_5494),
.B(n_5487),
.Y(n_7798)
);

OAI21x1_ASAP7_75t_L g7799 ( 
.A1(n_6541),
.A2(n_6069),
.B(n_6027),
.Y(n_7799)
);

AOI222xp33_ASAP7_75t_L g7800 ( 
.A1(n_6225),
.A2(n_5142),
.B1(n_5563),
.B2(n_5499),
.C1(n_6040),
.C2(n_6033),
.Y(n_7800)
);

AOI21xp5_ASAP7_75t_L g7801 ( 
.A1(n_6942),
.A2(n_5730),
.B(n_5721),
.Y(n_7801)
);

O2A1O1Ixp33_ASAP7_75t_SL g7802 ( 
.A1(n_7118),
.A2(n_5580),
.B(n_5578),
.C(n_5205),
.Y(n_7802)
);

INVx2_ASAP7_75t_L g7803 ( 
.A(n_6268),
.Y(n_7803)
);

OAI21x1_ASAP7_75t_L g7804 ( 
.A1(n_6541),
.A2(n_6111),
.B(n_6069),
.Y(n_7804)
);

AND2x4_ASAP7_75t_L g7805 ( 
.A(n_6389),
.B(n_5365),
.Y(n_7805)
);

AOI22xp33_ASAP7_75t_L g7806 ( 
.A1(n_7009),
.A2(n_5576),
.B1(n_4595),
.B2(n_4621),
.Y(n_7806)
);

INVx1_ASAP7_75t_L g7807 ( 
.A(n_6342),
.Y(n_7807)
);

NOR2x1_ASAP7_75t_R g7808 ( 
.A(n_6785),
.B(n_4159),
.Y(n_7808)
);

INVx1_ASAP7_75t_SL g7809 ( 
.A(n_6413),
.Y(n_7809)
);

CKINVDCx20_ASAP7_75t_R g7810 ( 
.A(n_6346),
.Y(n_7810)
);

OAI22xp5_ASAP7_75t_L g7811 ( 
.A1(n_6539),
.A2(n_5631),
.B1(n_5205),
.B2(n_5837),
.Y(n_7811)
);

INVx1_ASAP7_75t_L g7812 ( 
.A(n_6349),
.Y(n_7812)
);

OA21x2_ASAP7_75t_L g7813 ( 
.A1(n_7107),
.A2(n_5521),
.B(n_5494),
.Y(n_7813)
);

BUFx3_ASAP7_75t_L g7814 ( 
.A(n_6405),
.Y(n_7814)
);

CKINVDCx6p67_ASAP7_75t_R g7815 ( 
.A(n_6182),
.Y(n_7815)
);

AO31x2_ASAP7_75t_L g7816 ( 
.A1(n_6620),
.A2(n_5695),
.A3(n_5701),
.B(n_5693),
.Y(n_7816)
);

AOI22xp33_ASAP7_75t_L g7817 ( 
.A1(n_7009),
.A2(n_5576),
.B1(n_4595),
.B2(n_4621),
.Y(n_7817)
);

AND2x2_ASAP7_75t_L g7818 ( 
.A(n_6877),
.B(n_5171),
.Y(n_7818)
);

INVx1_ASAP7_75t_L g7819 ( 
.A(n_6349),
.Y(n_7819)
);

AOI22xp33_ASAP7_75t_L g7820 ( 
.A1(n_6841),
.A2(n_5576),
.B1(n_4595),
.B2(n_4621),
.Y(n_7820)
);

BUFx2_ASAP7_75t_L g7821 ( 
.A(n_6389),
.Y(n_7821)
);

OAI21x1_ASAP7_75t_L g7822 ( 
.A1(n_7064),
.A2(n_6111),
.B(n_6069),
.Y(n_7822)
);

O2A1O1Ixp33_ASAP7_75t_L g7823 ( 
.A1(n_6391),
.A2(n_5733),
.B(n_5766),
.C(n_5731),
.Y(n_7823)
);

BUFx3_ASAP7_75t_L g7824 ( 
.A(n_6405),
.Y(n_7824)
);

NAND2x1p5_ASAP7_75t_L g7825 ( 
.A(n_6679),
.B(n_4795),
.Y(n_7825)
);

AOI21xp5_ASAP7_75t_L g7826 ( 
.A1(n_6942),
.A2(n_5733),
.B(n_5731),
.Y(n_7826)
);

OAI21x1_ASAP7_75t_L g7827 ( 
.A1(n_7064),
.A2(n_6111),
.B(n_6069),
.Y(n_7827)
);

OAI21x1_ASAP7_75t_L g7828 ( 
.A1(n_6589),
.A2(n_6111),
.B(n_6069),
.Y(n_7828)
);

NAND2xp5_ASAP7_75t_L g7829 ( 
.A(n_6437),
.B(n_6442),
.Y(n_7829)
);

INVxp67_ASAP7_75t_L g7830 ( 
.A(n_7019),
.Y(n_7830)
);

INVx1_ASAP7_75t_L g7831 ( 
.A(n_6349),
.Y(n_7831)
);

BUFx3_ASAP7_75t_L g7832 ( 
.A(n_6405),
.Y(n_7832)
);

AND2x2_ASAP7_75t_L g7833 ( 
.A(n_6877),
.B(n_5171),
.Y(n_7833)
);

OAI22xp5_ASAP7_75t_L g7834 ( 
.A1(n_6160),
.A2(n_5631),
.B1(n_5837),
.B2(n_6019),
.Y(n_7834)
);

AO31x2_ASAP7_75t_L g7835 ( 
.A1(n_6391),
.A2(n_6584),
.A3(n_6634),
.B(n_6497),
.Y(n_7835)
);

NOR2xp33_ASAP7_75t_L g7836 ( 
.A(n_6165),
.B(n_6046),
.Y(n_7836)
);

BUFx6f_ASAP7_75t_L g7837 ( 
.A(n_6149),
.Y(n_7837)
);

OAI21xp5_ASAP7_75t_L g7838 ( 
.A1(n_6538),
.A2(n_5775),
.B(n_5766),
.Y(n_7838)
);

INVx1_ASAP7_75t_L g7839 ( 
.A(n_6365),
.Y(n_7839)
);

INVx2_ASAP7_75t_L g7840 ( 
.A(n_6286),
.Y(n_7840)
);

INVx2_ASAP7_75t_SL g7841 ( 
.A(n_6405),
.Y(n_7841)
);

BUFx8_ASAP7_75t_L g7842 ( 
.A(n_6785),
.Y(n_7842)
);

INVx1_ASAP7_75t_SL g7843 ( 
.A(n_6418),
.Y(n_7843)
);

AOI22xp33_ASAP7_75t_L g7844 ( 
.A1(n_6841),
.A2(n_4595),
.B1(n_4621),
.B2(n_4501),
.Y(n_7844)
);

AO21x2_ASAP7_75t_L g7845 ( 
.A1(n_6996),
.A2(n_5522),
.B(n_5521),
.Y(n_7845)
);

INVx2_ASAP7_75t_L g7846 ( 
.A(n_6286),
.Y(n_7846)
);

OAI21x1_ASAP7_75t_L g7847 ( 
.A1(n_6589),
.A2(n_7107),
.B(n_6681),
.Y(n_7847)
);

NAND2xp5_ASAP7_75t_L g7848 ( 
.A(n_6437),
.B(n_5775),
.Y(n_7848)
);

OAI21x1_ASAP7_75t_L g7849 ( 
.A1(n_6589),
.A2(n_6681),
.B(n_6597),
.Y(n_7849)
);

INVx2_ASAP7_75t_L g7850 ( 
.A(n_6286),
.Y(n_7850)
);

OAI21x1_ASAP7_75t_L g7851 ( 
.A1(n_6589),
.A2(n_6116),
.B(n_6111),
.Y(n_7851)
);

AO31x2_ASAP7_75t_L g7852 ( 
.A1(n_6584),
.A2(n_5701),
.A3(n_5711),
.B(n_5695),
.Y(n_7852)
);

OAI21x1_ASAP7_75t_L g7853 ( 
.A1(n_6589),
.A2(n_6681),
.B(n_6597),
.Y(n_7853)
);

INVx1_ASAP7_75t_L g7854 ( 
.A(n_6365),
.Y(n_7854)
);

CKINVDCx11_ASAP7_75t_R g7855 ( 
.A(n_6428),
.Y(n_7855)
);

INVx1_ASAP7_75t_L g7856 ( 
.A(n_6365),
.Y(n_7856)
);

INVx1_ASAP7_75t_L g7857 ( 
.A(n_6368),
.Y(n_7857)
);

INVx1_ASAP7_75t_L g7858 ( 
.A(n_6368),
.Y(n_7858)
);

INVx1_ASAP7_75t_SL g7859 ( 
.A(n_6418),
.Y(n_7859)
);

AOI22xp5_ASAP7_75t_L g7860 ( 
.A1(n_6169),
.A2(n_5913),
.B1(n_5877),
.B2(n_5563),
.Y(n_7860)
);

NOR2xp67_ASAP7_75t_L g7861 ( 
.A(n_6430),
.B(n_5365),
.Y(n_7861)
);

BUFx6f_ASAP7_75t_L g7862 ( 
.A(n_6149),
.Y(n_7862)
);

NOR2x1_ASAP7_75t_SL g7863 ( 
.A(n_6920),
.B(n_5760),
.Y(n_7863)
);

OAI21x1_ASAP7_75t_L g7864 ( 
.A1(n_6543),
.A2(n_6856),
.B(n_7134),
.Y(n_7864)
);

OAI21x1_ASAP7_75t_L g7865 ( 
.A1(n_6543),
.A2(n_6116),
.B(n_6016),
.Y(n_7865)
);

OAI21x1_ASAP7_75t_L g7866 ( 
.A1(n_6856),
.A2(n_6116),
.B(n_6016),
.Y(n_7866)
);

AO21x2_ASAP7_75t_L g7867 ( 
.A1(n_6996),
.A2(n_6113),
.B(n_6110),
.Y(n_7867)
);

OAI22xp5_ASAP7_75t_L g7868 ( 
.A1(n_6160),
.A2(n_6024),
.B1(n_5199),
.B2(n_5209),
.Y(n_7868)
);

OA21x2_ASAP7_75t_L g7869 ( 
.A1(n_6950),
.A2(n_5522),
.B(n_5521),
.Y(n_7869)
);

NAND2x1p5_ASAP7_75t_L g7870 ( 
.A(n_6679),
.B(n_4795),
.Y(n_7870)
);

INVx1_ASAP7_75t_L g7871 ( 
.A(n_6368),
.Y(n_7871)
);

OAI21x1_ASAP7_75t_SL g7872 ( 
.A1(n_6950),
.A2(n_6063),
.B(n_6025),
.Y(n_7872)
);

BUFx4f_ASAP7_75t_SL g7873 ( 
.A(n_6840),
.Y(n_7873)
);

NOR2xp33_ASAP7_75t_SL g7874 ( 
.A(n_6988),
.B(n_5365),
.Y(n_7874)
);

INVx2_ASAP7_75t_L g7875 ( 
.A(n_6286),
.Y(n_7875)
);

OAI21xp5_ASAP7_75t_L g7876 ( 
.A1(n_6538),
.A2(n_5790),
.B(n_5782),
.Y(n_7876)
);

INVx1_ASAP7_75t_L g7877 ( 
.A(n_6376),
.Y(n_7877)
);

O2A1O1Ixp33_ASAP7_75t_L g7878 ( 
.A1(n_7094),
.A2(n_5790),
.B(n_5793),
.C(n_5782),
.Y(n_7878)
);

CKINVDCx20_ASAP7_75t_R g7879 ( 
.A(n_6346),
.Y(n_7879)
);

AOI21x1_ASAP7_75t_L g7880 ( 
.A1(n_6451),
.A2(n_5148),
.B(n_5105),
.Y(n_7880)
);

AOI22xp33_ASAP7_75t_L g7881 ( 
.A1(n_6253),
.A2(n_4595),
.B1(n_4621),
.B2(n_4501),
.Y(n_7881)
);

AND2x2_ASAP7_75t_L g7882 ( 
.A(n_6877),
.B(n_5245),
.Y(n_7882)
);

NOR2xp33_ASAP7_75t_L g7883 ( 
.A(n_6166),
.B(n_6033),
.Y(n_7883)
);

OAI21xp5_ASAP7_75t_L g7884 ( 
.A1(n_6533),
.A2(n_5803),
.B(n_5793),
.Y(n_7884)
);

OAI21x1_ASAP7_75t_L g7885 ( 
.A1(n_7134),
.A2(n_6102),
.B(n_5981),
.Y(n_7885)
);

OAI21xp5_ASAP7_75t_L g7886 ( 
.A1(n_6169),
.A2(n_5821),
.B(n_5803),
.Y(n_7886)
);

AO21x2_ASAP7_75t_L g7887 ( 
.A1(n_7099),
.A2(n_5525),
.B(n_5522),
.Y(n_7887)
);

INVx2_ASAP7_75t_L g7888 ( 
.A(n_6288),
.Y(n_7888)
);

BUFx3_ASAP7_75t_L g7889 ( 
.A(n_6495),
.Y(n_7889)
);

OA21x2_ASAP7_75t_L g7890 ( 
.A1(n_6240),
.A2(n_6461),
.B(n_6574),
.Y(n_7890)
);

CKINVDCx9p33_ASAP7_75t_R g7891 ( 
.A(n_6782),
.Y(n_7891)
);

INVx4_ASAP7_75t_L g7892 ( 
.A(n_6185),
.Y(n_7892)
);

AOI22xp5_ASAP7_75t_L g7893 ( 
.A1(n_6253),
.A2(n_5563),
.B1(n_5499),
.B2(n_4595),
.Y(n_7893)
);

OAI21x1_ASAP7_75t_L g7894 ( 
.A1(n_7134),
.A2(n_7153),
.B(n_6209),
.Y(n_7894)
);

AOI21xp5_ASAP7_75t_L g7895 ( 
.A1(n_6240),
.A2(n_5827),
.B(n_5821),
.Y(n_7895)
);

AND2x4_ASAP7_75t_L g7896 ( 
.A(n_6495),
.B(n_5389),
.Y(n_7896)
);

BUFx2_ASAP7_75t_L g7897 ( 
.A(n_6479),
.Y(n_7897)
);

INVx1_ASAP7_75t_L g7898 ( 
.A(n_6376),
.Y(n_7898)
);

BUFx3_ASAP7_75t_L g7899 ( 
.A(n_6479),
.Y(n_7899)
);

AND2x4_ASAP7_75t_L g7900 ( 
.A(n_6495),
.B(n_5389),
.Y(n_7900)
);

INVx3_ASAP7_75t_L g7901 ( 
.A(n_6479),
.Y(n_7901)
);

INVx2_ASAP7_75t_L g7902 ( 
.A(n_6288),
.Y(n_7902)
);

OAI21x1_ASAP7_75t_L g7903 ( 
.A1(n_7153),
.A2(n_6102),
.B(n_5981),
.Y(n_7903)
);

BUFx8_ASAP7_75t_SL g7904 ( 
.A(n_6259),
.Y(n_7904)
);

OAI21xp5_ASAP7_75t_L g7905 ( 
.A1(n_7031),
.A2(n_5835),
.B(n_5827),
.Y(n_7905)
);

BUFx6f_ASAP7_75t_L g7906 ( 
.A(n_6149),
.Y(n_7906)
);

OAI21x1_ASAP7_75t_L g7907 ( 
.A1(n_7153),
.A2(n_6102),
.B(n_5981),
.Y(n_7907)
);

AND2x4_ASAP7_75t_L g7908 ( 
.A(n_6479),
.B(n_5389),
.Y(n_7908)
);

INVx2_ASAP7_75t_L g7909 ( 
.A(n_6288),
.Y(n_7909)
);

OA21x2_ASAP7_75t_L g7910 ( 
.A1(n_6461),
.A2(n_5552),
.B(n_5525),
.Y(n_7910)
);

AND2x4_ASAP7_75t_L g7911 ( 
.A(n_6495),
.B(n_5389),
.Y(n_7911)
);

INVx1_ASAP7_75t_L g7912 ( 
.A(n_6376),
.Y(n_7912)
);

AOI22xp33_ASAP7_75t_L g7913 ( 
.A1(n_7099),
.A2(n_4621),
.B1(n_4753),
.B2(n_4501),
.Y(n_7913)
);

NAND2x1p5_ASAP7_75t_L g7914 ( 
.A(n_6412),
.B(n_4795),
.Y(n_7914)
);

BUFx2_ASAP7_75t_L g7915 ( 
.A(n_6430),
.Y(n_7915)
);

INVx2_ASAP7_75t_L g7916 ( 
.A(n_6288),
.Y(n_7916)
);

OAI21x1_ASAP7_75t_L g7917 ( 
.A1(n_7153),
.A2(n_6102),
.B(n_5981),
.Y(n_7917)
);

AO21x2_ASAP7_75t_L g7918 ( 
.A1(n_7114),
.A2(n_6115),
.B(n_6113),
.Y(n_7918)
);

AND2x2_ASAP7_75t_L g7919 ( 
.A(n_6778),
.B(n_7038),
.Y(n_7919)
);

INVx6_ASAP7_75t_L g7920 ( 
.A(n_6430),
.Y(n_7920)
);

NAND2xp5_ASAP7_75t_L g7921 ( 
.A(n_6442),
.B(n_5835),
.Y(n_7921)
);

OAI21xp5_ASAP7_75t_L g7922 ( 
.A1(n_7031),
.A2(n_6789),
.B(n_6465),
.Y(n_7922)
);

AO32x2_ASAP7_75t_L g7923 ( 
.A1(n_6129),
.A2(n_5185),
.A3(n_5305),
.B1(n_5148),
.B2(n_5105),
.Y(n_7923)
);

INVx1_ASAP7_75t_L g7924 ( 
.A(n_6381),
.Y(n_7924)
);

AND2x4_ASAP7_75t_L g7925 ( 
.A(n_6430),
.B(n_5389),
.Y(n_7925)
);

AND2x2_ASAP7_75t_L g7926 ( 
.A(n_6778),
.B(n_5245),
.Y(n_7926)
);

AND2x4_ASAP7_75t_L g7927 ( 
.A(n_6430),
.B(n_5394),
.Y(n_7927)
);

OAI21x1_ASAP7_75t_L g7928 ( 
.A1(n_6209),
.A2(n_6817),
.B(n_6806),
.Y(n_7928)
);

AOI21xp5_ASAP7_75t_L g7929 ( 
.A1(n_6574),
.A2(n_5849),
.B(n_5841),
.Y(n_7929)
);

AO31x2_ASAP7_75t_L g7930 ( 
.A1(n_6634),
.A2(n_5716),
.A3(n_5728),
.B(n_5711),
.Y(n_7930)
);

OAI21xp5_ASAP7_75t_L g7931 ( 
.A1(n_6465),
.A2(n_5849),
.B(n_5841),
.Y(n_7931)
);

NOR2xp33_ASAP7_75t_L g7932 ( 
.A(n_6166),
.B(n_6518),
.Y(n_7932)
);

NAND2xp5_ASAP7_75t_L g7933 ( 
.A(n_6448),
.B(n_5853),
.Y(n_7933)
);

OR2x2_ASAP7_75t_L g7934 ( 
.A(n_6756),
.B(n_6768),
.Y(n_7934)
);

AND2x2_ASAP7_75t_L g7935 ( 
.A(n_6778),
.B(n_5245),
.Y(n_7935)
);

INVx2_ASAP7_75t_L g7936 ( 
.A(n_6301),
.Y(n_7936)
);

NAND2xp5_ASAP7_75t_L g7937 ( 
.A(n_6448),
.B(n_5853),
.Y(n_7937)
);

CKINVDCx20_ASAP7_75t_R g7938 ( 
.A(n_6507),
.Y(n_7938)
);

AO21x2_ASAP7_75t_L g7939 ( 
.A1(n_7114),
.A2(n_7115),
.B(n_6451),
.Y(n_7939)
);

INVx2_ASAP7_75t_L g7940 ( 
.A(n_6301),
.Y(n_7940)
);

INVx3_ASAP7_75t_L g7941 ( 
.A(n_6569),
.Y(n_7941)
);

INVx1_ASAP7_75t_L g7942 ( 
.A(n_6381),
.Y(n_7942)
);

BUFx3_ASAP7_75t_L g7943 ( 
.A(n_6273),
.Y(n_7943)
);

NOR2xp33_ASAP7_75t_L g7944 ( 
.A(n_6518),
.B(n_6040),
.Y(n_7944)
);

OAI21x1_ASAP7_75t_L g7945 ( 
.A1(n_6209),
.A2(n_5423),
.B(n_5335),
.Y(n_7945)
);

OAI21x1_ASAP7_75t_L g7946 ( 
.A1(n_6806),
.A2(n_5423),
.B(n_5335),
.Y(n_7946)
);

NAND2xp5_ASAP7_75t_L g7947 ( 
.A(n_7024),
.B(n_5859),
.Y(n_7947)
);

NAND2xp5_ASAP7_75t_L g7948 ( 
.A(n_7024),
.B(n_5859),
.Y(n_7948)
);

OR2x6_ASAP7_75t_L g7949 ( 
.A(n_6222),
.B(n_5760),
.Y(n_7949)
);

AND2x2_ASAP7_75t_L g7950 ( 
.A(n_7038),
.B(n_5279),
.Y(n_7950)
);

NAND2xp33_ASAP7_75t_L g7951 ( 
.A(n_6615),
.B(n_5952),
.Y(n_7951)
);

OAI22xp5_ASAP7_75t_L g7952 ( 
.A1(n_6261),
.A2(n_5227),
.B1(n_5246),
.B2(n_5166),
.Y(n_7952)
);

NAND2xp5_ASAP7_75t_L g7953 ( 
.A(n_7050),
.B(n_5894),
.Y(n_7953)
);

OAI21x1_ASAP7_75t_SL g7954 ( 
.A1(n_6156),
.A2(n_6063),
.B(n_5989),
.Y(n_7954)
);

BUFx6f_ASAP7_75t_L g7955 ( 
.A(n_6149),
.Y(n_7955)
);

NAND2xp5_ASAP7_75t_L g7956 ( 
.A(n_7050),
.B(n_5894),
.Y(n_7956)
);

OAI21x1_ASAP7_75t_L g7957 ( 
.A1(n_6817),
.A2(n_5423),
.B(n_5335),
.Y(n_7957)
);

OA21x2_ASAP7_75t_L g7958 ( 
.A1(n_6605),
.A2(n_5552),
.B(n_5525),
.Y(n_7958)
);

OAI21x1_ASAP7_75t_L g7959 ( 
.A1(n_6173),
.A2(n_6175),
.B(n_6140),
.Y(n_7959)
);

OAI22xp5_ASAP7_75t_L g7960 ( 
.A1(n_6261),
.A2(n_5246),
.B1(n_5266),
.B2(n_5227),
.Y(n_7960)
);

OAI21xp5_ASAP7_75t_L g7961 ( 
.A1(n_6183),
.A2(n_6452),
.B(n_6514),
.Y(n_7961)
);

INVx2_ASAP7_75t_L g7962 ( 
.A(n_6301),
.Y(n_7962)
);

AND2x4_ASAP7_75t_L g7963 ( 
.A(n_6569),
.B(n_5394),
.Y(n_7963)
);

INVx2_ASAP7_75t_SL g7964 ( 
.A(n_6766),
.Y(n_7964)
);

CKINVDCx20_ASAP7_75t_R g7965 ( 
.A(n_6507),
.Y(n_7965)
);

INVx1_ASAP7_75t_L g7966 ( 
.A(n_6381),
.Y(n_7966)
);

AOI21x1_ASAP7_75t_L g7967 ( 
.A1(n_6981),
.A2(n_5148),
.B(n_5105),
.Y(n_7967)
);

OAI21x1_ASAP7_75t_L g7968 ( 
.A1(n_6173),
.A2(n_5565),
.B(n_5447),
.Y(n_7968)
);

INVxp67_ASAP7_75t_SL g7969 ( 
.A(n_7072),
.Y(n_7969)
);

NOR2xp33_ASAP7_75t_L g7970 ( 
.A(n_7135),
.B(n_4719),
.Y(n_7970)
);

AOI22xp33_ASAP7_75t_SL g7971 ( 
.A1(n_6792),
.A2(n_5760),
.B1(n_5874),
.B2(n_5822),
.Y(n_7971)
);

OAI22xp5_ASAP7_75t_L g7972 ( 
.A1(n_6452),
.A2(n_5274),
.B1(n_5286),
.B2(n_5266),
.Y(n_7972)
);

INVx1_ASAP7_75t_L g7973 ( 
.A(n_6390),
.Y(n_7973)
);

A2O1A1Ixp33_ASAP7_75t_L g7974 ( 
.A1(n_7040),
.A2(n_5282),
.B(n_5544),
.C(n_5517),
.Y(n_7974)
);

AND2x4_ASAP7_75t_L g7975 ( 
.A(n_6569),
.B(n_5394),
.Y(n_7975)
);

OAI21x1_ASAP7_75t_L g7976 ( 
.A1(n_6175),
.A2(n_5565),
.B(n_5447),
.Y(n_7976)
);

OAI21x1_ASAP7_75t_SL g7977 ( 
.A1(n_6156),
.A2(n_5989),
.B(n_5958),
.Y(n_7977)
);

A2O1A1Ixp33_ASAP7_75t_L g7978 ( 
.A1(n_7040),
.A2(n_5544),
.B(n_5517),
.C(n_5112),
.Y(n_7978)
);

BUFx3_ASAP7_75t_L g7979 ( 
.A(n_6273),
.Y(n_7979)
);

INVx1_ASAP7_75t_L g7980 ( 
.A(n_6390),
.Y(n_7980)
);

BUFx2_ASAP7_75t_L g7981 ( 
.A(n_6266),
.Y(n_7981)
);

AOI22xp33_ASAP7_75t_L g7982 ( 
.A1(n_7115),
.A2(n_4621),
.B1(n_4753),
.B2(n_4501),
.Y(n_7982)
);

BUFx2_ASAP7_75t_L g7983 ( 
.A(n_6266),
.Y(n_7983)
);

AO31x2_ASAP7_75t_L g7984 ( 
.A1(n_6497),
.A2(n_5728),
.A3(n_5742),
.B(n_5716),
.Y(n_7984)
);

BUFx12f_ASAP7_75t_L g7985 ( 
.A(n_6380),
.Y(n_7985)
);

O2A1O1Ixp33_ASAP7_75t_L g7986 ( 
.A1(n_6183),
.A2(n_5907),
.B(n_6122),
.C(n_6121),
.Y(n_7986)
);

BUFx3_ASAP7_75t_L g7987 ( 
.A(n_6273),
.Y(n_7987)
);

AO21x2_ASAP7_75t_L g7988 ( 
.A1(n_7019),
.A2(n_6110),
.B(n_6105),
.Y(n_7988)
);

AO31x2_ASAP7_75t_L g7989 ( 
.A1(n_6665),
.A2(n_5743),
.A3(n_5754),
.B(n_5742),
.Y(n_7989)
);

AND2x2_ASAP7_75t_L g7990 ( 
.A(n_7038),
.B(n_5279),
.Y(n_7990)
);

AO31x2_ASAP7_75t_L g7991 ( 
.A1(n_6665),
.A2(n_5754),
.A3(n_5764),
.B(n_5743),
.Y(n_7991)
);

NAND2xp5_ASAP7_75t_L g7992 ( 
.A(n_7058),
.B(n_5907),
.Y(n_7992)
);

AOI221xp5_ASAP7_75t_L g7993 ( 
.A1(n_6129),
.A2(n_6122),
.B1(n_6127),
.B2(n_6121),
.C(n_5499),
.Y(n_7993)
);

NAND2xp5_ASAP7_75t_L g7994 ( 
.A(n_7058),
.B(n_5648),
.Y(n_7994)
);

NOR2xp33_ASAP7_75t_L g7995 ( 
.A(n_7135),
.B(n_4719),
.Y(n_7995)
);

BUFx3_ASAP7_75t_L g7996 ( 
.A(n_6273),
.Y(n_7996)
);

NAND2xp5_ASAP7_75t_L g7997 ( 
.A(n_7084),
.B(n_5648),
.Y(n_7997)
);

INVx2_ASAP7_75t_L g7998 ( 
.A(n_6301),
.Y(n_7998)
);

OAI22xp5_ASAP7_75t_L g7999 ( 
.A1(n_7052),
.A2(n_5286),
.B1(n_5318),
.B2(n_5274),
.Y(n_7999)
);

AO21x2_ASAP7_75t_L g8000 ( 
.A1(n_7022),
.A2(n_7072),
.B(n_7075),
.Y(n_8000)
);

BUFx8_ASAP7_75t_L g8001 ( 
.A(n_6434),
.Y(n_8001)
);

BUFx6f_ASAP7_75t_L g8002 ( 
.A(n_6149),
.Y(n_8002)
);

BUFx4f_ASAP7_75t_L g8003 ( 
.A(n_6185),
.Y(n_8003)
);

INVx1_ASAP7_75t_L g8004 ( 
.A(n_6390),
.Y(n_8004)
);

AO21x2_ASAP7_75t_L g8005 ( 
.A1(n_7022),
.A2(n_5553),
.B(n_5552),
.Y(n_8005)
);

INVx6_ASAP7_75t_L g8006 ( 
.A(n_6422),
.Y(n_8006)
);

OA21x2_ASAP7_75t_L g8007 ( 
.A1(n_6605),
.A2(n_5567),
.B(n_5553),
.Y(n_8007)
);

OAI21x1_ASAP7_75t_L g8008 ( 
.A1(n_6140),
.A2(n_6159),
.B(n_6147),
.Y(n_8008)
);

OAI21x1_ASAP7_75t_SL g8009 ( 
.A1(n_6153),
.A2(n_5989),
.B(n_5958),
.Y(n_8009)
);

INVx2_ASAP7_75t_L g8010 ( 
.A(n_6318),
.Y(n_8010)
);

HB1xp67_ASAP7_75t_L g8011 ( 
.A(n_6133),
.Y(n_8011)
);

BUFx2_ASAP7_75t_L g8012 ( 
.A(n_6266),
.Y(n_8012)
);

OA21x2_ASAP7_75t_L g8013 ( 
.A1(n_6818),
.A2(n_5567),
.B(n_5553),
.Y(n_8013)
);

INVx5_ASAP7_75t_L g8014 ( 
.A(n_6920),
.Y(n_8014)
);

NAND2xp5_ASAP7_75t_L g8015 ( 
.A(n_7084),
.B(n_5648),
.Y(n_8015)
);

AOI22xp5_ASAP7_75t_L g8016 ( 
.A1(n_6293),
.A2(n_4621),
.B1(n_4753),
.B2(n_4501),
.Y(n_8016)
);

OA21x2_ASAP7_75t_L g8017 ( 
.A1(n_6818),
.A2(n_6768),
.B(n_6756),
.Y(n_8017)
);

OAI22xp33_ASAP7_75t_L g8018 ( 
.A1(n_7052),
.A2(n_5822),
.B1(n_5874),
.B2(n_5760),
.Y(n_8018)
);

NAND2xp5_ASAP7_75t_SL g8019 ( 
.A(n_7001),
.B(n_6036),
.Y(n_8019)
);

AOI21x1_ASAP7_75t_L g8020 ( 
.A1(n_6981),
.A2(n_5305),
.B(n_5185),
.Y(n_8020)
);

NOR2xp33_ASAP7_75t_L g8021 ( 
.A(n_6586),
.B(n_4735),
.Y(n_8021)
);

OA21x2_ASAP7_75t_L g8022 ( 
.A1(n_6791),
.A2(n_5573),
.B(n_5567),
.Y(n_8022)
);

AND2x4_ASAP7_75t_SL g8023 ( 
.A(n_6422),
.B(n_5765),
.Y(n_8023)
);

NOR2xp33_ASAP7_75t_L g8024 ( 
.A(n_6586),
.B(n_4812),
.Y(n_8024)
);

OA21x2_ASAP7_75t_L g8025 ( 
.A1(n_6791),
.A2(n_5579),
.B(n_5573),
.Y(n_8025)
);

OA21x2_ASAP7_75t_L g8026 ( 
.A1(n_6807),
.A2(n_5579),
.B(n_5573),
.Y(n_8026)
);

AND2x2_ASAP7_75t_L g8027 ( 
.A(n_7091),
.B(n_6178),
.Y(n_8027)
);

AND2x2_ASAP7_75t_L g8028 ( 
.A(n_7091),
.B(n_5279),
.Y(n_8028)
);

CKINVDCx5p33_ASAP7_75t_R g8029 ( 
.A(n_6893),
.Y(n_8029)
);

AOI21x1_ASAP7_75t_L g8030 ( 
.A1(n_6981),
.A2(n_5305),
.B(n_5185),
.Y(n_8030)
);

OAI21x1_ASAP7_75t_L g8031 ( 
.A1(n_6159),
.A2(n_4637),
.B(n_5419),
.Y(n_8031)
);

AOI21xp5_ASAP7_75t_L g8032 ( 
.A1(n_7143),
.A2(n_5773),
.B(n_5770),
.Y(n_8032)
);

OAI21x1_ASAP7_75t_SL g8033 ( 
.A1(n_6230),
.A2(n_5989),
.B(n_5958),
.Y(n_8033)
);

CKINVDCx16_ASAP7_75t_R g8034 ( 
.A(n_6815),
.Y(n_8034)
);

AO21x1_ASAP7_75t_L g8035 ( 
.A1(n_7075),
.A2(n_6127),
.B(n_4641),
.Y(n_8035)
);

OAI21x1_ASAP7_75t_L g8036 ( 
.A1(n_6161),
.A2(n_4637),
.B(n_5419),
.Y(n_8036)
);

AO21x2_ASAP7_75t_L g8037 ( 
.A1(n_6318),
.A2(n_5583),
.B(n_5582),
.Y(n_8037)
);

INVx2_ASAP7_75t_L g8038 ( 
.A(n_6318),
.Y(n_8038)
);

AOI21xp5_ASAP7_75t_SL g8039 ( 
.A1(n_6245),
.A2(n_5924),
.B(n_5915),
.Y(n_8039)
);

NOR2xp33_ASAP7_75t_L g8040 ( 
.A(n_6592),
.B(n_4812),
.Y(n_8040)
);

AO21x2_ASAP7_75t_L g8041 ( 
.A1(n_6318),
.A2(n_6110),
.B(n_6105),
.Y(n_8041)
);

CKINVDCx11_ASAP7_75t_R g8042 ( 
.A(n_6428),
.Y(n_8042)
);

AOI21xp5_ASAP7_75t_L g8043 ( 
.A1(n_7143),
.A2(n_5773),
.B(n_5770),
.Y(n_8043)
);

OAI21xp5_ASAP7_75t_L g8044 ( 
.A1(n_6514),
.A2(n_5358),
.B(n_5318),
.Y(n_8044)
);

AOI22xp33_ASAP7_75t_L g8045 ( 
.A1(n_6466),
.A2(n_4753),
.B1(n_4801),
.B2(n_4501),
.Y(n_8045)
);

AO31x2_ASAP7_75t_L g8046 ( 
.A1(n_6652),
.A2(n_5768),
.A3(n_5778),
.B(n_5764),
.Y(n_8046)
);

HB1xp67_ASAP7_75t_L g8047 ( 
.A(n_6133),
.Y(n_8047)
);

OR2x2_ASAP7_75t_L g8048 ( 
.A(n_6807),
.B(n_6810),
.Y(n_8048)
);

AO21x2_ASAP7_75t_L g8049 ( 
.A1(n_6321),
.A2(n_6115),
.B(n_6113),
.Y(n_8049)
);

NAND2xp5_ASAP7_75t_L g8050 ( 
.A(n_6934),
.B(n_6945),
.Y(n_8050)
);

AND2x4_ASAP7_75t_SL g8051 ( 
.A(n_6422),
.B(n_5770),
.Y(n_8051)
);

CKINVDCx9p33_ASAP7_75t_R g8052 ( 
.A(n_6782),
.Y(n_8052)
);

AO31x2_ASAP7_75t_L g8053 ( 
.A1(n_6652),
.A2(n_5778),
.A3(n_5779),
.B(n_5768),
.Y(n_8053)
);

NAND2xp5_ASAP7_75t_L g8054 ( 
.A(n_6934),
.B(n_5648),
.Y(n_8054)
);

INVx2_ASAP7_75t_SL g8055 ( 
.A(n_6766),
.Y(n_8055)
);

NAND2xp5_ASAP7_75t_L g8056 ( 
.A(n_6945),
.B(n_5648),
.Y(n_8056)
);

INVx2_ASAP7_75t_L g8057 ( 
.A(n_6321),
.Y(n_8057)
);

HB1xp67_ASAP7_75t_L g8058 ( 
.A(n_6176),
.Y(n_8058)
);

INVxp67_ASAP7_75t_L g8059 ( 
.A(n_6948),
.Y(n_8059)
);

NAND2xp5_ASAP7_75t_L g8060 ( 
.A(n_6948),
.B(n_5648),
.Y(n_8060)
);

AOI21xp5_ASAP7_75t_L g8061 ( 
.A1(n_7148),
.A2(n_5773),
.B(n_5770),
.Y(n_8061)
);

NAND2xp5_ASAP7_75t_L g8062 ( 
.A(n_6972),
.B(n_5648),
.Y(n_8062)
);

OAI21x1_ASAP7_75t_L g8063 ( 
.A1(n_6200),
.A2(n_6227),
.B(n_6208),
.Y(n_8063)
);

AND2x4_ASAP7_75t_L g8064 ( 
.A(n_6569),
.B(n_5394),
.Y(n_8064)
);

HB1xp67_ASAP7_75t_L g8065 ( 
.A(n_6176),
.Y(n_8065)
);

BUFx3_ASAP7_75t_L g8066 ( 
.A(n_6871),
.Y(n_8066)
);

OAI21x1_ASAP7_75t_SL g8067 ( 
.A1(n_6153),
.A2(n_5989),
.B(n_5958),
.Y(n_8067)
);

INVx1_ASAP7_75t_L g8068 ( 
.A(n_6397),
.Y(n_8068)
);

OAI21xp5_ASAP7_75t_L g8069 ( 
.A1(n_6982),
.A2(n_5363),
.B(n_5358),
.Y(n_8069)
);

HB1xp67_ASAP7_75t_L g8070 ( 
.A(n_6231),
.Y(n_8070)
);

NOR2xp33_ASAP7_75t_L g8071 ( 
.A(n_6592),
.B(n_5026),
.Y(n_8071)
);

AOI21xp5_ASAP7_75t_L g8072 ( 
.A1(n_7148),
.A2(n_5773),
.B(n_5770),
.Y(n_8072)
);

AOI21xp5_ASAP7_75t_L g8073 ( 
.A1(n_6835),
.A2(n_5794),
.B(n_5773),
.Y(n_8073)
);

INVx1_ASAP7_75t_L g8074 ( 
.A(n_6397),
.Y(n_8074)
);

BUFx2_ASAP7_75t_L g8075 ( 
.A(n_6871),
.Y(n_8075)
);

OAI21x1_ASAP7_75t_L g8076 ( 
.A1(n_6200),
.A2(n_6120),
.B(n_6090),
.Y(n_8076)
);

HB1xp67_ASAP7_75t_L g8077 ( 
.A(n_6231),
.Y(n_8077)
);

INVx1_ASAP7_75t_L g8078 ( 
.A(n_6397),
.Y(n_8078)
);

INVx1_ASAP7_75t_L g8079 ( 
.A(n_6404),
.Y(n_8079)
);

OAI22xp33_ASAP7_75t_L g8080 ( 
.A1(n_7052),
.A2(n_5822),
.B1(n_5874),
.B2(n_5760),
.Y(n_8080)
);

BUFx12f_ASAP7_75t_L g8081 ( 
.A(n_6394),
.Y(n_8081)
);

CKINVDCx5p33_ASAP7_75t_R g8082 ( 
.A(n_6893),
.Y(n_8082)
);

AND2x2_ASAP7_75t_L g8083 ( 
.A(n_7091),
.B(n_5288),
.Y(n_8083)
);

INVx1_ASAP7_75t_L g8084 ( 
.A(n_6404),
.Y(n_8084)
);

INVx1_ASAP7_75t_L g8085 ( 
.A(n_6404),
.Y(n_8085)
);

AOI22xp5_ASAP7_75t_L g8086 ( 
.A1(n_6293),
.A2(n_4801),
.B1(n_4901),
.B2(n_4753),
.Y(n_8086)
);

INVx1_ASAP7_75t_L g8087 ( 
.A(n_6415),
.Y(n_8087)
);

BUFx2_ASAP7_75t_R g8088 ( 
.A(n_6154),
.Y(n_8088)
);

INVx1_ASAP7_75t_L g8089 ( 
.A(n_6415),
.Y(n_8089)
);

AOI22xp33_ASAP7_75t_L g8090 ( 
.A1(n_6466),
.A2(n_4801),
.B1(n_4901),
.B2(n_4753),
.Y(n_8090)
);

OAI21x1_ASAP7_75t_L g8091 ( 
.A1(n_6200),
.A2(n_6120),
.B(n_6090),
.Y(n_8091)
);

OAI21x1_ASAP7_75t_L g8092 ( 
.A1(n_6208),
.A2(n_6235),
.B(n_6227),
.Y(n_8092)
);

OAI21xp5_ASAP7_75t_L g8093 ( 
.A1(n_6982),
.A2(n_5380),
.B(n_5363),
.Y(n_8093)
);

OAI21x1_ASAP7_75t_L g8094 ( 
.A1(n_6208),
.A2(n_5583),
.B(n_5582),
.Y(n_8094)
);

OAI21x1_ASAP7_75t_L g8095 ( 
.A1(n_6208),
.A2(n_5583),
.B(n_5582),
.Y(n_8095)
);

INVx3_ASAP7_75t_L g8096 ( 
.A(n_6578),
.Y(n_8096)
);

OR2x6_ASAP7_75t_L g8097 ( 
.A(n_6222),
.B(n_5822),
.Y(n_8097)
);

OAI21xp5_ASAP7_75t_L g8098 ( 
.A1(n_6314),
.A2(n_5413),
.B(n_5380),
.Y(n_8098)
);

OR2x2_ASAP7_75t_L g8099 ( 
.A(n_6810),
.B(n_5476),
.Y(n_8099)
);

OAI22xp5_ASAP7_75t_L g8100 ( 
.A1(n_6558),
.A2(n_5413),
.B1(n_5465),
.B2(n_5412),
.Y(n_8100)
);

INVx1_ASAP7_75t_L g8101 ( 
.A(n_6415),
.Y(n_8101)
);

INVx2_ASAP7_75t_L g8102 ( 
.A(n_6321),
.Y(n_8102)
);

O2A1O1Ixp33_ASAP7_75t_SL g8103 ( 
.A1(n_7118),
.A2(n_5700),
.B(n_5808),
.C(n_5600),
.Y(n_8103)
);

A2O1A1Ixp33_ASAP7_75t_L g8104 ( 
.A1(n_6748),
.A2(n_5112),
.B(n_5160),
.C(n_5144),
.Y(n_8104)
);

NAND2xp5_ASAP7_75t_L g8105 ( 
.A(n_6972),
.B(n_5587),
.Y(n_8105)
);

INVx1_ASAP7_75t_L g8106 ( 
.A(n_6416),
.Y(n_8106)
);

CKINVDCx6p67_ASAP7_75t_R g8107 ( 
.A(n_6185),
.Y(n_8107)
);

INVx1_ASAP7_75t_L g8108 ( 
.A(n_6416),
.Y(n_8108)
);

A2O1A1Ixp33_ASAP7_75t_L g8109 ( 
.A1(n_6748),
.A2(n_5112),
.B(n_5160),
.C(n_5144),
.Y(n_8109)
);

NAND2xp33_ASAP7_75t_R g8110 ( 
.A(n_6394),
.B(n_6050),
.Y(n_8110)
);

NAND2xp5_ASAP7_75t_L g8111 ( 
.A(n_6984),
.B(n_5587),
.Y(n_8111)
);

OAI21xp5_ASAP7_75t_L g8112 ( 
.A1(n_6314),
.A2(n_6068),
.B(n_6036),
.Y(n_8112)
);

INVx1_ASAP7_75t_L g8113 ( 
.A(n_6416),
.Y(n_8113)
);

OAI21x1_ASAP7_75t_SL g8114 ( 
.A1(n_6153),
.A2(n_6041),
.B(n_6029),
.Y(n_8114)
);

O2A1O1Ixp33_ASAP7_75t_SL g8115 ( 
.A1(n_6815),
.A2(n_5700),
.B(n_5808),
.C(n_5600),
.Y(n_8115)
);

NAND2xp5_ASAP7_75t_L g8116 ( 
.A(n_6984),
.B(n_5587),
.Y(n_8116)
);

AOI21xp5_ASAP7_75t_L g8117 ( 
.A1(n_6835),
.A2(n_5823),
.B(n_5794),
.Y(n_8117)
);

NAND2xp5_ASAP7_75t_L g8118 ( 
.A(n_7003),
.B(n_5779),
.Y(n_8118)
);

INVx1_ASAP7_75t_L g8119 ( 
.A(n_6420),
.Y(n_8119)
);

OAI21xp5_ASAP7_75t_L g8120 ( 
.A1(n_6489),
.A2(n_6754),
.B(n_6740),
.Y(n_8120)
);

OR2x6_ASAP7_75t_L g8121 ( 
.A(n_6402),
.B(n_5874),
.Y(n_8121)
);

AOI22xp33_ASAP7_75t_L g8122 ( 
.A1(n_6792),
.A2(n_4801),
.B1(n_4901),
.B2(n_4753),
.Y(n_8122)
);

OA21x2_ASAP7_75t_L g8123 ( 
.A1(n_6854),
.A2(n_5609),
.B(n_5604),
.Y(n_8123)
);

AND2x2_ASAP7_75t_L g8124 ( 
.A(n_6178),
.B(n_5288),
.Y(n_8124)
);

BUFx6f_ASAP7_75t_L g8125 ( 
.A(n_6149),
.Y(n_8125)
);

AND2x4_ASAP7_75t_L g8126 ( 
.A(n_6578),
.B(n_5394),
.Y(n_8126)
);

AO31x2_ASAP7_75t_L g8127 ( 
.A1(n_6738),
.A2(n_5788),
.A3(n_5792),
.B(n_5784),
.Y(n_8127)
);

INVx1_ASAP7_75t_L g8128 ( 
.A(n_6420),
.Y(n_8128)
);

INVx1_ASAP7_75t_L g8129 ( 
.A(n_6420),
.Y(n_8129)
);

BUFx3_ASAP7_75t_L g8130 ( 
.A(n_6871),
.Y(n_8130)
);

NAND2xp5_ASAP7_75t_L g8131 ( 
.A(n_7003),
.B(n_6660),
.Y(n_8131)
);

AOI22xp33_ASAP7_75t_L g8132 ( 
.A1(n_6792),
.A2(n_4801),
.B1(n_4901),
.B2(n_4753),
.Y(n_8132)
);

INVx1_ASAP7_75t_L g8133 ( 
.A(n_6421),
.Y(n_8133)
);

INVx4_ASAP7_75t_L g8134 ( 
.A(n_6434),
.Y(n_8134)
);

INVx1_ASAP7_75t_L g8135 ( 
.A(n_6421),
.Y(n_8135)
);

AND2x2_ASAP7_75t_L g8136 ( 
.A(n_6178),
.B(n_6184),
.Y(n_8136)
);

OAI21xp5_ASAP7_75t_L g8137 ( 
.A1(n_6754),
.A2(n_6083),
.B(n_6068),
.Y(n_8137)
);

INVx2_ASAP7_75t_L g8138 ( 
.A(n_6321),
.Y(n_8138)
);

INVx6_ASAP7_75t_L g8139 ( 
.A(n_6422),
.Y(n_8139)
);

HB1xp67_ASAP7_75t_L g8140 ( 
.A(n_6239),
.Y(n_8140)
);

OA21x2_ASAP7_75t_L g8141 ( 
.A1(n_6854),
.A2(n_5686),
.B(n_5669),
.Y(n_8141)
);

BUFx8_ASAP7_75t_L g8142 ( 
.A(n_6434),
.Y(n_8142)
);

OAI21xp5_ASAP7_75t_L g8143 ( 
.A1(n_6740),
.A2(n_6112),
.B(n_6083),
.Y(n_8143)
);

AND2x2_ASAP7_75t_L g8144 ( 
.A(n_6184),
.B(n_5288),
.Y(n_8144)
);

INVx2_ASAP7_75t_L g8145 ( 
.A(n_6324),
.Y(n_8145)
);

OAI21x1_ASAP7_75t_L g8146 ( 
.A1(n_6254),
.A2(n_6276),
.B(n_6265),
.Y(n_8146)
);

OAI21xp5_ASAP7_75t_L g8147 ( 
.A1(n_7017),
.A2(n_6112),
.B(n_6058),
.Y(n_8147)
);

AO31x2_ASAP7_75t_L g8148 ( 
.A1(n_6738),
.A2(n_6565),
.A3(n_6396),
.B(n_6936),
.Y(n_8148)
);

AND2x2_ASAP7_75t_L g8149 ( 
.A(n_6184),
.B(n_5307),
.Y(n_8149)
);

INVx1_ASAP7_75t_L g8150 ( 
.A(n_6421),
.Y(n_8150)
);

AND2x4_ASAP7_75t_L g8151 ( 
.A(n_6578),
.B(n_5399),
.Y(n_8151)
);

INVxp67_ASAP7_75t_L g8152 ( 
.A(n_7076),
.Y(n_8152)
);

OR2x2_ASAP7_75t_L g8153 ( 
.A(n_6868),
.B(n_5476),
.Y(n_8153)
);

AO21x2_ASAP7_75t_L g8154 ( 
.A1(n_6324),
.A2(n_5692),
.B(n_5686),
.Y(n_8154)
);

BUFx3_ASAP7_75t_L g8155 ( 
.A(n_6871),
.Y(n_8155)
);

BUFx4f_ASAP7_75t_L g8156 ( 
.A(n_6412),
.Y(n_8156)
);

AOI21x1_ASAP7_75t_L g8157 ( 
.A1(n_6549),
.A2(n_6606),
.B(n_6557),
.Y(n_8157)
);

INVx1_ASAP7_75t_L g8158 ( 
.A(n_6447),
.Y(n_8158)
);

BUFx2_ASAP7_75t_L g8159 ( 
.A(n_6882),
.Y(n_8159)
);

INVx1_ASAP7_75t_L g8160 ( 
.A(n_6447),
.Y(n_8160)
);

AOI22xp33_ASAP7_75t_L g8161 ( 
.A1(n_6792),
.A2(n_6761),
.B1(n_6752),
.B2(n_6780),
.Y(n_8161)
);

OAI21xp5_ASAP7_75t_L g8162 ( 
.A1(n_7017),
.A2(n_6058),
.B(n_6050),
.Y(n_8162)
);

NAND2x1p5_ASAP7_75t_L g8163 ( 
.A(n_6412),
.B(n_4809),
.Y(n_8163)
);

AND2x4_ASAP7_75t_L g8164 ( 
.A(n_6578),
.B(n_5399),
.Y(n_8164)
);

INVx2_ASAP7_75t_L g8165 ( 
.A(n_6324),
.Y(n_8165)
);

AOI22xp5_ASAP7_75t_L g8166 ( 
.A1(n_6558),
.A2(n_4901),
.B1(n_4911),
.B2(n_4801),
.Y(n_8166)
);

INVx2_ASAP7_75t_L g8167 ( 
.A(n_6324),
.Y(n_8167)
);

OAI222xp33_ASAP7_75t_L g8168 ( 
.A1(n_6580),
.A2(n_5882),
.B1(n_5874),
.B2(n_5047),
.C1(n_4801),
.C2(n_4911),
.Y(n_8168)
);

OR2x6_ASAP7_75t_L g8169 ( 
.A(n_6402),
.B(n_5882),
.Y(n_8169)
);

BUFx6f_ASAP7_75t_L g8170 ( 
.A(n_6149),
.Y(n_8170)
);

NOR2xp33_ASAP7_75t_SL g8171 ( 
.A(n_6724),
.B(n_5399),
.Y(n_8171)
);

INVx2_ASAP7_75t_L g8172 ( 
.A(n_6337),
.Y(n_8172)
);

INVxp67_ASAP7_75t_L g8173 ( 
.A(n_7076),
.Y(n_8173)
);

OR2x2_ASAP7_75t_L g8174 ( 
.A(n_6868),
.B(n_5476),
.Y(n_8174)
);

OR2x2_ASAP7_75t_L g8175 ( 
.A(n_6869),
.B(n_5412),
.Y(n_8175)
);

INVx1_ASAP7_75t_L g8176 ( 
.A(n_6447),
.Y(n_8176)
);

INVx1_ASAP7_75t_L g8177 ( 
.A(n_6456),
.Y(n_8177)
);

INVx2_ASAP7_75t_SL g8178 ( 
.A(n_6766),
.Y(n_8178)
);

AND2x2_ASAP7_75t_L g8179 ( 
.A(n_6189),
.B(n_5307),
.Y(n_8179)
);

HB1xp67_ASAP7_75t_L g8180 ( 
.A(n_6239),
.Y(n_8180)
);

INVx3_ASAP7_75t_L g8181 ( 
.A(n_6585),
.Y(n_8181)
);

INVx4_ASAP7_75t_SL g8182 ( 
.A(n_6753),
.Y(n_8182)
);

AND2x4_ASAP7_75t_SL g8183 ( 
.A(n_6422),
.B(n_5794),
.Y(n_8183)
);

OAI22xp5_ASAP7_75t_L g8184 ( 
.A1(n_6580),
.A2(n_5465),
.B1(n_5412),
.B2(n_5128),
.Y(n_8184)
);

OR2x6_ASAP7_75t_L g8185 ( 
.A(n_6402),
.B(n_5882),
.Y(n_8185)
);

OAI22xp5_ASAP7_75t_L g8186 ( 
.A1(n_6946),
.A2(n_5465),
.B1(n_5128),
.B2(n_5182),
.Y(n_8186)
);

AOI21xp5_ASAP7_75t_L g8187 ( 
.A1(n_6407),
.A2(n_5823),
.B(n_5794),
.Y(n_8187)
);

INVx2_ASAP7_75t_L g8188 ( 
.A(n_6337),
.Y(n_8188)
);

NOR2xp33_ASAP7_75t_L g8189 ( 
.A(n_6865),
.B(n_6077),
.Y(n_8189)
);

INVx1_ASAP7_75t_L g8190 ( 
.A(n_6456),
.Y(n_8190)
);

INVx2_ASAP7_75t_SL g8191 ( 
.A(n_6766),
.Y(n_8191)
);

OR2x2_ASAP7_75t_L g8192 ( 
.A(n_6869),
.B(n_5468),
.Y(n_8192)
);

INVx2_ASAP7_75t_L g8193 ( 
.A(n_6337),
.Y(n_8193)
);

OR2x2_ASAP7_75t_L g8194 ( 
.A(n_6701),
.B(n_5468),
.Y(n_8194)
);

AOI21xp5_ASAP7_75t_L g8195 ( 
.A1(n_6407),
.A2(n_5823),
.B(n_5794),
.Y(n_8195)
);

INVx2_ASAP7_75t_SL g8196 ( 
.A(n_6882),
.Y(n_8196)
);

AND2x4_ASAP7_75t_L g8197 ( 
.A(n_6585),
.B(n_5399),
.Y(n_8197)
);

AND2x4_ASAP7_75t_L g8198 ( 
.A(n_6585),
.B(n_5399),
.Y(n_8198)
);

AOI21xp5_ASAP7_75t_L g8199 ( 
.A1(n_6453),
.A2(n_5826),
.B(n_5823),
.Y(n_8199)
);

INVx3_ASAP7_75t_L g8200 ( 
.A(n_6585),
.Y(n_8200)
);

AOI22xp33_ASAP7_75t_L g8201 ( 
.A1(n_6752),
.A2(n_4901),
.B1(n_4911),
.B2(n_4801),
.Y(n_8201)
);

AO21x2_ASAP7_75t_L g8202 ( 
.A1(n_6337),
.A2(n_5725),
.B(n_5706),
.Y(n_8202)
);

INVx3_ASAP7_75t_L g8203 ( 
.A(n_6598),
.Y(n_8203)
);

INVx1_ASAP7_75t_L g8204 ( 
.A(n_6456),
.Y(n_8204)
);

INVx2_ASAP7_75t_L g8205 ( 
.A(n_6341),
.Y(n_8205)
);

INVx3_ASAP7_75t_L g8206 ( 
.A(n_6598),
.Y(n_8206)
);

CKINVDCx5p33_ASAP7_75t_R g8207 ( 
.A(n_6911),
.Y(n_8207)
);

INVx2_ASAP7_75t_L g8208 ( 
.A(n_6341),
.Y(n_8208)
);

OA21x2_ASAP7_75t_L g8209 ( 
.A1(n_6831),
.A2(n_5725),
.B(n_5706),
.Y(n_8209)
);

AOI22xp33_ASAP7_75t_L g8210 ( 
.A1(n_6761),
.A2(n_4911),
.B1(n_5047),
.B2(n_4901),
.Y(n_8210)
);

AO31x2_ASAP7_75t_L g8211 ( 
.A1(n_6565),
.A2(n_5788),
.A3(n_5792),
.B(n_5784),
.Y(n_8211)
);

INVx2_ASAP7_75t_L g8212 ( 
.A(n_6341),
.Y(n_8212)
);

OAI22xp5_ASAP7_75t_L g8213 ( 
.A1(n_6946),
.A2(n_5128),
.B1(n_5182),
.B2(n_5107),
.Y(n_8213)
);

INVx1_ASAP7_75t_L g8214 ( 
.A(n_6460),
.Y(n_8214)
);

AO21x2_ASAP7_75t_L g8215 ( 
.A1(n_6341),
.A2(n_5761),
.B(n_5756),
.Y(n_8215)
);

NAND2xp5_ASAP7_75t_L g8216 ( 
.A(n_6660),
.B(n_6087),
.Y(n_8216)
);

INVx1_ASAP7_75t_L g8217 ( 
.A(n_6460),
.Y(n_8217)
);

AOI22xp5_ASAP7_75t_L g8218 ( 
.A1(n_6724),
.A2(n_4911),
.B1(n_5047),
.B2(n_4901),
.Y(n_8218)
);

INVx1_ASAP7_75t_L g8219 ( 
.A(n_6460),
.Y(n_8219)
);

INVx2_ASAP7_75t_L g8220 ( 
.A(n_6357),
.Y(n_8220)
);

NOR2xp33_ASAP7_75t_L g8221 ( 
.A(n_7090),
.B(n_6077),
.Y(n_8221)
);

CKINVDCx11_ASAP7_75t_R g8222 ( 
.A(n_6428),
.Y(n_8222)
);

OR2x2_ASAP7_75t_L g8223 ( 
.A(n_6701),
.B(n_5498),
.Y(n_8223)
);

OA21x2_ASAP7_75t_L g8224 ( 
.A1(n_6831),
.A2(n_5761),
.B(n_5756),
.Y(n_8224)
);

INVx1_ASAP7_75t_L g8225 ( 
.A(n_6467),
.Y(n_8225)
);

O2A1O1Ixp33_ASAP7_75t_SL g8226 ( 
.A1(n_6221),
.A2(n_5926),
.B(n_5939),
.C(n_5893),
.Y(n_8226)
);

OAI21xp5_ASAP7_75t_L g8227 ( 
.A1(n_6641),
.A2(n_5926),
.B(n_5893),
.Y(n_8227)
);

HB1xp67_ASAP7_75t_L g8228 ( 
.A(n_6279),
.Y(n_8228)
);

OA21x2_ASAP7_75t_L g8229 ( 
.A1(n_7044),
.A2(n_5763),
.B(n_5756),
.Y(n_8229)
);

NOR2xp33_ASAP7_75t_L g8230 ( 
.A(n_7090),
.B(n_4879),
.Y(n_8230)
);

A2O1A1Ixp33_ASAP7_75t_L g8231 ( 
.A1(n_6882),
.A2(n_5112),
.B(n_5160),
.C(n_5144),
.Y(n_8231)
);

NAND2xp5_ASAP7_75t_L g8232 ( 
.A(n_6907),
.B(n_6117),
.Y(n_8232)
);

AND2x2_ASAP7_75t_L g8233 ( 
.A(n_6189),
.B(n_5307),
.Y(n_8233)
);

INVx1_ASAP7_75t_L g8234 ( 
.A(n_6467),
.Y(n_8234)
);

BUFx2_ASAP7_75t_L g8235 ( 
.A(n_6882),
.Y(n_8235)
);

OAI21xp5_ASAP7_75t_L g8236 ( 
.A1(n_6641),
.A2(n_5963),
.B(n_5939),
.Y(n_8236)
);

HB1xp67_ASAP7_75t_L g8237 ( 
.A(n_6279),
.Y(n_8237)
);

AOI21x1_ASAP7_75t_L g8238 ( 
.A1(n_6549),
.A2(n_5420),
.B(n_5336),
.Y(n_8238)
);

INVx1_ASAP7_75t_L g8239 ( 
.A(n_6467),
.Y(n_8239)
);

AO21x2_ASAP7_75t_L g8240 ( 
.A1(n_6357),
.A2(n_5774),
.B(n_5763),
.Y(n_8240)
);

INVx1_ASAP7_75t_L g8241 ( 
.A(n_6471),
.Y(n_8241)
);

INVx1_ASAP7_75t_L g8242 ( 
.A(n_6471),
.Y(n_8242)
);

BUFx12f_ASAP7_75t_L g8243 ( 
.A(n_6399),
.Y(n_8243)
);

AND2x4_ASAP7_75t_L g8244 ( 
.A(n_6598),
.B(n_5493),
.Y(n_8244)
);

INVx2_ASAP7_75t_SL g8245 ( 
.A(n_6903),
.Y(n_8245)
);

NAND2xp5_ASAP7_75t_L g8246 ( 
.A(n_6907),
.B(n_5798),
.Y(n_8246)
);

O2A1O1Ixp33_ASAP7_75t_SL g8247 ( 
.A1(n_6221),
.A2(n_5963),
.B(n_5456),
.C(n_5608),
.Y(n_8247)
);

INVx2_ASAP7_75t_L g8248 ( 
.A(n_6357),
.Y(n_8248)
);

AOI21xp5_ASAP7_75t_L g8249 ( 
.A1(n_6453),
.A2(n_5826),
.B(n_5823),
.Y(n_8249)
);

OR2x2_ASAP7_75t_L g8250 ( 
.A(n_6701),
.B(n_5498),
.Y(n_8250)
);

NAND2xp5_ASAP7_75t_L g8251 ( 
.A(n_6205),
.B(n_6087),
.Y(n_8251)
);

INVx1_ASAP7_75t_L g8252 ( 
.A(n_6471),
.Y(n_8252)
);

INVx1_ASAP7_75t_L g8253 ( 
.A(n_6472),
.Y(n_8253)
);

NAND2x1p5_ASAP7_75t_L g8254 ( 
.A(n_6412),
.B(n_4809),
.Y(n_8254)
);

BUFx8_ASAP7_75t_SL g8255 ( 
.A(n_6188),
.Y(n_8255)
);

CKINVDCx5p33_ASAP7_75t_R g8256 ( 
.A(n_6911),
.Y(n_8256)
);

NAND2xp5_ASAP7_75t_L g8257 ( 
.A(n_6205),
.B(n_6099),
.Y(n_8257)
);

NAND2xp5_ASAP7_75t_L g8258 ( 
.A(n_6333),
.B(n_6099),
.Y(n_8258)
);

NAND3xp33_ASAP7_75t_SL g8259 ( 
.A(n_6483),
.B(n_5702),
.C(n_5547),
.Y(n_8259)
);

AOI221xp5_ASAP7_75t_L g8260 ( 
.A1(n_7079),
.A2(n_5551),
.B1(n_5548),
.B2(n_5543),
.C(n_6107),
.Y(n_8260)
);

BUFx2_ASAP7_75t_L g8261 ( 
.A(n_6903),
.Y(n_8261)
);

INVx1_ASAP7_75t_L g8262 ( 
.A(n_6472),
.Y(n_8262)
);

BUFx3_ASAP7_75t_L g8263 ( 
.A(n_6903),
.Y(n_8263)
);

AO21x2_ASAP7_75t_L g8264 ( 
.A1(n_6357),
.A2(n_5816),
.B(n_5814),
.Y(n_8264)
);

AND2x2_ASAP7_75t_L g8265 ( 
.A(n_6189),
.B(n_5325),
.Y(n_8265)
);

OA21x2_ASAP7_75t_L g8266 ( 
.A1(n_7044),
.A2(n_5816),
.B(n_5814),
.Y(n_8266)
);

INVx1_ASAP7_75t_L g8267 ( 
.A(n_6472),
.Y(n_8267)
);

OR2x2_ASAP7_75t_L g8268 ( 
.A(n_6721),
.B(n_5526),
.Y(n_8268)
);

NAND2x1p5_ASAP7_75t_L g8269 ( 
.A(n_6170),
.B(n_4809),
.Y(n_8269)
);

HB1xp67_ASAP7_75t_L g8270 ( 
.A(n_6295),
.Y(n_8270)
);

INVx4_ASAP7_75t_L g8271 ( 
.A(n_6434),
.Y(n_8271)
);

INVx1_ASAP7_75t_L g8272 ( 
.A(n_6474),
.Y(n_8272)
);

NAND3xp33_ASAP7_75t_SL g8273 ( 
.A(n_6483),
.B(n_5702),
.C(n_5547),
.Y(n_8273)
);

NAND2x1p5_ASAP7_75t_L g8274 ( 
.A(n_6170),
.B(n_4809),
.Y(n_8274)
);

INVx2_ASAP7_75t_L g8275 ( 
.A(n_6369),
.Y(n_8275)
);

OA21x2_ASAP7_75t_L g8276 ( 
.A1(n_6549),
.A2(n_6606),
.B(n_6557),
.Y(n_8276)
);

INVx1_ASAP7_75t_L g8277 ( 
.A(n_6474),
.Y(n_8277)
);

AOI22xp33_ASAP7_75t_L g8278 ( 
.A1(n_6780),
.A2(n_5047),
.B1(n_4911),
.B2(n_5882),
.Y(n_8278)
);

INVx3_ASAP7_75t_L g8279 ( 
.A(n_6598),
.Y(n_8279)
);

INVx1_ASAP7_75t_L g8280 ( 
.A(n_6474),
.Y(n_8280)
);

AOI21xp5_ASAP7_75t_L g8281 ( 
.A1(n_6698),
.A2(n_5854),
.B(n_5826),
.Y(n_8281)
);

AOI21xp5_ASAP7_75t_L g8282 ( 
.A1(n_6698),
.A2(n_6739),
.B(n_6645),
.Y(n_8282)
);

A2O1A1Ixp33_ASAP7_75t_L g8283 ( 
.A1(n_6903),
.A2(n_5112),
.B(n_5160),
.C(n_5144),
.Y(n_8283)
);

INVx1_ASAP7_75t_SL g8284 ( 
.A(n_6470),
.Y(n_8284)
);

INVx1_ASAP7_75t_SL g8285 ( 
.A(n_6470),
.Y(n_8285)
);

NOR2xp33_ASAP7_75t_L g8286 ( 
.A(n_6151),
.B(n_4879),
.Y(n_8286)
);

NAND2xp5_ASAP7_75t_L g8287 ( 
.A(n_6333),
.B(n_5798),
.Y(n_8287)
);

AOI21xp5_ASAP7_75t_L g8288 ( 
.A1(n_6739),
.A2(n_5854),
.B(n_5826),
.Y(n_8288)
);

AOI21xp33_ASAP7_75t_SL g8289 ( 
.A1(n_6164),
.A2(n_4164),
.B(n_4159),
.Y(n_8289)
);

AND2x4_ASAP7_75t_L g8290 ( 
.A(n_6599),
.B(n_5493),
.Y(n_8290)
);

AND2x2_ASAP7_75t_L g8291 ( 
.A(n_6902),
.B(n_5325),
.Y(n_8291)
);

INVx1_ASAP7_75t_L g8292 ( 
.A(n_6477),
.Y(n_8292)
);

NOR2xp33_ASAP7_75t_L g8293 ( 
.A(n_6151),
.B(n_5526),
.Y(n_8293)
);

AOI22xp33_ASAP7_75t_L g8294 ( 
.A1(n_6795),
.A2(n_5047),
.B1(n_4911),
.B2(n_5882),
.Y(n_8294)
);

OA21x2_ASAP7_75t_L g8295 ( 
.A1(n_6557),
.A2(n_5845),
.B(n_5834),
.Y(n_8295)
);

AND2x4_ASAP7_75t_L g8296 ( 
.A(n_6599),
.B(n_5493),
.Y(n_8296)
);

OAI22xp5_ASAP7_75t_SL g8297 ( 
.A1(n_6360),
.A2(n_5608),
.B1(n_5456),
.B2(n_5897),
.Y(n_8297)
);

INVx2_ASAP7_75t_L g8298 ( 
.A(n_6369),
.Y(n_8298)
);

AO21x2_ASAP7_75t_L g8299 ( 
.A1(n_6369),
.A2(n_5850),
.B(n_5847),
.Y(n_8299)
);

NOR2xp33_ASAP7_75t_L g8300 ( 
.A(n_6162),
.B(n_5533),
.Y(n_8300)
);

AO21x2_ASAP7_75t_L g8301 ( 
.A1(n_6369),
.A2(n_6375),
.B(n_6373),
.Y(n_8301)
);

NOR2x1_ASAP7_75t_SL g8302 ( 
.A(n_6920),
.B(n_6029),
.Y(n_8302)
);

AND2x2_ASAP7_75t_L g8303 ( 
.A(n_6902),
.B(n_5325),
.Y(n_8303)
);

CKINVDCx14_ASAP7_75t_R g8304 ( 
.A(n_6615),
.Y(n_8304)
);

INVx2_ASAP7_75t_L g8305 ( 
.A(n_8295),
.Y(n_8305)
);

AOI22xp5_ASAP7_75t_SL g8306 ( 
.A1(n_7166),
.A2(n_6427),
.B1(n_6399),
.B2(n_6938),
.Y(n_8306)
);

INVx1_ASAP7_75t_L g8307 ( 
.A(n_7156),
.Y(n_8307)
);

INVx2_ASAP7_75t_L g8308 ( 
.A(n_8295),
.Y(n_8308)
);

BUFx8_ASAP7_75t_L g8309 ( 
.A(n_7283),
.Y(n_8309)
);

INVx1_ASAP7_75t_L g8310 ( 
.A(n_7156),
.Y(n_8310)
);

BUFx10_ASAP7_75t_L g8311 ( 
.A(n_7262),
.Y(n_8311)
);

OAI21xp5_ASAP7_75t_L g8312 ( 
.A1(n_7227),
.A2(n_6230),
.B(n_6156),
.Y(n_8312)
);

INVx1_ASAP7_75t_L g8313 ( 
.A(n_7189),
.Y(n_8313)
);

AO21x1_ASAP7_75t_L g8314 ( 
.A1(n_7194),
.A2(n_7049),
.B(n_6396),
.Y(n_8314)
);

OAI22xp33_ASAP7_75t_L g8315 ( 
.A1(n_7256),
.A2(n_6758),
.B1(n_6760),
.B2(n_6682),
.Y(n_8315)
);

AO21x1_ASAP7_75t_SL g8316 ( 
.A1(n_7259),
.A2(n_7577),
.B(n_7286),
.Y(n_8316)
);

OAI21xp5_ASAP7_75t_L g8317 ( 
.A1(n_7227),
.A2(n_6230),
.B(n_7097),
.Y(n_8317)
);

HB1xp67_ASAP7_75t_L g8318 ( 
.A(n_7176),
.Y(n_8318)
);

CKINVDCx5p33_ASAP7_75t_R g8319 ( 
.A(n_7245),
.Y(n_8319)
);

CKINVDCx20_ASAP7_75t_R g8320 ( 
.A(n_7375),
.Y(n_8320)
);

AOI22xp5_ASAP7_75t_L g8321 ( 
.A1(n_7166),
.A2(n_6722),
.B1(n_6993),
.B2(n_6493),
.Y(n_8321)
);

INVx2_ASAP7_75t_L g8322 ( 
.A(n_8295),
.Y(n_8322)
);

INVx2_ASAP7_75t_L g8323 ( 
.A(n_8295),
.Y(n_8323)
);

INVx1_ASAP7_75t_L g8324 ( 
.A(n_7189),
.Y(n_8324)
);

OAI21x1_ASAP7_75t_SL g8325 ( 
.A1(n_7604),
.A2(n_6395),
.B(n_6335),
.Y(n_8325)
);

INVx1_ASAP7_75t_L g8326 ( 
.A(n_7192),
.Y(n_8326)
);

BUFx6f_ASAP7_75t_L g8327 ( 
.A(n_7283),
.Y(n_8327)
);

INVx1_ASAP7_75t_L g8328 ( 
.A(n_7192),
.Y(n_8328)
);

BUFx8_ASAP7_75t_L g8329 ( 
.A(n_7283),
.Y(n_8329)
);

INVx1_ASAP7_75t_L g8330 ( 
.A(n_7204),
.Y(n_8330)
);

HB1xp67_ASAP7_75t_L g8331 ( 
.A(n_7176),
.Y(n_8331)
);

INVx1_ASAP7_75t_L g8332 ( 
.A(n_7204),
.Y(n_8332)
);

INVx2_ASAP7_75t_L g8333 ( 
.A(n_8295),
.Y(n_8333)
);

CKINVDCx16_ASAP7_75t_R g8334 ( 
.A(n_8034),
.Y(n_8334)
);

OAI22xp5_ASAP7_75t_L g8335 ( 
.A1(n_7515),
.A2(n_6870),
.B1(n_6715),
.B2(n_6845),
.Y(n_8335)
);

AOI22xp33_ASAP7_75t_L g8336 ( 
.A1(n_7394),
.A2(n_6417),
.B1(n_6795),
.B2(n_7014),
.Y(n_8336)
);

INVx3_ASAP7_75t_L g8337 ( 
.A(n_7182),
.Y(n_8337)
);

OAI21xp5_ASAP7_75t_L g8338 ( 
.A1(n_7604),
.A2(n_7097),
.B(n_7147),
.Y(n_8338)
);

OAI22xp5_ASAP7_75t_L g8339 ( 
.A1(n_7515),
.A2(n_6870),
.B1(n_6715),
.B2(n_6845),
.Y(n_8339)
);

BUFx8_ASAP7_75t_SL g8340 ( 
.A(n_7904),
.Y(n_8340)
);

BUFx3_ASAP7_75t_L g8341 ( 
.A(n_7842),
.Y(n_8341)
);

BUFx12f_ASAP7_75t_L g8342 ( 
.A(n_7245),
.Y(n_8342)
);

CKINVDCx6p67_ASAP7_75t_R g8343 ( 
.A(n_7283),
.Y(n_8343)
);

INVx3_ASAP7_75t_L g8344 ( 
.A(n_7182),
.Y(n_8344)
);

BUFx6f_ASAP7_75t_L g8345 ( 
.A(n_7339),
.Y(n_8345)
);

BUFx3_ASAP7_75t_L g8346 ( 
.A(n_7842),
.Y(n_8346)
);

OA21x2_ASAP7_75t_L g8347 ( 
.A1(n_7170),
.A2(n_6607),
.B(n_6606),
.Y(n_8347)
);

INVx1_ASAP7_75t_L g8348 ( 
.A(n_7208),
.Y(n_8348)
);

BUFx3_ASAP7_75t_L g8349 ( 
.A(n_7842),
.Y(n_8349)
);

BUFx3_ASAP7_75t_L g8350 ( 
.A(n_7842),
.Y(n_8350)
);

INVx1_ASAP7_75t_L g8351 ( 
.A(n_7208),
.Y(n_8351)
);

AOI21x1_ASAP7_75t_L g8352 ( 
.A1(n_7194),
.A2(n_6617),
.B(n_6607),
.Y(n_8352)
);

INVx1_ASAP7_75t_L g8353 ( 
.A(n_7214),
.Y(n_8353)
);

BUFx3_ASAP7_75t_L g8354 ( 
.A(n_7842),
.Y(n_8354)
);

CKINVDCx11_ASAP7_75t_R g8355 ( 
.A(n_7314),
.Y(n_8355)
);

INVx2_ASAP7_75t_L g8356 ( 
.A(n_8295),
.Y(n_8356)
);

AND2x2_ASAP7_75t_L g8357 ( 
.A(n_7712),
.B(n_6335),
.Y(n_8357)
);

AOI22xp33_ASAP7_75t_L g8358 ( 
.A1(n_7394),
.A2(n_6417),
.B1(n_7014),
.B2(n_6720),
.Y(n_8358)
);

INVx2_ASAP7_75t_L g8359 ( 
.A(n_7910),
.Y(n_8359)
);

INVx2_ASAP7_75t_L g8360 ( 
.A(n_7910),
.Y(n_8360)
);

AOI22xp33_ASAP7_75t_L g8361 ( 
.A1(n_7652),
.A2(n_7165),
.B1(n_7302),
.B2(n_7301),
.Y(n_8361)
);

HB1xp67_ASAP7_75t_L g8362 ( 
.A(n_7202),
.Y(n_8362)
);

INVx1_ASAP7_75t_L g8363 ( 
.A(n_7214),
.Y(n_8363)
);

AO21x1_ASAP7_75t_L g8364 ( 
.A1(n_7244),
.A2(n_7049),
.B(n_6993),
.Y(n_8364)
);

CKINVDCx8_ASAP7_75t_R g8365 ( 
.A(n_7521),
.Y(n_8365)
);

INVx1_ASAP7_75t_L g8366 ( 
.A(n_7216),
.Y(n_8366)
);

INVx1_ASAP7_75t_L g8367 ( 
.A(n_7216),
.Y(n_8367)
);

INVx2_ASAP7_75t_L g8368 ( 
.A(n_7910),
.Y(n_8368)
);

HB1xp67_ASAP7_75t_L g8369 ( 
.A(n_7202),
.Y(n_8369)
);

AOI22xp5_ASAP7_75t_L g8370 ( 
.A1(n_7561),
.A2(n_6722),
.B1(n_6493),
.B2(n_6733),
.Y(n_8370)
);

BUFx12f_ASAP7_75t_L g8371 ( 
.A(n_7639),
.Y(n_8371)
);

NOR2xp33_ASAP7_75t_L g8372 ( 
.A(n_7378),
.B(n_6583),
.Y(n_8372)
);

INVx2_ASAP7_75t_SL g8373 ( 
.A(n_7265),
.Y(n_8373)
);

NAND2x1p5_ASAP7_75t_L g8374 ( 
.A(n_8156),
.B(n_6245),
.Y(n_8374)
);

BUFx4_ASAP7_75t_SL g8375 ( 
.A(n_7314),
.Y(n_8375)
);

HB1xp67_ASAP7_75t_L g8376 ( 
.A(n_7322),
.Y(n_8376)
);

BUFx2_ASAP7_75t_R g8377 ( 
.A(n_7904),
.Y(n_8377)
);

INVx2_ASAP7_75t_L g8378 ( 
.A(n_7910),
.Y(n_8378)
);

OAI21x1_ASAP7_75t_L g8379 ( 
.A1(n_7967),
.A2(n_8030),
.B(n_8020),
.Y(n_8379)
);

INVx1_ASAP7_75t_L g8380 ( 
.A(n_7217),
.Y(n_8380)
);

INVx2_ASAP7_75t_L g8381 ( 
.A(n_7910),
.Y(n_8381)
);

INVx1_ASAP7_75t_L g8382 ( 
.A(n_7217),
.Y(n_8382)
);

INVx5_ASAP7_75t_L g8383 ( 
.A(n_7339),
.Y(n_8383)
);

BUFx3_ASAP7_75t_L g8384 ( 
.A(n_7339),
.Y(n_8384)
);

OAI21x1_ASAP7_75t_L g8385 ( 
.A1(n_7967),
.A2(n_6329),
.B(n_6325),
.Y(n_8385)
);

INVx2_ASAP7_75t_L g8386 ( 
.A(n_7910),
.Y(n_8386)
);

INVx2_ASAP7_75t_SL g8387 ( 
.A(n_7265),
.Y(n_8387)
);

AND2x4_ASAP7_75t_L g8388 ( 
.A(n_7299),
.B(n_6599),
.Y(n_8388)
);

OAI21xp5_ASAP7_75t_L g8389 ( 
.A1(n_7259),
.A2(n_7150),
.B(n_7147),
.Y(n_8389)
);

OA21x2_ASAP7_75t_L g8390 ( 
.A1(n_7170),
.A2(n_6617),
.B(n_6607),
.Y(n_8390)
);

NAND2x1p5_ASAP7_75t_L g8391 ( 
.A(n_8156),
.B(n_6245),
.Y(n_8391)
);

INVx6_ASAP7_75t_L g8392 ( 
.A(n_8001),
.Y(n_8392)
);

AOI22xp33_ASAP7_75t_L g8393 ( 
.A1(n_7652),
.A2(n_7165),
.B1(n_7302),
.B2(n_7301),
.Y(n_8393)
);

INVx1_ASAP7_75t_L g8394 ( 
.A(n_7223),
.Y(n_8394)
);

INVx2_ASAP7_75t_L g8395 ( 
.A(n_7869),
.Y(n_8395)
);

INVx1_ASAP7_75t_L g8396 ( 
.A(n_7223),
.Y(n_8396)
);

CKINVDCx6p67_ASAP7_75t_R g8397 ( 
.A(n_7339),
.Y(n_8397)
);

AOI21x1_ASAP7_75t_L g8398 ( 
.A1(n_7244),
.A2(n_7146),
.B(n_6646),
.Y(n_8398)
);

OR2x2_ASAP7_75t_L g8399 ( 
.A(n_7502),
.B(n_6364),
.Y(n_8399)
);

INVx1_ASAP7_75t_L g8400 ( 
.A(n_7228),
.Y(n_8400)
);

INVx4_ASAP7_75t_L g8401 ( 
.A(n_7694),
.Y(n_8401)
);

BUFx10_ASAP7_75t_L g8402 ( 
.A(n_7262),
.Y(n_8402)
);

INVx1_ASAP7_75t_L g8403 ( 
.A(n_7228),
.Y(n_8403)
);

AOI22xp5_ASAP7_75t_L g8404 ( 
.A1(n_7561),
.A2(n_6733),
.B1(n_6760),
.B2(n_6758),
.Y(n_8404)
);

INVx1_ASAP7_75t_L g8405 ( 
.A(n_7236),
.Y(n_8405)
);

BUFx6f_ASAP7_75t_L g8406 ( 
.A(n_7387),
.Y(n_8406)
);

INVx3_ASAP7_75t_L g8407 ( 
.A(n_7182),
.Y(n_8407)
);

BUFx5_ASAP7_75t_L g8408 ( 
.A(n_7661),
.Y(n_8408)
);

CKINVDCx11_ASAP7_75t_R g8409 ( 
.A(n_7600),
.Y(n_8409)
);

INVx2_ASAP7_75t_L g8410 ( 
.A(n_7869),
.Y(n_8410)
);

INVx4_ASAP7_75t_L g8411 ( 
.A(n_7694),
.Y(n_8411)
);

BUFx10_ASAP7_75t_L g8412 ( 
.A(n_7323),
.Y(n_8412)
);

CKINVDCx11_ASAP7_75t_R g8413 ( 
.A(n_7600),
.Y(n_8413)
);

INVx1_ASAP7_75t_L g8414 ( 
.A(n_7236),
.Y(n_8414)
);

INVx3_ASAP7_75t_L g8415 ( 
.A(n_7182),
.Y(n_8415)
);

INVx1_ASAP7_75t_L g8416 ( 
.A(n_7237),
.Y(n_8416)
);

INVx3_ASAP7_75t_L g8417 ( 
.A(n_7182),
.Y(n_8417)
);

OAI21x1_ASAP7_75t_L g8418 ( 
.A1(n_7967),
.A2(n_6329),
.B(n_6325),
.Y(n_8418)
);

AOI22xp33_ASAP7_75t_SL g8419 ( 
.A1(n_7165),
.A2(n_6938),
.B1(n_7008),
.B2(n_6944),
.Y(n_8419)
);

INVx1_ASAP7_75t_L g8420 ( 
.A(n_7237),
.Y(n_8420)
);

BUFx6f_ASAP7_75t_L g8421 ( 
.A(n_7387),
.Y(n_8421)
);

INVx1_ASAP7_75t_L g8422 ( 
.A(n_7250),
.Y(n_8422)
);

AND2x4_ASAP7_75t_L g8423 ( 
.A(n_7299),
.B(n_6599),
.Y(n_8423)
);

INVx1_ASAP7_75t_L g8424 ( 
.A(n_7250),
.Y(n_8424)
);

INVx1_ASAP7_75t_L g8425 ( 
.A(n_7252),
.Y(n_8425)
);

AOI22xp33_ASAP7_75t_L g8426 ( 
.A1(n_7652),
.A2(n_6417),
.B1(n_6720),
.B2(n_6670),
.Y(n_8426)
);

OAI21x1_ASAP7_75t_L g8427 ( 
.A1(n_8020),
.A2(n_6345),
.B(n_6329),
.Y(n_8427)
);

INVx2_ASAP7_75t_L g8428 ( 
.A(n_7741),
.Y(n_8428)
);

OAI21xp5_ASAP7_75t_L g8429 ( 
.A1(n_7399),
.A2(n_7286),
.B(n_7172),
.Y(n_8429)
);

INVx1_ASAP7_75t_L g8430 ( 
.A(n_7252),
.Y(n_8430)
);

INVx2_ASAP7_75t_L g8431 ( 
.A(n_7741),
.Y(n_8431)
);

INVx1_ASAP7_75t_L g8432 ( 
.A(n_7253),
.Y(n_8432)
);

NAND2xp5_ASAP7_75t_L g8433 ( 
.A(n_7415),
.B(n_6162),
.Y(n_8433)
);

OAI21x1_ASAP7_75t_L g8434 ( 
.A1(n_8020),
.A2(n_6345),
.B(n_6329),
.Y(n_8434)
);

INVx6_ASAP7_75t_L g8435 ( 
.A(n_8001),
.Y(n_8435)
);

INVx1_ASAP7_75t_L g8436 ( 
.A(n_7253),
.Y(n_8436)
);

INVx1_ASAP7_75t_L g8437 ( 
.A(n_7304),
.Y(n_8437)
);

CKINVDCx5p33_ASAP7_75t_R g8438 ( 
.A(n_7375),
.Y(n_8438)
);

INVx2_ASAP7_75t_SL g8439 ( 
.A(n_7265),
.Y(n_8439)
);

INVx2_ASAP7_75t_L g8440 ( 
.A(n_7741),
.Y(n_8440)
);

INVx1_ASAP7_75t_SL g8441 ( 
.A(n_7378),
.Y(n_8441)
);

INVx1_ASAP7_75t_L g8442 ( 
.A(n_7304),
.Y(n_8442)
);

AOI22xp33_ASAP7_75t_SL g8443 ( 
.A1(n_7190),
.A2(n_6938),
.B1(n_7008),
.B2(n_6944),
.Y(n_8443)
);

AOI22xp33_ASAP7_75t_L g8444 ( 
.A1(n_7939),
.A2(n_6417),
.B1(n_6670),
.B2(n_7010),
.Y(n_8444)
);

NAND2x1p5_ASAP7_75t_L g8445 ( 
.A(n_8156),
.B(n_7661),
.Y(n_8445)
);

INVx4_ASAP7_75t_L g8446 ( 
.A(n_7694),
.Y(n_8446)
);

BUFx12f_ASAP7_75t_L g8447 ( 
.A(n_7639),
.Y(n_8447)
);

INVx1_ASAP7_75t_L g8448 ( 
.A(n_7306),
.Y(n_8448)
);

AOI22xp33_ASAP7_75t_L g8449 ( 
.A1(n_7939),
.A2(n_6417),
.B1(n_7010),
.B2(n_6919),
.Y(n_8449)
);

INVx1_ASAP7_75t_L g8450 ( 
.A(n_7306),
.Y(n_8450)
);

INVx1_ASAP7_75t_L g8451 ( 
.A(n_7327),
.Y(n_8451)
);

AOI22xp33_ASAP7_75t_L g8452 ( 
.A1(n_7939),
.A2(n_6919),
.B1(n_6906),
.B2(n_6753),
.Y(n_8452)
);

BUFx2_ASAP7_75t_L g8453 ( 
.A(n_7891),
.Y(n_8453)
);

INVx1_ASAP7_75t_L g8454 ( 
.A(n_7327),
.Y(n_8454)
);

AOI21xp5_ASAP7_75t_L g8455 ( 
.A1(n_7222),
.A2(n_6473),
.B(n_6631),
.Y(n_8455)
);

INVx2_ASAP7_75t_L g8456 ( 
.A(n_7741),
.Y(n_8456)
);

INVx3_ASAP7_75t_L g8457 ( 
.A(n_7182),
.Y(n_8457)
);

AND2x2_ASAP7_75t_L g8458 ( 
.A(n_7712),
.B(n_6335),
.Y(n_8458)
);

INVx3_ASAP7_75t_L g8459 ( 
.A(n_7182),
.Y(n_8459)
);

AOI22xp33_ASAP7_75t_L g8460 ( 
.A1(n_7939),
.A2(n_6906),
.B1(n_6753),
.B2(n_7145),
.Y(n_8460)
);

INVx2_ASAP7_75t_L g8461 ( 
.A(n_7741),
.Y(n_8461)
);

INVx2_ASAP7_75t_L g8462 ( 
.A(n_7741),
.Y(n_8462)
);

OAI22xp5_ASAP7_75t_L g8463 ( 
.A1(n_7257),
.A2(n_6433),
.B1(n_6936),
.B2(n_6926),
.Y(n_8463)
);

AND2x4_ASAP7_75t_L g8464 ( 
.A(n_7299),
.B(n_6656),
.Y(n_8464)
);

INVx2_ASAP7_75t_L g8465 ( 
.A(n_7753),
.Y(n_8465)
);

NAND2xp5_ASAP7_75t_L g8466 ( 
.A(n_7415),
.B(n_6797),
.Y(n_8466)
);

AO21x1_ASAP7_75t_L g8467 ( 
.A1(n_7922),
.A2(n_6411),
.B(n_6401),
.Y(n_8467)
);

INVx2_ASAP7_75t_L g8468 ( 
.A(n_7753),
.Y(n_8468)
);

AOI22xp33_ASAP7_75t_L g8469 ( 
.A1(n_7939),
.A2(n_6753),
.B1(n_7145),
.B2(n_6944),
.Y(n_8469)
);

INVx1_ASAP7_75t_L g8470 ( 
.A(n_7336),
.Y(n_8470)
);

AOI22xp5_ASAP7_75t_SL g8471 ( 
.A1(n_7922),
.A2(n_6427),
.B1(n_6944),
.B2(n_6938),
.Y(n_8471)
);

AO21x2_ASAP7_75t_L g8472 ( 
.A1(n_8035),
.A2(n_7079),
.B(n_6411),
.Y(n_8472)
);

AOI22xp33_ASAP7_75t_SL g8473 ( 
.A1(n_7190),
.A2(n_7231),
.B1(n_7264),
.B2(n_7246),
.Y(n_8473)
);

INVx2_ASAP7_75t_SL g8474 ( 
.A(n_7265),
.Y(n_8474)
);

INVx1_ASAP7_75t_L g8475 ( 
.A(n_7336),
.Y(n_8475)
);

AOI22xp5_ASAP7_75t_SL g8476 ( 
.A1(n_7320),
.A2(n_7012),
.B1(n_7008),
.B2(n_6526),
.Y(n_8476)
);

INVx1_ASAP7_75t_L g8477 ( 
.A(n_7348),
.Y(n_8477)
);

INVx1_ASAP7_75t_L g8478 ( 
.A(n_7348),
.Y(n_8478)
);

CKINVDCx20_ASAP7_75t_R g8479 ( 
.A(n_7453),
.Y(n_8479)
);

INVx1_ASAP7_75t_L g8480 ( 
.A(n_7356),
.Y(n_8480)
);

NAND2x1p5_ASAP7_75t_L g8481 ( 
.A(n_8156),
.B(n_7661),
.Y(n_8481)
);

INVx2_ASAP7_75t_L g8482 ( 
.A(n_7753),
.Y(n_8482)
);

INVx1_ASAP7_75t_L g8483 ( 
.A(n_7356),
.Y(n_8483)
);

BUFx3_ASAP7_75t_L g8484 ( 
.A(n_8255),
.Y(n_8484)
);

AND2x2_ASAP7_75t_L g8485 ( 
.A(n_7712),
.B(n_6395),
.Y(n_8485)
);

INVx3_ASAP7_75t_L g8486 ( 
.A(n_7182),
.Y(n_8486)
);

INVx1_ASAP7_75t_L g8487 ( 
.A(n_7357),
.Y(n_8487)
);

BUFx3_ASAP7_75t_L g8488 ( 
.A(n_8255),
.Y(n_8488)
);

AOI22xp33_ASAP7_75t_L g8489 ( 
.A1(n_7287),
.A2(n_7008),
.B1(n_7012),
.B2(n_6619),
.Y(n_8489)
);

INVx1_ASAP7_75t_L g8490 ( 
.A(n_7357),
.Y(n_8490)
);

INVx2_ASAP7_75t_L g8491 ( 
.A(n_7753),
.Y(n_8491)
);

INVx6_ASAP7_75t_L g8492 ( 
.A(n_8001),
.Y(n_8492)
);

INVx2_ASAP7_75t_L g8493 ( 
.A(n_7753),
.Y(n_8493)
);

BUFx6f_ASAP7_75t_L g8494 ( 
.A(n_7387),
.Y(n_8494)
);

INVx1_ASAP7_75t_L g8495 ( 
.A(n_7361),
.Y(n_8495)
);

HB1xp67_ASAP7_75t_L g8496 ( 
.A(n_7322),
.Y(n_8496)
);

NOR2x1_ASAP7_75t_L g8497 ( 
.A(n_7694),
.B(n_6631),
.Y(n_8497)
);

INVxp33_ASAP7_75t_L g8498 ( 
.A(n_7808),
.Y(n_8498)
);

NAND2xp5_ASAP7_75t_L g8499 ( 
.A(n_7292),
.B(n_6797),
.Y(n_8499)
);

INVx2_ASAP7_75t_L g8500 ( 
.A(n_7753),
.Y(n_8500)
);

AOI222xp33_ASAP7_75t_L g8501 ( 
.A1(n_7480),
.A2(n_6401),
.B1(n_7012),
.B2(n_6834),
.C1(n_6755),
.C2(n_7119),
.Y(n_8501)
);

BUFx2_ASAP7_75t_L g8502 ( 
.A(n_7891),
.Y(n_8502)
);

INVx1_ASAP7_75t_L g8503 ( 
.A(n_7361),
.Y(n_8503)
);

INVx1_ASAP7_75t_L g8504 ( 
.A(n_7364),
.Y(n_8504)
);

NAND2x1p5_ASAP7_75t_L g8505 ( 
.A(n_8156),
.B(n_7661),
.Y(n_8505)
);

OR2x2_ASAP7_75t_L g8506 ( 
.A(n_7502),
.B(n_6364),
.Y(n_8506)
);

INVx1_ASAP7_75t_L g8507 ( 
.A(n_7364),
.Y(n_8507)
);

INVx2_ASAP7_75t_L g8508 ( 
.A(n_7266),
.Y(n_8508)
);

AOI22xp33_ASAP7_75t_SL g8509 ( 
.A1(n_7190),
.A2(n_7012),
.B1(n_6309),
.B2(n_6595),
.Y(n_8509)
);

INVx1_ASAP7_75t_L g8510 ( 
.A(n_7389),
.Y(n_8510)
);

INVx2_ASAP7_75t_L g8511 ( 
.A(n_7266),
.Y(n_8511)
);

INVx2_ASAP7_75t_L g8512 ( 
.A(n_7266),
.Y(n_8512)
);

AOI22xp5_ASAP7_75t_L g8513 ( 
.A1(n_7157),
.A2(n_6719),
.B1(n_6619),
.B2(n_6682),
.Y(n_8513)
);

BUFx2_ASAP7_75t_L g8514 ( 
.A(n_8052),
.Y(n_8514)
);

INVx2_ASAP7_75t_L g8515 ( 
.A(n_7869),
.Y(n_8515)
);

INVx1_ASAP7_75t_L g8516 ( 
.A(n_7389),
.Y(n_8516)
);

INVx1_ASAP7_75t_L g8517 ( 
.A(n_7416),
.Y(n_8517)
);

BUFx6f_ASAP7_75t_L g8518 ( 
.A(n_7387),
.Y(n_8518)
);

OAI22xp5_ASAP7_75t_L g8519 ( 
.A1(n_7257),
.A2(n_6433),
.B1(n_6937),
.B2(n_6926),
.Y(n_8519)
);

AO21x1_ASAP7_75t_L g8520 ( 
.A1(n_7562),
.A2(n_6755),
.B(n_6834),
.Y(n_8520)
);

NAND2xp5_ASAP7_75t_L g8521 ( 
.A(n_7292),
.B(n_6821),
.Y(n_8521)
);

INVx1_ASAP7_75t_L g8522 ( 
.A(n_7416),
.Y(n_8522)
);

AND2x2_ASAP7_75t_L g8523 ( 
.A(n_7732),
.B(n_6395),
.Y(n_8523)
);

INVx1_ASAP7_75t_L g8524 ( 
.A(n_7421),
.Y(n_8524)
);

INVx1_ASAP7_75t_L g8525 ( 
.A(n_7421),
.Y(n_8525)
);

INVx2_ASAP7_75t_L g8526 ( 
.A(n_7869),
.Y(n_8526)
);

INVx2_ASAP7_75t_L g8527 ( 
.A(n_7869),
.Y(n_8527)
);

BUFx3_ASAP7_75t_L g8528 ( 
.A(n_7648),
.Y(n_8528)
);

AND2x2_ASAP7_75t_L g8529 ( 
.A(n_7732),
.B(n_6425),
.Y(n_8529)
);

OAI21xp33_ASAP7_75t_L g8530 ( 
.A1(n_7629),
.A2(n_7150),
.B(n_6883),
.Y(n_8530)
);

HB1xp67_ASAP7_75t_L g8531 ( 
.A(n_7324),
.Y(n_8531)
);

INVx3_ASAP7_75t_L g8532 ( 
.A(n_7312),
.Y(n_8532)
);

BUFx2_ASAP7_75t_L g8533 ( 
.A(n_8052),
.Y(n_8533)
);

INVx1_ASAP7_75t_L g8534 ( 
.A(n_7427),
.Y(n_8534)
);

NOR2xp33_ASAP7_75t_L g8535 ( 
.A(n_7653),
.B(n_6583),
.Y(n_8535)
);

AOI22xp33_ASAP7_75t_L g8536 ( 
.A1(n_7287),
.A2(n_7011),
.B1(n_7070),
.B2(n_7059),
.Y(n_8536)
);

NAND2xp5_ASAP7_75t_L g8537 ( 
.A(n_7707),
.B(n_6821),
.Y(n_8537)
);

AOI22xp5_ASAP7_75t_L g8538 ( 
.A1(n_7157),
.A2(n_6719),
.B1(n_6526),
.B2(n_6608),
.Y(n_8538)
);

OAI22xp5_ASAP7_75t_L g8539 ( 
.A1(n_7257),
.A2(n_6937),
.B1(n_6979),
.B2(n_6873),
.Y(n_8539)
);

OAI21x1_ASAP7_75t_L g8540 ( 
.A1(n_8030),
.A2(n_6345),
.B(n_6329),
.Y(n_8540)
);

BUFx2_ASAP7_75t_R g8541 ( 
.A(n_7521),
.Y(n_8541)
);

HB1xp67_ASAP7_75t_L g8542 ( 
.A(n_7324),
.Y(n_8542)
);

AOI22xp33_ASAP7_75t_L g8543 ( 
.A1(n_7285),
.A2(n_7011),
.B1(n_7070),
.B2(n_7059),
.Y(n_8543)
);

INVx1_ASAP7_75t_L g8544 ( 
.A(n_7427),
.Y(n_8544)
);

INVx8_ASAP7_75t_L g8545 ( 
.A(n_7265),
.Y(n_8545)
);

INVx2_ASAP7_75t_L g8546 ( 
.A(n_7869),
.Y(n_8546)
);

NAND3xp33_ASAP7_75t_L g8547 ( 
.A(n_7172),
.B(n_6883),
.C(n_6881),
.Y(n_8547)
);

INVx1_ASAP7_75t_L g8548 ( 
.A(n_7434),
.Y(n_8548)
);

BUFx2_ASAP7_75t_L g8549 ( 
.A(n_7407),
.Y(n_8549)
);

AOI22xp33_ASAP7_75t_SL g8550 ( 
.A1(n_7190),
.A2(n_6309),
.B1(n_6595),
.B2(n_6236),
.Y(n_8550)
);

HB1xp67_ASAP7_75t_L g8551 ( 
.A(n_7351),
.Y(n_8551)
);

NOR2xp33_ASAP7_75t_L g8552 ( 
.A(n_7653),
.B(n_6567),
.Y(n_8552)
);

INVx2_ASAP7_75t_SL g8553 ( 
.A(n_7265),
.Y(n_8553)
);

INVx1_ASAP7_75t_L g8554 ( 
.A(n_7434),
.Y(n_8554)
);

CKINVDCx6p67_ASAP7_75t_R g8555 ( 
.A(n_7159),
.Y(n_8555)
);

BUFx6f_ASAP7_75t_L g8556 ( 
.A(n_7404),
.Y(n_8556)
);

INVx1_ASAP7_75t_L g8557 ( 
.A(n_7449),
.Y(n_8557)
);

OA21x2_ASAP7_75t_L g8558 ( 
.A1(n_7472),
.A2(n_6646),
.B(n_6617),
.Y(n_8558)
);

AND2x2_ASAP7_75t_L g8559 ( 
.A(n_7732),
.B(n_6425),
.Y(n_8559)
);

INVx2_ASAP7_75t_L g8560 ( 
.A(n_8022),
.Y(n_8560)
);

BUFx2_ASAP7_75t_SL g8561 ( 
.A(n_7453),
.Y(n_8561)
);

INVx1_ASAP7_75t_L g8562 ( 
.A(n_7449),
.Y(n_8562)
);

INVx1_ASAP7_75t_L g8563 ( 
.A(n_7455),
.Y(n_8563)
);

INVx2_ASAP7_75t_L g8564 ( 
.A(n_8022),
.Y(n_8564)
);

INVx2_ASAP7_75t_L g8565 ( 
.A(n_8022),
.Y(n_8565)
);

HB1xp67_ASAP7_75t_L g8566 ( 
.A(n_7351),
.Y(n_8566)
);

INVx2_ASAP7_75t_L g8567 ( 
.A(n_8022),
.Y(n_8567)
);

AO21x2_ASAP7_75t_L g8568 ( 
.A1(n_8035),
.A2(n_6881),
.B(n_6375),
.Y(n_8568)
);

BUFx2_ASAP7_75t_SL g8569 ( 
.A(n_7810),
.Y(n_8569)
);

INVx3_ASAP7_75t_L g8570 ( 
.A(n_7312),
.Y(n_8570)
);

INVx2_ASAP7_75t_L g8571 ( 
.A(n_8022),
.Y(n_8571)
);

OR2x2_ASAP7_75t_L g8572 ( 
.A(n_7502),
.B(n_6364),
.Y(n_8572)
);

INVx1_ASAP7_75t_L g8573 ( 
.A(n_7455),
.Y(n_8573)
);

AOI22xp33_ASAP7_75t_SL g8574 ( 
.A1(n_7231),
.A2(n_6309),
.B1(n_6595),
.B2(n_6236),
.Y(n_8574)
);

INVx1_ASAP7_75t_SL g8575 ( 
.A(n_7873),
.Y(n_8575)
);

BUFx2_ASAP7_75t_L g8576 ( 
.A(n_7407),
.Y(n_8576)
);

AOI22xp33_ASAP7_75t_L g8577 ( 
.A1(n_7285),
.A2(n_7011),
.B1(n_7070),
.B2(n_7059),
.Y(n_8577)
);

INVx2_ASAP7_75t_L g8578 ( 
.A(n_8022),
.Y(n_8578)
);

INVx2_ASAP7_75t_L g8579 ( 
.A(n_8025),
.Y(n_8579)
);

INVx2_ASAP7_75t_L g8580 ( 
.A(n_8025),
.Y(n_8580)
);

BUFx3_ASAP7_75t_L g8581 ( 
.A(n_7648),
.Y(n_8581)
);

INVx2_ASAP7_75t_L g8582 ( 
.A(n_8025),
.Y(n_8582)
);

INVx1_ASAP7_75t_L g8583 ( 
.A(n_7468),
.Y(n_8583)
);

AND2x2_ASAP7_75t_L g8584 ( 
.A(n_7756),
.B(n_6425),
.Y(n_8584)
);

AND2x4_ASAP7_75t_L g8585 ( 
.A(n_7316),
.B(n_6656),
.Y(n_8585)
);

AOI22xp33_ASAP7_75t_SL g8586 ( 
.A1(n_7231),
.A2(n_6309),
.B1(n_6595),
.B2(n_6236),
.Y(n_8586)
);

AOI22xp33_ASAP7_75t_L g8587 ( 
.A1(n_7406),
.A2(n_7282),
.B1(n_7330),
.B2(n_7497),
.Y(n_8587)
);

BUFx3_ASAP7_75t_L g8588 ( 
.A(n_7648),
.Y(n_8588)
);

BUFx2_ASAP7_75t_R g8589 ( 
.A(n_7743),
.Y(n_8589)
);

INVx2_ASAP7_75t_L g8590 ( 
.A(n_8025),
.Y(n_8590)
);

INVx2_ASAP7_75t_L g8591 ( 
.A(n_8025),
.Y(n_8591)
);

INVx2_ASAP7_75t_L g8592 ( 
.A(n_8025),
.Y(n_8592)
);

NAND2xp5_ASAP7_75t_L g8593 ( 
.A(n_7707),
.B(n_6828),
.Y(n_8593)
);

INVx1_ASAP7_75t_L g8594 ( 
.A(n_7468),
.Y(n_8594)
);

NAND2x1p5_ASAP7_75t_L g8595 ( 
.A(n_7645),
.B(n_6170),
.Y(n_8595)
);

INVx1_ASAP7_75t_L g8596 ( 
.A(n_7481),
.Y(n_8596)
);

AOI22xp33_ASAP7_75t_L g8597 ( 
.A1(n_7406),
.A2(n_7011),
.B1(n_7070),
.B2(n_7059),
.Y(n_8597)
);

INVx1_ASAP7_75t_L g8598 ( 
.A(n_7481),
.Y(n_8598)
);

INVx1_ASAP7_75t_SL g8599 ( 
.A(n_7873),
.Y(n_8599)
);

AND2x2_ASAP7_75t_L g8600 ( 
.A(n_7756),
.B(n_6440),
.Y(n_8600)
);

CKINVDCx11_ASAP7_75t_R g8601 ( 
.A(n_7810),
.Y(n_8601)
);

BUFx12f_ASAP7_75t_L g8602 ( 
.A(n_7855),
.Y(n_8602)
);

INVx1_ASAP7_75t_L g8603 ( 
.A(n_7482),
.Y(n_8603)
);

INVx1_ASAP7_75t_L g8604 ( 
.A(n_7482),
.Y(n_8604)
);

BUFx6f_ASAP7_75t_L g8605 ( 
.A(n_7404),
.Y(n_8605)
);

INVx3_ASAP7_75t_L g8606 ( 
.A(n_7312),
.Y(n_8606)
);

NAND2x1p5_ASAP7_75t_L g8607 ( 
.A(n_7645),
.B(n_6170),
.Y(n_8607)
);

HB1xp67_ASAP7_75t_L g8608 ( 
.A(n_7367),
.Y(n_8608)
);

NAND2xp5_ASAP7_75t_L g8609 ( 
.A(n_7750),
.B(n_6828),
.Y(n_8609)
);

INVx2_ASAP7_75t_L g8610 ( 
.A(n_8026),
.Y(n_8610)
);

AO21x1_ASAP7_75t_L g8611 ( 
.A1(n_7562),
.A2(n_6317),
.B(n_6979),
.Y(n_8611)
);

INVx1_ASAP7_75t_L g8612 ( 
.A(n_7490),
.Y(n_8612)
);

NAND2x1p5_ASAP7_75t_L g8613 ( 
.A(n_7694),
.B(n_6334),
.Y(n_8613)
);

INVx2_ASAP7_75t_L g8614 ( 
.A(n_8026),
.Y(n_8614)
);

OAI22xp33_ASAP7_75t_L g8615 ( 
.A1(n_7256),
.A2(n_7001),
.B1(n_6582),
.B2(n_6645),
.Y(n_8615)
);

OAI21xp5_ASAP7_75t_L g8616 ( 
.A1(n_7399),
.A2(n_6825),
.B(n_6677),
.Y(n_8616)
);

AO21x2_ASAP7_75t_L g8617 ( 
.A1(n_8035),
.A2(n_6375),
.B(n_6373),
.Y(n_8617)
);

OAI21x1_ASAP7_75t_L g8618 ( 
.A1(n_8030),
.A2(n_6361),
.B(n_6345),
.Y(n_8618)
);

INVx11_ASAP7_75t_L g8619 ( 
.A(n_7648),
.Y(n_8619)
);

INVx2_ASAP7_75t_L g8620 ( 
.A(n_8026),
.Y(n_8620)
);

INVx1_ASAP7_75t_L g8621 ( 
.A(n_7490),
.Y(n_8621)
);

AND2x2_ASAP7_75t_L g8622 ( 
.A(n_7756),
.B(n_6440),
.Y(n_8622)
);

AO21x1_ASAP7_75t_L g8623 ( 
.A1(n_7650),
.A2(n_6317),
.B(n_6228),
.Y(n_8623)
);

INVx2_ASAP7_75t_SL g8624 ( 
.A(n_7265),
.Y(n_8624)
);

INVx2_ASAP7_75t_L g8625 ( 
.A(n_8026),
.Y(n_8625)
);

AOI22xp33_ASAP7_75t_L g8626 ( 
.A1(n_7282),
.A2(n_7011),
.B1(n_7070),
.B2(n_7059),
.Y(n_8626)
);

INVx1_ASAP7_75t_L g8627 ( 
.A(n_7499),
.Y(n_8627)
);

INVx3_ASAP7_75t_L g8628 ( 
.A(n_7312),
.Y(n_8628)
);

OAI21x1_ASAP7_75t_L g8629 ( 
.A1(n_7880),
.A2(n_6361),
.B(n_6345),
.Y(n_8629)
);

INVx1_ASAP7_75t_L g8630 ( 
.A(n_7499),
.Y(n_8630)
);

OAI21x1_ASAP7_75t_L g8631 ( 
.A1(n_7880),
.A2(n_6367),
.B(n_6361),
.Y(n_8631)
);

BUFx12f_ASAP7_75t_L g8632 ( 
.A(n_7855),
.Y(n_8632)
);

INVx3_ASAP7_75t_L g8633 ( 
.A(n_7312),
.Y(n_8633)
);

BUFx3_ASAP7_75t_L g8634 ( 
.A(n_7985),
.Y(n_8634)
);

OAI21x1_ASAP7_75t_L g8635 ( 
.A1(n_7880),
.A2(n_6367),
.B(n_6361),
.Y(n_8635)
);

AND2x2_ASAP7_75t_L g8636 ( 
.A(n_7919),
.B(n_6440),
.Y(n_8636)
);

AND2x4_ASAP7_75t_L g8637 ( 
.A(n_7316),
.B(n_6656),
.Y(n_8637)
);

AOI22xp5_ASAP7_75t_L g8638 ( 
.A1(n_7716),
.A2(n_6608),
.B1(n_6643),
.B2(n_6563),
.Y(n_8638)
);

AND2x4_ASAP7_75t_L g8639 ( 
.A(n_7316),
.B(n_6656),
.Y(n_8639)
);

BUFx2_ASAP7_75t_R g8640 ( 
.A(n_7743),
.Y(n_8640)
);

INVx2_ASAP7_75t_L g8641 ( 
.A(n_8026),
.Y(n_8641)
);

HB1xp67_ASAP7_75t_L g8642 ( 
.A(n_7367),
.Y(n_8642)
);

INVx2_ASAP7_75t_SL g8643 ( 
.A(n_7726),
.Y(n_8643)
);

INVx3_ASAP7_75t_L g8644 ( 
.A(n_7312),
.Y(n_8644)
);

INVx1_ASAP7_75t_L g8645 ( 
.A(n_7524),
.Y(n_8645)
);

INVx2_ASAP7_75t_SL g8646 ( 
.A(n_7726),
.Y(n_8646)
);

INVx2_ASAP7_75t_L g8647 ( 
.A(n_8026),
.Y(n_8647)
);

INVx1_ASAP7_75t_L g8648 ( 
.A(n_7524),
.Y(n_8648)
);

BUFx6f_ASAP7_75t_L g8649 ( 
.A(n_7404),
.Y(n_8649)
);

INVx3_ASAP7_75t_L g8650 ( 
.A(n_7665),
.Y(n_8650)
);

AOI22xp33_ASAP7_75t_L g8651 ( 
.A1(n_7330),
.A2(n_7011),
.B1(n_7070),
.B2(n_7059),
.Y(n_8651)
);

OAI21xp5_ASAP7_75t_L g8652 ( 
.A1(n_7172),
.A2(n_6825),
.B(n_6677),
.Y(n_8652)
);

INVx2_ASAP7_75t_L g8653 ( 
.A(n_8123),
.Y(n_8653)
);

AOI22xp33_ASAP7_75t_L g8654 ( 
.A1(n_7497),
.A2(n_7011),
.B1(n_7070),
.B2(n_7059),
.Y(n_8654)
);

NAND2xp5_ASAP7_75t_L g8655 ( 
.A(n_7750),
.B(n_6933),
.Y(n_8655)
);

AOI22xp5_ASAP7_75t_SL g8656 ( 
.A1(n_7320),
.A2(n_6643),
.B1(n_6563),
.B2(n_7080),
.Y(n_8656)
);

HB1xp67_ASAP7_75t_L g8657 ( 
.A(n_7379),
.Y(n_8657)
);

INVx4_ASAP7_75t_L g8658 ( 
.A(n_7726),
.Y(n_8658)
);

OAI21x1_ASAP7_75t_L g8659 ( 
.A1(n_7436),
.A2(n_6367),
.B(n_6361),
.Y(n_8659)
);

NAND2xp5_ASAP7_75t_L g8660 ( 
.A(n_7708),
.B(n_6933),
.Y(n_8660)
);

BUFx6f_ASAP7_75t_L g8661 ( 
.A(n_7404),
.Y(n_8661)
);

BUFx2_ASAP7_75t_R g8662 ( 
.A(n_7363),
.Y(n_8662)
);

BUFx3_ASAP7_75t_L g8663 ( 
.A(n_7985),
.Y(n_8663)
);

INVx1_ASAP7_75t_L g8664 ( 
.A(n_7527),
.Y(n_8664)
);

OR2x2_ASAP7_75t_L g8665 ( 
.A(n_7502),
.B(n_6721),
.Y(n_8665)
);

INVx2_ASAP7_75t_L g8666 ( 
.A(n_8123),
.Y(n_8666)
);

INVx2_ASAP7_75t_L g8667 ( 
.A(n_8229),
.Y(n_8667)
);

INVx2_ASAP7_75t_L g8668 ( 
.A(n_8229),
.Y(n_8668)
);

INVx1_ASAP7_75t_L g8669 ( 
.A(n_7527),
.Y(n_8669)
);

HB1xp67_ASAP7_75t_L g8670 ( 
.A(n_7379),
.Y(n_8670)
);

INVx3_ASAP7_75t_L g8671 ( 
.A(n_7665),
.Y(n_8671)
);

INVx2_ASAP7_75t_L g8672 ( 
.A(n_8229),
.Y(n_8672)
);

INVx2_ASAP7_75t_L g8673 ( 
.A(n_8229),
.Y(n_8673)
);

INVx2_ASAP7_75t_L g8674 ( 
.A(n_8229),
.Y(n_8674)
);

AOI22xp33_ASAP7_75t_L g8675 ( 
.A1(n_7401),
.A2(n_7103),
.B1(n_6803),
.B2(n_7119),
.Y(n_8675)
);

OAI22xp5_ASAP7_75t_L g8676 ( 
.A1(n_7257),
.A2(n_6873),
.B1(n_6837),
.B2(n_6772),
.Y(n_8676)
);

AOI22xp33_ASAP7_75t_L g8677 ( 
.A1(n_7401),
.A2(n_7103),
.B1(n_6803),
.B2(n_6309),
.Y(n_8677)
);

INVx1_ASAP7_75t_L g8678 ( 
.A(n_7528),
.Y(n_8678)
);

BUFx6f_ASAP7_75t_L g8679 ( 
.A(n_7433),
.Y(n_8679)
);

INVx2_ASAP7_75t_SL g8680 ( 
.A(n_7726),
.Y(n_8680)
);

AOI21x1_ASAP7_75t_L g8681 ( 
.A1(n_7981),
.A2(n_8012),
.B(n_7983),
.Y(n_8681)
);

AOI22xp33_ASAP7_75t_L g8682 ( 
.A1(n_7573),
.A2(n_7103),
.B1(n_6803),
.B2(n_6309),
.Y(n_8682)
);

OA21x2_ASAP7_75t_L g8683 ( 
.A1(n_7472),
.A2(n_6667),
.B(n_6646),
.Y(n_8683)
);

INVx3_ASAP7_75t_L g8684 ( 
.A(n_7665),
.Y(n_8684)
);

BUFx3_ASAP7_75t_L g8685 ( 
.A(n_7985),
.Y(n_8685)
);

INVx1_ASAP7_75t_L g8686 ( 
.A(n_7528),
.Y(n_8686)
);

HB1xp67_ASAP7_75t_L g8687 ( 
.A(n_7400),
.Y(n_8687)
);

INVx2_ASAP7_75t_L g8688 ( 
.A(n_8123),
.Y(n_8688)
);

INVx1_ASAP7_75t_L g8689 ( 
.A(n_7537),
.Y(n_8689)
);

INVx1_ASAP7_75t_L g8690 ( 
.A(n_7537),
.Y(n_8690)
);

AND2x2_ASAP7_75t_L g8691 ( 
.A(n_7919),
.B(n_6459),
.Y(n_8691)
);

INVx1_ASAP7_75t_L g8692 ( 
.A(n_7556),
.Y(n_8692)
);

BUFx2_ASAP7_75t_L g8693 ( 
.A(n_7407),
.Y(n_8693)
);

BUFx10_ASAP7_75t_L g8694 ( 
.A(n_7323),
.Y(n_8694)
);

INVx3_ASAP7_75t_L g8695 ( 
.A(n_7665),
.Y(n_8695)
);

BUFx2_ASAP7_75t_SL g8696 ( 
.A(n_7879),
.Y(n_8696)
);

INVx1_ASAP7_75t_L g8697 ( 
.A(n_7556),
.Y(n_8697)
);

INVx2_ASAP7_75t_L g8698 ( 
.A(n_8123),
.Y(n_8698)
);

INVx6_ASAP7_75t_L g8699 ( 
.A(n_8001),
.Y(n_8699)
);

AOI22xp5_ASAP7_75t_L g8700 ( 
.A1(n_7716),
.A2(n_7001),
.B1(n_6582),
.B2(n_7041),
.Y(n_8700)
);

INVx1_ASAP7_75t_L g8701 ( 
.A(n_7558),
.Y(n_8701)
);

AOI22xp5_ASAP7_75t_L g8702 ( 
.A1(n_7736),
.A2(n_7222),
.B1(n_7699),
.B2(n_7332),
.Y(n_8702)
);

AND2x2_ASAP7_75t_L g8703 ( 
.A(n_7919),
.B(n_6459),
.Y(n_8703)
);

INVx3_ASAP7_75t_L g8704 ( 
.A(n_7835),
.Y(n_8704)
);

HB1xp67_ASAP7_75t_L g8705 ( 
.A(n_7400),
.Y(n_8705)
);

BUFx3_ASAP7_75t_L g8706 ( 
.A(n_7985),
.Y(n_8706)
);

INVx3_ASAP7_75t_L g8707 ( 
.A(n_7835),
.Y(n_8707)
);

OAI22xp33_ASAP7_75t_L g8708 ( 
.A1(n_7573),
.A2(n_6309),
.B1(n_6595),
.B2(n_6236),
.Y(n_8708)
);

INVx1_ASAP7_75t_L g8709 ( 
.A(n_7558),
.Y(n_8709)
);

INVx4_ASAP7_75t_L g8710 ( 
.A(n_7726),
.Y(n_8710)
);

AOI22xp33_ASAP7_75t_L g8711 ( 
.A1(n_7480),
.A2(n_7103),
.B1(n_6803),
.B2(n_6309),
.Y(n_8711)
);

INVx1_ASAP7_75t_SL g8712 ( 
.A(n_8088),
.Y(n_8712)
);

AND2x2_ASAP7_75t_L g8713 ( 
.A(n_8027),
.B(n_6459),
.Y(n_8713)
);

OAI21x1_ASAP7_75t_L g8714 ( 
.A1(n_7436),
.A2(n_6400),
.B(n_6367),
.Y(n_8714)
);

BUFx6f_ASAP7_75t_L g8715 ( 
.A(n_7433),
.Y(n_8715)
);

INVx2_ASAP7_75t_L g8716 ( 
.A(n_8123),
.Y(n_8716)
);

BUFx6f_ASAP7_75t_L g8717 ( 
.A(n_7433),
.Y(n_8717)
);

NAND2xp5_ASAP7_75t_L g8718 ( 
.A(n_7708),
.B(n_7027),
.Y(n_8718)
);

INVx6_ASAP7_75t_L g8719 ( 
.A(n_8001),
.Y(n_8719)
);

INVx1_ASAP7_75t_L g8720 ( 
.A(n_7569),
.Y(n_8720)
);

NAND2x1p5_ASAP7_75t_L g8721 ( 
.A(n_8003),
.B(n_6334),
.Y(n_8721)
);

AOI22xp5_ASAP7_75t_L g8722 ( 
.A1(n_7736),
.A2(n_7117),
.B1(n_7041),
.B2(n_6454),
.Y(n_8722)
);

NAND2x1p5_ASAP7_75t_L g8723 ( 
.A(n_8003),
.B(n_6334),
.Y(n_8723)
);

INVx2_ASAP7_75t_L g8724 ( 
.A(n_8123),
.Y(n_8724)
);

INVx1_ASAP7_75t_SL g8725 ( 
.A(n_8088),
.Y(n_8725)
);

INVx4_ASAP7_75t_L g8726 ( 
.A(n_7159),
.Y(n_8726)
);

INVx2_ASAP7_75t_L g8727 ( 
.A(n_8141),
.Y(n_8727)
);

INVx2_ASAP7_75t_L g8728 ( 
.A(n_8141),
.Y(n_8728)
);

INVx2_ASAP7_75t_L g8729 ( 
.A(n_8141),
.Y(n_8729)
);

INVx1_ASAP7_75t_L g8730 ( 
.A(n_7569),
.Y(n_8730)
);

AO21x1_ASAP7_75t_L g8731 ( 
.A1(n_7650),
.A2(n_6228),
.B(n_6202),
.Y(n_8731)
);

HB1xp67_ASAP7_75t_L g8732 ( 
.A(n_7435),
.Y(n_8732)
);

INVx4_ASAP7_75t_R g8733 ( 
.A(n_7433),
.Y(n_8733)
);

CKINVDCx5p33_ASAP7_75t_R g8734 ( 
.A(n_7879),
.Y(n_8734)
);

AOI22xp33_ASAP7_75t_SL g8735 ( 
.A1(n_7231),
.A2(n_6236),
.B1(n_6595),
.B2(n_6309),
.Y(n_8735)
);

INVx2_ASAP7_75t_L g8736 ( 
.A(n_8141),
.Y(n_8736)
);

CKINVDCx5p33_ASAP7_75t_R g8737 ( 
.A(n_7938),
.Y(n_8737)
);

BUFx12f_ASAP7_75t_L g8738 ( 
.A(n_8042),
.Y(n_8738)
);

AND2x2_ASAP7_75t_L g8739 ( 
.A(n_8027),
.B(n_6481),
.Y(n_8739)
);

AND2x4_ASAP7_75t_L g8740 ( 
.A(n_7331),
.B(n_6674),
.Y(n_8740)
);

AOI22xp33_ASAP7_75t_SL g8741 ( 
.A1(n_7246),
.A2(n_6236),
.B1(n_6786),
.B2(n_6595),
.Y(n_8741)
);

AND2x2_ASAP7_75t_L g8742 ( 
.A(n_8027),
.B(n_6481),
.Y(n_8742)
);

INVx1_ASAP7_75t_L g8743 ( 
.A(n_7574),
.Y(n_8743)
);

INVx2_ASAP7_75t_L g8744 ( 
.A(n_8141),
.Y(n_8744)
);

NAND2x1p5_ASAP7_75t_L g8745 ( 
.A(n_8003),
.B(n_6334),
.Y(n_8745)
);

AOI22xp33_ASAP7_75t_L g8746 ( 
.A1(n_7246),
.A2(n_7103),
.B1(n_6803),
.B2(n_6595),
.Y(n_8746)
);

INVx2_ASAP7_75t_L g8747 ( 
.A(n_8141),
.Y(n_8747)
);

INVx1_ASAP7_75t_L g8748 ( 
.A(n_7574),
.Y(n_8748)
);

AOI22xp33_ASAP7_75t_SL g8749 ( 
.A1(n_7246),
.A2(n_6236),
.B1(n_6786),
.B2(n_6595),
.Y(n_8749)
);

INVx2_ASAP7_75t_L g8750 ( 
.A(n_7760),
.Y(n_8750)
);

AOI22xp33_ASAP7_75t_L g8751 ( 
.A1(n_7264),
.A2(n_7103),
.B1(n_6803),
.B2(n_6786),
.Y(n_8751)
);

INVx2_ASAP7_75t_L g8752 ( 
.A(n_7760),
.Y(n_8752)
);

INVx1_ASAP7_75t_L g8753 ( 
.A(n_7578),
.Y(n_8753)
);

INVx2_ASAP7_75t_SL g8754 ( 
.A(n_7489),
.Y(n_8754)
);

OAI22xp5_ASAP7_75t_L g8755 ( 
.A1(n_7395),
.A2(n_6837),
.B1(n_6772),
.B2(n_6985),
.Y(n_8755)
);

INVx1_ASAP7_75t_L g8756 ( 
.A(n_7578),
.Y(n_8756)
);

INVx1_ASAP7_75t_L g8757 ( 
.A(n_7672),
.Y(n_8757)
);

AOI22xp33_ASAP7_75t_L g8758 ( 
.A1(n_7264),
.A2(n_7103),
.B1(n_6786),
.B2(n_6823),
.Y(n_8758)
);

INVx2_ASAP7_75t_L g8759 ( 
.A(n_7760),
.Y(n_8759)
);

CKINVDCx5p33_ASAP7_75t_R g8760 ( 
.A(n_7938),
.Y(n_8760)
);

CKINVDCx11_ASAP7_75t_R g8761 ( 
.A(n_7965),
.Y(n_8761)
);

INVx1_ASAP7_75t_L g8762 ( 
.A(n_7672),
.Y(n_8762)
);

OA21x2_ASAP7_75t_L g8763 ( 
.A1(n_7472),
.A2(n_6683),
.B(n_6667),
.Y(n_8763)
);

INVxp67_ASAP7_75t_SL g8764 ( 
.A(n_7749),
.Y(n_8764)
);

NAND2xp5_ASAP7_75t_L g8765 ( 
.A(n_7597),
.B(n_7027),
.Y(n_8765)
);

INVx1_ASAP7_75t_L g8766 ( 
.A(n_7673),
.Y(n_8766)
);

HB1xp67_ASAP7_75t_L g8767 ( 
.A(n_7435),
.Y(n_8767)
);

CKINVDCx5p33_ASAP7_75t_R g8768 ( 
.A(n_7965),
.Y(n_8768)
);

INVx1_ASAP7_75t_L g8769 ( 
.A(n_7673),
.Y(n_8769)
);

INVx2_ASAP7_75t_SL g8770 ( 
.A(n_7489),
.Y(n_8770)
);

OR2x2_ASAP7_75t_L g8771 ( 
.A(n_7502),
.B(n_6721),
.Y(n_8771)
);

INVxp67_ASAP7_75t_L g8772 ( 
.A(n_8189),
.Y(n_8772)
);

BUFx2_ASAP7_75t_L g8773 ( 
.A(n_7407),
.Y(n_8773)
);

INVx4_ASAP7_75t_L g8774 ( 
.A(n_7159),
.Y(n_8774)
);

OA21x2_ASAP7_75t_L g8775 ( 
.A1(n_7409),
.A2(n_6683),
.B(n_6667),
.Y(n_8775)
);

AO21x1_ASAP7_75t_L g8776 ( 
.A1(n_7969),
.A2(n_6280),
.B(n_6202),
.Y(n_8776)
);

INVx2_ASAP7_75t_L g8777 ( 
.A(n_8229),
.Y(n_8777)
);

AO21x1_ASAP7_75t_SL g8778 ( 
.A1(n_7577),
.A2(n_6464),
.B(n_6455),
.Y(n_8778)
);

INVx1_ASAP7_75t_L g8779 ( 
.A(n_7684),
.Y(n_8779)
);

CKINVDCx20_ASAP7_75t_R g8780 ( 
.A(n_7476),
.Y(n_8780)
);

INVx1_ASAP7_75t_L g8781 ( 
.A(n_7684),
.Y(n_8781)
);

INVx2_ASAP7_75t_L g8782 ( 
.A(n_8266),
.Y(n_8782)
);

INVx6_ASAP7_75t_L g8783 ( 
.A(n_8142),
.Y(n_8783)
);

INVx1_ASAP7_75t_L g8784 ( 
.A(n_7703),
.Y(n_8784)
);

OAI22xp33_ASAP7_75t_L g8785 ( 
.A1(n_8282),
.A2(n_6786),
.B1(n_6823),
.B2(n_6236),
.Y(n_8785)
);

AND2x2_ASAP7_75t_L g8786 ( 
.A(n_8136),
.B(n_6481),
.Y(n_8786)
);

CKINVDCx16_ASAP7_75t_R g8787 ( 
.A(n_8034),
.Y(n_8787)
);

INVx5_ASAP7_75t_L g8788 ( 
.A(n_7158),
.Y(n_8788)
);

INVx1_ASAP7_75t_L g8789 ( 
.A(n_7703),
.Y(n_8789)
);

INVx1_ASAP7_75t_L g8790 ( 
.A(n_7714),
.Y(n_8790)
);

AND2x4_ASAP7_75t_L g8791 ( 
.A(n_7331),
.B(n_6674),
.Y(n_8791)
);

INVx2_ASAP7_75t_L g8792 ( 
.A(n_8266),
.Y(n_8792)
);

INVx2_ASAP7_75t_SL g8793 ( 
.A(n_7489),
.Y(n_8793)
);

INVx2_ASAP7_75t_L g8794 ( 
.A(n_8266),
.Y(n_8794)
);

BUFx2_ASAP7_75t_L g8795 ( 
.A(n_7407),
.Y(n_8795)
);

INVx1_ASAP7_75t_L g8796 ( 
.A(n_7714),
.Y(n_8796)
);

NAND2x1p5_ASAP7_75t_L g8797 ( 
.A(n_8003),
.B(n_6786),
.Y(n_8797)
);

OAI21xp5_ASAP7_75t_L g8798 ( 
.A1(n_7332),
.A2(n_6850),
.B(n_7152),
.Y(n_8798)
);

AOI22xp33_ASAP7_75t_L g8799 ( 
.A1(n_7264),
.A2(n_6786),
.B1(n_6949),
.B2(n_6823),
.Y(n_8799)
);

INVx1_ASAP7_75t_L g8800 ( 
.A(n_7729),
.Y(n_8800)
);

OAI21x1_ASAP7_75t_L g8801 ( 
.A1(n_7436),
.A2(n_6400),
.B(n_6367),
.Y(n_8801)
);

BUFx3_ASAP7_75t_L g8802 ( 
.A(n_8081),
.Y(n_8802)
);

BUFx12f_ASAP7_75t_L g8803 ( 
.A(n_8042),
.Y(n_8803)
);

INVx1_ASAP7_75t_L g8804 ( 
.A(n_7729),
.Y(n_8804)
);

HB1xp67_ASAP7_75t_L g8805 ( 
.A(n_7523),
.Y(n_8805)
);

AOI22xp33_ASAP7_75t_L g8806 ( 
.A1(n_7381),
.A2(n_6786),
.B1(n_6949),
.B2(n_6823),
.Y(n_8806)
);

INVx1_ASAP7_75t_L g8807 ( 
.A(n_7739),
.Y(n_8807)
);

INVx1_ASAP7_75t_SL g8808 ( 
.A(n_7790),
.Y(n_8808)
);

INVx2_ASAP7_75t_L g8809 ( 
.A(n_8266),
.Y(n_8809)
);

AOI22xp33_ASAP7_75t_L g8810 ( 
.A1(n_7381),
.A2(n_6786),
.B1(n_6949),
.B2(n_6823),
.Y(n_8810)
);

INVx1_ASAP7_75t_SL g8811 ( 
.A(n_7790),
.Y(n_8811)
);

INVx1_ASAP7_75t_L g8812 ( 
.A(n_7739),
.Y(n_8812)
);

INVx2_ASAP7_75t_L g8813 ( 
.A(n_8266),
.Y(n_8813)
);

AOI21x1_ASAP7_75t_L g8814 ( 
.A1(n_7981),
.A2(n_6697),
.B(n_6683),
.Y(n_8814)
);

BUFx2_ASAP7_75t_R g8815 ( 
.A(n_7363),
.Y(n_8815)
);

INVx2_ASAP7_75t_L g8816 ( 
.A(n_8266),
.Y(n_8816)
);

OAI21x1_ASAP7_75t_L g8817 ( 
.A1(n_7864),
.A2(n_6436),
.B(n_6400),
.Y(n_8817)
);

INVx2_ASAP7_75t_L g8818 ( 
.A(n_8301),
.Y(n_8818)
);

OAI21x1_ASAP7_75t_L g8819 ( 
.A1(n_7864),
.A2(n_6436),
.B(n_6400),
.Y(n_8819)
);

CKINVDCx20_ASAP7_75t_R g8820 ( 
.A(n_8029),
.Y(n_8820)
);

INVx1_ASAP7_75t_L g8821 ( 
.A(n_7745),
.Y(n_8821)
);

BUFx2_ASAP7_75t_R g8822 ( 
.A(n_7420),
.Y(n_8822)
);

INVx2_ASAP7_75t_SL g8823 ( 
.A(n_7489),
.Y(n_8823)
);

INVx2_ASAP7_75t_L g8824 ( 
.A(n_8301),
.Y(n_8824)
);

BUFx2_ASAP7_75t_L g8825 ( 
.A(n_7407),
.Y(n_8825)
);

AO21x2_ASAP7_75t_L g8826 ( 
.A1(n_7235),
.A2(n_7974),
.B(n_7619),
.Y(n_8826)
);

INVx2_ASAP7_75t_L g8827 ( 
.A(n_8301),
.Y(n_8827)
);

AO21x1_ASAP7_75t_SL g8828 ( 
.A1(n_7584),
.A2(n_6464),
.B(n_6455),
.Y(n_8828)
);

AND2x2_ASAP7_75t_L g8829 ( 
.A(n_8136),
.B(n_6519),
.Y(n_8829)
);

CKINVDCx20_ASAP7_75t_R g8830 ( 
.A(n_8029),
.Y(n_8830)
);

INVx1_ASAP7_75t_SL g8831 ( 
.A(n_8082),
.Y(n_8831)
);

INVx2_ASAP7_75t_L g8832 ( 
.A(n_8301),
.Y(n_8832)
);

CKINVDCx20_ASAP7_75t_R g8833 ( 
.A(n_8082),
.Y(n_8833)
);

CKINVDCx11_ASAP7_75t_R g8834 ( 
.A(n_8222),
.Y(n_8834)
);

INVx2_ASAP7_75t_L g8835 ( 
.A(n_8301),
.Y(n_8835)
);

INVx1_ASAP7_75t_L g8836 ( 
.A(n_7745),
.Y(n_8836)
);

AOI22xp33_ASAP7_75t_SL g8837 ( 
.A1(n_7381),
.A2(n_6966),
.B1(n_7083),
.B2(n_6949),
.Y(n_8837)
);

AOI21x1_ASAP7_75t_L g8838 ( 
.A1(n_7981),
.A2(n_6723),
.B(n_6697),
.Y(n_8838)
);

INVx2_ASAP7_75t_L g8839 ( 
.A(n_7760),
.Y(n_8839)
);

INVx2_ASAP7_75t_L g8840 ( 
.A(n_7760),
.Y(n_8840)
);

NAND2xp5_ASAP7_75t_L g8841 ( 
.A(n_7597),
.B(n_7028),
.Y(n_8841)
);

INVx1_ASAP7_75t_L g8842 ( 
.A(n_7748),
.Y(n_8842)
);

BUFx3_ASAP7_75t_L g8843 ( 
.A(n_8081),
.Y(n_8843)
);

OAI22xp5_ASAP7_75t_L g8844 ( 
.A1(n_7395),
.A2(n_6985),
.B1(n_7117),
.B2(n_7121),
.Y(n_8844)
);

INVx1_ASAP7_75t_L g8845 ( 
.A(n_7748),
.Y(n_8845)
);

HB1xp67_ASAP7_75t_L g8846 ( 
.A(n_7523),
.Y(n_8846)
);

CKINVDCx11_ASAP7_75t_R g8847 ( 
.A(n_8222),
.Y(n_8847)
);

HB1xp67_ASAP7_75t_L g8848 ( 
.A(n_7551),
.Y(n_8848)
);

OAI22xp5_ASAP7_75t_L g8849 ( 
.A1(n_7619),
.A2(n_7344),
.B1(n_7273),
.B2(n_7500),
.Y(n_8849)
);

AND2x2_ASAP7_75t_L g8850 ( 
.A(n_8136),
.B(n_7728),
.Y(n_8850)
);

INVx1_ASAP7_75t_L g8851 ( 
.A(n_7758),
.Y(n_8851)
);

OAI22xp5_ASAP7_75t_L g8852 ( 
.A1(n_7344),
.A2(n_7121),
.B1(n_7032),
.B2(n_7043),
.Y(n_8852)
);

INVx2_ASAP7_75t_L g8853 ( 
.A(n_7760),
.Y(n_8853)
);

INVx2_ASAP7_75t_L g8854 ( 
.A(n_7798),
.Y(n_8854)
);

AOI22xp33_ASAP7_75t_L g8855 ( 
.A1(n_7381),
.A2(n_6823),
.B1(n_6966),
.B2(n_6949),
.Y(n_8855)
);

INVx2_ASAP7_75t_L g8856 ( 
.A(n_7798),
.Y(n_8856)
);

OA21x2_ASAP7_75t_L g8857 ( 
.A1(n_7409),
.A2(n_6723),
.B(n_6697),
.Y(n_8857)
);

OAI21x1_ASAP7_75t_L g8858 ( 
.A1(n_7864),
.A2(n_6436),
.B(n_6400),
.Y(n_8858)
);

BUFx6f_ASAP7_75t_L g8859 ( 
.A(n_8081),
.Y(n_8859)
);

BUFx2_ASAP7_75t_SL g8860 ( 
.A(n_7158),
.Y(n_8860)
);

NOR2x1_ASAP7_75t_SL g8861 ( 
.A(n_7195),
.B(n_6947),
.Y(n_8861)
);

INVx1_ASAP7_75t_L g8862 ( 
.A(n_7758),
.Y(n_8862)
);

HB1xp67_ASAP7_75t_SL g8863 ( 
.A(n_7420),
.Y(n_8863)
);

INVx1_ASAP7_75t_L g8864 ( 
.A(n_7762),
.Y(n_8864)
);

INVx1_ASAP7_75t_L g8865 ( 
.A(n_7762),
.Y(n_8865)
);

INVx1_ASAP7_75t_L g8866 ( 
.A(n_7770),
.Y(n_8866)
);

BUFx6f_ASAP7_75t_L g8867 ( 
.A(n_8081),
.Y(n_8867)
);

AND2x4_ASAP7_75t_L g8868 ( 
.A(n_7331),
.B(n_8302),
.Y(n_8868)
);

AOI22xp33_ASAP7_75t_SL g8869 ( 
.A1(n_7383),
.A2(n_7083),
.B1(n_7087),
.B2(n_6823),
.Y(n_8869)
);

OAI21x1_ASAP7_75t_L g8870 ( 
.A1(n_7576),
.A2(n_6443),
.B(n_6436),
.Y(n_8870)
);

OR2x2_ASAP7_75t_L g8871 ( 
.A(n_7502),
.B(n_7934),
.Y(n_8871)
);

NAND2xp5_ASAP7_75t_L g8872 ( 
.A(n_7633),
.B(n_7028),
.Y(n_8872)
);

OAI21x1_ASAP7_75t_L g8873 ( 
.A1(n_7576),
.A2(n_7640),
.B(n_8238),
.Y(n_8873)
);

AOI21x1_ASAP7_75t_L g8874 ( 
.A1(n_7983),
.A2(n_7146),
.B(n_7144),
.Y(n_8874)
);

AOI22xp33_ASAP7_75t_L g8875 ( 
.A1(n_7383),
.A2(n_6823),
.B1(n_6966),
.B2(n_6949),
.Y(n_8875)
);

AND2x2_ASAP7_75t_L g8876 ( 
.A(n_7728),
.B(n_7761),
.Y(n_8876)
);

INVx3_ASAP7_75t_L g8877 ( 
.A(n_7835),
.Y(n_8877)
);

HB1xp67_ASAP7_75t_L g8878 ( 
.A(n_7551),
.Y(n_8878)
);

AOI22xp33_ASAP7_75t_L g8879 ( 
.A1(n_7383),
.A2(n_6823),
.B1(n_6966),
.B2(n_6949),
.Y(n_8879)
);

BUFx2_ASAP7_75t_R g8880 ( 
.A(n_7197),
.Y(n_8880)
);

AOI22xp33_ASAP7_75t_SL g8881 ( 
.A1(n_7383),
.A2(n_6966),
.B1(n_7083),
.B2(n_6949),
.Y(n_8881)
);

AO21x1_ASAP7_75t_L g8882 ( 
.A1(n_7969),
.A2(n_6284),
.B(n_6280),
.Y(n_8882)
);

INVx2_ASAP7_75t_L g8883 ( 
.A(n_7798),
.Y(n_8883)
);

BUFx3_ASAP7_75t_L g8884 ( 
.A(n_8243),
.Y(n_8884)
);

INVx1_ASAP7_75t_L g8885 ( 
.A(n_7770),
.Y(n_8885)
);

CKINVDCx11_ASAP7_75t_R g8886 ( 
.A(n_8243),
.Y(n_8886)
);

INVx2_ASAP7_75t_L g8887 ( 
.A(n_7798),
.Y(n_8887)
);

AO21x2_ASAP7_75t_L g8888 ( 
.A1(n_7235),
.A2(n_6375),
.B(n_6373),
.Y(n_8888)
);

CKINVDCx11_ASAP7_75t_R g8889 ( 
.A(n_8243),
.Y(n_8889)
);

INVx1_ASAP7_75t_SL g8890 ( 
.A(n_8207),
.Y(n_8890)
);

OAI22xp5_ASAP7_75t_L g8891 ( 
.A1(n_7273),
.A2(n_7032),
.B1(n_7043),
.B2(n_6666),
.Y(n_8891)
);

AO21x2_ASAP7_75t_L g8892 ( 
.A1(n_7235),
.A2(n_6392),
.B(n_6373),
.Y(n_8892)
);

NAND2x1p5_ASAP7_75t_L g8893 ( 
.A(n_8003),
.B(n_6949),
.Y(n_8893)
);

INVx3_ASAP7_75t_L g8894 ( 
.A(n_7835),
.Y(n_8894)
);

BUFx3_ASAP7_75t_L g8895 ( 
.A(n_8243),
.Y(n_8895)
);

INVx2_ASAP7_75t_L g8896 ( 
.A(n_7798),
.Y(n_8896)
);

OAI21xp5_ASAP7_75t_L g8897 ( 
.A1(n_7797),
.A2(n_6850),
.B(n_7152),
.Y(n_8897)
);

INVx1_ASAP7_75t_L g8898 ( 
.A(n_7771),
.Y(n_8898)
);

NAND2xp5_ASAP7_75t_L g8899 ( 
.A(n_7633),
.B(n_7830),
.Y(n_8899)
);

CKINVDCx20_ASAP7_75t_R g8900 ( 
.A(n_8207),
.Y(n_8900)
);

NAND2xp5_ASAP7_75t_L g8901 ( 
.A(n_7830),
.B(n_7045),
.Y(n_8901)
);

OAI22xp5_ASAP7_75t_L g8902 ( 
.A1(n_7500),
.A2(n_7410),
.B1(n_7471),
.B2(n_7463),
.Y(n_8902)
);

NAND2xp5_ASAP7_75t_L g8903 ( 
.A(n_8000),
.B(n_7045),
.Y(n_8903)
);

AOI22xp33_ASAP7_75t_SL g8904 ( 
.A1(n_7536),
.A2(n_7083),
.B1(n_7087),
.B2(n_6966),
.Y(n_8904)
);

AOI22xp33_ASAP7_75t_SL g8905 ( 
.A1(n_7536),
.A2(n_7083),
.B1(n_7087),
.B2(n_6966),
.Y(n_8905)
);

INVx6_ASAP7_75t_L g8906 ( 
.A(n_8142),
.Y(n_8906)
);

NAND2x1p5_ASAP7_75t_L g8907 ( 
.A(n_7438),
.B(n_6966),
.Y(n_8907)
);

CKINVDCx11_ASAP7_75t_R g8908 ( 
.A(n_7159),
.Y(n_8908)
);

CKINVDCx11_ASAP7_75t_R g8909 ( 
.A(n_7787),
.Y(n_8909)
);

OAI22xp5_ASAP7_75t_L g8910 ( 
.A1(n_7410),
.A2(n_7471),
.B1(n_7463),
.B2(n_7380),
.Y(n_8910)
);

INVx3_ASAP7_75t_L g8911 ( 
.A(n_7835),
.Y(n_8911)
);

NAND2x1p5_ASAP7_75t_L g8912 ( 
.A(n_7439),
.B(n_6966),
.Y(n_8912)
);

OAI21x1_ASAP7_75t_SL g8913 ( 
.A1(n_8069),
.A2(n_6520),
.B(n_6519),
.Y(n_8913)
);

INVx1_ASAP7_75t_L g8914 ( 
.A(n_7771),
.Y(n_8914)
);

BUFx12f_ASAP7_75t_L g8915 ( 
.A(n_7197),
.Y(n_8915)
);

INVx1_ASAP7_75t_L g8916 ( 
.A(n_7774),
.Y(n_8916)
);

INVx2_ASAP7_75t_L g8917 ( 
.A(n_7798),
.Y(n_8917)
);

INVx1_ASAP7_75t_L g8918 ( 
.A(n_7774),
.Y(n_8918)
);

INVx1_ASAP7_75t_L g8919 ( 
.A(n_7778),
.Y(n_8919)
);

INVx1_ASAP7_75t_L g8920 ( 
.A(n_7778),
.Y(n_8920)
);

AND2x4_ASAP7_75t_L g8921 ( 
.A(n_8302),
.B(n_6674),
.Y(n_8921)
);

INVx3_ASAP7_75t_L g8922 ( 
.A(n_7835),
.Y(n_8922)
);

INVx3_ASAP7_75t_L g8923 ( 
.A(n_7835),
.Y(n_8923)
);

INVx1_ASAP7_75t_L g8924 ( 
.A(n_7780),
.Y(n_8924)
);

OAI21x1_ASAP7_75t_L g8925 ( 
.A1(n_7576),
.A2(n_6443),
.B(n_6436),
.Y(n_8925)
);

OAI22xp33_ASAP7_75t_L g8926 ( 
.A1(n_8282),
.A2(n_7459),
.B1(n_7702),
.B2(n_7609),
.Y(n_8926)
);

AOI22xp33_ASAP7_75t_L g8927 ( 
.A1(n_7160),
.A2(n_7083),
.B1(n_7087),
.B2(n_6359),
.Y(n_8927)
);

OAI21x1_ASAP7_75t_L g8928 ( 
.A1(n_7640),
.A2(n_6445),
.B(n_6443),
.Y(n_8928)
);

BUFx3_ASAP7_75t_L g8929 ( 
.A(n_8142),
.Y(n_8929)
);

AO21x2_ASAP7_75t_L g8930 ( 
.A1(n_7974),
.A2(n_6439),
.B(n_6392),
.Y(n_8930)
);

NAND2xp5_ASAP7_75t_L g8931 ( 
.A(n_8000),
.B(n_7829),
.Y(n_8931)
);

AOI22xp33_ASAP7_75t_L g8932 ( 
.A1(n_7160),
.A2(n_7083),
.B1(n_7087),
.B2(n_6359),
.Y(n_8932)
);

AOI22xp33_ASAP7_75t_SL g8933 ( 
.A1(n_7536),
.A2(n_7087),
.B1(n_7083),
.B2(n_6674),
.Y(n_8933)
);

OA21x2_ASAP7_75t_L g8934 ( 
.A1(n_7409),
.A2(n_6759),
.B(n_6723),
.Y(n_8934)
);

OAI21xp5_ASAP7_75t_SL g8935 ( 
.A1(n_7584),
.A2(n_6896),
.B(n_6876),
.Y(n_8935)
);

HB1xp67_ASAP7_75t_L g8936 ( 
.A(n_7570),
.Y(n_8936)
);

INVx3_ASAP7_75t_L g8937 ( 
.A(n_7835),
.Y(n_8937)
);

INVx6_ASAP7_75t_L g8938 ( 
.A(n_8142),
.Y(n_8938)
);

INVx1_ASAP7_75t_L g8939 ( 
.A(n_7780),
.Y(n_8939)
);

OR2x2_ASAP7_75t_L g8940 ( 
.A(n_7502),
.B(n_6424),
.Y(n_8940)
);

BUFx8_ASAP7_75t_L g8941 ( 
.A(n_7983),
.Y(n_8941)
);

INVx1_ASAP7_75t_L g8942 ( 
.A(n_7791),
.Y(n_8942)
);

CKINVDCx5p33_ASAP7_75t_R g8943 ( 
.A(n_8256),
.Y(n_8943)
);

OAI21xp5_ASAP7_75t_L g8944 ( 
.A1(n_7797),
.A2(n_7101),
.B(n_7093),
.Y(n_8944)
);

OA21x2_ASAP7_75t_L g8945 ( 
.A1(n_7196),
.A2(n_6763),
.B(n_6759),
.Y(n_8945)
);

AOI21xp5_ASAP7_75t_L g8946 ( 
.A1(n_7230),
.A2(n_7000),
.B(n_6947),
.Y(n_8946)
);

OAI21x1_ASAP7_75t_L g8947 ( 
.A1(n_7640),
.A2(n_6445),
.B(n_6443),
.Y(n_8947)
);

INVx3_ASAP7_75t_L g8948 ( 
.A(n_7505),
.Y(n_8948)
);

INVx2_ASAP7_75t_L g8949 ( 
.A(n_7887),
.Y(n_8949)
);

INVx1_ASAP7_75t_L g8950 ( 
.A(n_7791),
.Y(n_8950)
);

INVx1_ASAP7_75t_L g8951 ( 
.A(n_7807),
.Y(n_8951)
);

OAI22xp5_ASAP7_75t_L g8952 ( 
.A1(n_7380),
.A2(n_7032),
.B1(n_7043),
.B2(n_6666),
.Y(n_8952)
);

AOI22xp33_ASAP7_75t_SL g8953 ( 
.A1(n_7540),
.A2(n_7083),
.B1(n_7087),
.B2(n_6700),
.Y(n_8953)
);

AOI22xp33_ASAP7_75t_SL g8954 ( 
.A1(n_7540),
.A2(n_7087),
.B1(n_6700),
.B2(n_6702),
.Y(n_8954)
);

INVx2_ASAP7_75t_L g8955 ( 
.A(n_7887),
.Y(n_8955)
);

BUFx2_ASAP7_75t_L g8956 ( 
.A(n_7407),
.Y(n_8956)
);

INVx1_ASAP7_75t_L g8957 ( 
.A(n_7807),
.Y(n_8957)
);

NAND2xp5_ASAP7_75t_L g8958 ( 
.A(n_8000),
.B(n_6530),
.Y(n_8958)
);

INVx3_ASAP7_75t_L g8959 ( 
.A(n_7505),
.Y(n_8959)
);

INVx1_ASAP7_75t_L g8960 ( 
.A(n_7839),
.Y(n_8960)
);

INVx1_ASAP7_75t_L g8961 ( 
.A(n_7839),
.Y(n_8961)
);

AOI22xp33_ASAP7_75t_SL g8962 ( 
.A1(n_7540),
.A2(n_7087),
.B1(n_6700),
.B2(n_6702),
.Y(n_8962)
);

INVx1_ASAP7_75t_L g8963 ( 
.A(n_7854),
.Y(n_8963)
);

INVx1_ASAP7_75t_L g8964 ( 
.A(n_7854),
.Y(n_8964)
);

AO21x1_ASAP7_75t_SL g8965 ( 
.A1(n_8069),
.A2(n_6486),
.B(n_6475),
.Y(n_8965)
);

AOI22xp5_ASAP7_75t_L g8966 ( 
.A1(n_7699),
.A2(n_6454),
.B1(n_6579),
.B2(n_6567),
.Y(n_8966)
);

NAND2xp5_ASAP7_75t_L g8967 ( 
.A(n_8000),
.B(n_6530),
.Y(n_8967)
);

INVx1_ASAP7_75t_L g8968 ( 
.A(n_7856),
.Y(n_8968)
);

AOI22xp33_ASAP7_75t_L g8969 ( 
.A1(n_7160),
.A2(n_6359),
.B1(n_6866),
.B2(n_6402),
.Y(n_8969)
);

BUFx3_ASAP7_75t_L g8970 ( 
.A(n_8142),
.Y(n_8970)
);

AO21x1_ASAP7_75t_SL g8971 ( 
.A1(n_8093),
.A2(n_6486),
.B(n_6475),
.Y(n_8971)
);

NAND2xp5_ASAP7_75t_SL g8972 ( 
.A(n_7370),
.B(n_7142),
.Y(n_8972)
);

AOI22xp33_ASAP7_75t_SL g8973 ( 
.A1(n_7547),
.A2(n_6700),
.B1(n_6702),
.B2(n_6920),
.Y(n_8973)
);

AOI22xp33_ASAP7_75t_L g8974 ( 
.A1(n_7629),
.A2(n_6359),
.B1(n_6866),
.B2(n_6402),
.Y(n_8974)
);

INVx2_ASAP7_75t_L g8975 ( 
.A(n_7887),
.Y(n_8975)
);

INVx4_ASAP7_75t_L g8976 ( 
.A(n_7242),
.Y(n_8976)
);

AO21x1_ASAP7_75t_SL g8977 ( 
.A1(n_8093),
.A2(n_6523),
.B(n_6509),
.Y(n_8977)
);

INVx2_ASAP7_75t_L g8978 ( 
.A(n_8037),
.Y(n_8978)
);

AOI22xp33_ASAP7_75t_L g8979 ( 
.A1(n_8161),
.A2(n_6359),
.B1(n_6866),
.B2(n_6402),
.Y(n_8979)
);

OAI22xp5_ASAP7_75t_L g8980 ( 
.A1(n_7525),
.A2(n_6666),
.B1(n_6520),
.B2(n_6525),
.Y(n_8980)
);

INVx2_ASAP7_75t_L g8981 ( 
.A(n_8037),
.Y(n_8981)
);

AOI22xp33_ASAP7_75t_L g8982 ( 
.A1(n_8161),
.A2(n_6359),
.B1(n_6866),
.B2(n_6402),
.Y(n_8982)
);

AOI22xp33_ASAP7_75t_SL g8983 ( 
.A1(n_7547),
.A2(n_6702),
.B1(n_6943),
.B2(n_6920),
.Y(n_8983)
);

INVx1_ASAP7_75t_L g8984 ( 
.A(n_7856),
.Y(n_8984)
);

AOI22xp33_ASAP7_75t_L g8985 ( 
.A1(n_7609),
.A2(n_6866),
.B1(n_5160),
.B2(n_5276),
.Y(n_8985)
);

INVx1_ASAP7_75t_L g8986 ( 
.A(n_7857),
.Y(n_8986)
);

BUFx2_ASAP7_75t_L g8987 ( 
.A(n_7407),
.Y(n_8987)
);

AOI22xp33_ASAP7_75t_L g8988 ( 
.A1(n_7459),
.A2(n_6866),
.B1(n_5276),
.B2(n_5292),
.Y(n_8988)
);

INVx2_ASAP7_75t_L g8989 ( 
.A(n_8037),
.Y(n_8989)
);

INVx1_ASAP7_75t_L g8990 ( 
.A(n_7857),
.Y(n_8990)
);

NAND2xp5_ASAP7_75t_L g8991 ( 
.A(n_8000),
.B(n_6694),
.Y(n_8991)
);

BUFx2_ASAP7_75t_L g8992 ( 
.A(n_7169),
.Y(n_8992)
);

AO21x1_ASAP7_75t_SL g8993 ( 
.A1(n_8120),
.A2(n_6523),
.B(n_6509),
.Y(n_8993)
);

AND2x4_ASAP7_75t_L g8994 ( 
.A(n_8302),
.B(n_6128),
.Y(n_8994)
);

INVx1_ASAP7_75t_L g8995 ( 
.A(n_7858),
.Y(n_8995)
);

INVx1_ASAP7_75t_L g8996 ( 
.A(n_7858),
.Y(n_8996)
);

INVx2_ASAP7_75t_L g8997 ( 
.A(n_8037),
.Y(n_8997)
);

CKINVDCx11_ASAP7_75t_R g8998 ( 
.A(n_7787),
.Y(n_8998)
);

OAI22xp33_ASAP7_75t_L g8999 ( 
.A1(n_7702),
.A2(n_7599),
.B1(n_8171),
.B2(n_7352),
.Y(n_8999)
);

OR2x2_ASAP7_75t_L g9000 ( 
.A(n_7502),
.B(n_6424),
.Y(n_9000)
);

AND2x2_ASAP7_75t_L g9001 ( 
.A(n_7728),
.B(n_6519),
.Y(n_9001)
);

INVx1_ASAP7_75t_L g9002 ( 
.A(n_7871),
.Y(n_9002)
);

OR2x2_ASAP7_75t_L g9003 ( 
.A(n_7934),
.B(n_8048),
.Y(n_9003)
);

INVx2_ASAP7_75t_L g9004 ( 
.A(n_7887),
.Y(n_9004)
);

OAI22xp33_ASAP7_75t_L g9005 ( 
.A1(n_7599),
.A2(n_6943),
.B1(n_6920),
.B2(n_6775),
.Y(n_9005)
);

HB1xp67_ASAP7_75t_L g9006 ( 
.A(n_7570),
.Y(n_9006)
);

AND2x2_ASAP7_75t_L g9007 ( 
.A(n_7761),
.B(n_6520),
.Y(n_9007)
);

INVx1_ASAP7_75t_L g9008 ( 
.A(n_7871),
.Y(n_9008)
);

INVx1_ASAP7_75t_L g9009 ( 
.A(n_7877),
.Y(n_9009)
);

AND2x2_ASAP7_75t_L g9010 ( 
.A(n_7761),
.B(n_6525),
.Y(n_9010)
);

INVx1_ASAP7_75t_L g9011 ( 
.A(n_7877),
.Y(n_9011)
);

OAI21x1_ASAP7_75t_L g9012 ( 
.A1(n_8238),
.A2(n_6445),
.B(n_6443),
.Y(n_9012)
);

BUFx3_ASAP7_75t_L g9013 ( 
.A(n_7229),
.Y(n_9013)
);

AOI22xp33_ASAP7_75t_SL g9014 ( 
.A1(n_7547),
.A2(n_7611),
.B1(n_7270),
.B2(n_7601),
.Y(n_9014)
);

INVx2_ASAP7_75t_L g9015 ( 
.A(n_7887),
.Y(n_9015)
);

AO21x2_ASAP7_75t_L g9016 ( 
.A1(n_7338),
.A2(n_6439),
.B(n_6392),
.Y(n_9016)
);

INVx1_ASAP7_75t_L g9017 ( 
.A(n_7898),
.Y(n_9017)
);

AND2x2_ASAP7_75t_L g9018 ( 
.A(n_8012),
.B(n_7277),
.Y(n_9018)
);

BUFx2_ASAP7_75t_L g9019 ( 
.A(n_7169),
.Y(n_9019)
);

INVx1_ASAP7_75t_SL g9020 ( 
.A(n_8256),
.Y(n_9020)
);

OAI22xp5_ASAP7_75t_L g9021 ( 
.A1(n_7525),
.A2(n_6556),
.B1(n_6611),
.B2(n_6525),
.Y(n_9021)
);

NOR2xp33_ASAP7_75t_L g9022 ( 
.A(n_7297),
.B(n_6567),
.Y(n_9022)
);

HB1xp67_ASAP7_75t_L g9023 ( 
.A(n_7625),
.Y(n_9023)
);

BUFx3_ASAP7_75t_L g9024 ( 
.A(n_7229),
.Y(n_9024)
);

NAND2xp5_ASAP7_75t_L g9025 ( 
.A(n_7829),
.B(n_7199),
.Y(n_9025)
);

BUFx2_ASAP7_75t_L g9026 ( 
.A(n_7169),
.Y(n_9026)
);

INVx1_ASAP7_75t_L g9027 ( 
.A(n_7898),
.Y(n_9027)
);

CKINVDCx11_ASAP7_75t_R g9028 ( 
.A(n_7787),
.Y(n_9028)
);

AOI21x1_ASAP7_75t_L g9029 ( 
.A1(n_8012),
.A2(n_7146),
.B(n_6763),
.Y(n_9029)
);

INVx4_ASAP7_75t_L g9030 ( 
.A(n_7242),
.Y(n_9030)
);

INVx1_ASAP7_75t_L g9031 ( 
.A(n_7912),
.Y(n_9031)
);

BUFx3_ASAP7_75t_L g9032 ( 
.A(n_7242),
.Y(n_9032)
);

INVx1_ASAP7_75t_L g9033 ( 
.A(n_7912),
.Y(n_9033)
);

INVx2_ASAP7_75t_L g9034 ( 
.A(n_7918),
.Y(n_9034)
);

INVx2_ASAP7_75t_L g9035 ( 
.A(n_7918),
.Y(n_9035)
);

INVx2_ASAP7_75t_L g9036 ( 
.A(n_7918),
.Y(n_9036)
);

INVx1_ASAP7_75t_L g9037 ( 
.A(n_7924),
.Y(n_9037)
);

INVx6_ASAP7_75t_L g9038 ( 
.A(n_7158),
.Y(n_9038)
);

BUFx2_ASAP7_75t_L g9039 ( 
.A(n_7169),
.Y(n_9039)
);

INVx1_ASAP7_75t_L g9040 ( 
.A(n_7924),
.Y(n_9040)
);

OAI21x1_ASAP7_75t_L g9041 ( 
.A1(n_8238),
.A2(n_6457),
.B(n_6445),
.Y(n_9041)
);

AND2x2_ASAP7_75t_L g9042 ( 
.A(n_7277),
.B(n_6556),
.Y(n_9042)
);

AOI22xp33_ASAP7_75t_L g9043 ( 
.A1(n_7717),
.A2(n_5276),
.B1(n_5292),
.B2(n_5144),
.Y(n_9043)
);

INVx8_ASAP7_75t_L g9044 ( 
.A(n_7271),
.Y(n_9044)
);

INVx2_ASAP7_75t_SL g9045 ( 
.A(n_7581),
.Y(n_9045)
);

AOI21x1_ASAP7_75t_L g9046 ( 
.A1(n_7310),
.A2(n_6763),
.B(n_6759),
.Y(n_9046)
);

INVx4_ASAP7_75t_L g9047 ( 
.A(n_7328),
.Y(n_9047)
);

INVx2_ASAP7_75t_SL g9048 ( 
.A(n_7581),
.Y(n_9048)
);

INVx2_ASAP7_75t_L g9049 ( 
.A(n_7918),
.Y(n_9049)
);

AND2x2_ASAP7_75t_L g9050 ( 
.A(n_7277),
.B(n_6556),
.Y(n_9050)
);

OAI21x1_ASAP7_75t_L g9051 ( 
.A1(n_8157),
.A2(n_6457),
.B(n_6445),
.Y(n_9051)
);

INVx1_ASAP7_75t_L g9052 ( 
.A(n_7942),
.Y(n_9052)
);

AOI22xp33_ASAP7_75t_L g9053 ( 
.A1(n_7717),
.A2(n_5292),
.B1(n_5276),
.B2(n_5047),
.Y(n_9053)
);

INVx3_ASAP7_75t_L g9054 ( 
.A(n_7505),
.Y(n_9054)
);

BUFx3_ASAP7_75t_L g9055 ( 
.A(n_7328),
.Y(n_9055)
);

NOR3xp33_ASAP7_75t_SL g9056 ( 
.A(n_8110),
.B(n_7088),
.C(n_7080),
.Y(n_9056)
);

INVx1_ASAP7_75t_L g9057 ( 
.A(n_7942),
.Y(n_9057)
);

INVx1_ASAP7_75t_L g9058 ( 
.A(n_7966),
.Y(n_9058)
);

BUFx3_ASAP7_75t_L g9059 ( 
.A(n_7328),
.Y(n_9059)
);

OR2x2_ASAP7_75t_L g9060 ( 
.A(n_7934),
.B(n_6424),
.Y(n_9060)
);

HB1xp67_ASAP7_75t_L g9061 ( 
.A(n_7625),
.Y(n_9061)
);

INVx1_ASAP7_75t_L g9062 ( 
.A(n_7966),
.Y(n_9062)
);

NAND2xp5_ASAP7_75t_SL g9063 ( 
.A(n_7370),
.B(n_7142),
.Y(n_9063)
);

OAI21x1_ASAP7_75t_L g9064 ( 
.A1(n_8157),
.A2(n_6469),
.B(n_6457),
.Y(n_9064)
);

BUFx3_ASAP7_75t_L g9065 ( 
.A(n_7815),
.Y(n_9065)
);

INVx2_ASAP7_75t_L g9066 ( 
.A(n_7918),
.Y(n_9066)
);

CKINVDCx11_ASAP7_75t_R g9067 ( 
.A(n_7815),
.Y(n_9067)
);

INVx1_ASAP7_75t_L g9068 ( 
.A(n_8068),
.Y(n_9068)
);

INVxp67_ASAP7_75t_L g9069 ( 
.A(n_8189),
.Y(n_9069)
);

OR2x2_ASAP7_75t_L g9070 ( 
.A(n_8048),
.B(n_6446),
.Y(n_9070)
);

BUFx2_ASAP7_75t_L g9071 ( 
.A(n_7169),
.Y(n_9071)
);

INVx1_ASAP7_75t_L g9072 ( 
.A(n_8068),
.Y(n_9072)
);

INVx1_ASAP7_75t_L g9073 ( 
.A(n_8074),
.Y(n_9073)
);

INVx2_ASAP7_75t_L g9074 ( 
.A(n_8211),
.Y(n_9074)
);

HB1xp67_ASAP7_75t_L g9075 ( 
.A(n_7767),
.Y(n_9075)
);

INVx1_ASAP7_75t_L g9076 ( 
.A(n_8074),
.Y(n_9076)
);

INVx4_ASAP7_75t_L g9077 ( 
.A(n_7158),
.Y(n_9077)
);

AO21x1_ASAP7_75t_L g9078 ( 
.A1(n_7310),
.A2(n_6287),
.B(n_6284),
.Y(n_9078)
);

BUFx2_ASAP7_75t_R g9079 ( 
.A(n_7366),
.Y(n_9079)
);

INVx1_ASAP7_75t_L g9080 ( 
.A(n_8078),
.Y(n_9080)
);

AOI22xp33_ASAP7_75t_L g9081 ( 
.A1(n_7603),
.A2(n_5292),
.B1(n_5276),
.B2(n_5047),
.Y(n_9081)
);

INVx2_ASAP7_75t_L g9082 ( 
.A(n_8211),
.Y(n_9082)
);

NAND2xp5_ASAP7_75t_L g9083 ( 
.A(n_7199),
.B(n_7219),
.Y(n_9083)
);

INVx1_ASAP7_75t_L g9084 ( 
.A(n_8078),
.Y(n_9084)
);

INVx2_ASAP7_75t_L g9085 ( 
.A(n_8211),
.Y(n_9085)
);

INVx1_ASAP7_75t_L g9086 ( 
.A(n_8079),
.Y(n_9086)
);

AND2x4_ASAP7_75t_L g9087 ( 
.A(n_8066),
.B(n_6128),
.Y(n_9087)
);

INVx1_ASAP7_75t_L g9088 ( 
.A(n_8079),
.Y(n_9088)
);

OAI22xp5_ASAP7_75t_L g9089 ( 
.A1(n_7403),
.A2(n_6651),
.B1(n_6737),
.B2(n_6611),
.Y(n_9089)
);

BUFx2_ASAP7_75t_L g9090 ( 
.A(n_7169),
.Y(n_9090)
);

BUFx2_ASAP7_75t_SL g9091 ( 
.A(n_7158),
.Y(n_9091)
);

OAI21x1_ASAP7_75t_L g9092 ( 
.A1(n_8157),
.A2(n_6469),
.B(n_6457),
.Y(n_9092)
);

INVx2_ASAP7_75t_L g9093 ( 
.A(n_8211),
.Y(n_9093)
);

INVx1_ASAP7_75t_L g9094 ( 
.A(n_8084),
.Y(n_9094)
);

INVx2_ASAP7_75t_L g9095 ( 
.A(n_8211),
.Y(n_9095)
);

HB1xp67_ASAP7_75t_L g9096 ( 
.A(n_7767),
.Y(n_9096)
);

AO21x2_ASAP7_75t_L g9097 ( 
.A1(n_7338),
.A2(n_6439),
.B(n_6392),
.Y(n_9097)
);

INVx1_ASAP7_75t_L g9098 ( 
.A(n_8084),
.Y(n_9098)
);

INVx1_ASAP7_75t_L g9099 ( 
.A(n_8087),
.Y(n_9099)
);

INVx2_ASAP7_75t_L g9100 ( 
.A(n_8211),
.Y(n_9100)
);

INVx1_ASAP7_75t_L g9101 ( 
.A(n_8087),
.Y(n_9101)
);

AOI22xp33_ASAP7_75t_SL g9102 ( 
.A1(n_7611),
.A2(n_7270),
.B1(n_7601),
.B2(n_7593),
.Y(n_9102)
);

OR2x6_ASAP7_75t_L g9103 ( 
.A(n_7504),
.B(n_6654),
.Y(n_9103)
);

INVx1_ASAP7_75t_L g9104 ( 
.A(n_8089),
.Y(n_9104)
);

AND2x2_ASAP7_75t_L g9105 ( 
.A(n_7298),
.B(n_6611),
.Y(n_9105)
);

NAND2xp5_ASAP7_75t_L g9106 ( 
.A(n_7219),
.B(n_6694),
.Y(n_9106)
);

INVx1_ASAP7_75t_L g9107 ( 
.A(n_8089),
.Y(n_9107)
);

HB1xp67_ASAP7_75t_SL g9108 ( 
.A(n_7276),
.Y(n_9108)
);

AO21x1_ASAP7_75t_L g9109 ( 
.A1(n_7349),
.A2(n_6322),
.B(n_6287),
.Y(n_9109)
);

AOI22xp33_ASAP7_75t_L g9110 ( 
.A1(n_7603),
.A2(n_5292),
.B1(n_5047),
.B2(n_4911),
.Y(n_9110)
);

HB1xp67_ASAP7_75t_L g9111 ( 
.A(n_7793),
.Y(n_9111)
);

NAND2xp5_ASAP7_75t_L g9112 ( 
.A(n_7243),
.B(n_7565),
.Y(n_9112)
);

AOI22xp33_ASAP7_75t_SL g9113 ( 
.A1(n_7611),
.A2(n_6943),
.B1(n_6775),
.B2(n_7112),
.Y(n_9113)
);

NOR2x1_ASAP7_75t_SL g9114 ( 
.A(n_7195),
.B(n_7000),
.Y(n_9114)
);

INVx1_ASAP7_75t_L g9115 ( 
.A(n_8101),
.Y(n_9115)
);

INVx1_ASAP7_75t_L g9116 ( 
.A(n_8101),
.Y(n_9116)
);

AOI22xp33_ASAP7_75t_L g9117 ( 
.A1(n_7268),
.A2(n_6943),
.B1(n_6838),
.B2(n_6859),
.Y(n_9117)
);

INVx1_ASAP7_75t_L g9118 ( 
.A(n_8106),
.Y(n_9118)
);

AOI22xp5_ASAP7_75t_L g9119 ( 
.A1(n_7598),
.A2(n_6579),
.B1(n_6614),
.B2(n_6567),
.Y(n_9119)
);

INVx1_ASAP7_75t_L g9120 ( 
.A(n_8106),
.Y(n_9120)
);

INVx2_ASAP7_75t_L g9121 ( 
.A(n_8211),
.Y(n_9121)
);

OAI21xp33_ASAP7_75t_SL g9122 ( 
.A1(n_8162),
.A2(n_7535),
.B(n_7491),
.Y(n_9122)
);

INVx2_ASAP7_75t_SL g9123 ( 
.A(n_7581),
.Y(n_9123)
);

INVx1_ASAP7_75t_L g9124 ( 
.A(n_8108),
.Y(n_9124)
);

HB1xp67_ASAP7_75t_L g9125 ( 
.A(n_7793),
.Y(n_9125)
);

AOI22xp33_ASAP7_75t_L g9126 ( 
.A1(n_7268),
.A2(n_6943),
.B1(n_6838),
.B2(n_6859),
.Y(n_9126)
);

BUFx2_ASAP7_75t_R g9127 ( 
.A(n_7366),
.Y(n_9127)
);

HB1xp67_ASAP7_75t_L g9128 ( 
.A(n_7796),
.Y(n_9128)
);

BUFx2_ASAP7_75t_L g9129 ( 
.A(n_7169),
.Y(n_9129)
);

AO21x2_ASAP7_75t_L g9130 ( 
.A1(n_7338),
.A2(n_6441),
.B(n_6439),
.Y(n_9130)
);

AND2x2_ASAP7_75t_L g9131 ( 
.A(n_7298),
.B(n_6651),
.Y(n_9131)
);

INVx1_ASAP7_75t_L g9132 ( 
.A(n_8108),
.Y(n_9132)
);

INVx2_ASAP7_75t_SL g9133 ( 
.A(n_7581),
.Y(n_9133)
);

INVx2_ASAP7_75t_L g9134 ( 
.A(n_8211),
.Y(n_9134)
);

INVx1_ASAP7_75t_L g9135 ( 
.A(n_8113),
.Y(n_9135)
);

INVx2_ASAP7_75t_L g9136 ( 
.A(n_7988),
.Y(n_9136)
);

INVx1_ASAP7_75t_L g9137 ( 
.A(n_8113),
.Y(n_9137)
);

INVx2_ASAP7_75t_L g9138 ( 
.A(n_7988),
.Y(n_9138)
);

OAI22xp5_ASAP7_75t_L g9139 ( 
.A1(n_7403),
.A2(n_6737),
.B1(n_6746),
.B2(n_6651),
.Y(n_9139)
);

CKINVDCx5p33_ASAP7_75t_R g9140 ( 
.A(n_7815),
.Y(n_9140)
);

INVx1_ASAP7_75t_L g9141 ( 
.A(n_8119),
.Y(n_9141)
);

INVx2_ASAP7_75t_SL g9142 ( 
.A(n_7582),
.Y(n_9142)
);

INVx2_ASAP7_75t_SL g9143 ( 
.A(n_7582),
.Y(n_9143)
);

BUFx3_ASAP7_75t_L g9144 ( 
.A(n_8107),
.Y(n_9144)
);

INVx2_ASAP7_75t_L g9145 ( 
.A(n_7988),
.Y(n_9145)
);

INVx1_ASAP7_75t_L g9146 ( 
.A(n_8119),
.Y(n_9146)
);

INVxp67_ASAP7_75t_L g9147 ( 
.A(n_8110),
.Y(n_9147)
);

INVx2_ASAP7_75t_L g9148 ( 
.A(n_7988),
.Y(n_9148)
);

NAND2xp5_ASAP7_75t_L g9149 ( 
.A(n_7243),
.B(n_6727),
.Y(n_9149)
);

INVx1_ASAP7_75t_L g9150 ( 
.A(n_8135),
.Y(n_9150)
);

AND2x2_ASAP7_75t_L g9151 ( 
.A(n_7298),
.B(n_6737),
.Y(n_9151)
);

INVx4_ASAP7_75t_L g9152 ( 
.A(n_7276),
.Y(n_9152)
);

BUFx3_ASAP7_75t_L g9153 ( 
.A(n_8107),
.Y(n_9153)
);

NAND2x1p5_ASAP7_75t_L g9154 ( 
.A(n_7438),
.B(n_7063),
.Y(n_9154)
);

BUFx12f_ASAP7_75t_L g9155 ( 
.A(n_7276),
.Y(n_9155)
);

BUFx6f_ASAP7_75t_L g9156 ( 
.A(n_7276),
.Y(n_9156)
);

INVx1_ASAP7_75t_L g9157 ( 
.A(n_8135),
.Y(n_9157)
);

NAND2x1p5_ASAP7_75t_L g9158 ( 
.A(n_7439),
.B(n_7063),
.Y(n_9158)
);

AND2x4_ASAP7_75t_L g9159 ( 
.A(n_8066),
.B(n_6128),
.Y(n_9159)
);

AND2x2_ASAP7_75t_L g9160 ( 
.A(n_7317),
.B(n_6746),
.Y(n_9160)
);

INVx1_ASAP7_75t_L g9161 ( 
.A(n_8150),
.Y(n_9161)
);

BUFx2_ASAP7_75t_SL g9162 ( 
.A(n_7276),
.Y(n_9162)
);

INVx2_ASAP7_75t_SL g9163 ( 
.A(n_7582),
.Y(n_9163)
);

AND2x4_ASAP7_75t_L g9164 ( 
.A(n_8066),
.B(n_6128),
.Y(n_9164)
);

AND2x2_ASAP7_75t_L g9165 ( 
.A(n_7317),
.B(n_6746),
.Y(n_9165)
);

OAI21x1_ASAP7_75t_L g9166 ( 
.A1(n_7613),
.A2(n_6469),
.B(n_6457),
.Y(n_9166)
);

INVx4_ASAP7_75t_L g9167 ( 
.A(n_7422),
.Y(n_9167)
);

OAI21x1_ASAP7_75t_L g9168 ( 
.A1(n_7613),
.A2(n_6491),
.B(n_6469),
.Y(n_9168)
);

INVx1_ASAP7_75t_SL g9169 ( 
.A(n_7742),
.Y(n_9169)
);

CKINVDCx11_ASAP7_75t_R g9170 ( 
.A(n_8107),
.Y(n_9170)
);

NAND2x1p5_ASAP7_75t_L g9171 ( 
.A(n_7442),
.B(n_7105),
.Y(n_9171)
);

BUFx2_ASAP7_75t_L g9172 ( 
.A(n_7169),
.Y(n_9172)
);

AOI22xp33_ASAP7_75t_SL g9173 ( 
.A1(n_7270),
.A2(n_6943),
.B1(n_7112),
.B2(n_6875),
.Y(n_9173)
);

INVx11_ASAP7_75t_L g9174 ( 
.A(n_7808),
.Y(n_9174)
);

BUFx3_ASAP7_75t_L g9175 ( 
.A(n_8297),
.Y(n_9175)
);

OA21x2_ASAP7_75t_L g9176 ( 
.A1(n_7196),
.A2(n_6805),
.B(n_6767),
.Y(n_9176)
);

OAI22xp5_ASAP7_75t_L g9177 ( 
.A1(n_7300),
.A2(n_6799),
.B1(n_6814),
.B2(n_6773),
.Y(n_9177)
);

INVx2_ASAP7_75t_L g9178 ( 
.A(n_7988),
.Y(n_9178)
);

INVx1_ASAP7_75t_L g9179 ( 
.A(n_8150),
.Y(n_9179)
);

AOI22xp5_ASAP7_75t_L g9180 ( 
.A1(n_7598),
.A2(n_6614),
.B1(n_6629),
.B2(n_6579),
.Y(n_9180)
);

AOI22xp33_ASAP7_75t_SL g9181 ( 
.A1(n_7593),
.A2(n_6943),
.B1(n_7112),
.B2(n_6875),
.Y(n_9181)
);

INVx1_ASAP7_75t_L g9182 ( 
.A(n_8158),
.Y(n_9182)
);

INVx1_ASAP7_75t_L g9183 ( 
.A(n_8158),
.Y(n_9183)
);

INVx1_ASAP7_75t_L g9184 ( 
.A(n_8160),
.Y(n_9184)
);

INVx1_ASAP7_75t_L g9185 ( 
.A(n_8160),
.Y(n_9185)
);

BUFx6f_ASAP7_75t_L g9186 ( 
.A(n_7422),
.Y(n_9186)
);

OAI21x1_ASAP7_75t_L g9187 ( 
.A1(n_7613),
.A2(n_6491),
.B(n_6469),
.Y(n_9187)
);

HB1xp67_ASAP7_75t_L g9188 ( 
.A(n_7796),
.Y(n_9188)
);

CKINVDCx11_ASAP7_75t_R g9189 ( 
.A(n_7422),
.Y(n_9189)
);

INVx1_ASAP7_75t_L g9190 ( 
.A(n_8176),
.Y(n_9190)
);

OAI22xp33_ASAP7_75t_SL g9191 ( 
.A1(n_7308),
.A2(n_7669),
.B1(n_7579),
.B2(n_7437),
.Y(n_9191)
);

OAI22xp5_ASAP7_75t_L g9192 ( 
.A1(n_7300),
.A2(n_6799),
.B1(n_6814),
.B2(n_6773),
.Y(n_9192)
);

INVx1_ASAP7_75t_L g9193 ( 
.A(n_8176),
.Y(n_9193)
);

INVx3_ASAP7_75t_L g9194 ( 
.A(n_7505),
.Y(n_9194)
);

INVx1_ASAP7_75t_L g9195 ( 
.A(n_8177),
.Y(n_9195)
);

INVx2_ASAP7_75t_L g9196 ( 
.A(n_8005),
.Y(n_9196)
);

INVx1_ASAP7_75t_L g9197 ( 
.A(n_8177),
.Y(n_9197)
);

INVx2_ASAP7_75t_L g9198 ( 
.A(n_8005),
.Y(n_9198)
);

BUFx10_ASAP7_75t_L g9199 ( 
.A(n_7836),
.Y(n_9199)
);

AOI22xp5_ASAP7_75t_SL g9200 ( 
.A1(n_8230),
.A2(n_7088),
.B1(n_6542),
.B2(n_6561),
.Y(n_9200)
);

INVx2_ASAP7_75t_L g9201 ( 
.A(n_8005),
.Y(n_9201)
);

INVx1_ASAP7_75t_L g9202 ( 
.A(n_8190),
.Y(n_9202)
);

BUFx2_ASAP7_75t_L g9203 ( 
.A(n_7923),
.Y(n_9203)
);

INVx1_ASAP7_75t_L g9204 ( 
.A(n_8190),
.Y(n_9204)
);

AO21x2_ASAP7_75t_L g9205 ( 
.A1(n_7338),
.A2(n_6444),
.B(n_6441),
.Y(n_9205)
);

INVx1_ASAP7_75t_L g9206 ( 
.A(n_8204),
.Y(n_9206)
);

AND2x2_ASAP7_75t_L g9207 ( 
.A(n_7317),
.B(n_6773),
.Y(n_9207)
);

INVx2_ASAP7_75t_L g9208 ( 
.A(n_8005),
.Y(n_9208)
);

INVx2_ASAP7_75t_L g9209 ( 
.A(n_8005),
.Y(n_9209)
);

AOI22xp5_ASAP7_75t_L g9210 ( 
.A1(n_7722),
.A2(n_7437),
.B1(n_7352),
.B2(n_7595),
.Y(n_9210)
);

INVx2_ASAP7_75t_L g9211 ( 
.A(n_7958),
.Y(n_9211)
);

BUFx2_ASAP7_75t_SL g9212 ( 
.A(n_7422),
.Y(n_9212)
);

AOI21x1_ASAP7_75t_L g9213 ( 
.A1(n_7315),
.A2(n_7144),
.B(n_6805),
.Y(n_9213)
);

AND2x2_ASAP7_75t_L g9214 ( 
.A(n_7345),
.B(n_6799),
.Y(n_9214)
);

INVxp67_ASAP7_75t_L g9215 ( 
.A(n_7932),
.Y(n_9215)
);

CKINVDCx11_ASAP7_75t_R g9216 ( 
.A(n_7422),
.Y(n_9216)
);

AND2x2_ASAP7_75t_L g9217 ( 
.A(n_7345),
.B(n_6814),
.Y(n_9217)
);

INVx2_ASAP7_75t_L g9218 ( 
.A(n_7958),
.Y(n_9218)
);

INVx1_ASAP7_75t_L g9219 ( 
.A(n_8204),
.Y(n_9219)
);

INVx2_ASAP7_75t_L g9220 ( 
.A(n_7958),
.Y(n_9220)
);

OAI22xp5_ASAP7_75t_L g9221 ( 
.A1(n_7961),
.A2(n_7020),
.B1(n_7053),
.B2(n_6952),
.Y(n_9221)
);

AND2x2_ASAP7_75t_L g9222 ( 
.A(n_7345),
.B(n_6952),
.Y(n_9222)
);

NAND2x1p5_ASAP7_75t_L g9223 ( 
.A(n_7442),
.B(n_7105),
.Y(n_9223)
);

AO21x1_ASAP7_75t_L g9224 ( 
.A1(n_7315),
.A2(n_7360),
.B(n_7349),
.Y(n_9224)
);

INVx1_ASAP7_75t_SL g9225 ( 
.A(n_7742),
.Y(n_9225)
);

INVx1_ASAP7_75t_L g9226 ( 
.A(n_8214),
.Y(n_9226)
);

AOI22xp33_ASAP7_75t_L g9227 ( 
.A1(n_7595),
.A2(n_7905),
.B1(n_7691),
.B2(n_7961),
.Y(n_9227)
);

BUFx3_ASAP7_75t_L g9228 ( 
.A(n_8297),
.Y(n_9228)
);

NAND2xp5_ASAP7_75t_L g9229 ( 
.A(n_7565),
.B(n_6727),
.Y(n_9229)
);

BUFx3_ASAP7_75t_L g9230 ( 
.A(n_7943),
.Y(n_9230)
);

BUFx12f_ASAP7_75t_L g9231 ( 
.A(n_8134),
.Y(n_9231)
);

INVx3_ASAP7_75t_L g9232 ( 
.A(n_7505),
.Y(n_9232)
);

INVx8_ASAP7_75t_L g9233 ( 
.A(n_7271),
.Y(n_9233)
);

INVx1_ASAP7_75t_L g9234 ( 
.A(n_8214),
.Y(n_9234)
);

INVx2_ASAP7_75t_L g9235 ( 
.A(n_7958),
.Y(n_9235)
);

INVx2_ASAP7_75t_L g9236 ( 
.A(n_7958),
.Y(n_9236)
);

NAND2xp5_ASAP7_75t_L g9237 ( 
.A(n_7583),
.B(n_6776),
.Y(n_9237)
);

INVx11_ASAP7_75t_L g9238 ( 
.A(n_7271),
.Y(n_9238)
);

INVx1_ASAP7_75t_L g9239 ( 
.A(n_8217),
.Y(n_9239)
);

AND2x2_ASAP7_75t_L g9240 ( 
.A(n_7347),
.B(n_6952),
.Y(n_9240)
);

INVx1_ASAP7_75t_L g9241 ( 
.A(n_8217),
.Y(n_9241)
);

INVx2_ASAP7_75t_L g9242 ( 
.A(n_7958),
.Y(n_9242)
);

HB1xp67_ASAP7_75t_L g9243 ( 
.A(n_8011),
.Y(n_9243)
);

INVx1_ASAP7_75t_L g9244 ( 
.A(n_8219),
.Y(n_9244)
);

INVx2_ASAP7_75t_L g9245 ( 
.A(n_8007),
.Y(n_9245)
);

HB1xp67_ASAP7_75t_L g9246 ( 
.A(n_8011),
.Y(n_9246)
);

INVx1_ASAP7_75t_L g9247 ( 
.A(n_8219),
.Y(n_9247)
);

OAI22xp5_ASAP7_75t_L g9248 ( 
.A1(n_7297),
.A2(n_7053),
.B1(n_7062),
.B2(n_7020),
.Y(n_9248)
);

INVx1_ASAP7_75t_L g9249 ( 
.A(n_8252),
.Y(n_9249)
);

INVx2_ASAP7_75t_L g9250 ( 
.A(n_8007),
.Y(n_9250)
);

INVx1_ASAP7_75t_L g9251 ( 
.A(n_8252),
.Y(n_9251)
);

AO21x1_ASAP7_75t_SL g9252 ( 
.A1(n_8120),
.A2(n_6602),
.B(n_6550),
.Y(n_9252)
);

INVx1_ASAP7_75t_L g9253 ( 
.A(n_8253),
.Y(n_9253)
);

INVx2_ASAP7_75t_L g9254 ( 
.A(n_8007),
.Y(n_9254)
);

INVx2_ASAP7_75t_L g9255 ( 
.A(n_8007),
.Y(n_9255)
);

INVx1_ASAP7_75t_L g9256 ( 
.A(n_8253),
.Y(n_9256)
);

INVx2_ASAP7_75t_L g9257 ( 
.A(n_8007),
.Y(n_9257)
);

INVx1_ASAP7_75t_L g9258 ( 
.A(n_8262),
.Y(n_9258)
);

INVx1_ASAP7_75t_L g9259 ( 
.A(n_8262),
.Y(n_9259)
);

INVx1_ASAP7_75t_L g9260 ( 
.A(n_8267),
.Y(n_9260)
);

INVx2_ASAP7_75t_L g9261 ( 
.A(n_8007),
.Y(n_9261)
);

AO21x1_ASAP7_75t_L g9262 ( 
.A1(n_7360),
.A2(n_6363),
.B(n_6322),
.Y(n_9262)
);

INVx1_ASAP7_75t_L g9263 ( 
.A(n_8267),
.Y(n_9263)
);

INVx2_ASAP7_75t_L g9264 ( 
.A(n_7733),
.Y(n_9264)
);

INVx2_ASAP7_75t_L g9265 ( 
.A(n_7733),
.Y(n_9265)
);

INVx2_ASAP7_75t_L g9266 ( 
.A(n_7733),
.Y(n_9266)
);

INVx1_ASAP7_75t_L g9267 ( 
.A(n_8272),
.Y(n_9267)
);

INVx1_ASAP7_75t_L g9268 ( 
.A(n_8272),
.Y(n_9268)
);

INVx3_ASAP7_75t_L g9269 ( 
.A(n_7505),
.Y(n_9269)
);

INVx2_ASAP7_75t_L g9270 ( 
.A(n_7733),
.Y(n_9270)
);

AOI21x1_ASAP7_75t_L g9271 ( 
.A1(n_8075),
.A2(n_6805),
.B(n_6767),
.Y(n_9271)
);

AOI21xp33_ASAP7_75t_L g9272 ( 
.A1(n_7583),
.A2(n_6372),
.B(n_6363),
.Y(n_9272)
);

AO21x1_ASAP7_75t_L g9273 ( 
.A1(n_8054),
.A2(n_6372),
.B(n_6550),
.Y(n_9273)
);

INVx1_ASAP7_75t_L g9274 ( 
.A(n_8277),
.Y(n_9274)
);

INVx2_ASAP7_75t_L g9275 ( 
.A(n_7733),
.Y(n_9275)
);

INVx2_ASAP7_75t_L g9276 ( 
.A(n_7733),
.Y(n_9276)
);

AOI21x1_ASAP7_75t_L g9277 ( 
.A1(n_8075),
.A2(n_8235),
.B(n_8159),
.Y(n_9277)
);

INVxp33_ASAP7_75t_L g9278 ( 
.A(n_8071),
.Y(n_9278)
);

BUFx6f_ASAP7_75t_L g9279 ( 
.A(n_7923),
.Y(n_9279)
);

OAI21x1_ASAP7_75t_L g9280 ( 
.A1(n_7680),
.A2(n_6502),
.B(n_6491),
.Y(n_9280)
);

INVx6_ASAP7_75t_L g9281 ( 
.A(n_7892),
.Y(n_9281)
);

OAI22xp33_ASAP7_75t_L g9282 ( 
.A1(n_8171),
.A2(n_6809),
.B1(n_6450),
.B2(n_6714),
.Y(n_9282)
);

AOI21x1_ASAP7_75t_L g9283 ( 
.A1(n_8075),
.A2(n_7144),
.B(n_6813),
.Y(n_9283)
);

HB1xp67_ASAP7_75t_L g9284 ( 
.A(n_8047),
.Y(n_9284)
);

OAI22xp5_ASAP7_75t_L g9285 ( 
.A1(n_7722),
.A2(n_7053),
.B1(n_7062),
.B2(n_7020),
.Y(n_9285)
);

INVx1_ASAP7_75t_L g9286 ( 
.A(n_8277),
.Y(n_9286)
);

INVx1_ASAP7_75t_SL g9287 ( 
.A(n_7809),
.Y(n_9287)
);

AOI22xp33_ASAP7_75t_L g9288 ( 
.A1(n_7905),
.A2(n_6838),
.B1(n_6859),
.B2(n_6714),
.Y(n_9288)
);

INVx4_ASAP7_75t_SL g9289 ( 
.A(n_7179),
.Y(n_9289)
);

INVx1_ASAP7_75t_L g9290 ( 
.A(n_8280),
.Y(n_9290)
);

INVx3_ASAP7_75t_L g9291 ( 
.A(n_7505),
.Y(n_9291)
);

AND2x4_ASAP7_75t_L g9292 ( 
.A(n_8066),
.B(n_6128),
.Y(n_9292)
);

OAI22xp33_ASAP7_75t_L g9293 ( 
.A1(n_7308),
.A2(n_6809),
.B1(n_6450),
.B2(n_6714),
.Y(n_9293)
);

OA21x2_ASAP7_75t_L g9294 ( 
.A1(n_7196),
.A2(n_6813),
.B(n_6767),
.Y(n_9294)
);

INVx6_ASAP7_75t_L g9295 ( 
.A(n_7892),
.Y(n_9295)
);

INVx1_ASAP7_75t_L g9296 ( 
.A(n_8280),
.Y(n_9296)
);

AND2x4_ASAP7_75t_L g9297 ( 
.A(n_8130),
.B(n_6128),
.Y(n_9297)
);

AOI21x1_ASAP7_75t_L g9298 ( 
.A1(n_8159),
.A2(n_6820),
.B(n_6813),
.Y(n_9298)
);

OR2x6_ASAP7_75t_L g9299 ( 
.A(n_7504),
.B(n_6654),
.Y(n_9299)
);

INVx2_ASAP7_75t_L g9300 ( 
.A(n_7226),
.Y(n_9300)
);

INVxp67_ASAP7_75t_L g9301 ( 
.A(n_7932),
.Y(n_9301)
);

INVx2_ASAP7_75t_L g9302 ( 
.A(n_7226),
.Y(n_9302)
);

AOI21x1_ASAP7_75t_L g9303 ( 
.A1(n_8159),
.A2(n_6824),
.B(n_6820),
.Y(n_9303)
);

AND2x2_ASAP7_75t_L g9304 ( 
.A(n_7347),
.B(n_7062),
.Y(n_9304)
);

BUFx2_ASAP7_75t_L g9305 ( 
.A(n_7923),
.Y(n_9305)
);

OAI21xp5_ASAP7_75t_L g9306 ( 
.A1(n_7749),
.A2(n_7101),
.B(n_7093),
.Y(n_9306)
);

NAND2xp5_ASAP7_75t_L g9307 ( 
.A(n_8131),
.B(n_6776),
.Y(n_9307)
);

OAI21x1_ASAP7_75t_L g9308 ( 
.A1(n_7680),
.A2(n_6502),
.B(n_6491),
.Y(n_9308)
);

AOI22xp33_ASAP7_75t_L g9309 ( 
.A1(n_7691),
.A2(n_6838),
.B1(n_6859),
.B2(n_6714),
.Y(n_9309)
);

INVx1_ASAP7_75t_L g9310 ( 
.A(n_8292),
.Y(n_9310)
);

INVx1_ASAP7_75t_L g9311 ( 
.A(n_8292),
.Y(n_9311)
);

BUFx2_ASAP7_75t_L g9312 ( 
.A(n_7923),
.Y(n_9312)
);

CKINVDCx5p33_ASAP7_75t_R g9313 ( 
.A(n_8071),
.Y(n_9313)
);

INVx3_ASAP7_75t_L g9314 ( 
.A(n_7505),
.Y(n_9314)
);

BUFx2_ASAP7_75t_L g9315 ( 
.A(n_7923),
.Y(n_9315)
);

INVx1_ASAP7_75t_L g9316 ( 
.A(n_7163),
.Y(n_9316)
);

AO21x2_ASAP7_75t_L g9317 ( 
.A1(n_7338),
.A2(n_6444),
.B(n_6441),
.Y(n_9317)
);

INVxp33_ASAP7_75t_L g9318 ( 
.A(n_7836),
.Y(n_9318)
);

INVx1_ASAP7_75t_L g9319 ( 
.A(n_7163),
.Y(n_9319)
);

HB1xp67_ASAP7_75t_L g9320 ( 
.A(n_8047),
.Y(n_9320)
);

INVx1_ASAP7_75t_L g9321 ( 
.A(n_7163),
.Y(n_9321)
);

OA21x2_ASAP7_75t_L g9322 ( 
.A1(n_7289),
.A2(n_6824),
.B(n_6820),
.Y(n_9322)
);

INVx4_ASAP7_75t_L g9323 ( 
.A(n_8134),
.Y(n_9323)
);

INVx2_ASAP7_75t_L g9324 ( 
.A(n_7226),
.Y(n_9324)
);

INVx1_ASAP7_75t_L g9325 ( 
.A(n_7258),
.Y(n_9325)
);

INVx3_ASAP7_75t_L g9326 ( 
.A(n_7890),
.Y(n_9326)
);

INVx2_ASAP7_75t_L g9327 ( 
.A(n_8037),
.Y(n_9327)
);

BUFx2_ASAP7_75t_L g9328 ( 
.A(n_7923),
.Y(n_9328)
);

OR2x2_ASAP7_75t_L g9329 ( 
.A(n_8048),
.B(n_6446),
.Y(n_9329)
);

INVx2_ASAP7_75t_L g9330 ( 
.A(n_8041),
.Y(n_9330)
);

INVx1_ASAP7_75t_SL g9331 ( 
.A(n_7809),
.Y(n_9331)
);

AOI22xp33_ASAP7_75t_L g9332 ( 
.A1(n_7763),
.A2(n_6838),
.B1(n_6859),
.B2(n_6714),
.Y(n_9332)
);

INVx2_ASAP7_75t_L g9333 ( 
.A(n_8041),
.Y(n_9333)
);

BUFx2_ASAP7_75t_L g9334 ( 
.A(n_7923),
.Y(n_9334)
);

INVx3_ASAP7_75t_L g9335 ( 
.A(n_7890),
.Y(n_9335)
);

INVx3_ASAP7_75t_L g9336 ( 
.A(n_7890),
.Y(n_9336)
);

AO21x1_ASAP7_75t_L g9337 ( 
.A1(n_8054),
.A2(n_6613),
.B(n_6602),
.Y(n_9337)
);

AOI222xp33_ASAP7_75t_L g9338 ( 
.A1(n_7886),
.A2(n_7089),
.B1(n_5584),
.B2(n_5548),
.C1(n_5551),
.C2(n_5543),
.Y(n_9338)
);

HB1xp67_ASAP7_75t_L g9339 ( 
.A(n_8058),
.Y(n_9339)
);

INVxp67_ASAP7_75t_SL g9340 ( 
.A(n_7823),
.Y(n_9340)
);

OA21x2_ASAP7_75t_L g9341 ( 
.A1(n_7289),
.A2(n_6839),
.B(n_6824),
.Y(n_9341)
);

AOI22xp33_ASAP7_75t_L g9342 ( 
.A1(n_7763),
.A2(n_6838),
.B1(n_6859),
.B2(n_6714),
.Y(n_9342)
);

INVxp67_ASAP7_75t_L g9343 ( 
.A(n_8286),
.Y(n_9343)
);

INVx1_ASAP7_75t_L g9344 ( 
.A(n_7258),
.Y(n_9344)
);

INVx1_ASAP7_75t_L g9345 ( 
.A(n_7258),
.Y(n_9345)
);

BUFx6f_ASAP7_75t_L g9346 ( 
.A(n_7923),
.Y(n_9346)
);

NAND2x1_ASAP7_75t_L g9347 ( 
.A(n_7586),
.B(n_7073),
.Y(n_9347)
);

INVx1_ASAP7_75t_L g9348 ( 
.A(n_7260),
.Y(n_9348)
);

OR2x2_ASAP7_75t_L g9349 ( 
.A(n_7414),
.B(n_6446),
.Y(n_9349)
);

INVx3_ASAP7_75t_L g9350 ( 
.A(n_7890),
.Y(n_9350)
);

HB1xp67_ASAP7_75t_L g9351 ( 
.A(n_8058),
.Y(n_9351)
);

INVx1_ASAP7_75t_L g9352 ( 
.A(n_7260),
.Y(n_9352)
);

INVx1_ASAP7_75t_SL g9353 ( 
.A(n_7843),
.Y(n_9353)
);

INVx2_ASAP7_75t_L g9354 ( 
.A(n_8041),
.Y(n_9354)
);

BUFx10_ASAP7_75t_L g9355 ( 
.A(n_8021),
.Y(n_9355)
);

BUFx2_ASAP7_75t_L g9356 ( 
.A(n_8148),
.Y(n_9356)
);

INVx1_ASAP7_75t_L g9357 ( 
.A(n_7260),
.Y(n_9357)
);

HB1xp67_ASAP7_75t_L g9358 ( 
.A(n_8065),
.Y(n_9358)
);

INVx1_ASAP7_75t_L g9359 ( 
.A(n_7274),
.Y(n_9359)
);

INVx1_ASAP7_75t_L g9360 ( 
.A(n_7274),
.Y(n_9360)
);

INVx2_ASAP7_75t_L g9361 ( 
.A(n_8041),
.Y(n_9361)
);

INVx3_ASAP7_75t_L g9362 ( 
.A(n_7890),
.Y(n_9362)
);

OA21x2_ASAP7_75t_L g9363 ( 
.A1(n_7289),
.A2(n_6852),
.B(n_6839),
.Y(n_9363)
);

OAI21x1_ASAP7_75t_L g9364 ( 
.A1(n_7508),
.A2(n_6502),
.B(n_6491),
.Y(n_9364)
);

AND2x4_ASAP7_75t_L g9365 ( 
.A(n_8130),
.B(n_6210),
.Y(n_9365)
);

AOI22xp33_ASAP7_75t_SL g9366 ( 
.A1(n_7593),
.A2(n_7601),
.B1(n_7535),
.B2(n_7491),
.Y(n_9366)
);

OAI22xp5_ASAP7_75t_L g9367 ( 
.A1(n_7860),
.A2(n_7096),
.B1(n_7108),
.B2(n_7073),
.Y(n_9367)
);

OAI21x1_ASAP7_75t_L g9368 ( 
.A1(n_7508),
.A2(n_6532),
.B(n_6502),
.Y(n_9368)
);

INVxp67_ASAP7_75t_L g9369 ( 
.A(n_8286),
.Y(n_9369)
);

INVx1_ASAP7_75t_L g9370 ( 
.A(n_7274),
.Y(n_9370)
);

INVx1_ASAP7_75t_L g9371 ( 
.A(n_7278),
.Y(n_9371)
);

AO21x1_ASAP7_75t_SL g9372 ( 
.A1(n_8044),
.A2(n_6616),
.B(n_6613),
.Y(n_9372)
);

OAI21x1_ASAP7_75t_L g9373 ( 
.A1(n_7509),
.A2(n_6532),
.B(n_6502),
.Y(n_9373)
);

HB1xp67_ASAP7_75t_L g9374 ( 
.A(n_8065),
.Y(n_9374)
);

INVx4_ASAP7_75t_L g9375 ( 
.A(n_8134),
.Y(n_9375)
);

OA21x2_ASAP7_75t_L g9376 ( 
.A1(n_7293),
.A2(n_6852),
.B(n_6839),
.Y(n_9376)
);

OAI21xp5_ASAP7_75t_L g9377 ( 
.A1(n_7230),
.A2(n_7123),
.B(n_7122),
.Y(n_9377)
);

INVx3_ASAP7_75t_L g9378 ( 
.A(n_7890),
.Y(n_9378)
);

OAI21x1_ASAP7_75t_L g9379 ( 
.A1(n_7509),
.A2(n_6536),
.B(n_6532),
.Y(n_9379)
);

AOI22xp33_ASAP7_75t_SL g9380 ( 
.A1(n_7593),
.A2(n_7112),
.B1(n_6630),
.B2(n_6450),
.Y(n_9380)
);

INVx2_ASAP7_75t_L g9381 ( 
.A(n_8041),
.Y(n_9381)
);

INVx2_ASAP7_75t_L g9382 ( 
.A(n_8049),
.Y(n_9382)
);

AOI21xp5_ASAP7_75t_L g9383 ( 
.A1(n_7430),
.A2(n_6627),
.B(n_6616),
.Y(n_9383)
);

INVx1_ASAP7_75t_L g9384 ( 
.A(n_7278),
.Y(n_9384)
);

OAI22xp33_ASAP7_75t_L g9385 ( 
.A1(n_7308),
.A2(n_6450),
.B1(n_6860),
.B2(n_6686),
.Y(n_9385)
);

AOI21xp5_ASAP7_75t_SL g9386 ( 
.A1(n_7769),
.A2(n_7111),
.B(n_6450),
.Y(n_9386)
);

INVx4_ASAP7_75t_L g9387 ( 
.A(n_8134),
.Y(n_9387)
);

AOI22xp33_ASAP7_75t_SL g9388 ( 
.A1(n_7593),
.A2(n_6630),
.B1(n_6135),
.B2(n_6516),
.Y(n_9388)
);

BUFx6f_ASAP7_75t_L g9389 ( 
.A(n_8134),
.Y(n_9389)
);

BUFx3_ASAP7_75t_L g9390 ( 
.A(n_7943),
.Y(n_9390)
);

CKINVDCx5p33_ASAP7_75t_R g9391 ( 
.A(n_8021),
.Y(n_9391)
);

HB1xp67_ASAP7_75t_L g9392 ( 
.A(n_8070),
.Y(n_9392)
);

INVx1_ASAP7_75t_L g9393 ( 
.A(n_7278),
.Y(n_9393)
);

INVx1_ASAP7_75t_L g9394 ( 
.A(n_7290),
.Y(n_9394)
);

INVx2_ASAP7_75t_L g9395 ( 
.A(n_8049),
.Y(n_9395)
);

AND2x2_ASAP7_75t_L g9396 ( 
.A(n_7347),
.B(n_7073),
.Y(n_9396)
);

AND2x2_ASAP7_75t_L g9397 ( 
.A(n_7350),
.B(n_7096),
.Y(n_9397)
);

INVx2_ASAP7_75t_L g9398 ( 
.A(n_8049),
.Y(n_9398)
);

AND2x4_ASAP7_75t_L g9399 ( 
.A(n_8130),
.B(n_6210),
.Y(n_9399)
);

INVx1_ASAP7_75t_L g9400 ( 
.A(n_7290),
.Y(n_9400)
);

INVx1_ASAP7_75t_L g9401 ( 
.A(n_7290),
.Y(n_9401)
);

INVx2_ASAP7_75t_L g9402 ( 
.A(n_8049),
.Y(n_9402)
);

AOI22xp33_ASAP7_75t_L g9403 ( 
.A1(n_7706),
.A2(n_7800),
.B1(n_7593),
.B2(n_7601),
.Y(n_9403)
);

INVx1_ASAP7_75t_L g9404 ( 
.A(n_7295),
.Y(n_9404)
);

AOI22xp33_ASAP7_75t_L g9405 ( 
.A1(n_7706),
.A2(n_6860),
.B1(n_4420),
.B2(n_4429),
.Y(n_9405)
);

BUFx4_ASAP7_75t_SL g9406 ( 
.A(n_7943),
.Y(n_9406)
);

INVx2_ASAP7_75t_L g9407 ( 
.A(n_8049),
.Y(n_9407)
);

INVx1_ASAP7_75t_L g9408 ( 
.A(n_7295),
.Y(n_9408)
);

AOI22xp33_ASAP7_75t_L g9409 ( 
.A1(n_7800),
.A2(n_7601),
.B1(n_7616),
.B2(n_7377),
.Y(n_9409)
);

OAI21x1_ASAP7_75t_L g9410 ( 
.A1(n_7509),
.A2(n_6536),
.B(n_6532),
.Y(n_9410)
);

AND2x2_ASAP7_75t_L g9411 ( 
.A(n_7350),
.B(n_7096),
.Y(n_9411)
);

AOI22xp33_ASAP7_75t_L g9412 ( 
.A1(n_7601),
.A2(n_6860),
.B1(n_4420),
.B2(n_4429),
.Y(n_9412)
);

INVx2_ASAP7_75t_L g9413 ( 
.A(n_8154),
.Y(n_9413)
);

INVx1_ASAP7_75t_L g9414 ( 
.A(n_7295),
.Y(n_9414)
);

INVx2_ASAP7_75t_L g9415 ( 
.A(n_8154),
.Y(n_9415)
);

BUFx3_ASAP7_75t_L g9416 ( 
.A(n_7943),
.Y(n_9416)
);

INVx1_ASAP7_75t_L g9417 ( 
.A(n_7446),
.Y(n_9417)
);

CKINVDCx11_ASAP7_75t_R g9418 ( 
.A(n_7892),
.Y(n_9418)
);

BUFx3_ASAP7_75t_L g9419 ( 
.A(n_7979),
.Y(n_9419)
);

CKINVDCx11_ASAP7_75t_R g9420 ( 
.A(n_7892),
.Y(n_9420)
);

INVx2_ASAP7_75t_SL g9421 ( 
.A(n_7582),
.Y(n_9421)
);

INVx2_ASAP7_75t_L g9422 ( 
.A(n_8154),
.Y(n_9422)
);

BUFx4f_ASAP7_75t_SL g9423 ( 
.A(n_7892),
.Y(n_9423)
);

INVx1_ASAP7_75t_L g9424 ( 
.A(n_7446),
.Y(n_9424)
);

INVx1_ASAP7_75t_L g9425 ( 
.A(n_7446),
.Y(n_9425)
);

INVx1_ASAP7_75t_L g9426 ( 
.A(n_7614),
.Y(n_9426)
);

INVx1_ASAP7_75t_L g9427 ( 
.A(n_7614),
.Y(n_9427)
);

CKINVDCx20_ASAP7_75t_R g9428 ( 
.A(n_7795),
.Y(n_9428)
);

BUFx2_ASAP7_75t_L g9429 ( 
.A(n_8148),
.Y(n_9429)
);

BUFx2_ASAP7_75t_L g9430 ( 
.A(n_8148),
.Y(n_9430)
);

OA21x2_ASAP7_75t_L g9431 ( 
.A1(n_7293),
.A2(n_6862),
.B(n_6852),
.Y(n_9431)
);

BUFx6f_ASAP7_75t_L g9432 ( 
.A(n_8271),
.Y(n_9432)
);

INVx1_ASAP7_75t_L g9433 ( 
.A(n_7614),
.Y(n_9433)
);

BUFx6f_ASAP7_75t_L g9434 ( 
.A(n_8271),
.Y(n_9434)
);

INVx1_ASAP7_75t_L g9435 ( 
.A(n_7617),
.Y(n_9435)
);

INVx2_ASAP7_75t_L g9436 ( 
.A(n_8154),
.Y(n_9436)
);

INVx2_ASAP7_75t_L g9437 ( 
.A(n_8395),
.Y(n_9437)
);

AOI22xp33_ASAP7_75t_L g9438 ( 
.A1(n_8587),
.A2(n_7377),
.B1(n_7355),
.B2(n_7470),
.Y(n_9438)
);

INVx1_ASAP7_75t_L g9439 ( 
.A(n_8307),
.Y(n_9439)
);

INVx2_ASAP7_75t_L g9440 ( 
.A(n_8395),
.Y(n_9440)
);

OR2x6_ASAP7_75t_L g9441 ( 
.A(n_8429),
.B(n_8271),
.Y(n_9441)
);

AOI21x1_ASAP7_75t_L g9442 ( 
.A1(n_8453),
.A2(n_8261),
.B(n_8235),
.Y(n_9442)
);

OAI21x1_ASAP7_75t_L g9443 ( 
.A1(n_8337),
.A2(n_7641),
.B(n_7269),
.Y(n_9443)
);

CKINVDCx5p33_ASAP7_75t_R g9444 ( 
.A(n_8340),
.Y(n_9444)
);

NOR2xp33_ASAP7_75t_L g9445 ( 
.A(n_8334),
.B(n_7970),
.Y(n_9445)
);

INVx1_ASAP7_75t_L g9446 ( 
.A(n_8307),
.Y(n_9446)
);

OAI21x1_ASAP7_75t_L g9447 ( 
.A1(n_8337),
.A2(n_7641),
.B(n_7269),
.Y(n_9447)
);

AND2x2_ASAP7_75t_L g9448 ( 
.A(n_8993),
.B(n_8148),
.Y(n_9448)
);

OAI21x1_ASAP7_75t_L g9449 ( 
.A1(n_8337),
.A2(n_7641),
.B(n_7615),
.Y(n_9449)
);

INVx1_ASAP7_75t_L g9450 ( 
.A(n_8310),
.Y(n_9450)
);

HB1xp67_ASAP7_75t_L g9451 ( 
.A(n_9169),
.Y(n_9451)
);

INVx2_ASAP7_75t_L g9452 ( 
.A(n_8395),
.Y(n_9452)
);

CKINVDCx16_ASAP7_75t_R g9453 ( 
.A(n_8334),
.Y(n_9453)
);

INVx2_ASAP7_75t_L g9454 ( 
.A(n_8410),
.Y(n_9454)
);

INVx3_ASAP7_75t_L g9455 ( 
.A(n_9279),
.Y(n_9455)
);

OA21x2_ASAP7_75t_L g9456 ( 
.A1(n_8873),
.A2(n_7319),
.B(n_7293),
.Y(n_9456)
);

BUFx2_ASAP7_75t_L g9457 ( 
.A(n_8371),
.Y(n_9457)
);

INVxp33_ASAP7_75t_L g9458 ( 
.A(n_8372),
.Y(n_9458)
);

HB1xp67_ASAP7_75t_L g9459 ( 
.A(n_9225),
.Y(n_9459)
);

INVx1_ASAP7_75t_L g9460 ( 
.A(n_8310),
.Y(n_9460)
);

INVx2_ASAP7_75t_L g9461 ( 
.A(n_8410),
.Y(n_9461)
);

INVx2_ASAP7_75t_L g9462 ( 
.A(n_8410),
.Y(n_9462)
);

AND2x2_ASAP7_75t_L g9463 ( 
.A(n_8993),
.B(n_8148),
.Y(n_9463)
);

HB1xp67_ASAP7_75t_L g9464 ( 
.A(n_9287),
.Y(n_9464)
);

CKINVDCx9p33_ASAP7_75t_R g9465 ( 
.A(n_8453),
.Y(n_9465)
);

INVx1_ASAP7_75t_SL g9466 ( 
.A(n_8355),
.Y(n_9466)
);

BUFx2_ASAP7_75t_L g9467 ( 
.A(n_8371),
.Y(n_9467)
);

INVx2_ASAP7_75t_L g9468 ( 
.A(n_8515),
.Y(n_9468)
);

AND2x2_ASAP7_75t_L g9469 ( 
.A(n_9252),
.B(n_8148),
.Y(n_9469)
);

INVx2_ASAP7_75t_L g9470 ( 
.A(n_8515),
.Y(n_9470)
);

INVx1_ASAP7_75t_L g9471 ( 
.A(n_8313),
.Y(n_9471)
);

INVx1_ASAP7_75t_L g9472 ( 
.A(n_8313),
.Y(n_9472)
);

BUFx12f_ASAP7_75t_L g9473 ( 
.A(n_8834),
.Y(n_9473)
);

INVx1_ASAP7_75t_L g9474 ( 
.A(n_8324),
.Y(n_9474)
);

INVx1_ASAP7_75t_L g9475 ( 
.A(n_8324),
.Y(n_9475)
);

INVxp67_ASAP7_75t_L g9476 ( 
.A(n_8316),
.Y(n_9476)
);

INVx1_ASAP7_75t_L g9477 ( 
.A(n_8326),
.Y(n_9477)
);

INVx1_ASAP7_75t_L g9478 ( 
.A(n_8326),
.Y(n_9478)
);

INVx2_ASAP7_75t_L g9479 ( 
.A(n_8526),
.Y(n_9479)
);

AND2x2_ASAP7_75t_L g9480 ( 
.A(n_9252),
.B(n_8148),
.Y(n_9480)
);

HB1xp67_ASAP7_75t_L g9481 ( 
.A(n_9331),
.Y(n_9481)
);

HB1xp67_ASAP7_75t_L g9482 ( 
.A(n_9353),
.Y(n_9482)
);

INVx3_ASAP7_75t_L g9483 ( 
.A(n_9279),
.Y(n_9483)
);

BUFx2_ASAP7_75t_L g9484 ( 
.A(n_8447),
.Y(n_9484)
);

INVx1_ASAP7_75t_L g9485 ( 
.A(n_8328),
.Y(n_9485)
);

BUFx2_ASAP7_75t_L g9486 ( 
.A(n_8447),
.Y(n_9486)
);

INVx4_ASAP7_75t_L g9487 ( 
.A(n_8602),
.Y(n_9487)
);

INVx2_ASAP7_75t_L g9488 ( 
.A(n_8526),
.Y(n_9488)
);

INVx4_ASAP7_75t_L g9489 ( 
.A(n_8602),
.Y(n_9489)
);

INVx1_ASAP7_75t_L g9490 ( 
.A(n_8328),
.Y(n_9490)
);

INVx2_ASAP7_75t_L g9491 ( 
.A(n_8527),
.Y(n_9491)
);

INVx1_ASAP7_75t_L g9492 ( 
.A(n_8330),
.Y(n_9492)
);

INVx2_ASAP7_75t_SL g9493 ( 
.A(n_8619),
.Y(n_9493)
);

INVx3_ASAP7_75t_L g9494 ( 
.A(n_9279),
.Y(n_9494)
);

AOI22xp33_ASAP7_75t_L g9495 ( 
.A1(n_8549),
.A2(n_8693),
.B1(n_8773),
.B2(n_8576),
.Y(n_9495)
);

NAND2x1p5_ASAP7_75t_L g9496 ( 
.A(n_8497),
.B(n_8271),
.Y(n_9496)
);

AOI22xp33_ASAP7_75t_L g9497 ( 
.A1(n_8549),
.A2(n_7377),
.B1(n_7355),
.B2(n_7470),
.Y(n_9497)
);

AND2x4_ASAP7_75t_L g9498 ( 
.A(n_8502),
.B(n_7179),
.Y(n_9498)
);

INVx4_ASAP7_75t_L g9499 ( 
.A(n_8632),
.Y(n_9499)
);

A2O1A1Ixp33_ASAP7_75t_L g9500 ( 
.A1(n_8576),
.A2(n_7752),
.B(n_7823),
.C(n_7735),
.Y(n_9500)
);

INVx2_ASAP7_75t_L g9501 ( 
.A(n_8527),
.Y(n_9501)
);

AND2x4_ASAP7_75t_L g9502 ( 
.A(n_8502),
.B(n_7179),
.Y(n_9502)
);

INVx2_ASAP7_75t_L g9503 ( 
.A(n_8546),
.Y(n_9503)
);

INVx2_ASAP7_75t_L g9504 ( 
.A(n_8546),
.Y(n_9504)
);

INVx1_ASAP7_75t_L g9505 ( 
.A(n_8330),
.Y(n_9505)
);

INVx1_ASAP7_75t_L g9506 ( 
.A(n_8332),
.Y(n_9506)
);

BUFx2_ASAP7_75t_L g9507 ( 
.A(n_8632),
.Y(n_9507)
);

BUFx6f_ASAP7_75t_L g9508 ( 
.A(n_8484),
.Y(n_9508)
);

AO21x2_ASAP7_75t_L g9509 ( 
.A1(n_8467),
.A2(n_8060),
.B(n_8056),
.Y(n_9509)
);

AO21x1_ASAP7_75t_L g9510 ( 
.A1(n_8849),
.A2(n_8926),
.B(n_9191),
.Y(n_9510)
);

INVx1_ASAP7_75t_L g9511 ( 
.A(n_8332),
.Y(n_9511)
);

INVx1_ASAP7_75t_L g9512 ( 
.A(n_8348),
.Y(n_9512)
);

OR2x6_ASAP7_75t_L g9513 ( 
.A(n_8467),
.B(n_8271),
.Y(n_9513)
);

INVx1_ASAP7_75t_L g9514 ( 
.A(n_8348),
.Y(n_9514)
);

INVx1_ASAP7_75t_L g9515 ( 
.A(n_8351),
.Y(n_9515)
);

INVx1_ASAP7_75t_L g9516 ( 
.A(n_8351),
.Y(n_9516)
);

AOI22xp33_ASAP7_75t_L g9517 ( 
.A1(n_8693),
.A2(n_8795),
.B1(n_8825),
.B2(n_8773),
.Y(n_9517)
);

OAI21x1_ASAP7_75t_L g9518 ( 
.A1(n_8337),
.A2(n_7615),
.B(n_7634),
.Y(n_9518)
);

NAND2xp5_ASAP7_75t_L g9519 ( 
.A(n_9340),
.B(n_8059),
.Y(n_9519)
);

AOI21xp5_ASAP7_75t_L g9520 ( 
.A1(n_8314),
.A2(n_7654),
.B(n_7802),
.Y(n_9520)
);

INVx1_ASAP7_75t_L g9521 ( 
.A(n_8353),
.Y(n_9521)
);

AND2x2_ASAP7_75t_L g9522 ( 
.A(n_8778),
.B(n_8148),
.Y(n_9522)
);

INVx1_ASAP7_75t_L g9523 ( 
.A(n_8353),
.Y(n_9523)
);

INVx1_ASAP7_75t_L g9524 ( 
.A(n_8363),
.Y(n_9524)
);

BUFx2_ASAP7_75t_L g9525 ( 
.A(n_8738),
.Y(n_9525)
);

INVx1_ASAP7_75t_L g9526 ( 
.A(n_8363),
.Y(n_9526)
);

BUFx3_ASAP7_75t_L g9527 ( 
.A(n_8342),
.Y(n_9527)
);

OAI21x1_ASAP7_75t_L g9528 ( 
.A1(n_8344),
.A2(n_7615),
.B(n_7634),
.Y(n_9528)
);

HB1xp67_ASAP7_75t_L g9529 ( 
.A(n_8466),
.Y(n_9529)
);

NAND2xp5_ASAP7_75t_L g9530 ( 
.A(n_9383),
.B(n_8059),
.Y(n_9530)
);

INVx1_ASAP7_75t_L g9531 ( 
.A(n_8366),
.Y(n_9531)
);

INVx1_ASAP7_75t_L g9532 ( 
.A(n_8366),
.Y(n_9532)
);

INVx1_ASAP7_75t_L g9533 ( 
.A(n_8367),
.Y(n_9533)
);

INVx2_ASAP7_75t_SL g9534 ( 
.A(n_8619),
.Y(n_9534)
);

INVx1_ASAP7_75t_L g9535 ( 
.A(n_8367),
.Y(n_9535)
);

INVx2_ASAP7_75t_L g9536 ( 
.A(n_8667),
.Y(n_9536)
);

OAI22xp5_ASAP7_75t_L g9537 ( 
.A1(n_8702),
.A2(n_7834),
.B1(n_7193),
.B2(n_8304),
.Y(n_9537)
);

BUFx3_ASAP7_75t_L g9538 ( 
.A(n_8342),
.Y(n_9538)
);

HB1xp67_ASAP7_75t_L g9539 ( 
.A(n_8765),
.Y(n_9539)
);

AO222x2_ASAP7_75t_L g9540 ( 
.A1(n_8316),
.A2(n_7535),
.B1(n_7491),
.B2(n_7180),
.C1(n_7203),
.C2(n_7291),
.Y(n_9540)
);

INVx1_ASAP7_75t_L g9541 ( 
.A(n_8380),
.Y(n_9541)
);

AO21x2_ASAP7_75t_L g9542 ( 
.A1(n_9224),
.A2(n_8060),
.B(n_8056),
.Y(n_9542)
);

CKINVDCx11_ASAP7_75t_R g9543 ( 
.A(n_8365),
.Y(n_9543)
);

INVx2_ASAP7_75t_L g9544 ( 
.A(n_8667),
.Y(n_9544)
);

INVx1_ASAP7_75t_L g9545 ( 
.A(n_8380),
.Y(n_9545)
);

INVx2_ASAP7_75t_SL g9546 ( 
.A(n_8311),
.Y(n_9546)
);

INVx1_ASAP7_75t_L g9547 ( 
.A(n_8382),
.Y(n_9547)
);

INVx2_ASAP7_75t_L g9548 ( 
.A(n_8667),
.Y(n_9548)
);

HB1xp67_ASAP7_75t_L g9549 ( 
.A(n_8841),
.Y(n_9549)
);

NAND2x1p5_ASAP7_75t_L g9550 ( 
.A(n_8497),
.B(n_7979),
.Y(n_9550)
);

AND2x2_ASAP7_75t_L g9551 ( 
.A(n_8778),
.B(n_7350),
.Y(n_9551)
);

INVx1_ASAP7_75t_L g9552 ( 
.A(n_8382),
.Y(n_9552)
);

AND2x2_ASAP7_75t_L g9553 ( 
.A(n_8828),
.B(n_8235),
.Y(n_9553)
);

INVx1_ASAP7_75t_L g9554 ( 
.A(n_8394),
.Y(n_9554)
);

BUFx6f_ASAP7_75t_L g9555 ( 
.A(n_8484),
.Y(n_9555)
);

BUFx6f_ASAP7_75t_L g9556 ( 
.A(n_8484),
.Y(n_9556)
);

AOI22xp33_ASAP7_75t_L g9557 ( 
.A1(n_8795),
.A2(n_7377),
.B1(n_7355),
.B2(n_7470),
.Y(n_9557)
);

INVx1_ASAP7_75t_L g9558 ( 
.A(n_8394),
.Y(n_9558)
);

INVx2_ASAP7_75t_L g9559 ( 
.A(n_8668),
.Y(n_9559)
);

INVx1_ASAP7_75t_L g9560 ( 
.A(n_8396),
.Y(n_9560)
);

INVx2_ASAP7_75t_L g9561 ( 
.A(n_8668),
.Y(n_9561)
);

AOI21xp33_ASAP7_75t_L g9562 ( 
.A1(n_8826),
.A2(n_7377),
.B(n_7247),
.Y(n_9562)
);

INVx1_ASAP7_75t_L g9563 ( 
.A(n_8396),
.Y(n_9563)
);

INVx2_ASAP7_75t_L g9564 ( 
.A(n_8668),
.Y(n_9564)
);

INVx1_ASAP7_75t_L g9565 ( 
.A(n_8400),
.Y(n_9565)
);

INVx1_ASAP7_75t_L g9566 ( 
.A(n_8400),
.Y(n_9566)
);

OAI21x1_ASAP7_75t_SL g9567 ( 
.A1(n_8314),
.A2(n_7586),
.B(n_7563),
.Y(n_9567)
);

BUFx2_ASAP7_75t_L g9568 ( 
.A(n_8738),
.Y(n_9568)
);

INVx1_ASAP7_75t_L g9569 ( 
.A(n_8403),
.Y(n_9569)
);

AND2x2_ASAP7_75t_L g9570 ( 
.A(n_8828),
.B(n_8261),
.Y(n_9570)
);

INVx1_ASAP7_75t_L g9571 ( 
.A(n_8403),
.Y(n_9571)
);

AOI22xp33_ASAP7_75t_L g9572 ( 
.A1(n_8825),
.A2(n_7355),
.B1(n_7470),
.B2(n_7458),
.Y(n_9572)
);

INVxp67_ASAP7_75t_L g9573 ( 
.A(n_8561),
.Y(n_9573)
);

INVx1_ASAP7_75t_L g9574 ( 
.A(n_8405),
.Y(n_9574)
);

INVx2_ASAP7_75t_L g9575 ( 
.A(n_8672),
.Y(n_9575)
);

INVx1_ASAP7_75t_L g9576 ( 
.A(n_8405),
.Y(n_9576)
);

INVx1_ASAP7_75t_L g9577 ( 
.A(n_8414),
.Y(n_9577)
);

INVx2_ASAP7_75t_L g9578 ( 
.A(n_8672),
.Y(n_9578)
);

O2A1O1Ixp33_ASAP7_75t_SL g9579 ( 
.A1(n_8935),
.A2(n_8273),
.B(n_8259),
.C(n_8230),
.Y(n_9579)
);

AO21x2_ASAP7_75t_L g9580 ( 
.A1(n_9224),
.A2(n_8062),
.B(n_7997),
.Y(n_9580)
);

OR2x2_ASAP7_75t_L g9581 ( 
.A(n_9003),
.B(n_7280),
.Y(n_9581)
);

AND2x4_ASAP7_75t_L g9582 ( 
.A(n_8514),
.B(n_7179),
.Y(n_9582)
);

AND2x2_ASAP7_75t_L g9583 ( 
.A(n_8514),
.B(n_8261),
.Y(n_9583)
);

AND2x4_ASAP7_75t_L g9584 ( 
.A(n_8533),
.B(n_9289),
.Y(n_9584)
);

INVx2_ASAP7_75t_L g9585 ( 
.A(n_8672),
.Y(n_9585)
);

INVx1_ASAP7_75t_L g9586 ( 
.A(n_8414),
.Y(n_9586)
);

AND2x2_ASAP7_75t_L g9587 ( 
.A(n_8533),
.B(n_7335),
.Y(n_9587)
);

INVx2_ASAP7_75t_L g9588 ( 
.A(n_8673),
.Y(n_9588)
);

AND2x4_ASAP7_75t_L g9589 ( 
.A(n_9289),
.B(n_7179),
.Y(n_9589)
);

INVx1_ASAP7_75t_L g9590 ( 
.A(n_8416),
.Y(n_9590)
);

BUFx2_ASAP7_75t_L g9591 ( 
.A(n_8803),
.Y(n_9591)
);

INVx4_ASAP7_75t_SL g9592 ( 
.A(n_8803),
.Y(n_9592)
);

INVx1_ASAP7_75t_L g9593 ( 
.A(n_8416),
.Y(n_9593)
);

AO21x2_ASAP7_75t_L g9594 ( 
.A1(n_8826),
.A2(n_8062),
.B(n_7997),
.Y(n_9594)
);

AND2x2_ASAP7_75t_L g9595 ( 
.A(n_8876),
.B(n_7335),
.Y(n_9595)
);

INVx1_ASAP7_75t_L g9596 ( 
.A(n_8420),
.Y(n_9596)
);

INVx3_ASAP7_75t_L g9597 ( 
.A(n_9279),
.Y(n_9597)
);

NAND2xp5_ASAP7_75t_L g9598 ( 
.A(n_8956),
.B(n_8152),
.Y(n_9598)
);

INVx2_ASAP7_75t_L g9599 ( 
.A(n_8673),
.Y(n_9599)
);

OAI21x1_ASAP7_75t_L g9600 ( 
.A1(n_8344),
.A2(n_7637),
.B(n_7634),
.Y(n_9600)
);

INVx2_ASAP7_75t_L g9601 ( 
.A(n_8673),
.Y(n_9601)
);

INVx2_ASAP7_75t_L g9602 ( 
.A(n_8674),
.Y(n_9602)
);

BUFx6f_ASAP7_75t_L g9603 ( 
.A(n_8488),
.Y(n_9603)
);

OR2x2_ASAP7_75t_L g9604 ( 
.A(n_9003),
.B(n_7280),
.Y(n_9604)
);

HB1xp67_ASAP7_75t_L g9605 ( 
.A(n_8872),
.Y(n_9605)
);

OAI21xp5_ASAP7_75t_L g9606 ( 
.A1(n_8702),
.A2(n_8162),
.B(n_7451),
.Y(n_9606)
);

INVx2_ASAP7_75t_L g9607 ( 
.A(n_8674),
.Y(n_9607)
);

INVx1_ASAP7_75t_SL g9608 ( 
.A(n_8601),
.Y(n_9608)
);

OA21x2_ASAP7_75t_L g9609 ( 
.A1(n_8873),
.A2(n_7333),
.B(n_7319),
.Y(n_9609)
);

INVx1_ASAP7_75t_L g9610 ( 
.A(n_8420),
.Y(n_9610)
);

INVx2_ASAP7_75t_L g9611 ( 
.A(n_8674),
.Y(n_9611)
);

INVx2_ASAP7_75t_L g9612 ( 
.A(n_8777),
.Y(n_9612)
);

INVx1_ASAP7_75t_L g9613 ( 
.A(n_8422),
.Y(n_9613)
);

OAI21xp5_ASAP7_75t_L g9614 ( 
.A1(n_8361),
.A2(n_7451),
.B(n_7986),
.Y(n_9614)
);

HB1xp67_ASAP7_75t_L g9615 ( 
.A(n_8660),
.Y(n_9615)
);

OR2x6_ASAP7_75t_L g9616 ( 
.A(n_9103),
.B(n_7677),
.Y(n_9616)
);

INVx2_ASAP7_75t_SL g9617 ( 
.A(n_8311),
.Y(n_9617)
);

OR2x2_ASAP7_75t_L g9618 ( 
.A(n_9349),
.B(n_8131),
.Y(n_9618)
);

AND2x4_ASAP7_75t_L g9619 ( 
.A(n_9289),
.B(n_8994),
.Y(n_9619)
);

OR2x2_ASAP7_75t_L g9620 ( 
.A(n_9349),
.B(n_7511),
.Y(n_9620)
);

INVx1_ASAP7_75t_L g9621 ( 
.A(n_8422),
.Y(n_9621)
);

INVx2_ASAP7_75t_L g9622 ( 
.A(n_8777),
.Y(n_9622)
);

AOI22xp33_ASAP7_75t_L g9623 ( 
.A1(n_8956),
.A2(n_7355),
.B1(n_7470),
.B2(n_7458),
.Y(n_9623)
);

OAI21x1_ASAP7_75t_L g9624 ( 
.A1(n_8344),
.A2(n_7637),
.B(n_7464),
.Y(n_9624)
);

BUFx3_ASAP7_75t_L g9625 ( 
.A(n_8915),
.Y(n_9625)
);

INVx1_ASAP7_75t_L g9626 ( 
.A(n_8424),
.Y(n_9626)
);

INVx3_ASAP7_75t_L g9627 ( 
.A(n_9279),
.Y(n_9627)
);

INVx1_ASAP7_75t_L g9628 ( 
.A(n_8424),
.Y(n_9628)
);

INVx1_ASAP7_75t_L g9629 ( 
.A(n_8425),
.Y(n_9629)
);

INVx1_ASAP7_75t_L g9630 ( 
.A(n_8425),
.Y(n_9630)
);

AND2x2_ASAP7_75t_L g9631 ( 
.A(n_8876),
.B(n_7335),
.Y(n_9631)
);

INVx1_ASAP7_75t_L g9632 ( 
.A(n_8430),
.Y(n_9632)
);

AND2x4_ASAP7_75t_L g9633 ( 
.A(n_9289),
.B(n_7179),
.Y(n_9633)
);

BUFx6f_ASAP7_75t_L g9634 ( 
.A(n_8488),
.Y(n_9634)
);

INVx2_ASAP7_75t_L g9635 ( 
.A(n_8777),
.Y(n_9635)
);

INVx2_ASAP7_75t_L g9636 ( 
.A(n_8782),
.Y(n_9636)
);

INVx1_ASAP7_75t_L g9637 ( 
.A(n_8430),
.Y(n_9637)
);

HB1xp67_ASAP7_75t_L g9638 ( 
.A(n_8718),
.Y(n_9638)
);

NAND2xp5_ASAP7_75t_SL g9639 ( 
.A(n_8364),
.B(n_7682),
.Y(n_9639)
);

INVx1_ASAP7_75t_SL g9640 ( 
.A(n_8761),
.Y(n_9640)
);

INVx1_ASAP7_75t_L g9641 ( 
.A(n_8432),
.Y(n_9641)
);

BUFx2_ASAP7_75t_L g9642 ( 
.A(n_8787),
.Y(n_9642)
);

AOI21x1_ASAP7_75t_L g9643 ( 
.A1(n_8681),
.A2(n_8077),
.B(n_8070),
.Y(n_9643)
);

OR2x6_ASAP7_75t_L g9644 ( 
.A(n_9103),
.B(n_9299),
.Y(n_9644)
);

INVx1_ASAP7_75t_L g9645 ( 
.A(n_8432),
.Y(n_9645)
);

INVx2_ASAP7_75t_L g9646 ( 
.A(n_8782),
.Y(n_9646)
);

CKINVDCx11_ASAP7_75t_R g9647 ( 
.A(n_8365),
.Y(n_9647)
);

INVx1_ASAP7_75t_L g9648 ( 
.A(n_8436),
.Y(n_9648)
);

AO21x2_ASAP7_75t_L g9649 ( 
.A1(n_8826),
.A2(n_8015),
.B(n_7994),
.Y(n_9649)
);

AND2x2_ASAP7_75t_L g9650 ( 
.A(n_9372),
.B(n_7371),
.Y(n_9650)
);

INVx2_ASAP7_75t_L g9651 ( 
.A(n_8782),
.Y(n_9651)
);

INVx1_ASAP7_75t_L g9652 ( 
.A(n_8436),
.Y(n_9652)
);

INVx2_ASAP7_75t_L g9653 ( 
.A(n_8792),
.Y(n_9653)
);

INVx1_ASAP7_75t_L g9654 ( 
.A(n_8437),
.Y(n_9654)
);

INVx1_ASAP7_75t_L g9655 ( 
.A(n_8437),
.Y(n_9655)
);

CKINVDCx20_ASAP7_75t_R g9656 ( 
.A(n_8320),
.Y(n_9656)
);

INVx1_ASAP7_75t_L g9657 ( 
.A(n_8442),
.Y(n_9657)
);

NAND2xp5_ASAP7_75t_L g9658 ( 
.A(n_8987),
.B(n_8152),
.Y(n_9658)
);

OAI21x1_ASAP7_75t_L g9659 ( 
.A1(n_8344),
.A2(n_7637),
.B(n_7464),
.Y(n_9659)
);

AOI22xp5_ASAP7_75t_L g9660 ( 
.A1(n_8987),
.A2(n_8992),
.B1(n_9026),
.B2(n_9019),
.Y(n_9660)
);

AOI21xp33_ASAP7_75t_SL g9661 ( 
.A1(n_8787),
.A2(n_8902),
.B(n_8910),
.Y(n_9661)
);

AND2x2_ASAP7_75t_L g9662 ( 
.A(n_9372),
.B(n_7371),
.Y(n_9662)
);

INVx2_ASAP7_75t_L g9663 ( 
.A(n_8792),
.Y(n_9663)
);

BUFx2_ASAP7_75t_L g9664 ( 
.A(n_8309),
.Y(n_9664)
);

INVx2_ASAP7_75t_L g9665 ( 
.A(n_8792),
.Y(n_9665)
);

INVx3_ASAP7_75t_L g9666 ( 
.A(n_9279),
.Y(n_9666)
);

INVx2_ASAP7_75t_L g9667 ( 
.A(n_8794),
.Y(n_9667)
);

INVxp67_ASAP7_75t_L g9668 ( 
.A(n_8561),
.Y(n_9668)
);

HB1xp67_ASAP7_75t_L g9669 ( 
.A(n_9215),
.Y(n_9669)
);

AO31x2_ASAP7_75t_L g9670 ( 
.A1(n_8992),
.A2(n_7209),
.A3(n_7210),
.B(n_7183),
.Y(n_9670)
);

INVx1_ASAP7_75t_L g9671 ( 
.A(n_8442),
.Y(n_9671)
);

AO21x2_ASAP7_75t_L g9672 ( 
.A1(n_8364),
.A2(n_8015),
.B(n_7994),
.Y(n_9672)
);

AO21x2_ASAP7_75t_L g9673 ( 
.A1(n_8312),
.A2(n_7720),
.B(n_7698),
.Y(n_9673)
);

OAI21x1_ASAP7_75t_L g9674 ( 
.A1(n_8407),
.A2(n_7464),
.B(n_7441),
.Y(n_9674)
);

BUFx2_ASAP7_75t_L g9675 ( 
.A(n_8309),
.Y(n_9675)
);

NOR2xp33_ASAP7_75t_L g9676 ( 
.A(n_8441),
.B(n_7970),
.Y(n_9676)
);

AND2x2_ASAP7_75t_L g9677 ( 
.A(n_8850),
.B(n_7371),
.Y(n_9677)
);

INVx2_ASAP7_75t_L g9678 ( 
.A(n_8794),
.Y(n_9678)
);

INVx1_ASAP7_75t_L g9679 ( 
.A(n_8448),
.Y(n_9679)
);

OAI21x1_ASAP7_75t_L g9680 ( 
.A1(n_8407),
.A2(n_8417),
.B(n_8415),
.Y(n_9680)
);

INVx2_ASAP7_75t_L g9681 ( 
.A(n_8794),
.Y(n_9681)
);

NOR2xp33_ASAP7_75t_L g9682 ( 
.A(n_8712),
.B(n_7995),
.Y(n_9682)
);

INVx2_ASAP7_75t_L g9683 ( 
.A(n_8809),
.Y(n_9683)
);

INVx2_ASAP7_75t_L g9684 ( 
.A(n_8809),
.Y(n_9684)
);

INVxp33_ASAP7_75t_L g9685 ( 
.A(n_9200),
.Y(n_9685)
);

BUFx6f_ASAP7_75t_L g9686 ( 
.A(n_8488),
.Y(n_9686)
);

INVx1_ASAP7_75t_L g9687 ( 
.A(n_8448),
.Y(n_9687)
);

NAND2xp33_ASAP7_75t_SL g9688 ( 
.A(n_9056),
.B(n_7212),
.Y(n_9688)
);

AND2x2_ASAP7_75t_L g9689 ( 
.A(n_8850),
.B(n_7374),
.Y(n_9689)
);

INVx1_ASAP7_75t_L g9690 ( 
.A(n_8450),
.Y(n_9690)
);

BUFx2_ASAP7_75t_L g9691 ( 
.A(n_8309),
.Y(n_9691)
);

BUFx2_ASAP7_75t_L g9692 ( 
.A(n_8309),
.Y(n_9692)
);

INVx1_ASAP7_75t_L g9693 ( 
.A(n_8450),
.Y(n_9693)
);

INVx1_ASAP7_75t_L g9694 ( 
.A(n_8451),
.Y(n_9694)
);

INVx1_ASAP7_75t_L g9695 ( 
.A(n_8451),
.Y(n_9695)
);

CKINVDCx6p67_ASAP7_75t_R g9696 ( 
.A(n_8915),
.Y(n_9696)
);

INVx2_ASAP7_75t_L g9697 ( 
.A(n_8809),
.Y(n_9697)
);

INVx1_ASAP7_75t_L g9698 ( 
.A(n_8454),
.Y(n_9698)
);

HB1xp67_ASAP7_75t_SL g9699 ( 
.A(n_8377),
.Y(n_9699)
);

INVx1_ASAP7_75t_L g9700 ( 
.A(n_8454),
.Y(n_9700)
);

INVx2_ASAP7_75t_L g9701 ( 
.A(n_8813),
.Y(n_9701)
);

INVx2_ASAP7_75t_L g9702 ( 
.A(n_8813),
.Y(n_9702)
);

NAND2xp5_ASAP7_75t_L g9703 ( 
.A(n_9019),
.B(n_8173),
.Y(n_9703)
);

AND2x2_ASAP7_75t_L g9704 ( 
.A(n_9014),
.B(n_7374),
.Y(n_9704)
);

INVx1_ASAP7_75t_L g9705 ( 
.A(n_8470),
.Y(n_9705)
);

INVx2_ASAP7_75t_L g9706 ( 
.A(n_8813),
.Y(n_9706)
);

OAI21x1_ASAP7_75t_L g9707 ( 
.A1(n_8407),
.A2(n_7441),
.B(n_7895),
.Y(n_9707)
);

HB1xp67_ASAP7_75t_L g9708 ( 
.A(n_9301),
.Y(n_9708)
);

AOI21x1_ASAP7_75t_L g9709 ( 
.A1(n_8681),
.A2(n_8140),
.B(n_8077),
.Y(n_9709)
);

INVx1_ASAP7_75t_L g9710 ( 
.A(n_8470),
.Y(n_9710)
);

INVx2_ASAP7_75t_L g9711 ( 
.A(n_8816),
.Y(n_9711)
);

INVx1_ASAP7_75t_L g9712 ( 
.A(n_8475),
.Y(n_9712)
);

AOI21xp5_ASAP7_75t_SL g9713 ( 
.A1(n_9026),
.A2(n_8273),
.B(n_8259),
.Y(n_9713)
);

INVx3_ASAP7_75t_L g9714 ( 
.A(n_9346),
.Y(n_9714)
);

AND2x4_ASAP7_75t_L g9715 ( 
.A(n_9289),
.B(n_7179),
.Y(n_9715)
);

AOI21x1_ASAP7_75t_L g9716 ( 
.A1(n_9277),
.A2(n_8180),
.B(n_8140),
.Y(n_9716)
);

INVx1_ASAP7_75t_L g9717 ( 
.A(n_8475),
.Y(n_9717)
);

AND2x2_ASAP7_75t_L g9718 ( 
.A(n_9039),
.B(n_7374),
.Y(n_9718)
);

INVx2_ASAP7_75t_L g9719 ( 
.A(n_8816),
.Y(n_9719)
);

OR2x2_ASAP7_75t_L g9720 ( 
.A(n_9060),
.B(n_7511),
.Y(n_9720)
);

AOI22xp33_ASAP7_75t_SL g9721 ( 
.A1(n_9039),
.A2(n_7638),
.B1(n_7662),
.B2(n_7660),
.Y(n_9721)
);

INVx1_ASAP7_75t_L g9722 ( 
.A(n_8477),
.Y(n_9722)
);

AND2x2_ASAP7_75t_L g9723 ( 
.A(n_9071),
.B(n_9090),
.Y(n_9723)
);

OAI21x1_ASAP7_75t_L g9724 ( 
.A1(n_8407),
.A2(n_7441),
.B(n_7895),
.Y(n_9724)
);

INVx2_ASAP7_75t_L g9725 ( 
.A(n_8816),
.Y(n_9725)
);

INVx1_ASAP7_75t_L g9726 ( 
.A(n_8477),
.Y(n_9726)
);

INVx2_ASAP7_75t_L g9727 ( 
.A(n_9346),
.Y(n_9727)
);

NAND2xp5_ASAP7_75t_L g9728 ( 
.A(n_9071),
.B(n_8173),
.Y(n_9728)
);

BUFx3_ASAP7_75t_L g9729 ( 
.A(n_8409),
.Y(n_9729)
);

INVx1_ASAP7_75t_L g9730 ( 
.A(n_8478),
.Y(n_9730)
);

BUFx2_ASAP7_75t_L g9731 ( 
.A(n_8329),
.Y(n_9731)
);

AO21x2_ASAP7_75t_L g9732 ( 
.A1(n_8764),
.A2(n_7720),
.B(n_7698),
.Y(n_9732)
);

AND2x2_ASAP7_75t_L g9733 ( 
.A(n_9090),
.B(n_7382),
.Y(n_9733)
);

INVx1_ASAP7_75t_L g9734 ( 
.A(n_8478),
.Y(n_9734)
);

BUFx4f_ASAP7_75t_L g9735 ( 
.A(n_8343),
.Y(n_9735)
);

INVx2_ASAP7_75t_L g9736 ( 
.A(n_9346),
.Y(n_9736)
);

INVx1_ASAP7_75t_L g9737 ( 
.A(n_8480),
.Y(n_9737)
);

INVx2_ASAP7_75t_L g9738 ( 
.A(n_9346),
.Y(n_9738)
);

INVx1_ASAP7_75t_L g9739 ( 
.A(n_8480),
.Y(n_9739)
);

INVx1_ASAP7_75t_SL g9740 ( 
.A(n_8375),
.Y(n_9740)
);

INVx1_ASAP7_75t_L g9741 ( 
.A(n_8483),
.Y(n_9741)
);

OAI21x1_ASAP7_75t_L g9742 ( 
.A1(n_8415),
.A2(n_7929),
.B(n_7804),
.Y(n_9742)
);

INVx2_ASAP7_75t_L g9743 ( 
.A(n_9346),
.Y(n_9743)
);

INVx3_ASAP7_75t_L g9744 ( 
.A(n_9346),
.Y(n_9744)
);

INVx1_ASAP7_75t_L g9745 ( 
.A(n_8483),
.Y(n_9745)
);

INVx2_ASAP7_75t_L g9746 ( 
.A(n_8428),
.Y(n_9746)
);

INVx1_ASAP7_75t_L g9747 ( 
.A(n_8487),
.Y(n_9747)
);

INVxp67_ASAP7_75t_L g9748 ( 
.A(n_8569),
.Y(n_9748)
);

AOI21x1_ASAP7_75t_L g9749 ( 
.A1(n_9277),
.A2(n_8228),
.B(n_8180),
.Y(n_9749)
);

INVx2_ASAP7_75t_L g9750 ( 
.A(n_8428),
.Y(n_9750)
);

AOI22xp33_ASAP7_75t_L g9751 ( 
.A1(n_9129),
.A2(n_9172),
.B1(n_8393),
.B2(n_9356),
.Y(n_9751)
);

BUFx3_ASAP7_75t_L g9752 ( 
.A(n_8413),
.Y(n_9752)
);

INVx1_ASAP7_75t_L g9753 ( 
.A(n_8487),
.Y(n_9753)
);

AOI21x1_ASAP7_75t_L g9754 ( 
.A1(n_8520),
.A2(n_8237),
.B(n_8228),
.Y(n_9754)
);

HB1xp67_ASAP7_75t_L g9755 ( 
.A(n_9307),
.Y(n_9755)
);

OAI22xp5_ASAP7_75t_L g9756 ( 
.A1(n_9129),
.A2(n_7834),
.B1(n_7193),
.B2(n_8304),
.Y(n_9756)
);

AOI22xp33_ASAP7_75t_L g9757 ( 
.A1(n_9172),
.A2(n_7458),
.B1(n_7638),
.B2(n_7234),
.Y(n_9757)
);

OAI21xp5_ASAP7_75t_SL g9758 ( 
.A1(n_9356),
.A2(n_7288),
.B(n_7185),
.Y(n_9758)
);

INVx1_ASAP7_75t_L g9759 ( 
.A(n_8490),
.Y(n_9759)
);

INVx1_ASAP7_75t_L g9760 ( 
.A(n_8490),
.Y(n_9760)
);

OR2x6_ASAP7_75t_L g9761 ( 
.A(n_9103),
.B(n_7677),
.Y(n_9761)
);

INVx1_ASAP7_75t_L g9762 ( 
.A(n_8495),
.Y(n_9762)
);

INVx3_ASAP7_75t_L g9763 ( 
.A(n_8347),
.Y(n_9763)
);

INVx2_ASAP7_75t_L g9764 ( 
.A(n_8431),
.Y(n_9764)
);

BUFx2_ASAP7_75t_L g9765 ( 
.A(n_8329),
.Y(n_9765)
);

AND2x2_ASAP7_75t_L g9766 ( 
.A(n_9018),
.B(n_7382),
.Y(n_9766)
);

INVx2_ASAP7_75t_L g9767 ( 
.A(n_8431),
.Y(n_9767)
);

INVx3_ASAP7_75t_L g9768 ( 
.A(n_8347),
.Y(n_9768)
);

OAI21x1_ASAP7_75t_L g9769 ( 
.A1(n_8415),
.A2(n_7929),
.B(n_7804),
.Y(n_9769)
);

BUFx6f_ASAP7_75t_L g9770 ( 
.A(n_8847),
.Y(n_9770)
);

OR2x2_ASAP7_75t_L g9771 ( 
.A(n_9060),
.B(n_7559),
.Y(n_9771)
);

INVx1_ASAP7_75t_L g9772 ( 
.A(n_8495),
.Y(n_9772)
);

AND2x2_ASAP7_75t_L g9773 ( 
.A(n_9018),
.B(n_7382),
.Y(n_9773)
);

INVx2_ASAP7_75t_L g9774 ( 
.A(n_8440),
.Y(n_9774)
);

INVx1_ASAP7_75t_L g9775 ( 
.A(n_8503),
.Y(n_9775)
);

INVx2_ASAP7_75t_L g9776 ( 
.A(n_8440),
.Y(n_9776)
);

OA21x2_ASAP7_75t_L g9777 ( 
.A1(n_8317),
.A2(n_7333),
.B(n_7319),
.Y(n_9777)
);

BUFx4f_ASAP7_75t_SL g9778 ( 
.A(n_8780),
.Y(n_9778)
);

NAND2xp5_ASAP7_75t_L g9779 ( 
.A(n_8899),
.B(n_7993),
.Y(n_9779)
);

NAND2xp5_ASAP7_75t_L g9780 ( 
.A(n_8499),
.B(n_7993),
.Y(n_9780)
);

INVx1_ASAP7_75t_L g9781 ( 
.A(n_8503),
.Y(n_9781)
);

INVx2_ASAP7_75t_L g9782 ( 
.A(n_8456),
.Y(n_9782)
);

INVx2_ASAP7_75t_L g9783 ( 
.A(n_8456),
.Y(n_9783)
);

INVx2_ASAP7_75t_L g9784 ( 
.A(n_8461),
.Y(n_9784)
);

AND2x4_ASAP7_75t_L g9785 ( 
.A(n_8994),
.B(n_7179),
.Y(n_9785)
);

OAI21x1_ASAP7_75t_L g9786 ( 
.A1(n_8415),
.A2(n_7804),
.B(n_7799),
.Y(n_9786)
);

INVx1_ASAP7_75t_L g9787 ( 
.A(n_8504),
.Y(n_9787)
);

OAI21x1_ASAP7_75t_L g9788 ( 
.A1(n_8417),
.A2(n_7799),
.B(n_7649),
.Y(n_9788)
);

INVx2_ASAP7_75t_SL g9789 ( 
.A(n_8311),
.Y(n_9789)
);

INVx2_ASAP7_75t_L g9790 ( 
.A(n_8461),
.Y(n_9790)
);

BUFx2_ASAP7_75t_L g9791 ( 
.A(n_8329),
.Y(n_9791)
);

AND2x2_ASAP7_75t_L g9792 ( 
.A(n_8994),
.B(n_8861),
.Y(n_9792)
);

INVx2_ASAP7_75t_L g9793 ( 
.A(n_8462),
.Y(n_9793)
);

NAND2xp5_ASAP7_75t_L g9794 ( 
.A(n_8521),
.B(n_7883),
.Y(n_9794)
);

OAI22xp5_ASAP7_75t_L g9795 ( 
.A1(n_8538),
.A2(n_7579),
.B1(n_7669),
.B2(n_7860),
.Y(n_9795)
);

AO21x2_ASAP7_75t_L g9796 ( 
.A1(n_8520),
.A2(n_7720),
.B(n_7698),
.Y(n_9796)
);

AND2x2_ASAP7_75t_L g9797 ( 
.A(n_8994),
.B(n_7413),
.Y(n_9797)
);

INVx2_ASAP7_75t_L g9798 ( 
.A(n_8462),
.Y(n_9798)
);

INVx1_ASAP7_75t_L g9799 ( 
.A(n_8504),
.Y(n_9799)
);

OAI21x1_ASAP7_75t_L g9800 ( 
.A1(n_8417),
.A2(n_7799),
.B(n_7649),
.Y(n_9800)
);

INVx1_ASAP7_75t_L g9801 ( 
.A(n_8507),
.Y(n_9801)
);

AND2x2_ASAP7_75t_L g9802 ( 
.A(n_8861),
.B(n_7413),
.Y(n_9802)
);

AO21x2_ASAP7_75t_L g9803 ( 
.A1(n_8611),
.A2(n_7720),
.B(n_7698),
.Y(n_9803)
);

AOI21xp5_ASAP7_75t_L g9804 ( 
.A1(n_8999),
.A2(n_7654),
.B(n_7802),
.Y(n_9804)
);

INVx1_ASAP7_75t_L g9805 ( 
.A(n_8507),
.Y(n_9805)
);

AOI22xp33_ASAP7_75t_SL g9806 ( 
.A1(n_9429),
.A2(n_7638),
.B1(n_7662),
.B2(n_7660),
.Y(n_9806)
);

OR2x2_ASAP7_75t_L g9807 ( 
.A(n_9070),
.B(n_7559),
.Y(n_9807)
);

BUFx2_ASAP7_75t_L g9808 ( 
.A(n_8329),
.Y(n_9808)
);

INVx1_ASAP7_75t_L g9809 ( 
.A(n_8510),
.Y(n_9809)
);

NOR2xp33_ASAP7_75t_L g9810 ( 
.A(n_8725),
.B(n_9013),
.Y(n_9810)
);

INVx2_ASAP7_75t_L g9811 ( 
.A(n_8465),
.Y(n_9811)
);

OAI21x1_ASAP7_75t_L g9812 ( 
.A1(n_8417),
.A2(n_7649),
.B(n_7644),
.Y(n_9812)
);

INVx1_ASAP7_75t_L g9813 ( 
.A(n_8510),
.Y(n_9813)
);

INVx1_ASAP7_75t_SL g9814 ( 
.A(n_8662),
.Y(n_9814)
);

HB1xp67_ASAP7_75t_L g9815 ( 
.A(n_8901),
.Y(n_9815)
);

OAI22xp5_ASAP7_75t_L g9816 ( 
.A1(n_8538),
.A2(n_7579),
.B1(n_7669),
.B2(n_7978),
.Y(n_9816)
);

HB1xp67_ASAP7_75t_L g9817 ( 
.A(n_9106),
.Y(n_9817)
);

INVx2_ASAP7_75t_L g9818 ( 
.A(n_8465),
.Y(n_9818)
);

INVx1_ASAP7_75t_L g9819 ( 
.A(n_8516),
.Y(n_9819)
);

INVx2_ASAP7_75t_SL g9820 ( 
.A(n_8311),
.Y(n_9820)
);

OR2x2_ASAP7_75t_L g9821 ( 
.A(n_9070),
.B(n_7590),
.Y(n_9821)
);

HB1xp67_ASAP7_75t_L g9822 ( 
.A(n_9149),
.Y(n_9822)
);

INVx2_ASAP7_75t_L g9823 ( 
.A(n_8468),
.Y(n_9823)
);

INVx1_ASAP7_75t_L g9824 ( 
.A(n_8516),
.Y(n_9824)
);

BUFx6f_ASAP7_75t_L g9825 ( 
.A(n_9013),
.Y(n_9825)
);

INVx1_ASAP7_75t_L g9826 ( 
.A(n_8517),
.Y(n_9826)
);

INVx3_ASAP7_75t_L g9827 ( 
.A(n_8347),
.Y(n_9827)
);

INVx1_ASAP7_75t_L g9828 ( 
.A(n_8517),
.Y(n_9828)
);

INVx2_ASAP7_75t_L g9829 ( 
.A(n_8468),
.Y(n_9829)
);

INVx2_ASAP7_75t_L g9830 ( 
.A(n_8482),
.Y(n_9830)
);

INVx1_ASAP7_75t_L g9831 ( 
.A(n_8522),
.Y(n_9831)
);

OR2x2_ASAP7_75t_L g9832 ( 
.A(n_9329),
.B(n_7590),
.Y(n_9832)
);

AND2x2_ASAP7_75t_L g9833 ( 
.A(n_9114),
.B(n_7413),
.Y(n_9833)
);

INVx2_ASAP7_75t_L g9834 ( 
.A(n_8482),
.Y(n_9834)
);

INVx2_ASAP7_75t_SL g9835 ( 
.A(n_8402),
.Y(n_9835)
);

INVx2_ASAP7_75t_L g9836 ( 
.A(n_8491),
.Y(n_9836)
);

A2O1A1Ixp33_ASAP7_75t_L g9837 ( 
.A1(n_8656),
.A2(n_7752),
.B(n_7735),
.C(n_7769),
.Y(n_9837)
);

AND2x2_ASAP7_75t_SL g9838 ( 
.A(n_9429),
.B(n_7682),
.Y(n_9838)
);

HB1xp67_ASAP7_75t_L g9839 ( 
.A(n_9229),
.Y(n_9839)
);

INVxp33_ASAP7_75t_L g9840 ( 
.A(n_9200),
.Y(n_9840)
);

AND2x2_ASAP7_75t_L g9841 ( 
.A(n_9114),
.B(n_7964),
.Y(n_9841)
);

INVx1_ASAP7_75t_L g9842 ( 
.A(n_8522),
.Y(n_9842)
);

INVx2_ASAP7_75t_L g9843 ( 
.A(n_8491),
.Y(n_9843)
);

INVx2_ASAP7_75t_L g9844 ( 
.A(n_8493),
.Y(n_9844)
);

NAND2xp5_ASAP7_75t_L g9845 ( 
.A(n_9025),
.B(n_8537),
.Y(n_9845)
);

NOR2xp33_ASAP7_75t_L g9846 ( 
.A(n_9013),
.B(n_9024),
.Y(n_9846)
);

INVx2_ASAP7_75t_L g9847 ( 
.A(n_8493),
.Y(n_9847)
);

INVx1_ASAP7_75t_L g9848 ( 
.A(n_8524),
.Y(n_9848)
);

AO21x2_ASAP7_75t_L g9849 ( 
.A1(n_8611),
.A2(n_7720),
.B(n_7698),
.Y(n_9849)
);

OR2x6_ASAP7_75t_L g9850 ( 
.A(n_9103),
.B(n_7677),
.Y(n_9850)
);

NAND2xp5_ASAP7_75t_L g9851 ( 
.A(n_8593),
.B(n_7883),
.Y(n_9851)
);

INVx2_ASAP7_75t_SL g9852 ( 
.A(n_8402),
.Y(n_9852)
);

BUFx2_ASAP7_75t_L g9853 ( 
.A(n_8941),
.Y(n_9853)
);

AOI21x1_ASAP7_75t_L g9854 ( 
.A1(n_8972),
.A2(n_8270),
.B(n_8237),
.Y(n_9854)
);

INVx1_ASAP7_75t_L g9855 ( 
.A(n_8524),
.Y(n_9855)
);

INVx1_ASAP7_75t_L g9856 ( 
.A(n_8525),
.Y(n_9856)
);

INVx2_ASAP7_75t_L g9857 ( 
.A(n_8500),
.Y(n_9857)
);

INVx2_ASAP7_75t_L g9858 ( 
.A(n_8500),
.Y(n_9858)
);

HB1xp67_ASAP7_75t_L g9859 ( 
.A(n_9237),
.Y(n_9859)
);

BUFx12f_ASAP7_75t_L g9860 ( 
.A(n_8886),
.Y(n_9860)
);

INVx2_ASAP7_75t_L g9861 ( 
.A(n_8472),
.Y(n_9861)
);

INVx1_ASAP7_75t_L g9862 ( 
.A(n_8525),
.Y(n_9862)
);

INVx1_ASAP7_75t_SL g9863 ( 
.A(n_8815),
.Y(n_9863)
);

INVx1_ASAP7_75t_L g9864 ( 
.A(n_8534),
.Y(n_9864)
);

INVx2_ASAP7_75t_L g9865 ( 
.A(n_8472),
.Y(n_9865)
);

INVx1_ASAP7_75t_L g9866 ( 
.A(n_8534),
.Y(n_9866)
);

INVx1_ASAP7_75t_L g9867 ( 
.A(n_8544),
.Y(n_9867)
);

AND2x2_ASAP7_75t_L g9868 ( 
.A(n_9087),
.B(n_7964),
.Y(n_9868)
);

INVx1_ASAP7_75t_L g9869 ( 
.A(n_8544),
.Y(n_9869)
);

INVx1_ASAP7_75t_L g9870 ( 
.A(n_8548),
.Y(n_9870)
);

INVx2_ASAP7_75t_L g9871 ( 
.A(n_8472),
.Y(n_9871)
);

INVx1_ASAP7_75t_L g9872 ( 
.A(n_8548),
.Y(n_9872)
);

HB1xp67_ASAP7_75t_L g9873 ( 
.A(n_9112),
.Y(n_9873)
);

OAI22xp5_ASAP7_75t_SL g9874 ( 
.A1(n_8638),
.A2(n_6614),
.B1(n_6629),
.B2(n_6579),
.Y(n_9874)
);

NAND2xp5_ASAP7_75t_L g9875 ( 
.A(n_8404),
.B(n_7944),
.Y(n_9875)
);

INVx1_ASAP7_75t_L g9876 ( 
.A(n_8554),
.Y(n_9876)
);

AND2x4_ASAP7_75t_L g9877 ( 
.A(n_9087),
.B(n_8130),
.Y(n_9877)
);

INVx8_ASAP7_75t_L g9878 ( 
.A(n_8545),
.Y(n_9878)
);

AND2x2_ASAP7_75t_L g9879 ( 
.A(n_9087),
.B(n_7964),
.Y(n_9879)
);

CKINVDCx5p33_ASAP7_75t_R g9880 ( 
.A(n_8319),
.Y(n_9880)
);

INVx1_ASAP7_75t_L g9881 ( 
.A(n_8554),
.Y(n_9881)
);

INVx2_ASAP7_75t_L g9882 ( 
.A(n_8457),
.Y(n_9882)
);

INVx1_ASAP7_75t_L g9883 ( 
.A(n_8557),
.Y(n_9883)
);

INVx2_ASAP7_75t_L g9884 ( 
.A(n_8457),
.Y(n_9884)
);

HB1xp67_ASAP7_75t_L g9885 ( 
.A(n_8318),
.Y(n_9885)
);

INVx2_ASAP7_75t_L g9886 ( 
.A(n_8457),
.Y(n_9886)
);

INVx1_ASAP7_75t_L g9887 ( 
.A(n_8557),
.Y(n_9887)
);

INVx1_ASAP7_75t_L g9888 ( 
.A(n_8562),
.Y(n_9888)
);

BUFx2_ASAP7_75t_L g9889 ( 
.A(n_8941),
.Y(n_9889)
);

INVx2_ASAP7_75t_L g9890 ( 
.A(n_8457),
.Y(n_9890)
);

OAI21x1_ASAP7_75t_L g9891 ( 
.A1(n_8459),
.A2(n_7644),
.B(n_7866),
.Y(n_9891)
);

OAI21x1_ASAP7_75t_L g9892 ( 
.A1(n_8459),
.A2(n_8486),
.B(n_8532),
.Y(n_9892)
);

INVx1_ASAP7_75t_L g9893 ( 
.A(n_8562),
.Y(n_9893)
);

HB1xp67_ASAP7_75t_L g9894 ( 
.A(n_8331),
.Y(n_9894)
);

INVx1_ASAP7_75t_L g9895 ( 
.A(n_8563),
.Y(n_9895)
);

BUFx3_ASAP7_75t_L g9896 ( 
.A(n_9024),
.Y(n_9896)
);

INVx1_ASAP7_75t_L g9897 ( 
.A(n_8563),
.Y(n_9897)
);

INVx2_ASAP7_75t_L g9898 ( 
.A(n_8459),
.Y(n_9898)
);

AND2x2_ASAP7_75t_L g9899 ( 
.A(n_9087),
.B(n_8055),
.Y(n_9899)
);

INVx1_ASAP7_75t_L g9900 ( 
.A(n_8573),
.Y(n_9900)
);

BUFx3_ASAP7_75t_L g9901 ( 
.A(n_9024),
.Y(n_9901)
);

BUFx3_ASAP7_75t_L g9902 ( 
.A(n_8820),
.Y(n_9902)
);

INVx3_ASAP7_75t_SL g9903 ( 
.A(n_8863),
.Y(n_9903)
);

AND2x2_ASAP7_75t_L g9904 ( 
.A(n_9159),
.B(n_8055),
.Y(n_9904)
);

INVx1_ASAP7_75t_L g9905 ( 
.A(n_8573),
.Y(n_9905)
);

INVx1_ASAP7_75t_L g9906 ( 
.A(n_8583),
.Y(n_9906)
);

NOR2xp33_ASAP7_75t_L g9907 ( 
.A(n_9278),
.B(n_7995),
.Y(n_9907)
);

INVx1_ASAP7_75t_L g9908 ( 
.A(n_8583),
.Y(n_9908)
);

INVx2_ASAP7_75t_SL g9909 ( 
.A(n_8402),
.Y(n_9909)
);

AND2x2_ASAP7_75t_L g9910 ( 
.A(n_9159),
.B(n_8055),
.Y(n_9910)
);

INVx1_ASAP7_75t_L g9911 ( 
.A(n_8594),
.Y(n_9911)
);

INVx1_ASAP7_75t_L g9912 ( 
.A(n_8594),
.Y(n_9912)
);

INVx1_ASAP7_75t_L g9913 ( 
.A(n_8596),
.Y(n_9913)
);

INVx2_ASAP7_75t_L g9914 ( 
.A(n_8459),
.Y(n_9914)
);

AND2x4_ASAP7_75t_L g9915 ( 
.A(n_9159),
.B(n_8155),
.Y(n_9915)
);

INVx2_ASAP7_75t_L g9916 ( 
.A(n_8486),
.Y(n_9916)
);

INVx1_ASAP7_75t_L g9917 ( 
.A(n_8596),
.Y(n_9917)
);

INVx2_ASAP7_75t_SL g9918 ( 
.A(n_8402),
.Y(n_9918)
);

INVx1_ASAP7_75t_SL g9919 ( 
.A(n_8822),
.Y(n_9919)
);

INVx1_ASAP7_75t_L g9920 ( 
.A(n_8598),
.Y(n_9920)
);

HB1xp67_ASAP7_75t_L g9921 ( 
.A(n_8362),
.Y(n_9921)
);

INVx2_ASAP7_75t_L g9922 ( 
.A(n_8486),
.Y(n_9922)
);

AOI21xp5_ASAP7_75t_L g9923 ( 
.A1(n_8455),
.A2(n_8050),
.B(n_7341),
.Y(n_9923)
);

INVx1_ASAP7_75t_L g9924 ( 
.A(n_8598),
.Y(n_9924)
);

NAND2xp5_ASAP7_75t_L g9925 ( 
.A(n_8404),
.B(n_7944),
.Y(n_9925)
);

BUFx3_ASAP7_75t_L g9926 ( 
.A(n_8830),
.Y(n_9926)
);

AND2x2_ASAP7_75t_L g9927 ( 
.A(n_9159),
.B(n_9164),
.Y(n_9927)
);

HB1xp67_ASAP7_75t_L g9928 ( 
.A(n_8369),
.Y(n_9928)
);

INVx1_ASAP7_75t_L g9929 ( 
.A(n_8603),
.Y(n_9929)
);

INVx2_ASAP7_75t_L g9930 ( 
.A(n_8486),
.Y(n_9930)
);

INVx1_ASAP7_75t_L g9931 ( 
.A(n_8603),
.Y(n_9931)
);

OAI21x1_ASAP7_75t_L g9932 ( 
.A1(n_8532),
.A2(n_7644),
.B(n_7866),
.Y(n_9932)
);

INVx1_ASAP7_75t_L g9933 ( 
.A(n_8604),
.Y(n_9933)
);

OR2x2_ASAP7_75t_L g9934 ( 
.A(n_9329),
.B(n_7628),
.Y(n_9934)
);

INVx1_ASAP7_75t_L g9935 ( 
.A(n_8604),
.Y(n_9935)
);

AND2x4_ASAP7_75t_L g9936 ( 
.A(n_9164),
.B(n_8155),
.Y(n_9936)
);

INVx2_ASAP7_75t_SL g9937 ( 
.A(n_8412),
.Y(n_9937)
);

OR2x2_ASAP7_75t_L g9938 ( 
.A(n_8940),
.B(n_7628),
.Y(n_9938)
);

INVx1_ASAP7_75t_L g9939 ( 
.A(n_8612),
.Y(n_9939)
);

AND2x2_ASAP7_75t_L g9940 ( 
.A(n_9164),
.B(n_8178),
.Y(n_9940)
);

INVx3_ASAP7_75t_L g9941 ( 
.A(n_8347),
.Y(n_9941)
);

OAI21x1_ASAP7_75t_L g9942 ( 
.A1(n_8532),
.A2(n_7866),
.B(n_8044),
.Y(n_9942)
);

INVx2_ASAP7_75t_SL g9943 ( 
.A(n_8412),
.Y(n_9943)
);

INVx2_ASAP7_75t_L g9944 ( 
.A(n_8948),
.Y(n_9944)
);

INVx2_ASAP7_75t_L g9945 ( 
.A(n_8948),
.Y(n_9945)
);

BUFx6f_ASAP7_75t_L g9946 ( 
.A(n_8889),
.Y(n_9946)
);

INVx1_ASAP7_75t_L g9947 ( 
.A(n_8612),
.Y(n_9947)
);

AO21x1_ASAP7_75t_L g9948 ( 
.A1(n_9191),
.A2(n_7878),
.B(n_8050),
.Y(n_9948)
);

AO21x2_ASAP7_75t_L g9949 ( 
.A1(n_9078),
.A2(n_7751),
.B(n_7724),
.Y(n_9949)
);

BUFx2_ASAP7_75t_L g9950 ( 
.A(n_8941),
.Y(n_9950)
);

INVx2_ASAP7_75t_L g9951 ( 
.A(n_8948),
.Y(n_9951)
);

INVx1_ASAP7_75t_L g9952 ( 
.A(n_8621),
.Y(n_9952)
);

INVx3_ASAP7_75t_L g9953 ( 
.A(n_8390),
.Y(n_9953)
);

BUFx2_ASAP7_75t_L g9954 ( 
.A(n_8941),
.Y(n_9954)
);

BUFx3_ASAP7_75t_L g9955 ( 
.A(n_8833),
.Y(n_9955)
);

INVx1_ASAP7_75t_L g9956 ( 
.A(n_8621),
.Y(n_9956)
);

INVx2_ASAP7_75t_L g9957 ( 
.A(n_8948),
.Y(n_9957)
);

INVx2_ASAP7_75t_L g9958 ( 
.A(n_8959),
.Y(n_9958)
);

INVx2_ASAP7_75t_L g9959 ( 
.A(n_8959),
.Y(n_9959)
);

INVx2_ASAP7_75t_L g9960 ( 
.A(n_8959),
.Y(n_9960)
);

INVx1_ASAP7_75t_L g9961 ( 
.A(n_8627),
.Y(n_9961)
);

INVx2_ASAP7_75t_L g9962 ( 
.A(n_8959),
.Y(n_9962)
);

INVx1_ASAP7_75t_L g9963 ( 
.A(n_8627),
.Y(n_9963)
);

INVx2_ASAP7_75t_L g9964 ( 
.A(n_9054),
.Y(n_9964)
);

INVx2_ASAP7_75t_L g9965 ( 
.A(n_9054),
.Y(n_9965)
);

AO21x1_ASAP7_75t_SL g9966 ( 
.A1(n_9119),
.A2(n_8137),
.B(n_8098),
.Y(n_9966)
);

INVx1_ASAP7_75t_L g9967 ( 
.A(n_8630),
.Y(n_9967)
);

INVx2_ASAP7_75t_L g9968 ( 
.A(n_9054),
.Y(n_9968)
);

INVxp67_ASAP7_75t_L g9969 ( 
.A(n_8569),
.Y(n_9969)
);

INVx3_ASAP7_75t_L g9970 ( 
.A(n_8390),
.Y(n_9970)
);

OAI21x1_ASAP7_75t_L g9971 ( 
.A1(n_8532),
.A2(n_7602),
.B(n_7585),
.Y(n_9971)
);

INVx2_ASAP7_75t_SL g9972 ( 
.A(n_8412),
.Y(n_9972)
);

INVx2_ASAP7_75t_L g9973 ( 
.A(n_9054),
.Y(n_9973)
);

INVx1_ASAP7_75t_L g9974 ( 
.A(n_8630),
.Y(n_9974)
);

OAI21x1_ASAP7_75t_L g9975 ( 
.A1(n_8570),
.A2(n_7602),
.B(n_7585),
.Y(n_9975)
);

OAI21x1_ASAP7_75t_L g9976 ( 
.A1(n_8570),
.A2(n_7602),
.B(n_7585),
.Y(n_9976)
);

INVx1_ASAP7_75t_L g9977 ( 
.A(n_8645),
.Y(n_9977)
);

INVxp67_ASAP7_75t_L g9978 ( 
.A(n_8696),
.Y(n_9978)
);

BUFx2_ASAP7_75t_L g9979 ( 
.A(n_9140),
.Y(n_9979)
);

INVx1_ASAP7_75t_L g9980 ( 
.A(n_8645),
.Y(n_9980)
);

INVx2_ASAP7_75t_L g9981 ( 
.A(n_9194),
.Y(n_9981)
);

OR2x6_ASAP7_75t_L g9982 ( 
.A(n_9103),
.B(n_7677),
.Y(n_9982)
);

INVx1_ASAP7_75t_L g9983 ( 
.A(n_8648),
.Y(n_9983)
);

OR2x2_ASAP7_75t_L g9984 ( 
.A(n_8940),
.B(n_7679),
.Y(n_9984)
);

INVx1_ASAP7_75t_L g9985 ( 
.A(n_8648),
.Y(n_9985)
);

INVx2_ASAP7_75t_L g9986 ( 
.A(n_9194),
.Y(n_9986)
);

INVx3_ASAP7_75t_L g9987 ( 
.A(n_8390),
.Y(n_9987)
);

INVx1_ASAP7_75t_L g9988 ( 
.A(n_8664),
.Y(n_9988)
);

OR2x2_ASAP7_75t_L g9989 ( 
.A(n_9000),
.B(n_7679),
.Y(n_9989)
);

AND2x2_ASAP7_75t_L g9990 ( 
.A(n_9164),
.B(n_8178),
.Y(n_9990)
);

AND2x2_ASAP7_75t_L g9991 ( 
.A(n_9292),
.B(n_8178),
.Y(n_9991)
);

AND2x4_ASAP7_75t_L g9992 ( 
.A(n_9292),
.B(n_9297),
.Y(n_9992)
);

BUFx2_ASAP7_75t_L g9993 ( 
.A(n_8341),
.Y(n_9993)
);

INVx1_ASAP7_75t_L g9994 ( 
.A(n_8664),
.Y(n_9994)
);

BUFx2_ASAP7_75t_L g9995 ( 
.A(n_8341),
.Y(n_9995)
);

INVx1_ASAP7_75t_L g9996 ( 
.A(n_8669),
.Y(n_9996)
);

INVx2_ASAP7_75t_L g9997 ( 
.A(n_9194),
.Y(n_9997)
);

INVx1_ASAP7_75t_L g9998 ( 
.A(n_8669),
.Y(n_9998)
);

INVx1_ASAP7_75t_L g9999 ( 
.A(n_8678),
.Y(n_9999)
);

INVx1_ASAP7_75t_SL g10000 ( 
.A(n_8880),
.Y(n_10000)
);

INVx1_ASAP7_75t_L g10001 ( 
.A(n_8678),
.Y(n_10001)
);

AND2x2_ASAP7_75t_L g10002 ( 
.A(n_9292),
.B(n_8191),
.Y(n_10002)
);

INVx1_ASAP7_75t_L g10003 ( 
.A(n_8686),
.Y(n_10003)
);

INVx3_ASAP7_75t_L g10004 ( 
.A(n_8390),
.Y(n_10004)
);

INVx1_ASAP7_75t_L g10005 ( 
.A(n_8686),
.Y(n_10005)
);

INVx1_ASAP7_75t_L g10006 ( 
.A(n_8689),
.Y(n_10006)
);

OAI21x1_ASAP7_75t_L g10007 ( 
.A1(n_8570),
.A2(n_7872),
.B(n_7494),
.Y(n_10007)
);

INVx2_ASAP7_75t_L g10008 ( 
.A(n_9194),
.Y(n_10008)
);

AND2x2_ASAP7_75t_L g10009 ( 
.A(n_9292),
.B(n_8191),
.Y(n_10009)
);

BUFx2_ASAP7_75t_L g10010 ( 
.A(n_8341),
.Y(n_10010)
);

INVx1_ASAP7_75t_L g10011 ( 
.A(n_8689),
.Y(n_10011)
);

CKINVDCx5p33_ASAP7_75t_R g10012 ( 
.A(n_8479),
.Y(n_10012)
);

INVx2_ASAP7_75t_L g10013 ( 
.A(n_9232),
.Y(n_10013)
);

INVx1_ASAP7_75t_L g10014 ( 
.A(n_8690),
.Y(n_10014)
);

INVx2_ASAP7_75t_L g10015 ( 
.A(n_9232),
.Y(n_10015)
);

NAND2xp5_ASAP7_75t_L g10016 ( 
.A(n_8609),
.B(n_7786),
.Y(n_10016)
);

INVx1_ASAP7_75t_L g10017 ( 
.A(n_8690),
.Y(n_10017)
);

BUFx3_ASAP7_75t_L g10018 ( 
.A(n_8900),
.Y(n_10018)
);

INVx6_ASAP7_75t_L g10019 ( 
.A(n_8412),
.Y(n_10019)
);

INVx1_ASAP7_75t_L g10020 ( 
.A(n_8692),
.Y(n_10020)
);

INVx1_ASAP7_75t_L g10021 ( 
.A(n_8692),
.Y(n_10021)
);

AND2x2_ASAP7_75t_L g10022 ( 
.A(n_9297),
.B(n_9365),
.Y(n_10022)
);

INVx2_ASAP7_75t_SL g10023 ( 
.A(n_8694),
.Y(n_10023)
);

INVx2_ASAP7_75t_L g10024 ( 
.A(n_9232),
.Y(n_10024)
);

INVx2_ASAP7_75t_L g10025 ( 
.A(n_9232),
.Y(n_10025)
);

BUFx2_ASAP7_75t_L g10026 ( 
.A(n_8346),
.Y(n_10026)
);

AOI21x1_ASAP7_75t_L g10027 ( 
.A1(n_9063),
.A2(n_8270),
.B(n_7494),
.Y(n_10027)
);

INVx1_ASAP7_75t_L g10028 ( 
.A(n_8697),
.Y(n_10028)
);

OAI22xp5_ASAP7_75t_L g10029 ( 
.A1(n_9210),
.A2(n_7978),
.B1(n_7430),
.B2(n_7486),
.Y(n_10029)
);

INVx2_ASAP7_75t_L g10030 ( 
.A(n_9269),
.Y(n_10030)
);

BUFx2_ASAP7_75t_L g10031 ( 
.A(n_8346),
.Y(n_10031)
);

HB1xp67_ASAP7_75t_L g10032 ( 
.A(n_8376),
.Y(n_10032)
);

INVx2_ASAP7_75t_L g10033 ( 
.A(n_9269),
.Y(n_10033)
);

AOI21x1_ASAP7_75t_L g10034 ( 
.A1(n_8814),
.A2(n_7414),
.B(n_7747),
.Y(n_10034)
);

INVx2_ASAP7_75t_L g10035 ( 
.A(n_9269),
.Y(n_10035)
);

INVx1_ASAP7_75t_L g10036 ( 
.A(n_8697),
.Y(n_10036)
);

AND2x2_ASAP7_75t_L g10037 ( 
.A(n_9297),
.B(n_8191),
.Y(n_10037)
);

OA21x2_ASAP7_75t_L g10038 ( 
.A1(n_9074),
.A2(n_7333),
.B(n_7457),
.Y(n_10038)
);

INVx4_ASAP7_75t_L g10039 ( 
.A(n_8383),
.Y(n_10039)
);

INVx3_ASAP7_75t_L g10040 ( 
.A(n_9238),
.Y(n_10040)
);

INVx2_ASAP7_75t_L g10041 ( 
.A(n_9269),
.Y(n_10041)
);

AND2x2_ASAP7_75t_L g10042 ( 
.A(n_9297),
.B(n_7408),
.Y(n_10042)
);

NAND2xp5_ASAP7_75t_L g10043 ( 
.A(n_8655),
.B(n_7786),
.Y(n_10043)
);

INVx1_ASAP7_75t_L g10044 ( 
.A(n_8701),
.Y(n_10044)
);

AOI21x1_ASAP7_75t_L g10045 ( 
.A1(n_8814),
.A2(n_7747),
.B(n_7999),
.Y(n_10045)
);

INVxp67_ASAP7_75t_L g10046 ( 
.A(n_8696),
.Y(n_10046)
);

INVx1_ASAP7_75t_L g10047 ( 
.A(n_8701),
.Y(n_10047)
);

INVx2_ASAP7_75t_L g10048 ( 
.A(n_9291),
.Y(n_10048)
);

INVx2_ASAP7_75t_L g10049 ( 
.A(n_9291),
.Y(n_10049)
);

INVx1_ASAP7_75t_L g10050 ( 
.A(n_8709),
.Y(n_10050)
);

INVx2_ASAP7_75t_SL g10051 ( 
.A(n_8694),
.Y(n_10051)
);

BUFx3_ASAP7_75t_L g10052 ( 
.A(n_8694),
.Y(n_10052)
);

AO21x2_ASAP7_75t_L g10053 ( 
.A1(n_9078),
.A2(n_7751),
.B(n_7724),
.Y(n_10053)
);

BUFx2_ASAP7_75t_L g10054 ( 
.A(n_8346),
.Y(n_10054)
);

INVx1_ASAP7_75t_L g10055 ( 
.A(n_8709),
.Y(n_10055)
);

OAI21x1_ASAP7_75t_L g10056 ( 
.A1(n_8570),
.A2(n_7872),
.B(n_7885),
.Y(n_10056)
);

AOI22xp33_ASAP7_75t_SL g10057 ( 
.A1(n_9430),
.A2(n_7638),
.B1(n_7662),
.B2(n_7660),
.Y(n_10057)
);

INVx1_ASAP7_75t_L g10058 ( 
.A(n_8720),
.Y(n_10058)
);

OA21x2_ASAP7_75t_L g10059 ( 
.A1(n_9074),
.A2(n_7457),
.B(n_7232),
.Y(n_10059)
);

CKINVDCx20_ASAP7_75t_R g10060 ( 
.A(n_8438),
.Y(n_10060)
);

HB1xp67_ASAP7_75t_L g10061 ( 
.A(n_8496),
.Y(n_10061)
);

OR2x6_ASAP7_75t_L g10062 ( 
.A(n_9299),
.B(n_7713),
.Y(n_10062)
);

CKINVDCx20_ASAP7_75t_R g10063 ( 
.A(n_8734),
.Y(n_10063)
);

INVx2_ASAP7_75t_L g10064 ( 
.A(n_9291),
.Y(n_10064)
);

INVx2_ASAP7_75t_L g10065 ( 
.A(n_9291),
.Y(n_10065)
);

INVx1_ASAP7_75t_L g10066 ( 
.A(n_8720),
.Y(n_10066)
);

OA21x2_ASAP7_75t_L g10067 ( 
.A1(n_9082),
.A2(n_7457),
.B(n_7232),
.Y(n_10067)
);

NAND2xp5_ASAP7_75t_L g10068 ( 
.A(n_9210),
.B(n_7986),
.Y(n_10068)
);

INVx2_ASAP7_75t_L g10069 ( 
.A(n_9314),
.Y(n_10069)
);

HB1xp67_ASAP7_75t_L g10070 ( 
.A(n_8531),
.Y(n_10070)
);

OAI21xp5_ASAP7_75t_L g10071 ( 
.A1(n_9227),
.A2(n_7931),
.B(n_7878),
.Y(n_10071)
);

BUFx6f_ASAP7_75t_L g10072 ( 
.A(n_8327),
.Y(n_10072)
);

HB1xp67_ASAP7_75t_L g10073 ( 
.A(n_8542),
.Y(n_10073)
);

AND2x2_ASAP7_75t_L g10074 ( 
.A(n_9365),
.B(n_9399),
.Y(n_10074)
);

INVx2_ASAP7_75t_L g10075 ( 
.A(n_9314),
.Y(n_10075)
);

INVx2_ASAP7_75t_L g10076 ( 
.A(n_9314),
.Y(n_10076)
);

INVx1_ASAP7_75t_L g10077 ( 
.A(n_8730),
.Y(n_10077)
);

HB1xp67_ASAP7_75t_L g10078 ( 
.A(n_8551),
.Y(n_10078)
);

INVx1_ASAP7_75t_L g10079 ( 
.A(n_8730),
.Y(n_10079)
);

BUFx4f_ASAP7_75t_SL g10080 ( 
.A(n_8343),
.Y(n_10080)
);

INVx2_ASAP7_75t_L g10081 ( 
.A(n_9314),
.Y(n_10081)
);

INVx2_ASAP7_75t_L g10082 ( 
.A(n_8617),
.Y(n_10082)
);

HB1xp67_ASAP7_75t_L g10083 ( 
.A(n_8566),
.Y(n_10083)
);

INVx3_ASAP7_75t_L g10084 ( 
.A(n_9238),
.Y(n_10084)
);

INVx2_ASAP7_75t_L g10085 ( 
.A(n_8617),
.Y(n_10085)
);

INVx1_ASAP7_75t_L g10086 ( 
.A(n_8743),
.Y(n_10086)
);

AOI22xp5_ASAP7_75t_L g10087 ( 
.A1(n_9430),
.A2(n_7715),
.B1(n_7893),
.B2(n_7234),
.Y(n_10087)
);

INVx1_ASAP7_75t_L g10088 ( 
.A(n_8743),
.Y(n_10088)
);

INVx1_ASAP7_75t_L g10089 ( 
.A(n_8748),
.Y(n_10089)
);

CKINVDCx11_ASAP7_75t_R g10090 ( 
.A(n_8694),
.Y(n_10090)
);

AO21x2_ASAP7_75t_L g10091 ( 
.A1(n_9109),
.A2(n_7751),
.B(n_7724),
.Y(n_10091)
);

OA21x2_ASAP7_75t_L g10092 ( 
.A1(n_9082),
.A2(n_9093),
.B(n_9085),
.Y(n_10092)
);

INVx1_ASAP7_75t_L g10093 ( 
.A(n_8748),
.Y(n_10093)
);

INVx1_ASAP7_75t_L g10094 ( 
.A(n_8753),
.Y(n_10094)
);

INVx1_ASAP7_75t_L g10095 ( 
.A(n_8753),
.Y(n_10095)
);

HB1xp67_ASAP7_75t_L g10096 ( 
.A(n_8608),
.Y(n_10096)
);

INVx1_ASAP7_75t_L g10097 ( 
.A(n_8756),
.Y(n_10097)
);

HB1xp67_ASAP7_75t_L g10098 ( 
.A(n_8642),
.Y(n_10098)
);

INVx2_ASAP7_75t_L g10099 ( 
.A(n_8617),
.Y(n_10099)
);

OAI21x1_ASAP7_75t_L g10100 ( 
.A1(n_8606),
.A2(n_7872),
.B(n_7885),
.Y(n_10100)
);

INVx1_ASAP7_75t_L g10101 ( 
.A(n_8756),
.Y(n_10101)
);

NAND2x1p5_ASAP7_75t_L g10102 ( 
.A(n_8788),
.B(n_7979),
.Y(n_10102)
);

BUFx3_ASAP7_75t_L g10103 ( 
.A(n_8909),
.Y(n_10103)
);

INVx1_ASAP7_75t_L g10104 ( 
.A(n_8757),
.Y(n_10104)
);

INVx1_ASAP7_75t_L g10105 ( 
.A(n_8757),
.Y(n_10105)
);

INVx1_ASAP7_75t_L g10106 ( 
.A(n_8762),
.Y(n_10106)
);

AND2x2_ASAP7_75t_L g10107 ( 
.A(n_9365),
.B(n_7408),
.Y(n_10107)
);

INVx2_ASAP7_75t_L g10108 ( 
.A(n_9203),
.Y(n_10108)
);

AOI22xp33_ASAP7_75t_L g10109 ( 
.A1(n_8704),
.A2(n_7458),
.B1(n_7638),
.B2(n_7234),
.Y(n_10109)
);

INVx1_ASAP7_75t_L g10110 ( 
.A(n_8762),
.Y(n_10110)
);

OAI21x1_ASAP7_75t_L g10111 ( 
.A1(n_8606),
.A2(n_7903),
.B(n_7885),
.Y(n_10111)
);

INVx1_ASAP7_75t_L g10112 ( 
.A(n_8766),
.Y(n_10112)
);

INVx3_ASAP7_75t_L g10113 ( 
.A(n_8606),
.Y(n_10113)
);

OAI21xp5_ASAP7_75t_L g10114 ( 
.A1(n_8547),
.A2(n_7931),
.B(n_7288),
.Y(n_10114)
);

INVx1_ASAP7_75t_L g10115 ( 
.A(n_8766),
.Y(n_10115)
);

INVx2_ASAP7_75t_L g10116 ( 
.A(n_9203),
.Y(n_10116)
);

INVx2_ASAP7_75t_L g10117 ( 
.A(n_9305),
.Y(n_10117)
);

INVxp67_ASAP7_75t_L g10118 ( 
.A(n_8656),
.Y(n_10118)
);

INVx1_ASAP7_75t_L g10119 ( 
.A(n_8769),
.Y(n_10119)
);

NAND2xp5_ASAP7_75t_L g10120 ( 
.A(n_8433),
.B(n_7886),
.Y(n_10120)
);

INVx3_ASAP7_75t_L g10121 ( 
.A(n_8606),
.Y(n_10121)
);

INVx3_ASAP7_75t_L g10122 ( 
.A(n_8628),
.Y(n_10122)
);

AND2x2_ASAP7_75t_L g10123 ( 
.A(n_9365),
.B(n_7408),
.Y(n_10123)
);

INVx2_ASAP7_75t_L g10124 ( 
.A(n_9305),
.Y(n_10124)
);

INVx1_ASAP7_75t_L g10125 ( 
.A(n_8769),
.Y(n_10125)
);

BUFx6f_ASAP7_75t_L g10126 ( 
.A(n_8327),
.Y(n_10126)
);

INVx2_ASAP7_75t_SL g10127 ( 
.A(n_9406),
.Y(n_10127)
);

BUFx10_ASAP7_75t_L g10128 ( 
.A(n_8859),
.Y(n_10128)
);

HB1xp67_ASAP7_75t_L g10129 ( 
.A(n_8657),
.Y(n_10129)
);

INVx1_ASAP7_75t_L g10130 ( 
.A(n_8779),
.Y(n_10130)
);

BUFx3_ASAP7_75t_L g10131 ( 
.A(n_8998),
.Y(n_10131)
);

AOI22xp33_ASAP7_75t_L g10132 ( 
.A1(n_8704),
.A2(n_7458),
.B1(n_7638),
.B2(n_7234),
.Y(n_10132)
);

AND2x2_ASAP7_75t_L g10133 ( 
.A(n_9399),
.B(n_8306),
.Y(n_10133)
);

AND2x2_ASAP7_75t_L g10134 ( 
.A(n_9399),
.B(n_7452),
.Y(n_10134)
);

INVx2_ASAP7_75t_SL g10135 ( 
.A(n_9174),
.Y(n_10135)
);

INVx2_ASAP7_75t_L g10136 ( 
.A(n_9312),
.Y(n_10136)
);

OAI22xp5_ASAP7_75t_SL g10137 ( 
.A1(n_8638),
.A2(n_6629),
.B1(n_6637),
.B2(n_6614),
.Y(n_10137)
);

INVx1_ASAP7_75t_L g10138 ( 
.A(n_8779),
.Y(n_10138)
);

OAI21x1_ASAP7_75t_L g10139 ( 
.A1(n_8628),
.A2(n_7907),
.B(n_7903),
.Y(n_10139)
);

INVx1_ASAP7_75t_L g10140 ( 
.A(n_8781),
.Y(n_10140)
);

OAI21x1_ASAP7_75t_L g10141 ( 
.A1(n_8628),
.A2(n_8644),
.B(n_8633),
.Y(n_10141)
);

AND2x2_ASAP7_75t_L g10142 ( 
.A(n_9399),
.B(n_8306),
.Y(n_10142)
);

OR2x2_ASAP7_75t_L g10143 ( 
.A(n_9000),
.B(n_8871),
.Y(n_10143)
);

INVx2_ASAP7_75t_L g10144 ( 
.A(n_9312),
.Y(n_10144)
);

OAI21x1_ASAP7_75t_L g10145 ( 
.A1(n_8628),
.A2(n_7907),
.B(n_7903),
.Y(n_10145)
);

INVx2_ASAP7_75t_SL g10146 ( 
.A(n_9174),
.Y(n_10146)
);

INVx2_ASAP7_75t_L g10147 ( 
.A(n_9315),
.Y(n_10147)
);

INVx1_ASAP7_75t_L g10148 ( 
.A(n_8781),
.Y(n_10148)
);

INVx1_ASAP7_75t_L g10149 ( 
.A(n_8784),
.Y(n_10149)
);

AND2x2_ASAP7_75t_L g10150 ( 
.A(n_8965),
.B(n_7452),
.Y(n_10150)
);

INVx1_ASAP7_75t_L g10151 ( 
.A(n_8784),
.Y(n_10151)
);

INVx1_ASAP7_75t_L g10152 ( 
.A(n_8789),
.Y(n_10152)
);

HB1xp67_ASAP7_75t_L g10153 ( 
.A(n_8670),
.Y(n_10153)
);

INVx3_ASAP7_75t_L g10154 ( 
.A(n_8633),
.Y(n_10154)
);

INVx1_ASAP7_75t_L g10155 ( 
.A(n_8789),
.Y(n_10155)
);

INVx2_ASAP7_75t_L g10156 ( 
.A(n_9315),
.Y(n_10156)
);

NAND2xp5_ASAP7_75t_L g10157 ( 
.A(n_9083),
.B(n_7479),
.Y(n_10157)
);

INVx3_ASAP7_75t_L g10158 ( 
.A(n_8633),
.Y(n_10158)
);

BUFx2_ASAP7_75t_L g10159 ( 
.A(n_8349),
.Y(n_10159)
);

HB1xp67_ASAP7_75t_L g10160 ( 
.A(n_8687),
.Y(n_10160)
);

INVx2_ASAP7_75t_L g10161 ( 
.A(n_9328),
.Y(n_10161)
);

OAI21x1_ASAP7_75t_L g10162 ( 
.A1(n_8633),
.A2(n_7917),
.B(n_7907),
.Y(n_10162)
);

INVx1_ASAP7_75t_L g10163 ( 
.A(n_8790),
.Y(n_10163)
);

AND2x2_ASAP7_75t_L g10164 ( 
.A(n_8965),
.B(n_8971),
.Y(n_10164)
);

AND2x2_ASAP7_75t_L g10165 ( 
.A(n_8971),
.B(n_7452),
.Y(n_10165)
);

BUFx3_ASAP7_75t_L g10166 ( 
.A(n_9028),
.Y(n_10166)
);

NAND2x1p5_ASAP7_75t_L g10167 ( 
.A(n_8788),
.B(n_7979),
.Y(n_10167)
);

INVx1_ASAP7_75t_L g10168 ( 
.A(n_8790),
.Y(n_10168)
);

INVx2_ASAP7_75t_L g10169 ( 
.A(n_9328),
.Y(n_10169)
);

BUFx2_ASAP7_75t_L g10170 ( 
.A(n_8349),
.Y(n_10170)
);

INVx3_ASAP7_75t_L g10171 ( 
.A(n_8644),
.Y(n_10171)
);

INVx2_ASAP7_75t_L g10172 ( 
.A(n_9334),
.Y(n_10172)
);

AND2x2_ASAP7_75t_L g10173 ( 
.A(n_8977),
.B(n_7466),
.Y(n_10173)
);

NAND2x1_ASAP7_75t_L g10174 ( 
.A(n_8325),
.B(n_7586),
.Y(n_10174)
);

OAI22xp5_ASAP7_75t_L g10175 ( 
.A1(n_8513),
.A2(n_8370),
.B1(n_8707),
.B2(n_8704),
.Y(n_10175)
);

INVx2_ASAP7_75t_L g10176 ( 
.A(n_9334),
.Y(n_10176)
);

INVx1_ASAP7_75t_L g10177 ( 
.A(n_8796),
.Y(n_10177)
);

HB1xp67_ASAP7_75t_L g10178 ( 
.A(n_8705),
.Y(n_10178)
);

OR2x2_ASAP7_75t_L g10179 ( 
.A(n_8871),
.B(n_7718),
.Y(n_10179)
);

AND2x4_ASAP7_75t_L g10180 ( 
.A(n_9230),
.B(n_8155),
.Y(n_10180)
);

HB1xp67_ASAP7_75t_L g10181 ( 
.A(n_8732),
.Y(n_10181)
);

INVx2_ASAP7_75t_L g10182 ( 
.A(n_9085),
.Y(n_10182)
);

INVx3_ASAP7_75t_L g10183 ( 
.A(n_8644),
.Y(n_10183)
);

INVx3_ASAP7_75t_L g10184 ( 
.A(n_8644),
.Y(n_10184)
);

NOR2x1_ASAP7_75t_R g10185 ( 
.A(n_9067),
.B(n_6629),
.Y(n_10185)
);

INVx3_ASAP7_75t_L g10186 ( 
.A(n_9044),
.Y(n_10186)
);

INVx2_ASAP7_75t_L g10187 ( 
.A(n_9093),
.Y(n_10187)
);

OAI21x1_ASAP7_75t_L g10188 ( 
.A1(n_8352),
.A2(n_7917),
.B(n_7692),
.Y(n_10188)
);

INVx2_ASAP7_75t_L g10189 ( 
.A(n_9095),
.Y(n_10189)
);

BUFx2_ASAP7_75t_L g10190 ( 
.A(n_8349),
.Y(n_10190)
);

INVx1_ASAP7_75t_SL g10191 ( 
.A(n_8541),
.Y(n_10191)
);

INVx2_ASAP7_75t_L g10192 ( 
.A(n_9095),
.Y(n_10192)
);

OAI21x1_ASAP7_75t_L g10193 ( 
.A1(n_8352),
.A2(n_7917),
.B(n_7692),
.Y(n_10193)
);

NOR2xp33_ASAP7_75t_L g10194 ( 
.A(n_9391),
.B(n_7479),
.Y(n_10194)
);

BUFx6f_ASAP7_75t_L g10195 ( 
.A(n_8327),
.Y(n_10195)
);

INVx1_ASAP7_75t_L g10196 ( 
.A(n_8796),
.Y(n_10196)
);

INVx1_ASAP7_75t_L g10197 ( 
.A(n_8800),
.Y(n_10197)
);

OAI21x1_ASAP7_75t_L g10198 ( 
.A1(n_8379),
.A2(n_7692),
.B(n_7687),
.Y(n_10198)
);

OR2x2_ASAP7_75t_L g10199 ( 
.A(n_8399),
.B(n_7718),
.Y(n_10199)
);

INVx1_ASAP7_75t_L g10200 ( 
.A(n_8800),
.Y(n_10200)
);

INVx1_ASAP7_75t_L g10201 ( 
.A(n_8804),
.Y(n_10201)
);

OAI21x1_ASAP7_75t_L g10202 ( 
.A1(n_8379),
.A2(n_7693),
.B(n_7687),
.Y(n_10202)
);

CKINVDCx5p33_ASAP7_75t_R g10203 ( 
.A(n_8589),
.Y(n_10203)
);

AND2x6_ASAP7_75t_L g10204 ( 
.A(n_8350),
.B(n_7987),
.Y(n_10204)
);

INVx1_ASAP7_75t_L g10205 ( 
.A(n_8804),
.Y(n_10205)
);

INVx1_ASAP7_75t_L g10206 ( 
.A(n_8807),
.Y(n_10206)
);

OR2x2_ASAP7_75t_L g10207 ( 
.A(n_8399),
.B(n_7718),
.Y(n_10207)
);

AND2x4_ASAP7_75t_L g10208 ( 
.A(n_9230),
.B(n_8155),
.Y(n_10208)
);

INVx2_ASAP7_75t_L g10209 ( 
.A(n_9100),
.Y(n_10209)
);

INVx1_ASAP7_75t_L g10210 ( 
.A(n_8807),
.Y(n_10210)
);

OA21x2_ASAP7_75t_L g10211 ( 
.A1(n_9100),
.A2(n_7232),
.B(n_7343),
.Y(n_10211)
);

INVx2_ASAP7_75t_SL g10212 ( 
.A(n_8859),
.Y(n_10212)
);

INVx1_ASAP7_75t_L g10213 ( 
.A(n_8812),
.Y(n_10213)
);

INVx3_ASAP7_75t_L g10214 ( 
.A(n_9044),
.Y(n_10214)
);

INVx2_ASAP7_75t_L g10215 ( 
.A(n_9121),
.Y(n_10215)
);

INVx1_ASAP7_75t_L g10216 ( 
.A(n_8812),
.Y(n_10216)
);

OAI21x1_ASAP7_75t_L g10217 ( 
.A1(n_9271),
.A2(n_7693),
.B(n_7687),
.Y(n_10217)
);

INVx2_ASAP7_75t_L g10218 ( 
.A(n_9121),
.Y(n_10218)
);

AOI22xp5_ASAP7_75t_L g10219 ( 
.A1(n_8704),
.A2(n_8707),
.B1(n_8894),
.B2(n_8877),
.Y(n_10219)
);

AND2x2_ASAP7_75t_L g10220 ( 
.A(n_8977),
.B(n_7466),
.Y(n_10220)
);

HB1xp67_ASAP7_75t_L g10221 ( 
.A(n_8767),
.Y(n_10221)
);

INVx1_ASAP7_75t_L g10222 ( 
.A(n_8821),
.Y(n_10222)
);

INVx3_ASAP7_75t_L g10223 ( 
.A(n_9044),
.Y(n_10223)
);

AND2x2_ASAP7_75t_L g10224 ( 
.A(n_8707),
.B(n_8877),
.Y(n_10224)
);

INVx1_ASAP7_75t_L g10225 ( 
.A(n_8821),
.Y(n_10225)
);

AOI22xp33_ASAP7_75t_L g10226 ( 
.A1(n_8707),
.A2(n_7234),
.B1(n_8017),
.B2(n_7632),
.Y(n_10226)
);

INVx1_ASAP7_75t_L g10227 ( 
.A(n_8836),
.Y(n_10227)
);

INVx1_ASAP7_75t_L g10228 ( 
.A(n_8836),
.Y(n_10228)
);

OR2x6_ASAP7_75t_L g10229 ( 
.A(n_9299),
.B(n_7713),
.Y(n_10229)
);

INVx1_ASAP7_75t_L g10230 ( 
.A(n_8842),
.Y(n_10230)
);

INVx2_ASAP7_75t_L g10231 ( 
.A(n_9134),
.Y(n_10231)
);

NAND2xp5_ASAP7_75t_L g10232 ( 
.A(n_8877),
.B(n_7486),
.Y(n_10232)
);

INVx1_ASAP7_75t_L g10233 ( 
.A(n_8842),
.Y(n_10233)
);

BUFx2_ASAP7_75t_L g10234 ( 
.A(n_8350),
.Y(n_10234)
);

AND2x2_ASAP7_75t_L g10235 ( 
.A(n_8877),
.B(n_7466),
.Y(n_10235)
);

INVx1_ASAP7_75t_L g10236 ( 
.A(n_8845),
.Y(n_10236)
);

BUFx6f_ASAP7_75t_L g10237 ( 
.A(n_8327),
.Y(n_10237)
);

INVx1_ASAP7_75t_L g10238 ( 
.A(n_8845),
.Y(n_10238)
);

INVx1_ASAP7_75t_L g10239 ( 
.A(n_8851),
.Y(n_10239)
);

INVx1_ASAP7_75t_L g10240 ( 
.A(n_8851),
.Y(n_10240)
);

INVx3_ASAP7_75t_L g10241 ( 
.A(n_9044),
.Y(n_10241)
);

INVx2_ASAP7_75t_L g10242 ( 
.A(n_9134),
.Y(n_10242)
);

INVx2_ASAP7_75t_SL g10243 ( 
.A(n_8859),
.Y(n_10243)
);

OAI22xp5_ASAP7_75t_L g10244 ( 
.A1(n_8513),
.A2(n_7612),
.B1(n_7868),
.B2(n_7398),
.Y(n_10244)
);

HB1xp67_ASAP7_75t_L g10245 ( 
.A(n_8805),
.Y(n_10245)
);

INVx1_ASAP7_75t_L g10246 ( 
.A(n_8862),
.Y(n_10246)
);

INVx1_ASAP7_75t_L g10247 ( 
.A(n_8862),
.Y(n_10247)
);

INVx3_ASAP7_75t_L g10248 ( 
.A(n_9044),
.Y(n_10248)
);

HB1xp67_ASAP7_75t_L g10249 ( 
.A(n_8846),
.Y(n_10249)
);

INVx2_ASAP7_75t_L g10250 ( 
.A(n_9326),
.Y(n_10250)
);

INVx2_ASAP7_75t_L g10251 ( 
.A(n_9326),
.Y(n_10251)
);

AO21x1_ASAP7_75t_SL g10252 ( 
.A1(n_9119),
.A2(n_8137),
.B(n_8098),
.Y(n_10252)
);

HB1xp67_ASAP7_75t_L g10253 ( 
.A(n_8848),
.Y(n_10253)
);

INVx2_ASAP7_75t_L g10254 ( 
.A(n_9326),
.Y(n_10254)
);

INVx2_ASAP7_75t_L g10255 ( 
.A(n_9326),
.Y(n_10255)
);

NOR2xp33_ASAP7_75t_L g10256 ( 
.A(n_9313),
.B(n_7612),
.Y(n_10256)
);

AND2x4_ASAP7_75t_L g10257 ( 
.A(n_9230),
.B(n_9390),
.Y(n_10257)
);

INVx3_ASAP7_75t_L g10258 ( 
.A(n_9233),
.Y(n_10258)
);

INVx1_ASAP7_75t_L g10259 ( 
.A(n_8864),
.Y(n_10259)
);

INVx1_ASAP7_75t_L g10260 ( 
.A(n_8864),
.Y(n_10260)
);

OA21x2_ASAP7_75t_L g10261 ( 
.A1(n_8652),
.A2(n_9218),
.B(n_9211),
.Y(n_10261)
);

INVx2_ASAP7_75t_L g10262 ( 
.A(n_9335),
.Y(n_10262)
);

AOI21x1_ASAP7_75t_L g10263 ( 
.A1(n_8838),
.A2(n_7999),
.B(n_8196),
.Y(n_10263)
);

AOI21xp33_ASAP7_75t_SL g10264 ( 
.A1(n_9147),
.A2(n_6223),
.B(n_7795),
.Y(n_10264)
);

BUFx3_ASAP7_75t_L g10265 ( 
.A(n_9170),
.Y(n_10265)
);

INVx1_ASAP7_75t_L g10266 ( 
.A(n_8865),
.Y(n_10266)
);

INVx1_ASAP7_75t_L g10267 ( 
.A(n_8865),
.Y(n_10267)
);

INVx2_ASAP7_75t_L g10268 ( 
.A(n_9335),
.Y(n_10268)
);

INVx1_ASAP7_75t_L g10269 ( 
.A(n_8866),
.Y(n_10269)
);

BUFx10_ASAP7_75t_L g10270 ( 
.A(n_8859),
.Y(n_10270)
);

HB1xp67_ASAP7_75t_L g10271 ( 
.A(n_8878),
.Y(n_10271)
);

AND2x2_ASAP7_75t_L g10272 ( 
.A(n_8894),
.B(n_7469),
.Y(n_10272)
);

AND2x4_ASAP7_75t_L g10273 ( 
.A(n_9390),
.B(n_9416),
.Y(n_10273)
);

INVx1_ASAP7_75t_L g10274 ( 
.A(n_8866),
.Y(n_10274)
);

BUFx6f_ASAP7_75t_L g10275 ( 
.A(n_8327),
.Y(n_10275)
);

INVx2_ASAP7_75t_L g10276 ( 
.A(n_9335),
.Y(n_10276)
);

INVx1_ASAP7_75t_L g10277 ( 
.A(n_8885),
.Y(n_10277)
);

OAI22xp5_ASAP7_75t_L g10278 ( 
.A1(n_8370),
.A2(n_7868),
.B1(n_7398),
.B2(n_7477),
.Y(n_10278)
);

INVx1_ASAP7_75t_L g10279 ( 
.A(n_8885),
.Y(n_10279)
);

AOI222xp33_ASAP7_75t_L g10280 ( 
.A1(n_9122),
.A2(n_7876),
.B1(n_7838),
.B2(n_7591),
.C1(n_8147),
.C2(n_8260),
.Y(n_10280)
);

INVx3_ASAP7_75t_L g10281 ( 
.A(n_9233),
.Y(n_10281)
);

AOI22xp33_ASAP7_75t_L g10282 ( 
.A1(n_8894),
.A2(n_8017),
.B1(n_7632),
.B2(n_7168),
.Y(n_10282)
);

INVx1_ASAP7_75t_L g10283 ( 
.A(n_8898),
.Y(n_10283)
);

OAI21x1_ASAP7_75t_L g10284 ( 
.A1(n_9271),
.A2(n_7695),
.B(n_7693),
.Y(n_10284)
);

INVxp67_ASAP7_75t_L g10285 ( 
.A(n_8535),
.Y(n_10285)
);

INVxp67_ASAP7_75t_L g10286 ( 
.A(n_8640),
.Y(n_10286)
);

AOI22xp33_ASAP7_75t_SL g10287 ( 
.A1(n_8894),
.A2(n_7662),
.B1(n_7660),
.B2(n_7632),
.Y(n_10287)
);

INVx1_ASAP7_75t_L g10288 ( 
.A(n_8898),
.Y(n_10288)
);

INVx4_ASAP7_75t_SL g10289 ( 
.A(n_8392),
.Y(n_10289)
);

INVx1_ASAP7_75t_L g10290 ( 
.A(n_8914),
.Y(n_10290)
);

INVx2_ASAP7_75t_L g10291 ( 
.A(n_9335),
.Y(n_10291)
);

INVxp67_ASAP7_75t_L g10292 ( 
.A(n_9022),
.Y(n_10292)
);

HB1xp67_ASAP7_75t_L g10293 ( 
.A(n_8936),
.Y(n_10293)
);

INVx2_ASAP7_75t_L g10294 ( 
.A(n_9336),
.Y(n_10294)
);

INVx1_ASAP7_75t_L g10295 ( 
.A(n_8914),
.Y(n_10295)
);

BUFx2_ASAP7_75t_L g10296 ( 
.A(n_8350),
.Y(n_10296)
);

INVx2_ASAP7_75t_L g10297 ( 
.A(n_9336),
.Y(n_10297)
);

BUFx2_ASAP7_75t_L g10298 ( 
.A(n_8354),
.Y(n_10298)
);

OAI21x1_ASAP7_75t_L g10299 ( 
.A1(n_9283),
.A2(n_7695),
.B(n_7658),
.Y(n_10299)
);

INVx1_ASAP7_75t_L g10300 ( 
.A(n_8916),
.Y(n_10300)
);

AND2x2_ASAP7_75t_L g10301 ( 
.A(n_8911),
.B(n_7469),
.Y(n_10301)
);

INVx2_ASAP7_75t_L g10302 ( 
.A(n_9336),
.Y(n_10302)
);

INVx1_ASAP7_75t_L g10303 ( 
.A(n_8916),
.Y(n_10303)
);

INVx1_ASAP7_75t_L g10304 ( 
.A(n_8918),
.Y(n_10304)
);

OR2x2_ASAP7_75t_L g10305 ( 
.A(n_8506),
.B(n_7718),
.Y(n_10305)
);

INVx1_ASAP7_75t_L g10306 ( 
.A(n_8918),
.Y(n_10306)
);

INVx1_ASAP7_75t_L g10307 ( 
.A(n_8919),
.Y(n_10307)
);

INVx2_ASAP7_75t_SL g10308 ( 
.A(n_8859),
.Y(n_10308)
);

OAI22xp5_ASAP7_75t_L g10309 ( 
.A1(n_8911),
.A2(n_7477),
.B1(n_7811),
.B2(n_8263),
.Y(n_10309)
);

INVx1_ASAP7_75t_L g10310 ( 
.A(n_8919),
.Y(n_10310)
);

INVx2_ASAP7_75t_L g10311 ( 
.A(n_9336),
.Y(n_10311)
);

INVx1_ASAP7_75t_L g10312 ( 
.A(n_8920),
.Y(n_10312)
);

BUFx3_ASAP7_75t_L g10313 ( 
.A(n_8354),
.Y(n_10313)
);

INVx2_ASAP7_75t_L g10314 ( 
.A(n_9350),
.Y(n_10314)
);

INVx1_ASAP7_75t_L g10315 ( 
.A(n_8920),
.Y(n_10315)
);

INVx1_ASAP7_75t_SL g10316 ( 
.A(n_8737),
.Y(n_10316)
);

OR2x6_ASAP7_75t_L g10317 ( 
.A(n_9299),
.B(n_7185),
.Y(n_10317)
);

BUFx6f_ASAP7_75t_L g10318 ( 
.A(n_8327),
.Y(n_10318)
);

INVx3_ASAP7_75t_L g10319 ( 
.A(n_9233),
.Y(n_10319)
);

AOI22xp5_ASAP7_75t_L g10320 ( 
.A1(n_8911),
.A2(n_8923),
.B1(n_8937),
.B2(n_8922),
.Y(n_10320)
);

INVx2_ASAP7_75t_SL g10321 ( 
.A(n_8859),
.Y(n_10321)
);

INVx2_ASAP7_75t_SL g10322 ( 
.A(n_8867),
.Y(n_10322)
);

AO21x2_ASAP7_75t_L g10323 ( 
.A1(n_9109),
.A2(n_7751),
.B(n_7724),
.Y(n_10323)
);

INVx1_ASAP7_75t_SL g10324 ( 
.A(n_8760),
.Y(n_10324)
);

INVx2_ASAP7_75t_L g10325 ( 
.A(n_9350),
.Y(n_10325)
);

AOI21xp5_ASAP7_75t_L g10326 ( 
.A1(n_8389),
.A2(n_7341),
.B(n_7567),
.Y(n_10326)
);

BUFx2_ASAP7_75t_L g10327 ( 
.A(n_8354),
.Y(n_10327)
);

INVx1_ASAP7_75t_L g10328 ( 
.A(n_8924),
.Y(n_10328)
);

INVx2_ASAP7_75t_L g10329 ( 
.A(n_9350),
.Y(n_10329)
);

INVx2_ASAP7_75t_L g10330 ( 
.A(n_9350),
.Y(n_10330)
);

INVx2_ASAP7_75t_L g10331 ( 
.A(n_9362),
.Y(n_10331)
);

HB1xp67_ASAP7_75t_L g10332 ( 
.A(n_9006),
.Y(n_10332)
);

BUFx2_ASAP7_75t_L g10333 ( 
.A(n_8528),
.Y(n_10333)
);

INVx1_ASAP7_75t_L g10334 ( 
.A(n_8924),
.Y(n_10334)
);

INVx1_ASAP7_75t_L g10335 ( 
.A(n_8939),
.Y(n_10335)
);

INVx3_ASAP7_75t_L g10336 ( 
.A(n_9233),
.Y(n_10336)
);

INVx2_ASAP7_75t_L g10337 ( 
.A(n_9362),
.Y(n_10337)
);

INVx2_ASAP7_75t_L g10338 ( 
.A(n_9362),
.Y(n_10338)
);

NOR2xp33_ASAP7_75t_L g10339 ( 
.A(n_9343),
.B(n_8024),
.Y(n_10339)
);

INVx2_ASAP7_75t_L g10340 ( 
.A(n_9362),
.Y(n_10340)
);

OR2x2_ASAP7_75t_L g10341 ( 
.A(n_8506),
.B(n_7718),
.Y(n_10341)
);

OAI21x1_ASAP7_75t_L g10342 ( 
.A1(n_9283),
.A2(n_7695),
.B(n_7658),
.Y(n_10342)
);

OAI21x1_ASAP7_75t_L g10343 ( 
.A1(n_9298),
.A2(n_7658),
.B(n_7657),
.Y(n_10343)
);

AOI22xp33_ASAP7_75t_L g10344 ( 
.A1(n_8911),
.A2(n_8017),
.B1(n_7632),
.B2(n_7168),
.Y(n_10344)
);

INVx1_ASAP7_75t_L g10345 ( 
.A(n_8939),
.Y(n_10345)
);

INVx2_ASAP7_75t_L g10346 ( 
.A(n_9378),
.Y(n_10346)
);

INVx1_ASAP7_75t_L g10347 ( 
.A(n_8942),
.Y(n_10347)
);

INVx1_ASAP7_75t_L g10348 ( 
.A(n_8942),
.Y(n_10348)
);

INVx1_ASAP7_75t_L g10349 ( 
.A(n_8950),
.Y(n_10349)
);

INVx3_ASAP7_75t_L g10350 ( 
.A(n_9233),
.Y(n_10350)
);

INVx1_ASAP7_75t_L g10351 ( 
.A(n_8950),
.Y(n_10351)
);

AOI21x1_ASAP7_75t_L g10352 ( 
.A1(n_8838),
.A2(n_8245),
.B(n_8196),
.Y(n_10352)
);

AOI21xp5_ASAP7_75t_L g10353 ( 
.A1(n_8335),
.A2(n_7567),
.B(n_7440),
.Y(n_10353)
);

OAI21xp5_ASAP7_75t_L g10354 ( 
.A1(n_8547),
.A2(n_7440),
.B(n_8147),
.Y(n_10354)
);

INVx1_ASAP7_75t_L g10355 ( 
.A(n_8951),
.Y(n_10355)
);

INVx1_ASAP7_75t_L g10356 ( 
.A(n_8951),
.Y(n_10356)
);

OAI21x1_ASAP7_75t_L g10357 ( 
.A1(n_9298),
.A2(n_7667),
.B(n_7657),
.Y(n_10357)
);

BUFx2_ASAP7_75t_L g10358 ( 
.A(n_8528),
.Y(n_10358)
);

BUFx2_ASAP7_75t_L g10359 ( 
.A(n_8528),
.Y(n_10359)
);

AND2x4_ASAP7_75t_L g10360 ( 
.A(n_9390),
.B(n_8263),
.Y(n_10360)
);

INVx1_ASAP7_75t_L g10361 ( 
.A(n_8957),
.Y(n_10361)
);

BUFx3_ASAP7_75t_L g10362 ( 
.A(n_8908),
.Y(n_10362)
);

BUFx2_ASAP7_75t_L g10363 ( 
.A(n_8581),
.Y(n_10363)
);

INVx1_ASAP7_75t_L g10364 ( 
.A(n_8957),
.Y(n_10364)
);

BUFx3_ASAP7_75t_L g10365 ( 
.A(n_8867),
.Y(n_10365)
);

AND2x2_ASAP7_75t_L g10366 ( 
.A(n_8922),
.B(n_7469),
.Y(n_10366)
);

BUFx2_ASAP7_75t_SL g10367 ( 
.A(n_9175),
.Y(n_10367)
);

INVx2_ASAP7_75t_L g10368 ( 
.A(n_9378),
.Y(n_10368)
);

INVxp67_ASAP7_75t_L g10369 ( 
.A(n_8552),
.Y(n_10369)
);

NAND2xp5_ASAP7_75t_L g10370 ( 
.A(n_8922),
.B(n_7838),
.Y(n_10370)
);

INVx2_ASAP7_75t_L g10371 ( 
.A(n_9378),
.Y(n_10371)
);

INVx1_ASAP7_75t_L g10372 ( 
.A(n_8960),
.Y(n_10372)
);

INVx1_ASAP7_75t_L g10373 ( 
.A(n_8960),
.Y(n_10373)
);

INVx1_ASAP7_75t_L g10374 ( 
.A(n_8961),
.Y(n_10374)
);

OAI21x1_ASAP7_75t_L g10375 ( 
.A1(n_9303),
.A2(n_7667),
.B(n_7657),
.Y(n_10375)
);

OAI21x1_ASAP7_75t_L g10376 ( 
.A1(n_9303),
.A2(n_7675),
.B(n_7667),
.Y(n_10376)
);

BUFx3_ASAP7_75t_L g10377 ( 
.A(n_8867),
.Y(n_10377)
);

INVx2_ASAP7_75t_L g10378 ( 
.A(n_9378),
.Y(n_10378)
);

INVx1_ASAP7_75t_L g10379 ( 
.A(n_8961),
.Y(n_10379)
);

INVx2_ASAP7_75t_L g10380 ( 
.A(n_9211),
.Y(n_10380)
);

OAI21x1_ASAP7_75t_L g10381 ( 
.A1(n_8398),
.A2(n_7675),
.B(n_7594),
.Y(n_10381)
);

INVx2_ASAP7_75t_L g10382 ( 
.A(n_9218),
.Y(n_10382)
);

AND2x2_ASAP7_75t_L g10383 ( 
.A(n_8922),
.B(n_7492),
.Y(n_10383)
);

INVxp67_ASAP7_75t_L g10384 ( 
.A(n_8754),
.Y(n_10384)
);

OAI21x1_ASAP7_75t_L g10385 ( 
.A1(n_8398),
.A2(n_7675),
.B(n_7594),
.Y(n_10385)
);

AO21x2_ASAP7_75t_L g10386 ( 
.A1(n_9262),
.A2(n_7751),
.B(n_7724),
.Y(n_10386)
);

AOI21xp33_ASAP7_75t_L g10387 ( 
.A1(n_8476),
.A2(n_7247),
.B(n_7588),
.Y(n_10387)
);

INVx2_ASAP7_75t_L g10388 ( 
.A(n_9220),
.Y(n_10388)
);

INVx1_ASAP7_75t_L g10389 ( 
.A(n_8963),
.Y(n_10389)
);

AO21x2_ASAP7_75t_L g10390 ( 
.A1(n_9262),
.A2(n_7167),
.B(n_7845),
.Y(n_10390)
);

INVxp67_ASAP7_75t_L g10391 ( 
.A(n_8754),
.Y(n_10391)
);

NAND2xp5_ASAP7_75t_L g10392 ( 
.A(n_8923),
.B(n_7876),
.Y(n_10392)
);

AO21x1_ASAP7_75t_L g10393 ( 
.A1(n_8665),
.A2(n_7392),
.B(n_7376),
.Y(n_10393)
);

AND2x2_ASAP7_75t_L g10394 ( 
.A(n_8923),
.B(n_7492),
.Y(n_10394)
);

AND2x2_ASAP7_75t_L g10395 ( 
.A(n_8923),
.B(n_7492),
.Y(n_10395)
);

INVx4_ASAP7_75t_SL g10396 ( 
.A(n_8392),
.Y(n_10396)
);

INVx1_ASAP7_75t_L g10397 ( 
.A(n_8963),
.Y(n_10397)
);

AND2x2_ASAP7_75t_L g10398 ( 
.A(n_8937),
.B(n_7522),
.Y(n_10398)
);

INVx1_ASAP7_75t_L g10399 ( 
.A(n_8964),
.Y(n_10399)
);

INVx2_ASAP7_75t_L g10400 ( 
.A(n_9220),
.Y(n_10400)
);

INVx1_ASAP7_75t_L g10401 ( 
.A(n_8964),
.Y(n_10401)
);

INVx2_ASAP7_75t_SL g10402 ( 
.A(n_8867),
.Y(n_10402)
);

OAI21xp5_ASAP7_75t_L g10403 ( 
.A1(n_9122),
.A2(n_7392),
.B(n_7376),
.Y(n_10403)
);

INVx3_ASAP7_75t_L g10404 ( 
.A(n_8558),
.Y(n_10404)
);

AND2x2_ASAP7_75t_L g10405 ( 
.A(n_8937),
.B(n_7522),
.Y(n_10405)
);

BUFx6f_ASAP7_75t_L g10406 ( 
.A(n_8345),
.Y(n_10406)
);

INVx3_ASAP7_75t_L g10407 ( 
.A(n_8558),
.Y(n_10407)
);

AOI21x1_ASAP7_75t_L g10408 ( 
.A1(n_8874),
.A2(n_8245),
.B(n_8196),
.Y(n_10408)
);

INVx2_ASAP7_75t_L g10409 ( 
.A(n_9235),
.Y(n_10409)
);

INVx2_ASAP7_75t_L g10410 ( 
.A(n_9235),
.Y(n_10410)
);

NAND2xp5_ASAP7_75t_L g10411 ( 
.A(n_8937),
.B(n_8293),
.Y(n_10411)
);

AND2x2_ASAP7_75t_L g10412 ( 
.A(n_9045),
.B(n_7522),
.Y(n_10412)
);

OAI211xp5_ASAP7_75t_L g10413 ( 
.A1(n_9661),
.A2(n_9366),
.B(n_9175),
.C(n_9228),
.Y(n_10413)
);

INVx2_ASAP7_75t_L g10414 ( 
.A(n_9642),
.Y(n_10414)
);

AOI221xp5_ASAP7_75t_L g10415 ( 
.A1(n_9510),
.A2(n_9409),
.B1(n_9403),
.B2(n_9102),
.C(n_9337),
.Y(n_10415)
);

INVx2_ASAP7_75t_L g10416 ( 
.A(n_9583),
.Y(n_10416)
);

OAI22xp5_ASAP7_75t_L g10417 ( 
.A1(n_9837),
.A2(n_8419),
.B1(n_8321),
.B2(n_8572),
.Y(n_10417)
);

INVx1_ASAP7_75t_L g10418 ( 
.A(n_9669),
.Y(n_10418)
);

AND2x4_ASAP7_75t_L g10419 ( 
.A(n_9584),
.B(n_10313),
.Y(n_10419)
);

NAND2xp5_ASAP7_75t_L g10420 ( 
.A(n_10068),
.B(n_8772),
.Y(n_10420)
);

AOI22xp33_ASAP7_75t_L g10421 ( 
.A1(n_9510),
.A2(n_9948),
.B1(n_9606),
.B2(n_10280),
.Y(n_10421)
);

INVx1_ASAP7_75t_L g10422 ( 
.A(n_9708),
.Y(n_10422)
);

OAI21xp5_ASAP7_75t_L g10423 ( 
.A1(n_9639),
.A2(n_8471),
.B(n_8476),
.Y(n_10423)
);

AOI22xp5_ASAP7_75t_L g10424 ( 
.A1(n_9948),
.A2(n_8930),
.B1(n_8844),
.B2(n_8426),
.Y(n_10424)
);

AOI221xp5_ASAP7_75t_L g10425 ( 
.A1(n_9562),
.A2(n_9337),
.B1(n_9273),
.B2(n_8530),
.C(n_8572),
.Y(n_10425)
);

AOI211xp5_ASAP7_75t_L g10426 ( 
.A1(n_9713),
.A2(n_8771),
.B(n_8665),
.C(n_8623),
.Y(n_10426)
);

AOI221xp5_ASAP7_75t_L g10427 ( 
.A1(n_10354),
.A2(n_9273),
.B1(n_8530),
.B2(n_8771),
.C(n_8776),
.Y(n_10427)
);

HB1xp67_ASAP7_75t_L g10428 ( 
.A(n_9451),
.Y(n_10428)
);

OAI22xp33_ASAP7_75t_L g10429 ( 
.A1(n_9780),
.A2(n_9299),
.B1(n_8700),
.B2(n_8321),
.Y(n_10429)
);

INVx2_ASAP7_75t_L g10430 ( 
.A(n_9583),
.Y(n_10430)
);

OAI211xp5_ASAP7_75t_L g10431 ( 
.A1(n_9579),
.A2(n_9228),
.B(n_9175),
.C(n_8338),
.Y(n_10431)
);

OAI221xp5_ASAP7_75t_L g10432 ( 
.A1(n_9500),
.A2(n_8473),
.B1(n_8982),
.B2(n_8979),
.C(n_9380),
.Y(n_10432)
);

INVx1_ASAP7_75t_L g10433 ( 
.A(n_9439),
.Y(n_10433)
);

OR2x2_ASAP7_75t_L g10434 ( 
.A(n_9598),
.B(n_7718),
.Y(n_10434)
);

OAI21x1_ASAP7_75t_L g10435 ( 
.A1(n_9754),
.A2(n_9442),
.B(n_10352),
.Y(n_10435)
);

BUFx5_ASAP7_75t_L g10436 ( 
.A(n_9860),
.Y(n_10436)
);

AND2x2_ASAP7_75t_L g10437 ( 
.A(n_9453),
.B(n_8555),
.Y(n_10437)
);

INVx1_ASAP7_75t_L g10438 ( 
.A(n_9446),
.Y(n_10438)
);

AO21x2_ASAP7_75t_L g10439 ( 
.A1(n_9639),
.A2(n_8776),
.B(n_8731),
.Y(n_10439)
);

INVx2_ASAP7_75t_L g10440 ( 
.A(n_9680),
.Y(n_10440)
);

OR2x6_ASAP7_75t_SL g10441 ( 
.A(n_10203),
.B(n_8768),
.Y(n_10441)
);

AOI21xp5_ASAP7_75t_L g10442 ( 
.A1(n_9579),
.A2(n_8471),
.B(n_8798),
.Y(n_10442)
);

BUFx4f_ASAP7_75t_SL g10443 ( 
.A(n_9473),
.Y(n_10443)
);

INVx2_ASAP7_75t_L g10444 ( 
.A(n_9680),
.Y(n_10444)
);

BUFx3_ASAP7_75t_L g10445 ( 
.A(n_9473),
.Y(n_10445)
);

AND2x2_ASAP7_75t_L g10446 ( 
.A(n_9587),
.B(n_8555),
.Y(n_10446)
);

INVx1_ASAP7_75t_L g10447 ( 
.A(n_9450),
.Y(n_10447)
);

AO31x2_ASAP7_75t_L g10448 ( 
.A1(n_10175),
.A2(n_8731),
.A3(n_8882),
.B(n_8623),
.Y(n_10448)
);

OAI22xp33_ASAP7_75t_L g10449 ( 
.A1(n_9520),
.A2(n_8700),
.B1(n_8722),
.B2(n_8966),
.Y(n_10449)
);

AOI21xp33_ASAP7_75t_SL g10450 ( 
.A1(n_9903),
.A2(n_8498),
.B(n_8952),
.Y(n_10450)
);

AOI22xp33_ASAP7_75t_L g10451 ( 
.A1(n_9448),
.A2(n_8930),
.B1(n_8452),
.B2(n_8460),
.Y(n_10451)
);

AOI22xp33_ASAP7_75t_L g10452 ( 
.A1(n_9448),
.A2(n_8930),
.B1(n_8469),
.B2(n_8444),
.Y(n_10452)
);

OR2x6_ASAP7_75t_L g10453 ( 
.A(n_9860),
.B(n_9946),
.Y(n_10453)
);

AOI22xp33_ASAP7_75t_SL g10454 ( 
.A1(n_9463),
.A2(n_9236),
.B1(n_9245),
.B2(n_9242),
.Y(n_10454)
);

AOI22xp33_ASAP7_75t_L g10455 ( 
.A1(n_9463),
.A2(n_8449),
.B1(n_8501),
.B2(n_9236),
.Y(n_10455)
);

AOI22xp33_ASAP7_75t_SL g10456 ( 
.A1(n_9480),
.A2(n_9242),
.B1(n_9250),
.B2(n_9245),
.Y(n_10456)
);

AOI22xp33_ASAP7_75t_L g10457 ( 
.A1(n_9469),
.A2(n_9250),
.B1(n_9255),
.B2(n_9254),
.Y(n_10457)
);

AOI22xp33_ASAP7_75t_L g10458 ( 
.A1(n_9469),
.A2(n_9254),
.B1(n_9257),
.B2(n_9255),
.Y(n_10458)
);

AOI22xp33_ASAP7_75t_L g10459 ( 
.A1(n_9480),
.A2(n_9257),
.B1(n_9261),
.B2(n_8755),
.Y(n_10459)
);

OAI22xp33_ASAP7_75t_L g10460 ( 
.A1(n_10114),
.A2(n_8722),
.B1(n_8966),
.B2(n_9180),
.Y(n_10460)
);

AOI22xp33_ASAP7_75t_L g10461 ( 
.A1(n_10393),
.A2(n_9261),
.B1(n_8336),
.B2(n_8443),
.Y(n_10461)
);

INVx1_ASAP7_75t_L g10462 ( 
.A(n_9460),
.Y(n_10462)
);

AOI21xp5_ASAP7_75t_L g10463 ( 
.A1(n_9713),
.A2(n_9377),
.B(n_8339),
.Y(n_10463)
);

AOI22xp33_ASAP7_75t_L g10464 ( 
.A1(n_10393),
.A2(n_9723),
.B1(n_9589),
.B2(n_9715),
.Y(n_10464)
);

AND2x2_ASAP7_75t_L g10465 ( 
.A(n_9587),
.B(n_8581),
.Y(n_10465)
);

NAND2xp5_ASAP7_75t_L g10466 ( 
.A(n_10071),
.B(n_9069),
.Y(n_10466)
);

AOI21xp5_ASAP7_75t_L g10467 ( 
.A1(n_10326),
.A2(n_8616),
.B(n_8931),
.Y(n_10467)
);

INVx1_ASAP7_75t_L g10468 ( 
.A(n_9471),
.Y(n_10468)
);

OAI211xp5_ASAP7_75t_SL g10469 ( 
.A1(n_10353),
.A2(n_9758),
.B(n_9476),
.C(n_10118),
.Y(n_10469)
);

INVx1_ASAP7_75t_L g10470 ( 
.A(n_9472),
.Y(n_10470)
);

NAND2xp5_ASAP7_75t_L g10471 ( 
.A(n_9614),
.B(n_7718),
.Y(n_10471)
);

AOI22xp33_ASAP7_75t_L g10472 ( 
.A1(n_9723),
.A2(n_9589),
.B1(n_9715),
.B2(n_9633),
.Y(n_10472)
);

OAI22xp5_ASAP7_75t_L g10473 ( 
.A1(n_9837),
.A2(n_9079),
.B1(n_9127),
.B2(n_8489),
.Y(n_10473)
);

AND2x2_ASAP7_75t_L g10474 ( 
.A(n_9853),
.B(n_8581),
.Y(n_10474)
);

OAI221xp5_ASAP7_75t_L g10475 ( 
.A1(n_9500),
.A2(n_9180),
.B1(n_9388),
.B2(n_8969),
.C(n_8927),
.Y(n_10475)
);

AOI221xp5_ASAP7_75t_SL g10476 ( 
.A1(n_9537),
.A2(n_8980),
.B1(n_9369),
.B2(n_8539),
.C(n_9285),
.Y(n_10476)
);

AO221x2_ASAP7_75t_L g10477 ( 
.A1(n_9540),
.A2(n_8852),
.B1(n_8891),
.B2(n_8676),
.C(n_8944),
.Y(n_10477)
);

INVx1_ASAP7_75t_L g10478 ( 
.A(n_9474),
.Y(n_10478)
);

OAI21xp5_ASAP7_75t_SL g10479 ( 
.A1(n_9685),
.A2(n_8723),
.B(n_8721),
.Y(n_10479)
);

OAI22xp5_ASAP7_75t_L g10480 ( 
.A1(n_9804),
.A2(n_8607),
.B1(n_8595),
.B2(n_8946),
.Y(n_10480)
);

INVx5_ASAP7_75t_SL g10481 ( 
.A(n_9770),
.Y(n_10481)
);

OAI22xp33_ASAP7_75t_L g10482 ( 
.A1(n_10087),
.A2(n_8263),
.B1(n_7704),
.B2(n_7893),
.Y(n_10482)
);

AND2x4_ASAP7_75t_L g10483 ( 
.A(n_9584),
.B(n_8588),
.Y(n_10483)
);

AOI221xp5_ASAP7_75t_L g10484 ( 
.A1(n_9572),
.A2(n_8882),
.B1(n_8903),
.B2(n_8967),
.C(n_8958),
.Y(n_10484)
);

HB1xp67_ASAP7_75t_L g10485 ( 
.A(n_9459),
.Y(n_10485)
);

OAI221xp5_ASAP7_75t_SL g10486 ( 
.A1(n_9757),
.A2(n_8315),
.B1(n_7337),
.B2(n_9386),
.C(n_8597),
.Y(n_10486)
);

AOI22xp33_ASAP7_75t_L g10487 ( 
.A1(n_9589),
.A2(n_8675),
.B1(n_8017),
.B2(n_8358),
.Y(n_10487)
);

AOI21xp5_ASAP7_75t_L g10488 ( 
.A1(n_10029),
.A2(n_8897),
.B(n_8325),
.Y(n_10488)
);

OAI211xp5_ASAP7_75t_L g10489 ( 
.A1(n_10403),
.A2(n_9228),
.B(n_7643),
.C(n_8774),
.Y(n_10489)
);

OAI22xp5_ASAP7_75t_L g10490 ( 
.A1(n_9875),
.A2(n_9925),
.B1(n_10244),
.B2(n_9794),
.Y(n_10490)
);

BUFx6f_ASAP7_75t_L g10491 ( 
.A(n_9770),
.Y(n_10491)
);

AOI22xp33_ASAP7_75t_L g10492 ( 
.A1(n_9633),
.A2(n_8017),
.B1(n_8677),
.B2(n_9005),
.Y(n_10492)
);

INVx1_ASAP7_75t_L g10493 ( 
.A(n_9475),
.Y(n_10493)
);

OAI22xp5_ASAP7_75t_SL g10494 ( 
.A1(n_9685),
.A2(n_9428),
.B1(n_6647),
.B2(n_6649),
.Y(n_10494)
);

INVx3_ASAP7_75t_L g10495 ( 
.A(n_9770),
.Y(n_10495)
);

AOI22xp33_ASAP7_75t_L g10496 ( 
.A1(n_9633),
.A2(n_8017),
.B1(n_9338),
.B2(n_7660),
.Y(n_10496)
);

INVx2_ASAP7_75t_SL g10497 ( 
.A(n_9778),
.Y(n_10497)
);

INVx3_ASAP7_75t_L g10498 ( 
.A(n_9770),
.Y(n_10498)
);

NOR2xp33_ASAP7_75t_L g10499 ( 
.A(n_9778),
.B(n_8575),
.Y(n_10499)
);

OAI321xp33_ASAP7_75t_L g10500 ( 
.A1(n_9438),
.A2(n_8615),
.A3(n_8708),
.B1(n_8785),
.B2(n_8463),
.C(n_8932),
.Y(n_10500)
);

OAI211xp5_ASAP7_75t_L g10501 ( 
.A1(n_9522),
.A2(n_7643),
.B(n_8774),
.C(n_8726),
.Y(n_10501)
);

HB1xp67_ASAP7_75t_L g10502 ( 
.A(n_9464),
.Y(n_10502)
);

AOI21xp33_ASAP7_75t_L g10503 ( 
.A1(n_9458),
.A2(n_7247),
.B(n_8991),
.Y(n_10503)
);

INVx1_ASAP7_75t_L g10504 ( 
.A(n_9477),
.Y(n_10504)
);

OAI22xp33_ASAP7_75t_SL g10505 ( 
.A1(n_10199),
.A2(n_8263),
.B1(n_8308),
.B2(n_8305),
.Y(n_10505)
);

AOI22xp33_ASAP7_75t_L g10506 ( 
.A1(n_9715),
.A2(n_9522),
.B1(n_9751),
.B2(n_9517),
.Y(n_10506)
);

NAND2xp5_ASAP7_75t_L g10507 ( 
.A(n_9530),
.B(n_7718),
.Y(n_10507)
);

OAI22xp33_ASAP7_75t_L g10508 ( 
.A1(n_10143),
.A2(n_9644),
.B1(n_9660),
.B2(n_9779),
.Y(n_10508)
);

BUFx6f_ASAP7_75t_L g10509 ( 
.A(n_9729),
.Y(n_10509)
);

INVx2_ASAP7_75t_L g10510 ( 
.A(n_9797),
.Y(n_10510)
);

OAI22xp5_ASAP7_75t_L g10511 ( 
.A1(n_9495),
.A2(n_8607),
.B1(n_8595),
.B2(n_8481),
.Y(n_10511)
);

NOR2xp33_ASAP7_75t_L g10512 ( 
.A(n_9699),
.B(n_8599),
.Y(n_10512)
);

OAI22xp33_ASAP7_75t_L g10513 ( 
.A1(n_9644),
.A2(n_7704),
.B1(n_9021),
.B2(n_8481),
.Y(n_10513)
);

AOI22xp33_ASAP7_75t_L g10514 ( 
.A1(n_9751),
.A2(n_7660),
.B1(n_7662),
.B2(n_7632),
.Y(n_10514)
);

AOI21xp5_ASAP7_75t_L g10515 ( 
.A1(n_10016),
.A2(n_9318),
.B(n_7450),
.Y(n_10515)
);

A2O1A1Ixp33_ASAP7_75t_L g10516 ( 
.A1(n_10387),
.A2(n_7461),
.B(n_7444),
.C(n_7337),
.Y(n_10516)
);

NAND2xp5_ASAP7_75t_L g10517 ( 
.A(n_9851),
.B(n_7674),
.Y(n_10517)
);

OAI21x1_ASAP7_75t_L g10518 ( 
.A1(n_10408),
.A2(n_9709),
.B(n_9643),
.Y(n_10518)
);

AOI21xp5_ASAP7_75t_L g10519 ( 
.A1(n_10043),
.A2(n_7450),
.B(n_9386),
.Y(n_10519)
);

HB1xp67_ASAP7_75t_L g10520 ( 
.A(n_9481),
.Y(n_10520)
);

OAI22xp5_ASAP7_75t_L g10521 ( 
.A1(n_9495),
.A2(n_8607),
.B1(n_8595),
.B2(n_8445),
.Y(n_10521)
);

INVx1_ASAP7_75t_L g10522 ( 
.A(n_9478),
.Y(n_10522)
);

AOI22xp33_ASAP7_75t_L g10523 ( 
.A1(n_9517),
.A2(n_7662),
.B1(n_7632),
.B2(n_7325),
.Y(n_10523)
);

AND2x2_ASAP7_75t_L g10524 ( 
.A(n_9889),
.B(n_9950),
.Y(n_10524)
);

AOI22xp33_ASAP7_75t_SL g10525 ( 
.A1(n_9838),
.A2(n_8408),
.B1(n_7529),
.B2(n_7688),
.Y(n_10525)
);

OAI221xp5_ASAP7_75t_L g10526 ( 
.A1(n_9438),
.A2(n_9181),
.B1(n_8983),
.B2(n_8974),
.C(n_9173),
.Y(n_10526)
);

NAND2xp5_ASAP7_75t_SL g10527 ( 
.A(n_9445),
.B(n_8408),
.Y(n_10527)
);

AOI22xp33_ASAP7_75t_L g10528 ( 
.A1(n_9838),
.A2(n_7325),
.B1(n_7688),
.B2(n_7588),
.Y(n_10528)
);

BUFx3_ASAP7_75t_L g10529 ( 
.A(n_9656),
.Y(n_10529)
);

OAI22xp5_ASAP7_75t_L g10530 ( 
.A1(n_10278),
.A2(n_8445),
.B1(n_8505),
.B2(n_8481),
.Y(n_10530)
);

NOR2xp33_ASAP7_75t_L g10531 ( 
.A(n_10203),
.B(n_9729),
.Y(n_10531)
);

OAI22xp33_ASAP7_75t_L g10532 ( 
.A1(n_9644),
.A2(n_10229),
.B1(n_10062),
.B2(n_10317),
.Y(n_10532)
);

OAI21x1_ASAP7_75t_L g10533 ( 
.A1(n_10263),
.A2(n_9029),
.B(n_8874),
.Y(n_10533)
);

OAI221xp5_ASAP7_75t_L g10534 ( 
.A1(n_9757),
.A2(n_8839),
.B1(n_8840),
.B2(n_8962),
.C(n_8954),
.Y(n_10534)
);

INVx2_ASAP7_75t_L g10535 ( 
.A(n_9797),
.Y(n_10535)
);

AOI22xp33_ASAP7_75t_L g10536 ( 
.A1(n_9816),
.A2(n_7688),
.B1(n_7588),
.B2(n_8519),
.Y(n_10536)
);

OAI221xp5_ASAP7_75t_L g10537 ( 
.A1(n_9572),
.A2(n_8839),
.B1(n_8840),
.B2(n_8509),
.C(n_8682),
.Y(n_10537)
);

AOI22xp33_ASAP7_75t_L g10538 ( 
.A1(n_9721),
.A2(n_7688),
.B1(n_7588),
.B2(n_8626),
.Y(n_10538)
);

OR2x2_ASAP7_75t_L g10539 ( 
.A(n_9658),
.B(n_7605),
.Y(n_10539)
);

AND2x2_ASAP7_75t_L g10540 ( 
.A(n_9954),
.B(n_8588),
.Y(n_10540)
);

OR2x2_ASAP7_75t_L g10541 ( 
.A(n_9703),
.B(n_7605),
.Y(n_10541)
);

OR2x2_ASAP7_75t_L g10542 ( 
.A(n_9728),
.B(n_7605),
.Y(n_10542)
);

INVx1_ASAP7_75t_SL g10543 ( 
.A(n_9656),
.Y(n_10543)
);

BUFx3_ASAP7_75t_L g10544 ( 
.A(n_10060),
.Y(n_10544)
);

INVx3_ASAP7_75t_L g10545 ( 
.A(n_9752),
.Y(n_10545)
);

BUFx6f_ASAP7_75t_L g10546 ( 
.A(n_9752),
.Y(n_10546)
);

INVx1_ASAP7_75t_L g10547 ( 
.A(n_9485),
.Y(n_10547)
);

AOI22xp33_ASAP7_75t_L g10548 ( 
.A1(n_10207),
.A2(n_7688),
.B1(n_7588),
.B2(n_8650),
.Y(n_10548)
);

AO21x2_ASAP7_75t_L g10549 ( 
.A1(n_9861),
.A2(n_8511),
.B(n_8508),
.Y(n_10549)
);

OAI22xp5_ASAP7_75t_L g10550 ( 
.A1(n_10282),
.A2(n_8445),
.B1(n_8505),
.B2(n_9309),
.Y(n_10550)
);

AO221x1_ASAP7_75t_L g10551 ( 
.A1(n_9567),
.A2(n_8913),
.B1(n_8684),
.B2(n_8695),
.C(n_8671),
.Y(n_10551)
);

OAI22xp33_ASAP7_75t_L g10552 ( 
.A1(n_9644),
.A2(n_7704),
.B1(n_8505),
.B2(n_7461),
.Y(n_10552)
);

INVx2_ASAP7_75t_L g10553 ( 
.A(n_10235),
.Y(n_10553)
);

OAI22xp5_ASAP7_75t_L g10554 ( 
.A1(n_10282),
.A2(n_9117),
.B1(n_9126),
.B2(n_8613),
.Y(n_10554)
);

OAI22xp5_ASAP7_75t_L g10555 ( 
.A1(n_10344),
.A2(n_9623),
.B1(n_9704),
.B2(n_10317),
.Y(n_10555)
);

AND2x4_ASAP7_75t_L g10556 ( 
.A(n_9584),
.B(n_8588),
.Y(n_10556)
);

AOI221xp5_ASAP7_75t_L g10557 ( 
.A1(n_9623),
.A2(n_8565),
.B1(n_8567),
.B2(n_8564),
.C(n_8560),
.Y(n_10557)
);

OAI22xp5_ASAP7_75t_L g10558 ( 
.A1(n_10344),
.A2(n_8613),
.B1(n_9342),
.B2(n_9332),
.Y(n_10558)
);

OAI22xp5_ASAP7_75t_L g10559 ( 
.A1(n_9704),
.A2(n_8613),
.B1(n_9288),
.B2(n_8985),
.Y(n_10559)
);

AND2x2_ASAP7_75t_L g10560 ( 
.A(n_9445),
.B(n_8634),
.Y(n_10560)
);

AOI221xp5_ASAP7_75t_L g10561 ( 
.A1(n_9497),
.A2(n_8565),
.B1(n_8567),
.B2(n_8564),
.C(n_8560),
.Y(n_10561)
);

AOI22xp33_ASAP7_75t_L g10562 ( 
.A1(n_10305),
.A2(n_7688),
.B1(n_8671),
.B2(n_8650),
.Y(n_10562)
);

OAI22xp5_ASAP7_75t_L g10563 ( 
.A1(n_10317),
.A2(n_8721),
.B1(n_8745),
.B2(n_8723),
.Y(n_10563)
);

INVx2_ASAP7_75t_L g10564 ( 
.A(n_10235),
.Y(n_10564)
);

INVx1_ASAP7_75t_L g10565 ( 
.A(n_9490),
.Y(n_10565)
);

AND2x4_ASAP7_75t_L g10566 ( 
.A(n_10313),
.B(n_8634),
.Y(n_10566)
);

OAI221xp5_ASAP7_75t_L g10567 ( 
.A1(n_9497),
.A2(n_8840),
.B1(n_8839),
.B2(n_9265),
.C(n_9264),
.Y(n_10567)
);

OAI22xp5_ASAP7_75t_L g10568 ( 
.A1(n_10317),
.A2(n_8721),
.B1(n_8745),
.B2(n_8723),
.Y(n_10568)
);

AND2x2_ASAP7_75t_L g10569 ( 
.A(n_10289),
.B(n_8634),
.Y(n_10569)
);

HB1xp67_ASAP7_75t_L g10570 ( 
.A(n_9482),
.Y(n_10570)
);

AND2x2_ASAP7_75t_L g10571 ( 
.A(n_10289),
.B(n_8663),
.Y(n_10571)
);

INVx3_ASAP7_75t_L g10572 ( 
.A(n_10362),
.Y(n_10572)
);

AOI22xp33_ASAP7_75t_L g10573 ( 
.A1(n_10341),
.A2(n_8650),
.B1(n_8684),
.B2(n_8671),
.Y(n_10573)
);

INVx1_ASAP7_75t_L g10574 ( 
.A(n_9492),
.Y(n_10574)
);

OAI22xp5_ASAP7_75t_L g10575 ( 
.A1(n_9840),
.A2(n_8745),
.B1(n_8973),
.B2(n_8245),
.Y(n_10575)
);

OA21x2_ASAP7_75t_L g10576 ( 
.A1(n_9557),
.A2(n_8511),
.B(n_8508),
.Y(n_10576)
);

BUFx6f_ASAP7_75t_L g10577 ( 
.A(n_9527),
.Y(n_10577)
);

AND2x4_ASAP7_75t_L g10578 ( 
.A(n_10289),
.B(n_8663),
.Y(n_10578)
);

AOI22xp33_ASAP7_75t_L g10579 ( 
.A1(n_10179),
.A2(n_9795),
.B1(n_10116),
.B2(n_10108),
.Y(n_10579)
);

INVx1_ASAP7_75t_L g10580 ( 
.A(n_9505),
.Y(n_10580)
);

AOI22xp33_ASAP7_75t_L g10581 ( 
.A1(n_10108),
.A2(n_8650),
.B1(n_8684),
.B2(n_8671),
.Y(n_10581)
);

BUFx2_ASAP7_75t_L g10582 ( 
.A(n_10103),
.Y(n_10582)
);

OAI211xp5_ASAP7_75t_L g10583 ( 
.A1(n_9923),
.A2(n_8774),
.B(n_8726),
.C(n_9306),
.Y(n_10583)
);

AOI221xp5_ASAP7_75t_L g10584 ( 
.A1(n_9557),
.A2(n_10226),
.B1(n_10132),
.B2(n_10109),
.C(n_10370),
.Y(n_10584)
);

OAI22xp5_ASAP7_75t_L g10585 ( 
.A1(n_9840),
.A2(n_9756),
.B1(n_9513),
.B2(n_10226),
.Y(n_10585)
);

AOI22xp5_ASAP7_75t_L g10586 ( 
.A1(n_9806),
.A2(n_7715),
.B1(n_9081),
.B2(n_9110),
.Y(n_10586)
);

AOI22xp33_ASAP7_75t_L g10587 ( 
.A1(n_10116),
.A2(n_8684),
.B1(n_8695),
.B2(n_7560),
.Y(n_10587)
);

NAND2xp5_ASAP7_75t_L g10588 ( 
.A(n_9519),
.B(n_7674),
.Y(n_10588)
);

INVx3_ASAP7_75t_L g10589 ( 
.A(n_10362),
.Y(n_10589)
);

OR2x2_ASAP7_75t_L g10590 ( 
.A(n_9618),
.B(n_7783),
.Y(n_10590)
);

OAI22xp5_ASAP7_75t_L g10591 ( 
.A1(n_9513),
.A2(n_8988),
.B1(n_8695),
.B2(n_7721),
.Y(n_10591)
);

OA21x2_ASAP7_75t_L g10592 ( 
.A1(n_10141),
.A2(n_8512),
.B(n_8949),
.Y(n_10592)
);

OAI21xp5_ASAP7_75t_L g10593 ( 
.A1(n_9513),
.A2(n_7444),
.B(n_9364),
.Y(n_10593)
);

INVx2_ASAP7_75t_L g10594 ( 
.A(n_10272),
.Y(n_10594)
);

AOI22xp33_ASAP7_75t_L g10595 ( 
.A1(n_10117),
.A2(n_8695),
.B1(n_7560),
.B2(n_7820),
.Y(n_10595)
);

AOI22xp33_ASAP7_75t_L g10596 ( 
.A1(n_10117),
.A2(n_10136),
.B1(n_10144),
.B2(n_10124),
.Y(n_10596)
);

AOI22xp33_ASAP7_75t_SL g10597 ( 
.A1(n_10164),
.A2(n_8408),
.B1(n_7529),
.B2(n_7549),
.Y(n_10597)
);

AOI22xp33_ASAP7_75t_L g10598 ( 
.A1(n_10124),
.A2(n_7560),
.B1(n_7820),
.B2(n_7529),
.Y(n_10598)
);

OA21x2_ASAP7_75t_L g10599 ( 
.A1(n_10141),
.A2(n_8512),
.B(n_8949),
.Y(n_10599)
);

OAI211xp5_ASAP7_75t_L g10600 ( 
.A1(n_10027),
.A2(n_8774),
.B(n_8726),
.C(n_7247),
.Y(n_10600)
);

AOI221xp5_ASAP7_75t_L g10601 ( 
.A1(n_10109),
.A2(n_8579),
.B1(n_8580),
.B2(n_8578),
.C(n_8571),
.Y(n_10601)
);

OAI22xp33_ASAP7_75t_L g10602 ( 
.A1(n_10062),
.A2(n_8086),
.B1(n_8016),
.B2(n_8166),
.Y(n_10602)
);

INVx2_ASAP7_75t_L g10603 ( 
.A(n_10272),
.Y(n_10603)
);

OAI22xp5_ASAP7_75t_L g10604 ( 
.A1(n_9513),
.A2(n_7721),
.B1(n_7782),
.B2(n_7781),
.Y(n_10604)
);

AOI221xp5_ASAP7_75t_L g10605 ( 
.A1(n_10132),
.A2(n_10392),
.B1(n_10057),
.B2(n_10287),
.C(n_10136),
.Y(n_10605)
);

AOI22xp33_ASAP7_75t_L g10606 ( 
.A1(n_10144),
.A2(n_10156),
.B1(n_10161),
.B2(n_10147),
.Y(n_10606)
);

O2A1O1Ixp33_ASAP7_75t_L g10607 ( 
.A1(n_9441),
.A2(n_8913),
.B(n_9221),
.C(n_9192),
.Y(n_10607)
);

INVx1_ASAP7_75t_L g10608 ( 
.A(n_9506),
.Y(n_10608)
);

OAI22xp5_ASAP7_75t_L g10609 ( 
.A1(n_9498),
.A2(n_7721),
.B1(n_7782),
.B2(n_7781),
.Y(n_10609)
);

INVx1_ASAP7_75t_L g10610 ( 
.A(n_9511),
.Y(n_10610)
);

OAI22xp5_ASAP7_75t_L g10611 ( 
.A1(n_9498),
.A2(n_7782),
.B1(n_7821),
.B2(n_7781),
.Y(n_10611)
);

BUFx12f_ASAP7_75t_L g10612 ( 
.A(n_9543),
.Y(n_10612)
);

NAND2xp5_ASAP7_75t_L g10613 ( 
.A(n_10157),
.B(n_7674),
.Y(n_10613)
);

AOI22xp33_ASAP7_75t_L g10614 ( 
.A1(n_10147),
.A2(n_7560),
.B1(n_7529),
.B2(n_8408),
.Y(n_10614)
);

AOI21xp33_ASAP7_75t_SL g10615 ( 
.A1(n_9903),
.A2(n_8545),
.B(n_9177),
.Y(n_10615)
);

INVx1_ASAP7_75t_L g10616 ( 
.A(n_9512),
.Y(n_10616)
);

OAI221xp5_ASAP7_75t_L g10617 ( 
.A1(n_9441),
.A2(n_9266),
.B1(n_9270),
.B2(n_9265),
.C(n_9264),
.Y(n_10617)
);

AND2x2_ASAP7_75t_L g10618 ( 
.A(n_10396),
.B(n_8663),
.Y(n_10618)
);

AOI22xp33_ASAP7_75t_L g10619 ( 
.A1(n_10156),
.A2(n_7560),
.B1(n_7529),
.B2(n_8408),
.Y(n_10619)
);

OAI321xp33_ASAP7_75t_L g10620 ( 
.A1(n_10062),
.A2(n_7591),
.A3(n_7757),
.B1(n_8143),
.B2(n_8391),
.C(n_8374),
.Y(n_10620)
);

AOI222xp33_ASAP7_75t_L g10621 ( 
.A1(n_10161),
.A2(n_9275),
.B1(n_9270),
.B2(n_9276),
.C1(n_9266),
.C2(n_8260),
.Y(n_10621)
);

OAI22xp5_ASAP7_75t_L g10622 ( 
.A1(n_9498),
.A2(n_7821),
.B1(n_7897),
.B2(n_8392),
.Y(n_10622)
);

AOI222xp33_ASAP7_75t_L g10623 ( 
.A1(n_10169),
.A2(n_9276),
.B1(n_9275),
.B2(n_8853),
.C1(n_8752),
.C2(n_8854),
.Y(n_10623)
);

AOI21xp33_ASAP7_75t_SL g10624 ( 
.A1(n_10127),
.A2(n_8545),
.B(n_9045),
.Y(n_10624)
);

AND2x2_ASAP7_75t_L g10625 ( 
.A(n_10396),
.B(n_8685),
.Y(n_10625)
);

AOI21xp5_ASAP7_75t_L g10626 ( 
.A1(n_9688),
.A2(n_9845),
.B(n_10194),
.Y(n_10626)
);

OR2x6_ASAP7_75t_L g10627 ( 
.A(n_9946),
.B(n_8867),
.Y(n_10627)
);

BUFx10_ASAP7_75t_L g10628 ( 
.A(n_9946),
.Y(n_10628)
);

OAI211xp5_ASAP7_75t_L g10629 ( 
.A1(n_9854),
.A2(n_9688),
.B(n_9465),
.C(n_10164),
.Y(n_10629)
);

INVx2_ASAP7_75t_L g10630 ( 
.A(n_10301),
.Y(n_10630)
);

OR2x2_ASAP7_75t_L g10631 ( 
.A(n_9581),
.B(n_7783),
.Y(n_10631)
);

INVx1_ASAP7_75t_L g10632 ( 
.A(n_9514),
.Y(n_10632)
);

O2A1O1Ixp33_ASAP7_75t_L g10633 ( 
.A1(n_9441),
.A2(n_7960),
.B(n_7952),
.C(n_8143),
.Y(n_10633)
);

AOI22xp5_ASAP7_75t_L g10634 ( 
.A1(n_9502),
.A2(n_8536),
.B1(n_8086),
.B2(n_8016),
.Y(n_10634)
);

AOI22xp33_ASAP7_75t_SL g10635 ( 
.A1(n_9502),
.A2(n_8408),
.B1(n_7529),
.B2(n_7549),
.Y(n_10635)
);

INVx2_ASAP7_75t_L g10636 ( 
.A(n_10301),
.Y(n_10636)
);

AOI222xp33_ASAP7_75t_L g10637 ( 
.A1(n_10169),
.A2(n_8853),
.B1(n_8752),
.B2(n_8854),
.C1(n_8759),
.C2(n_8750),
.Y(n_10637)
);

CKINVDCx11_ASAP7_75t_R g10638 ( 
.A(n_9543),
.Y(n_10638)
);

INVx3_ASAP7_75t_SL g10639 ( 
.A(n_9444),
.Y(n_10639)
);

OAI21x1_ASAP7_75t_L g10640 ( 
.A1(n_10045),
.A2(n_9029),
.B(n_9046),
.Y(n_10640)
);

HB1xp67_ASAP7_75t_L g10641 ( 
.A(n_9573),
.Y(n_10641)
);

BUFx2_ASAP7_75t_L g10642 ( 
.A(n_10103),
.Y(n_10642)
);

BUFx6f_ASAP7_75t_SL g10643 ( 
.A(n_9487),
.Y(n_10643)
);

BUFx3_ASAP7_75t_L g10644 ( 
.A(n_10060),
.Y(n_10644)
);

AOI222xp33_ASAP7_75t_L g10645 ( 
.A1(n_10172),
.A2(n_8883),
.B1(n_8759),
.B2(n_8887),
.C1(n_8856),
.C2(n_8750),
.Y(n_10645)
);

AO31x2_ASAP7_75t_L g10646 ( 
.A1(n_9861),
.A2(n_8975),
.A3(n_9004),
.B(n_8955),
.Y(n_10646)
);

INVx2_ASAP7_75t_L g10647 ( 
.A(n_10366),
.Y(n_10647)
);

AOI22xp33_ASAP7_75t_L g10648 ( 
.A1(n_10172),
.A2(n_8408),
.B1(n_8013),
.B2(n_7168),
.Y(n_10648)
);

INVx3_ASAP7_75t_L g10649 ( 
.A(n_10131),
.Y(n_10649)
);

AND2x2_ASAP7_75t_L g10650 ( 
.A(n_10396),
.B(n_8685),
.Y(n_10650)
);

OAI21x1_ASAP7_75t_L g10651 ( 
.A1(n_9716),
.A2(n_9213),
.B(n_9046),
.Y(n_10651)
);

OAI22xp5_ASAP7_75t_SL g10652 ( 
.A1(n_10367),
.A2(n_6647),
.B1(n_6649),
.B2(n_6637),
.Y(n_10652)
);

INVxp67_ASAP7_75t_L g10653 ( 
.A(n_9810),
.Y(n_10653)
);

AOI21xp5_ASAP7_75t_L g10654 ( 
.A1(n_10194),
.A2(n_8103),
.B(n_8115),
.Y(n_10654)
);

INVx4_ASAP7_75t_L g10655 ( 
.A(n_9592),
.Y(n_10655)
);

AOI21xp5_ASAP7_75t_L g10656 ( 
.A1(n_10256),
.A2(n_8103),
.B(n_8115),
.Y(n_10656)
);

AOI22xp33_ASAP7_75t_L g10657 ( 
.A1(n_10176),
.A2(n_8408),
.B1(n_8013),
.B2(n_7168),
.Y(n_10657)
);

OA21x2_ASAP7_75t_L g10658 ( 
.A1(n_9865),
.A2(n_8975),
.B(n_8955),
.Y(n_10658)
);

OR2x6_ASAP7_75t_L g10659 ( 
.A(n_9946),
.B(n_8867),
.Y(n_10659)
);

OAI21x1_ASAP7_75t_L g10660 ( 
.A1(n_9749),
.A2(n_9213),
.B(n_9347),
.Y(n_10660)
);

OAI21x1_ASAP7_75t_L g10661 ( 
.A1(n_10034),
.A2(n_9347),
.B(n_8714),
.Y(n_10661)
);

AND2x2_ASAP7_75t_L g10662 ( 
.A(n_9718),
.B(n_8685),
.Y(n_10662)
);

NAND2xp5_ASAP7_75t_L g10663 ( 
.A(n_9539),
.B(n_7674),
.Y(n_10663)
);

NAND2xp5_ASAP7_75t_L g10664 ( 
.A(n_9549),
.B(n_7674),
.Y(n_10664)
);

INVx2_ASAP7_75t_L g10665 ( 
.A(n_10366),
.Y(n_10665)
);

AOI322xp5_ASAP7_75t_L g10666 ( 
.A1(n_9718),
.A2(n_9733),
.A3(n_9540),
.B1(n_10176),
.B2(n_9582),
.C1(n_9502),
.C2(n_9871),
.Y(n_10666)
);

OAI22xp33_ASAP7_75t_L g10667 ( 
.A1(n_10062),
.A2(n_8166),
.B1(n_8391),
.B2(n_8374),
.Y(n_10667)
);

AND2x2_ASAP7_75t_L g10668 ( 
.A(n_9733),
.B(n_8706),
.Y(n_10668)
);

AOI22xp33_ASAP7_75t_L g10669 ( 
.A1(n_9594),
.A2(n_8408),
.B1(n_8013),
.B2(n_7168),
.Y(n_10669)
);

INVx2_ASAP7_75t_L g10670 ( 
.A(n_10383),
.Y(n_10670)
);

INVx1_ASAP7_75t_L g10671 ( 
.A(n_9515),
.Y(n_10671)
);

NAND2xp5_ASAP7_75t_L g10672 ( 
.A(n_9605),
.B(n_7674),
.Y(n_10672)
);

INVx2_ASAP7_75t_L g10673 ( 
.A(n_10383),
.Y(n_10673)
);

OAI22xp33_ASAP7_75t_L g10674 ( 
.A1(n_10229),
.A2(n_8391),
.B1(n_8374),
.B2(n_7765),
.Y(n_10674)
);

AOI22xp33_ASAP7_75t_L g10675 ( 
.A1(n_9594),
.A2(n_8013),
.B1(n_7168),
.B2(n_8654),
.Y(n_10675)
);

OAI221xp5_ASAP7_75t_SL g10676 ( 
.A1(n_9441),
.A2(n_7580),
.B1(n_8578),
.B2(n_8579),
.C(n_8571),
.Y(n_10676)
);

OA21x2_ASAP7_75t_L g10677 ( 
.A1(n_9865),
.A2(n_9015),
.B(n_9004),
.Y(n_10677)
);

OAI21xp5_ASAP7_75t_L g10678 ( 
.A1(n_9707),
.A2(n_9368),
.B(n_9364),
.Y(n_10678)
);

INVx1_ASAP7_75t_L g10679 ( 
.A(n_9516),
.Y(n_10679)
);

AOI22xp33_ASAP7_75t_L g10680 ( 
.A1(n_9649),
.A2(n_8013),
.B1(n_7309),
.B2(n_7616),
.Y(n_10680)
);

OAI22xp5_ASAP7_75t_L g10681 ( 
.A1(n_9582),
.A2(n_7821),
.B1(n_7897),
.B2(n_8392),
.Y(n_10681)
);

AOI21xp33_ASAP7_75t_L g10682 ( 
.A1(n_9458),
.A2(n_9582),
.B(n_9803),
.Y(n_10682)
);

AOI222xp33_ASAP7_75t_L g10683 ( 
.A1(n_10120),
.A2(n_8896),
.B1(n_8883),
.B2(n_8917),
.C1(n_8887),
.C2(n_8856),
.Y(n_10683)
);

AO21x2_ASAP7_75t_L g10684 ( 
.A1(n_9871),
.A2(n_8892),
.B(n_8888),
.Y(n_10684)
);

OAI22xp5_ASAP7_75t_L g10685 ( 
.A1(n_10256),
.A2(n_7897),
.B1(n_8492),
.B2(n_8435),
.Y(n_10685)
);

AND2x2_ASAP7_75t_L g10686 ( 
.A(n_10133),
.B(n_8706),
.Y(n_10686)
);

CKINVDCx5p33_ASAP7_75t_R g10687 ( 
.A(n_9444),
.Y(n_10687)
);

AOI22xp33_ASAP7_75t_SL g10688 ( 
.A1(n_9509),
.A2(n_7549),
.B1(n_8360),
.B2(n_8359),
.Y(n_10688)
);

OAI22xp5_ASAP7_75t_L g10689 ( 
.A1(n_10229),
.A2(n_8435),
.B1(n_8699),
.B2(n_8492),
.Y(n_10689)
);

AOI22xp33_ASAP7_75t_L g10690 ( 
.A1(n_9649),
.A2(n_8013),
.B1(n_7309),
.B2(n_8543),
.Y(n_10690)
);

AND2x2_ASAP7_75t_L g10691 ( 
.A(n_10133),
.B(n_8706),
.Y(n_10691)
);

HB1xp67_ASAP7_75t_L g10692 ( 
.A(n_9668),
.Y(n_10692)
);

AOI22xp33_ASAP7_75t_L g10693 ( 
.A1(n_9509),
.A2(n_7309),
.B1(n_8577),
.B2(n_7247),
.Y(n_10693)
);

CKINVDCx5p33_ASAP7_75t_R g10694 ( 
.A(n_10012),
.Y(n_10694)
);

AND2x2_ASAP7_75t_L g10695 ( 
.A(n_10142),
.B(n_8802),
.Y(n_10695)
);

A2O1A1Ixp33_ASAP7_75t_L g10696 ( 
.A1(n_9707),
.A2(n_7580),
.B(n_9368),
.C(n_8308),
.Y(n_10696)
);

AOI22xp33_ASAP7_75t_L g10697 ( 
.A1(n_9673),
.A2(n_7309),
.B1(n_7247),
.B2(n_7792),
.Y(n_10697)
);

AOI221xp5_ASAP7_75t_L g10698 ( 
.A1(n_9672),
.A2(n_9542),
.B1(n_9727),
.B2(n_9738),
.C(n_9736),
.Y(n_10698)
);

OAI22xp33_ASAP7_75t_L g10699 ( 
.A1(n_10229),
.A2(n_7765),
.B1(n_8014),
.B2(n_7686),
.Y(n_10699)
);

INVx1_ASAP7_75t_L g10700 ( 
.A(n_9521),
.Y(n_10700)
);

AOI21xp5_ASAP7_75t_L g10701 ( 
.A1(n_10232),
.A2(n_9907),
.B(n_10339),
.Y(n_10701)
);

AO21x2_ASAP7_75t_L g10702 ( 
.A1(n_10219),
.A2(n_10320),
.B(n_10085),
.Y(n_10702)
);

OAI22xp5_ASAP7_75t_L g10703 ( 
.A1(n_10309),
.A2(n_8435),
.B1(n_8699),
.B2(n_8492),
.Y(n_10703)
);

INVx1_ASAP7_75t_L g10704 ( 
.A(n_9523),
.Y(n_10704)
);

AOI22xp33_ASAP7_75t_L g10705 ( 
.A1(n_9673),
.A2(n_7309),
.B1(n_7792),
.B2(n_7544),
.Y(n_10705)
);

AOI22xp33_ASAP7_75t_L g10706 ( 
.A1(n_10261),
.A2(n_7544),
.B1(n_7844),
.B2(n_7215),
.Y(n_10706)
);

AOI22xp33_ASAP7_75t_L g10707 ( 
.A1(n_10261),
.A2(n_7544),
.B1(n_7844),
.B2(n_7215),
.Y(n_10707)
);

AOI21xp5_ASAP7_75t_L g10708 ( 
.A1(n_9907),
.A2(n_9272),
.B(n_9367),
.Y(n_10708)
);

AO21x1_ASAP7_75t_L g10709 ( 
.A1(n_9785),
.A2(n_8582),
.B(n_8580),
.Y(n_10709)
);

AOI21xp33_ASAP7_75t_L g10710 ( 
.A1(n_9803),
.A2(n_8892),
.B(n_8888),
.Y(n_10710)
);

AOI22xp5_ASAP7_75t_L g10711 ( 
.A1(n_9672),
.A2(n_9053),
.B1(n_7757),
.B2(n_8568),
.Y(n_10711)
);

OAI221xp5_ASAP7_75t_L g10712 ( 
.A1(n_9938),
.A2(n_8322),
.B1(n_8323),
.B2(n_8308),
.C(n_8305),
.Y(n_10712)
);

AOI22xp33_ASAP7_75t_L g10713 ( 
.A1(n_10261),
.A2(n_7544),
.B1(n_7215),
.B2(n_8651),
.Y(n_10713)
);

AND2x2_ASAP7_75t_L g10714 ( 
.A(n_10142),
.B(n_8802),
.Y(n_10714)
);

AOI22xp33_ASAP7_75t_SL g10715 ( 
.A1(n_9542),
.A2(n_7549),
.B1(n_8360),
.B2(n_8359),
.Y(n_10715)
);

AND2x2_ASAP7_75t_L g10716 ( 
.A(n_9993),
.B(n_8802),
.Y(n_10716)
);

BUFx2_ASAP7_75t_L g10717 ( 
.A(n_10131),
.Y(n_10717)
);

AND2x2_ASAP7_75t_L g10718 ( 
.A(n_9995),
.B(n_8843),
.Y(n_10718)
);

INVx2_ASAP7_75t_L g10719 ( 
.A(n_10394),
.Y(n_10719)
);

NOR2xp67_ASAP7_75t_L g10720 ( 
.A(n_9487),
.B(n_8726),
.Y(n_10720)
);

INVx3_ASAP7_75t_L g10721 ( 
.A(n_10166),
.Y(n_10721)
);

INVx2_ASAP7_75t_L g10722 ( 
.A(n_10394),
.Y(n_10722)
);

AND2x2_ASAP7_75t_L g10723 ( 
.A(n_10010),
.B(n_8843),
.Y(n_10723)
);

OAI22xp5_ASAP7_75t_L g10724 ( 
.A1(n_9785),
.A2(n_8435),
.B1(n_8699),
.B2(n_8492),
.Y(n_10724)
);

AOI222xp33_ASAP7_75t_L g10725 ( 
.A1(n_9873),
.A2(n_8917),
.B1(n_8896),
.B2(n_8592),
.C1(n_8590),
.C2(n_8610),
.Y(n_10725)
);

AOI22xp33_ASAP7_75t_L g10726 ( 
.A1(n_9966),
.A2(n_7544),
.B1(n_7215),
.B2(n_7806),
.Y(n_10726)
);

AOI22xp33_ASAP7_75t_L g10727 ( 
.A1(n_10252),
.A2(n_7215),
.B1(n_7817),
.B2(n_7806),
.Y(n_10727)
);

OAI22xp5_ASAP7_75t_L g10728 ( 
.A1(n_9785),
.A2(n_8699),
.B1(n_8783),
.B2(n_8719),
.Y(n_10728)
);

AOI221xp5_ASAP7_75t_L g10729 ( 
.A1(n_9727),
.A2(n_8591),
.B1(n_8592),
.B2(n_8590),
.C(n_8582),
.Y(n_10729)
);

INVx1_ASAP7_75t_L g10730 ( 
.A(n_9524),
.Y(n_10730)
);

AND2x2_ASAP7_75t_L g10731 ( 
.A(n_10026),
.B(n_8843),
.Y(n_10731)
);

BUFx6f_ASAP7_75t_L g10732 ( 
.A(n_9527),
.Y(n_10732)
);

AND2x2_ASAP7_75t_L g10733 ( 
.A(n_10031),
.B(n_8884),
.Y(n_10733)
);

NOR2xp67_ASAP7_75t_L g10734 ( 
.A(n_9487),
.B(n_9048),
.Y(n_10734)
);

INVx1_ASAP7_75t_L g10735 ( 
.A(n_9526),
.Y(n_10735)
);

INVx1_ASAP7_75t_L g10736 ( 
.A(n_9531),
.Y(n_10736)
);

AOI221xp5_ASAP7_75t_L g10737 ( 
.A1(n_9736),
.A2(n_9738),
.B1(n_9743),
.B2(n_10407),
.C(n_10404),
.Y(n_10737)
);

INVx2_ASAP7_75t_L g10738 ( 
.A(n_10395),
.Y(n_10738)
);

BUFx3_ASAP7_75t_L g10739 ( 
.A(n_10063),
.Y(n_10739)
);

AOI221xp5_ASAP7_75t_L g10740 ( 
.A1(n_9743),
.A2(n_8614),
.B1(n_8620),
.B2(n_8610),
.C(n_8591),
.Y(n_10740)
);

INVx1_ASAP7_75t_L g10741 ( 
.A(n_9532),
.Y(n_10741)
);

OAI211xp5_ASAP7_75t_SL g10742 ( 
.A1(n_10369),
.A2(n_9216),
.B(n_9189),
.C(n_9418),
.Y(n_10742)
);

NAND2xp5_ASAP7_75t_L g10743 ( 
.A(n_9615),
.B(n_7674),
.Y(n_10743)
);

AOI22xp33_ASAP7_75t_L g10744 ( 
.A1(n_9580),
.A2(n_7817),
.B1(n_7867),
.B2(n_7845),
.Y(n_10744)
);

AOI22xp33_ASAP7_75t_L g10745 ( 
.A1(n_9580),
.A2(n_7845),
.B1(n_7867),
.B2(n_7971),
.Y(n_10745)
);

O2A1O1Ixp33_ASAP7_75t_L g10746 ( 
.A1(n_9763),
.A2(n_7952),
.B(n_7960),
.C(n_8614),
.Y(n_10746)
);

AO222x2_ASAP7_75t_L g10747 ( 
.A1(n_9553),
.A2(n_7180),
.B1(n_7203),
.B2(n_7291),
.C1(n_8868),
.C2(n_7683),
.Y(n_10747)
);

AND2x2_ASAP7_75t_L g10748 ( 
.A(n_10054),
.B(n_8884),
.Y(n_10748)
);

OAI211xp5_ASAP7_75t_L g10749 ( 
.A1(n_9465),
.A2(n_8401),
.B(n_8446),
.C(n_8411),
.Y(n_10749)
);

AOI221xp5_ASAP7_75t_L g10750 ( 
.A1(n_10404),
.A2(n_8641),
.B1(n_8647),
.B2(n_8625),
.C(n_8620),
.Y(n_10750)
);

NOR2xp67_ASAP7_75t_L g10751 ( 
.A(n_9489),
.B(n_9048),
.Y(n_10751)
);

AOI21xp5_ASAP7_75t_L g10752 ( 
.A1(n_10339),
.A2(n_8226),
.B(n_7921),
.Y(n_10752)
);

OAI21xp33_ASAP7_75t_L g10753 ( 
.A1(n_10411),
.A2(n_9419),
.B(n_9416),
.Y(n_10753)
);

AOI22xp5_ASAP7_75t_L g10754 ( 
.A1(n_9849),
.A2(n_8568),
.B1(n_8186),
.B2(n_9405),
.Y(n_10754)
);

AOI22xp5_ASAP7_75t_L g10755 ( 
.A1(n_9849),
.A2(n_8568),
.B1(n_8186),
.B2(n_7845),
.Y(n_10755)
);

OAI22xp33_ASAP7_75t_L g10756 ( 
.A1(n_9616),
.A2(n_7765),
.B1(n_8014),
.B2(n_7686),
.Y(n_10756)
);

AOI221xp5_ASAP7_75t_L g10757 ( 
.A1(n_10404),
.A2(n_8647),
.B1(n_8653),
.B2(n_8641),
.C(n_8625),
.Y(n_10757)
);

AOI222xp33_ASAP7_75t_L g10758 ( 
.A1(n_10082),
.A2(n_8698),
.B1(n_8666),
.B2(n_8716),
.C1(n_8688),
.C2(n_8653),
.Y(n_10758)
);

OAI22xp33_ASAP7_75t_L g10759 ( 
.A1(n_9616),
.A2(n_7765),
.B1(n_8014),
.B2(n_7686),
.Y(n_10759)
);

AOI221xp5_ASAP7_75t_L g10760 ( 
.A1(n_10407),
.A2(n_8698),
.B1(n_8716),
.B2(n_8688),
.C(n_8666),
.Y(n_10760)
);

OA21x2_ASAP7_75t_L g10761 ( 
.A1(n_9971),
.A2(n_9976),
.B(n_9975),
.Y(n_10761)
);

AOI221xp5_ASAP7_75t_L g10762 ( 
.A1(n_10407),
.A2(n_8728),
.B1(n_8729),
.B2(n_8727),
.C(n_8724),
.Y(n_10762)
);

AOI22xp33_ASAP7_75t_L g10763 ( 
.A1(n_9796),
.A2(n_7845),
.B1(n_7867),
.B2(n_7971),
.Y(n_10763)
);

OA21x2_ASAP7_75t_L g10764 ( 
.A1(n_9971),
.A2(n_9034),
.B(n_9015),
.Y(n_10764)
);

OAI22xp5_ASAP7_75t_L g10765 ( 
.A1(n_9748),
.A2(n_8783),
.B1(n_8906),
.B2(n_8719),
.Y(n_10765)
);

INVx3_ASAP7_75t_L g10766 ( 
.A(n_10166),
.Y(n_10766)
);

AOI22xp33_ASAP7_75t_L g10767 ( 
.A1(n_9796),
.A2(n_7867),
.B1(n_9035),
.B2(n_9034),
.Y(n_10767)
);

AOI22xp33_ASAP7_75t_SL g10768 ( 
.A1(n_9763),
.A2(n_7549),
.B1(n_8360),
.B2(n_8359),
.Y(n_10768)
);

AO21x2_ASAP7_75t_L g10769 ( 
.A1(n_10082),
.A2(n_10099),
.B(n_10085),
.Y(n_10769)
);

INVx3_ASAP7_75t_L g10770 ( 
.A(n_10265),
.Y(n_10770)
);

AOI22xp33_ASAP7_75t_L g10771 ( 
.A1(n_9437),
.A2(n_7867),
.B1(n_9036),
.B2(n_9035),
.Y(n_10771)
);

AOI22xp33_ASAP7_75t_L g10772 ( 
.A1(n_9437),
.A2(n_9036),
.B1(n_9066),
.B2(n_9049),
.Y(n_10772)
);

AOI21xp5_ASAP7_75t_L g10773 ( 
.A1(n_9735),
.A2(n_8226),
.B(n_7921),
.Y(n_10773)
);

A2O1A1Ixp33_ASAP7_75t_L g10774 ( 
.A1(n_9724),
.A2(n_8322),
.B(n_8323),
.C(n_8305),
.Y(n_10774)
);

INVx1_ASAP7_75t_L g10775 ( 
.A(n_9533),
.Y(n_10775)
);

AOI22xp33_ASAP7_75t_SL g10776 ( 
.A1(n_9763),
.A2(n_7549),
.B1(n_8378),
.B2(n_8368),
.Y(n_10776)
);

OAI22xp5_ASAP7_75t_L g10777 ( 
.A1(n_9969),
.A2(n_8783),
.B1(n_8906),
.B2(n_8719),
.Y(n_10777)
);

AOI22xp33_ASAP7_75t_L g10778 ( 
.A1(n_9440),
.A2(n_9049),
.B1(n_9066),
.B2(n_7630),
.Y(n_10778)
);

OR2x2_ASAP7_75t_L g10779 ( 
.A(n_9604),
.B(n_7848),
.Y(n_10779)
);

CKINVDCx8_ASAP7_75t_R g10780 ( 
.A(n_10012),
.Y(n_10780)
);

OAI211xp5_ASAP7_75t_L g10781 ( 
.A1(n_9647),
.A2(n_8401),
.B(n_8446),
.C(n_8411),
.Y(n_10781)
);

NAND3xp33_ASAP7_75t_L g10782 ( 
.A(n_10384),
.B(n_7279),
.C(n_9077),
.Y(n_10782)
);

AND2x2_ASAP7_75t_L g10783 ( 
.A(n_10159),
.B(n_10170),
.Y(n_10783)
);

CKINVDCx5p33_ASAP7_75t_R g10784 ( 
.A(n_9647),
.Y(n_10784)
);

AOI211xp5_ASAP7_75t_L g10785 ( 
.A1(n_9724),
.A2(n_7779),
.B(n_7275),
.C(n_8227),
.Y(n_10785)
);

AOI22xp33_ASAP7_75t_L g10786 ( 
.A1(n_9440),
.A2(n_7630),
.B1(n_8294),
.B2(n_8278),
.Y(n_10786)
);

BUFx6f_ASAP7_75t_L g10787 ( 
.A(n_9538),
.Y(n_10787)
);

INVxp67_ASAP7_75t_L g10788 ( 
.A(n_9810),
.Y(n_10788)
);

AOI22xp33_ASAP7_75t_L g10789 ( 
.A1(n_9452),
.A2(n_8294),
.B1(n_8278),
.B2(n_8014),
.Y(n_10789)
);

INVx2_ASAP7_75t_SL g10790 ( 
.A(n_9902),
.Y(n_10790)
);

NAND2xp5_ASAP7_75t_L g10791 ( 
.A(n_9638),
.B(n_7674),
.Y(n_10791)
);

INVx1_ASAP7_75t_L g10792 ( 
.A(n_9535),
.Y(n_10792)
);

AOI21xp33_ASAP7_75t_L g10793 ( 
.A1(n_9732),
.A2(n_8892),
.B(n_8888),
.Y(n_10793)
);

AOI21xp5_ASAP7_75t_L g10794 ( 
.A1(n_9735),
.A2(n_7933),
.B(n_7848),
.Y(n_10794)
);

OAI221xp5_ASAP7_75t_L g10795 ( 
.A1(n_9984),
.A2(n_9989),
.B1(n_9768),
.B2(n_9953),
.C(n_9941),
.Y(n_10795)
);

NOR2xp33_ASAP7_75t_L g10796 ( 
.A(n_9814),
.B(n_8808),
.Y(n_10796)
);

OAI22xp5_ASAP7_75t_L g10797 ( 
.A1(n_9978),
.A2(n_8783),
.B1(n_8906),
.B2(n_8719),
.Y(n_10797)
);

OR2x6_ASAP7_75t_L g10798 ( 
.A(n_9489),
.B(n_8884),
.Y(n_10798)
);

AND2x2_ASAP7_75t_L g10799 ( 
.A(n_10190),
.B(n_8895),
.Y(n_10799)
);

NAND2xp5_ASAP7_75t_L g10800 ( 
.A(n_9815),
.B(n_7683),
.Y(n_10800)
);

OR2x6_ASAP7_75t_L g10801 ( 
.A(n_9489),
.B(n_8895),
.Y(n_10801)
);

AND2x2_ASAP7_75t_L g10802 ( 
.A(n_10234),
.B(n_8895),
.Y(n_10802)
);

NAND2x1_ASAP7_75t_L g10803 ( 
.A(n_9792),
.B(n_8733),
.Y(n_10803)
);

OAI211xp5_ASAP7_75t_SL g10804 ( 
.A1(n_10046),
.A2(n_9420),
.B(n_8831),
.C(n_8890),
.Y(n_10804)
);

INVx1_ASAP7_75t_L g10805 ( 
.A(n_9541),
.Y(n_10805)
);

OAI211xp5_ASAP7_75t_SL g10806 ( 
.A1(n_10292),
.A2(n_9020),
.B(n_8811),
.C(n_7251),
.Y(n_10806)
);

AND2x4_ASAP7_75t_L g10807 ( 
.A(n_10127),
.B(n_8384),
.Y(n_10807)
);

CKINVDCx20_ASAP7_75t_R g10808 ( 
.A(n_10063),
.Y(n_10808)
);

NOR2xp33_ASAP7_75t_L g10809 ( 
.A(n_9863),
.B(n_8397),
.Y(n_10809)
);

OAI22xp5_ASAP7_75t_L g10810 ( 
.A1(n_9676),
.A2(n_8938),
.B1(n_8906),
.B2(n_9108),
.Y(n_10810)
);

BUFx12f_ASAP7_75t_L g10811 ( 
.A(n_9499),
.Y(n_10811)
);

NOR2xp33_ASAP7_75t_L g10812 ( 
.A(n_9919),
.B(n_8397),
.Y(n_10812)
);

OAI22xp5_ASAP7_75t_L g10813 ( 
.A1(n_9676),
.A2(n_8938),
.B1(n_8104),
.B2(n_8109),
.Y(n_10813)
);

CKINVDCx5p33_ASAP7_75t_R g10814 ( 
.A(n_9880),
.Y(n_10814)
);

INVx2_ASAP7_75t_SL g10815 ( 
.A(n_9902),
.Y(n_10815)
);

AOI21xp5_ASAP7_75t_L g10816 ( 
.A1(n_9735),
.A2(n_7937),
.B(n_7933),
.Y(n_10816)
);

OAI22xp33_ASAP7_75t_L g10817 ( 
.A1(n_9616),
.A2(n_9850),
.B1(n_9982),
.B2(n_9761),
.Y(n_10817)
);

A2O1A1Ixp33_ASAP7_75t_L g10818 ( 
.A1(n_9768),
.A2(n_9827),
.B(n_9953),
.C(n_9941),
.Y(n_10818)
);

INVx1_ASAP7_75t_L g10819 ( 
.A(n_9545),
.Y(n_10819)
);

AOI22xp33_ASAP7_75t_L g10820 ( 
.A1(n_9452),
.A2(n_8014),
.B1(n_7765),
.B2(n_8368),
.Y(n_10820)
);

AOI221xp5_ASAP7_75t_L g10821 ( 
.A1(n_9768),
.A2(n_8728),
.B1(n_8729),
.B2(n_8727),
.C(n_8724),
.Y(n_10821)
);

OAI22xp5_ASAP7_75t_L g10822 ( 
.A1(n_9682),
.A2(n_8938),
.B1(n_8104),
.B2(n_8109),
.Y(n_10822)
);

OR2x6_ASAP7_75t_L g10823 ( 
.A(n_9499),
.B(n_6637),
.Y(n_10823)
);

AOI22xp33_ASAP7_75t_L g10824 ( 
.A1(n_9454),
.A2(n_8014),
.B1(n_7765),
.B2(n_8368),
.Y(n_10824)
);

A2O1A1Ixp33_ASAP7_75t_L g10825 ( 
.A1(n_9827),
.A2(n_8323),
.B(n_8333),
.C(n_8322),
.Y(n_10825)
);

INVx1_ASAP7_75t_L g10826 ( 
.A(n_9547),
.Y(n_10826)
);

AND2x2_ASAP7_75t_L g10827 ( 
.A(n_10296),
.B(n_9355),
.Y(n_10827)
);

AOI22xp33_ASAP7_75t_L g10828 ( 
.A1(n_9454),
.A2(n_8014),
.B1(n_7765),
.B2(n_8378),
.Y(n_10828)
);

OAI22xp5_ASAP7_75t_L g10829 ( 
.A1(n_9682),
.A2(n_8938),
.B1(n_8213),
.B2(n_9113),
.Y(n_10829)
);

AND2x2_ASAP7_75t_L g10830 ( 
.A(n_10298),
.B(n_9355),
.Y(n_10830)
);

AND2x2_ASAP7_75t_L g10831 ( 
.A(n_10327),
.B(n_9355),
.Y(n_10831)
);

AND2x2_ASAP7_75t_L g10832 ( 
.A(n_10180),
.B(n_9355),
.Y(n_10832)
);

AOI22xp33_ASAP7_75t_L g10833 ( 
.A1(n_9461),
.A2(n_8014),
.B1(n_7765),
.B2(n_8378),
.Y(n_10833)
);

AOI21xp33_ASAP7_75t_L g10834 ( 
.A1(n_9732),
.A2(n_7279),
.B(n_8770),
.Y(n_10834)
);

AOI22xp33_ASAP7_75t_L g10835 ( 
.A1(n_9461),
.A2(n_9462),
.B1(n_9544),
.B2(n_9536),
.Y(n_10835)
);

AOI22xp33_ASAP7_75t_L g10836 ( 
.A1(n_9462),
.A2(n_8014),
.B1(n_7765),
.B2(n_8381),
.Y(n_10836)
);

OAI221xp5_ASAP7_75t_L g10837 ( 
.A1(n_9827),
.A2(n_9970),
.B1(n_9987),
.B2(n_9953),
.C(n_9941),
.Y(n_10837)
);

OAI221xp5_ASAP7_75t_L g10838 ( 
.A1(n_9970),
.A2(n_8356),
.B1(n_8333),
.B2(n_8744),
.C(n_8736),
.Y(n_10838)
);

AOI22xp5_ASAP7_75t_L g10839 ( 
.A1(n_10285),
.A2(n_10053),
.B1(n_10091),
.B2(n_9949),
.Y(n_10839)
);

AOI22xp33_ASAP7_75t_SL g10840 ( 
.A1(n_9970),
.A2(n_8386),
.B1(n_8381),
.B2(n_8356),
.Y(n_10840)
);

OAI21x1_ASAP7_75t_L g10841 ( 
.A1(n_9892),
.A2(n_8714),
.B(n_8659),
.Y(n_10841)
);

OAI21xp5_ASAP7_75t_SL g10842 ( 
.A1(n_9550),
.A2(n_7811),
.B(n_8797),
.Y(n_10842)
);

INVx1_ASAP7_75t_L g10843 ( 
.A(n_9552),
.Y(n_10843)
);

INVx1_ASAP7_75t_L g10844 ( 
.A(n_9554),
.Y(n_10844)
);

AOI22xp33_ASAP7_75t_L g10845 ( 
.A1(n_9536),
.A2(n_8386),
.B1(n_8381),
.B2(n_7516),
.Y(n_10845)
);

OAI22xp33_ASAP7_75t_L g10846 ( 
.A1(n_9616),
.A2(n_7686),
.B1(n_7874),
.B2(n_7393),
.Y(n_10846)
);

OAI21x1_ASAP7_75t_L g10847 ( 
.A1(n_9892),
.A2(n_8801),
.B(n_8659),
.Y(n_10847)
);

NAND2xp5_ASAP7_75t_L g10848 ( 
.A(n_9817),
.B(n_7683),
.Y(n_10848)
);

AOI22xp33_ASAP7_75t_L g10849 ( 
.A1(n_9544),
.A2(n_8386),
.B1(n_7516),
.B2(n_7545),
.Y(n_10849)
);

OAI22xp33_ASAP7_75t_L g10850 ( 
.A1(n_9761),
.A2(n_7874),
.B1(n_7393),
.B2(n_7554),
.Y(n_10850)
);

OAI221xp5_ASAP7_75t_L g10851 ( 
.A1(n_9987),
.A2(n_8356),
.B1(n_8333),
.B2(n_8744),
.C(n_8736),
.Y(n_10851)
);

INVx1_ASAP7_75t_L g10852 ( 
.A(n_9558),
.Y(n_10852)
);

INVx1_ASAP7_75t_L g10853 ( 
.A(n_9560),
.Y(n_10853)
);

HB1xp67_ASAP7_75t_L g10854 ( 
.A(n_9885),
.Y(n_10854)
);

AOI22xp33_ASAP7_75t_L g10855 ( 
.A1(n_9548),
.A2(n_7516),
.B1(n_7545),
.B2(n_8747),
.Y(n_10855)
);

A2O1A1Ixp33_ASAP7_75t_L g10856 ( 
.A1(n_9987),
.A2(n_8747),
.B(n_7626),
.C(n_7928),
.Y(n_10856)
);

INVx1_ASAP7_75t_L g10857 ( 
.A(n_9563),
.Y(n_10857)
);

INVx2_ASAP7_75t_L g10858 ( 
.A(n_10395),
.Y(n_10858)
);

OAI221xp5_ASAP7_75t_L g10859 ( 
.A1(n_10004),
.A2(n_8953),
.B1(n_8933),
.B2(n_8905),
.C(n_8904),
.Y(n_10859)
);

BUFx6f_ASAP7_75t_L g10860 ( 
.A(n_9538),
.Y(n_10860)
);

AND2x4_ASAP7_75t_L g10861 ( 
.A(n_9896),
.B(n_8384),
.Y(n_10861)
);

INVx1_ASAP7_75t_L g10862 ( 
.A(n_9565),
.Y(n_10862)
);

INVxp67_ASAP7_75t_SL g10863 ( 
.A(n_9926),
.Y(n_10863)
);

OAI22xp5_ASAP7_75t_L g10864 ( 
.A1(n_9550),
.A2(n_8213),
.B1(n_8221),
.B2(n_9089),
.Y(n_10864)
);

AOI22xp33_ASAP7_75t_L g10865 ( 
.A1(n_9548),
.A2(n_9561),
.B1(n_9564),
.B2(n_9559),
.Y(n_10865)
);

AO22x1_ASAP7_75t_L g10866 ( 
.A1(n_10180),
.A2(n_8384),
.B1(n_8383),
.B2(n_8345),
.Y(n_10866)
);

AOI22xp33_ASAP7_75t_L g10867 ( 
.A1(n_9559),
.A2(n_7516),
.B1(n_7813),
.B2(n_7417),
.Y(n_10867)
);

NAND2xp5_ASAP7_75t_L g10868 ( 
.A(n_9822),
.B(n_7683),
.Y(n_10868)
);

AOI22xp33_ASAP7_75t_L g10869 ( 
.A1(n_9561),
.A2(n_7516),
.B1(n_7813),
.B2(n_7417),
.Y(n_10869)
);

A2O1A1Ixp33_ASAP7_75t_L g10870 ( 
.A1(n_10004),
.A2(n_9674),
.B(n_9570),
.C(n_9553),
.Y(n_10870)
);

INVx1_ASAP7_75t_L g10871 ( 
.A(n_9566),
.Y(n_10871)
);

AOI22xp33_ASAP7_75t_L g10872 ( 
.A1(n_9564),
.A2(n_7516),
.B1(n_7813),
.B2(n_7417),
.Y(n_10872)
);

AOI22xp33_ASAP7_75t_L g10873 ( 
.A1(n_9575),
.A2(n_7813),
.B1(n_7417),
.B2(n_8201),
.Y(n_10873)
);

NAND2xp5_ASAP7_75t_L g10874 ( 
.A(n_9839),
.B(n_7683),
.Y(n_10874)
);

OAI33xp33_ASAP7_75t_L g10875 ( 
.A1(n_10391),
.A2(n_9139),
.A3(n_7937),
.B1(n_9385),
.B2(n_7405),
.B3(n_9319),
.Y(n_10875)
);

AOI21xp5_ASAP7_75t_L g10876 ( 
.A1(n_10000),
.A2(n_8793),
.B(n_8770),
.Y(n_10876)
);

OR2x6_ASAP7_75t_L g10877 ( 
.A(n_9499),
.B(n_6637),
.Y(n_10877)
);

INVx1_ASAP7_75t_L g10878 ( 
.A(n_9569),
.Y(n_10878)
);

OAI22xp33_ASAP7_75t_L g10879 ( 
.A1(n_9761),
.A2(n_7393),
.B1(n_7554),
.B2(n_7225),
.Y(n_10879)
);

BUFx12f_ASAP7_75t_L g10880 ( 
.A(n_9880),
.Y(n_10880)
);

INVx4_ASAP7_75t_SL g10881 ( 
.A(n_10080),
.Y(n_10881)
);

OAI211xp5_ASAP7_75t_L g10882 ( 
.A1(n_9777),
.A2(n_8401),
.B(n_8446),
.C(n_8411),
.Y(n_10882)
);

AND2x2_ASAP7_75t_L g10883 ( 
.A(n_10180),
.B(n_9065),
.Y(n_10883)
);

OAI22xp5_ASAP7_75t_L g10884 ( 
.A1(n_10040),
.A2(n_8221),
.B1(n_8288),
.B2(n_8281),
.Y(n_10884)
);

INVx5_ASAP7_75t_SL g10885 ( 
.A(n_9696),
.Y(n_10885)
);

INVx1_ASAP7_75t_L g10886 ( 
.A(n_9571),
.Y(n_10886)
);

AOI222xp33_ASAP7_75t_L g10887 ( 
.A1(n_10099),
.A2(n_10004),
.B1(n_9597),
.B2(n_9483),
.C1(n_9627),
.C2(n_9494),
.Y(n_10887)
);

AOI22xp33_ASAP7_75t_L g10888 ( 
.A1(n_9575),
.A2(n_9585),
.B1(n_9588),
.B2(n_9578),
.Y(n_10888)
);

A2O1A1Ixp33_ASAP7_75t_L g10889 ( 
.A1(n_9674),
.A2(n_7626),
.B(n_7928),
.C(n_7546),
.Y(n_10889)
);

AOI22xp33_ASAP7_75t_L g10890 ( 
.A1(n_9578),
.A2(n_9588),
.B1(n_9599),
.B2(n_9585),
.Y(n_10890)
);

AOI22xp33_ASAP7_75t_L g10891 ( 
.A1(n_9599),
.A2(n_7813),
.B1(n_7417),
.B2(n_8201),
.Y(n_10891)
);

AOI22xp33_ASAP7_75t_L g10892 ( 
.A1(n_9601),
.A2(n_7813),
.B1(n_8210),
.B2(n_9016),
.Y(n_10892)
);

AOI22xp33_ASAP7_75t_L g10893 ( 
.A1(n_9601),
.A2(n_8210),
.B1(n_9097),
.B2(n_9016),
.Y(n_10893)
);

AOI22xp33_ASAP7_75t_L g10894 ( 
.A1(n_9602),
.A2(n_9097),
.B1(n_9130),
.B2(n_9016),
.Y(n_10894)
);

OR2x2_ASAP7_75t_L g10895 ( 
.A(n_9620),
.B(n_7225),
.Y(n_10895)
);

OAI21x1_ASAP7_75t_L g10896 ( 
.A1(n_10174),
.A2(n_8801),
.B(n_9373),
.Y(n_10896)
);

INVx2_ASAP7_75t_L g10897 ( 
.A(n_10398),
.Y(n_10897)
);

OAI22xp33_ASAP7_75t_L g10898 ( 
.A1(n_9761),
.A2(n_7554),
.B1(n_7225),
.B2(n_7689),
.Y(n_10898)
);

INVx3_ASAP7_75t_L g10899 ( 
.A(n_10265),
.Y(n_10899)
);

AOI21xp5_ASAP7_75t_L g10900 ( 
.A1(n_10191),
.A2(n_8823),
.B(n_8793),
.Y(n_10900)
);

NAND2xp5_ASAP7_75t_L g10901 ( 
.A(n_9859),
.B(n_7683),
.Y(n_10901)
);

AOI22xp33_ASAP7_75t_L g10902 ( 
.A1(n_9602),
.A2(n_9130),
.B1(n_9205),
.B2(n_9097),
.Y(n_10902)
);

AOI22xp5_ASAP7_75t_L g10903 ( 
.A1(n_9949),
.A2(n_8184),
.B1(n_8100),
.B2(n_9293),
.Y(n_10903)
);

NAND2xp5_ASAP7_75t_L g10904 ( 
.A(n_9755),
.B(n_7683),
.Y(n_10904)
);

AOI211xp5_ASAP7_75t_L g10905 ( 
.A1(n_9570),
.A2(n_7779),
.B(n_7275),
.C(n_8227),
.Y(n_10905)
);

AOI22xp33_ASAP7_75t_L g10906 ( 
.A1(n_9607),
.A2(n_9205),
.B1(n_9317),
.B2(n_9130),
.Y(n_10906)
);

INVx1_ASAP7_75t_L g10907 ( 
.A(n_9574),
.Y(n_10907)
);

NOR3xp33_ASAP7_75t_L g10908 ( 
.A(n_10333),
.B(n_8411),
.C(n_8401),
.Y(n_10908)
);

INVx2_ASAP7_75t_L g10909 ( 
.A(n_10398),
.Y(n_10909)
);

INVx2_ASAP7_75t_L g10910 ( 
.A(n_10405),
.Y(n_10910)
);

AOI33xp33_ASAP7_75t_L g10911 ( 
.A1(n_10150),
.A2(n_9143),
.A3(n_9133),
.B1(n_9163),
.B2(n_9142),
.B3(n_9123),
.Y(n_10911)
);

AO221x2_ASAP7_75t_L g10912 ( 
.A1(n_9874),
.A2(n_7972),
.B1(n_8100),
.B2(n_9248),
.C(n_8184),
.Y(n_10912)
);

BUFx4f_ASAP7_75t_SL g10913 ( 
.A(n_9696),
.Y(n_10913)
);

AND2x2_ASAP7_75t_L g10914 ( 
.A(n_10208),
.B(n_9065),
.Y(n_10914)
);

OR2x2_ASAP7_75t_L g10915 ( 
.A(n_9720),
.B(n_7683),
.Y(n_10915)
);

OAI22xp5_ASAP7_75t_L g10916 ( 
.A1(n_10040),
.A2(n_8288),
.B1(n_8281),
.B2(n_7730),
.Y(n_10916)
);

AOI22xp33_ASAP7_75t_SL g10917 ( 
.A1(n_9777),
.A2(n_7701),
.B1(n_7863),
.B2(n_8558),
.Y(n_10917)
);

BUFx2_ASAP7_75t_L g10918 ( 
.A(n_9457),
.Y(n_10918)
);

AOI22x1_ASAP7_75t_L g10919 ( 
.A1(n_9496),
.A2(n_8658),
.B1(n_8710),
.B2(n_8446),
.Y(n_10919)
);

OA21x2_ASAP7_75t_L g10920 ( 
.A1(n_9975),
.A2(n_8824),
.B(n_8818),
.Y(n_10920)
);

OAI22xp33_ASAP7_75t_L g10921 ( 
.A1(n_9850),
.A2(n_9982),
.B1(n_9483),
.B2(n_9494),
.Y(n_10921)
);

INVx1_ASAP7_75t_L g10922 ( 
.A(n_9576),
.Y(n_10922)
);

OAI22xp5_ASAP7_75t_L g10923 ( 
.A1(n_10040),
.A2(n_7730),
.B1(n_7755),
.B2(n_7531),
.Y(n_10923)
);

OR2x2_ASAP7_75t_L g10924 ( 
.A(n_9771),
.B(n_8175),
.Y(n_10924)
);

OAI22xp5_ASAP7_75t_L g10925 ( 
.A1(n_10084),
.A2(n_7730),
.B1(n_7755),
.B2(n_7531),
.Y(n_10925)
);

CKINVDCx20_ASAP7_75t_R g10926 ( 
.A(n_9926),
.Y(n_10926)
);

OAI22xp5_ASAP7_75t_L g10927 ( 
.A1(n_10084),
.A2(n_7755),
.B1(n_7841),
.B2(n_7531),
.Y(n_10927)
);

AOI21xp33_ASAP7_75t_R g10928 ( 
.A1(n_9455),
.A2(n_8733),
.B(n_9316),
.Y(n_10928)
);

AOI22xp33_ASAP7_75t_L g10929 ( 
.A1(n_9607),
.A2(n_9317),
.B1(n_9205),
.B2(n_7689),
.Y(n_10929)
);

NAND2xp5_ASAP7_75t_L g10930 ( 
.A(n_9529),
.B(n_9894),
.Y(n_10930)
);

BUFx12f_ASAP7_75t_L g10931 ( 
.A(n_9467),
.Y(n_10931)
);

AOI22xp5_ASAP7_75t_L g10932 ( 
.A1(n_10053),
.A2(n_9282),
.B1(n_9043),
.B2(n_8711),
.Y(n_10932)
);

BUFx6f_ASAP7_75t_L g10933 ( 
.A(n_9625),
.Y(n_10933)
);

HB1xp67_ASAP7_75t_L g10934 ( 
.A(n_9921),
.Y(n_10934)
);

HB1xp67_ASAP7_75t_L g10935 ( 
.A(n_9928),
.Y(n_10935)
);

OAI22xp33_ASAP7_75t_L g10936 ( 
.A1(n_9850),
.A2(n_7689),
.B1(n_7824),
.B2(n_7814),
.Y(n_10936)
);

AOI221xp5_ASAP7_75t_L g10937 ( 
.A1(n_10390),
.A2(n_9136),
.B1(n_9148),
.B2(n_9145),
.C(n_9138),
.Y(n_10937)
);

OA21x2_ASAP7_75t_L g10938 ( 
.A1(n_9976),
.A2(n_8824),
.B(n_8818),
.Y(n_10938)
);

NOR2xp67_ASAP7_75t_L g10939 ( 
.A(n_10286),
.B(n_9123),
.Y(n_10939)
);

INVx1_ASAP7_75t_L g10940 ( 
.A(n_9577),
.Y(n_10940)
);

NAND2xp5_ASAP7_75t_L g10941 ( 
.A(n_10032),
.B(n_8823),
.Y(n_10941)
);

AOI221xp5_ASAP7_75t_SL g10942 ( 
.A1(n_10264),
.A2(n_7731),
.B1(n_7884),
.B2(n_8112),
.C(n_7972),
.Y(n_10942)
);

OAI22xp5_ASAP7_75t_L g10943 ( 
.A1(n_10084),
.A2(n_9833),
.B1(n_9802),
.B2(n_9496),
.Y(n_10943)
);

AOI221xp5_ASAP7_75t_L g10944 ( 
.A1(n_10390),
.A2(n_9136),
.B1(n_9148),
.B2(n_9145),
.C(n_9138),
.Y(n_10944)
);

AND2x2_ASAP7_75t_L g10945 ( 
.A(n_10208),
.B(n_9065),
.Y(n_10945)
);

AOI22xp33_ASAP7_75t_L g10946 ( 
.A1(n_9611),
.A2(n_9317),
.B1(n_7689),
.B2(n_7824),
.Y(n_10946)
);

INVx2_ASAP7_75t_L g10947 ( 
.A(n_10405),
.Y(n_10947)
);

AND2x4_ASAP7_75t_L g10948 ( 
.A(n_9896),
.B(n_9144),
.Y(n_10948)
);

OAI22xp5_ASAP7_75t_L g10949 ( 
.A1(n_9802),
.A2(n_7841),
.B1(n_9142),
.B2(n_9133),
.Y(n_10949)
);

BUFx3_ASAP7_75t_L g10950 ( 
.A(n_9955),
.Y(n_10950)
);

OAI22xp5_ASAP7_75t_L g10951 ( 
.A1(n_9833),
.A2(n_7841),
.B1(n_9163),
.B2(n_9143),
.Y(n_10951)
);

INVx1_ASAP7_75t_L g10952 ( 
.A(n_9586),
.Y(n_10952)
);

OR2x2_ASAP7_75t_L g10953 ( 
.A(n_9807),
.B(n_8175),
.Y(n_10953)
);

OAI211xp5_ASAP7_75t_L g10954 ( 
.A1(n_9777),
.A2(n_9483),
.B(n_9494),
.C(n_9455),
.Y(n_10954)
);

AND2x4_ASAP7_75t_L g10955 ( 
.A(n_9901),
.B(n_9144),
.Y(n_10955)
);

INVx4_ASAP7_75t_L g10956 ( 
.A(n_9592),
.Y(n_10956)
);

AOI22xp33_ASAP7_75t_SL g10957 ( 
.A1(n_10091),
.A2(n_7701),
.B1(n_7863),
.B2(n_8558),
.Y(n_10957)
);

AOI22xp33_ASAP7_75t_SL g10958 ( 
.A1(n_10386),
.A2(n_7701),
.B1(n_7863),
.B2(n_8683),
.Y(n_10958)
);

NOR2xp33_ASAP7_75t_L g10959 ( 
.A(n_9740),
.B(n_8943),
.Y(n_10959)
);

NAND2xp5_ASAP7_75t_L g10960 ( 
.A(n_10061),
.B(n_8293),
.Y(n_10960)
);

OR2x2_ASAP7_75t_L g10961 ( 
.A(n_9821),
.B(n_8175),
.Y(n_10961)
);

AND2x2_ASAP7_75t_L g10962 ( 
.A(n_10208),
.B(n_9144),
.Y(n_10962)
);

INVx2_ASAP7_75t_L g10963 ( 
.A(n_10224),
.Y(n_10963)
);

INVx1_ASAP7_75t_L g10964 ( 
.A(n_9590),
.Y(n_10964)
);

AOI22xp33_ASAP7_75t_SL g10965 ( 
.A1(n_10323),
.A2(n_8683),
.B1(n_8763),
.B2(n_7279),
.Y(n_10965)
);

INVx1_ASAP7_75t_L g10966 ( 
.A(n_9593),
.Y(n_10966)
);

AOI22xp33_ASAP7_75t_L g10967 ( 
.A1(n_9611),
.A2(n_7814),
.B1(n_7832),
.B2(n_7824),
.Y(n_10967)
);

INVx1_ASAP7_75t_L g10968 ( 
.A(n_9596),
.Y(n_10968)
);

OR2x2_ASAP7_75t_L g10969 ( 
.A(n_9832),
.B(n_8192),
.Y(n_10969)
);

NAND3xp33_ASAP7_75t_L g10970 ( 
.A(n_10070),
.B(n_7279),
.C(n_9077),
.Y(n_10970)
);

AOI22xp33_ASAP7_75t_L g10971 ( 
.A1(n_9612),
.A2(n_7814),
.B1(n_7832),
.B2(n_7824),
.Y(n_10971)
);

BUFx3_ASAP7_75t_L g10972 ( 
.A(n_9955),
.Y(n_10972)
);

OAI22xp5_ASAP7_75t_L g10973 ( 
.A1(n_10186),
.A2(n_9421),
.B1(n_9412),
.B2(n_7832),
.Y(n_10973)
);

OAI22xp5_ASAP7_75t_L g10974 ( 
.A1(n_10186),
.A2(n_9421),
.B1(n_7832),
.B2(n_7889),
.Y(n_10974)
);

AOI222xp33_ASAP7_75t_L g10975 ( 
.A1(n_9455),
.A2(n_7884),
.B1(n_8236),
.B2(n_9198),
.C1(n_9196),
.C2(n_9178),
.Y(n_10975)
);

AOI21xp5_ASAP7_75t_L g10976 ( 
.A1(n_9846),
.A2(n_8646),
.B(n_8643),
.Y(n_10976)
);

AOI22xp33_ASAP7_75t_L g10977 ( 
.A1(n_9612),
.A2(n_7814),
.B1(n_7899),
.B2(n_7889),
.Y(n_10977)
);

INVx1_ASAP7_75t_L g10978 ( 
.A(n_9610),
.Y(n_10978)
);

OAI221xp5_ASAP7_75t_L g10979 ( 
.A1(n_9982),
.A2(n_8586),
.B1(n_8735),
.B2(n_8574),
.C(n_8550),
.Y(n_10979)
);

AOI21xp5_ASAP7_75t_L g10980 ( 
.A1(n_9846),
.A2(n_8646),
.B(n_8643),
.Y(n_10980)
);

INVx1_ASAP7_75t_L g10981 ( 
.A(n_9613),
.Y(n_10981)
);

CKINVDCx16_ASAP7_75t_R g10982 ( 
.A(n_10018),
.Y(n_10982)
);

AOI22xp33_ASAP7_75t_SL g10983 ( 
.A1(n_10386),
.A2(n_8683),
.B1(n_8763),
.B2(n_7279),
.Y(n_10983)
);

OAI33xp33_ASAP7_75t_L g10984 ( 
.A1(n_10137),
.A2(n_9629),
.A3(n_9626),
.B1(n_9630),
.B2(n_9628),
.B3(n_9621),
.Y(n_10984)
);

NAND2xp5_ASAP7_75t_L g10985 ( 
.A(n_10073),
.B(n_8300),
.Y(n_10985)
);

INVx1_ASAP7_75t_L g10986 ( 
.A(n_9632),
.Y(n_10986)
);

AOI22xp33_ASAP7_75t_L g10987 ( 
.A1(n_9622),
.A2(n_7889),
.B1(n_7899),
.B2(n_8388),
.Y(n_10987)
);

OR2x6_ASAP7_75t_L g10988 ( 
.A(n_9484),
.B(n_6647),
.Y(n_10988)
);

AOI22xp33_ASAP7_75t_SL g10989 ( 
.A1(n_10323),
.A2(n_8683),
.B1(n_8763),
.B2(n_7279),
.Y(n_10989)
);

NAND3xp33_ASAP7_75t_L g10990 ( 
.A(n_10078),
.B(n_9152),
.C(n_9077),
.Y(n_10990)
);

INVx1_ASAP7_75t_L g10991 ( 
.A(n_9637),
.Y(n_10991)
);

A2O1A1Ixp33_ASAP7_75t_L g10992 ( 
.A1(n_9942),
.A2(n_7928),
.B(n_7546),
.C(n_8921),
.Y(n_10992)
);

INVx3_ASAP7_75t_L g10993 ( 
.A(n_9508),
.Y(n_10993)
);

AOI221xp5_ASAP7_75t_L g10994 ( 
.A1(n_9744),
.A2(n_9196),
.B1(n_9201),
.B2(n_9198),
.C(n_9178),
.Y(n_10994)
);

INVx4_ASAP7_75t_L g10995 ( 
.A(n_9592),
.Y(n_10995)
);

OAI211xp5_ASAP7_75t_SL g10996 ( 
.A1(n_9597),
.A2(n_9666),
.B(n_9714),
.C(n_9627),
.Y(n_10996)
);

AOI22xp33_ASAP7_75t_L g10997 ( 
.A1(n_9622),
.A2(n_7889),
.B1(n_7899),
.B2(n_8388),
.Y(n_10997)
);

CKINVDCx5p33_ASAP7_75t_R g10998 ( 
.A(n_10090),
.Y(n_10998)
);

AOI22xp33_ASAP7_75t_L g10999 ( 
.A1(n_9635),
.A2(n_9646),
.B1(n_9651),
.B2(n_9636),
.Y(n_10999)
);

OAI22xp5_ASAP7_75t_L g11000 ( 
.A1(n_10186),
.A2(n_7899),
.B1(n_7212),
.B2(n_7915),
.Y(n_11000)
);

AOI22xp33_ASAP7_75t_L g11001 ( 
.A1(n_9635),
.A2(n_8388),
.B1(n_8464),
.B2(n_8423),
.Y(n_11001)
);

OR2x2_ASAP7_75t_L g11002 ( 
.A(n_9934),
.B(n_8192),
.Y(n_11002)
);

AOI221xp5_ASAP7_75t_L g11003 ( 
.A1(n_9714),
.A2(n_9208),
.B1(n_9209),
.B2(n_9201),
.C(n_8236),
.Y(n_11003)
);

AOI222xp33_ASAP7_75t_L g11004 ( 
.A1(n_9597),
.A2(n_9208),
.B1(n_9209),
.B2(n_7183),
.C1(n_7210),
.C2(n_7209),
.Y(n_11004)
);

AOI22xp33_ASAP7_75t_L g11005 ( 
.A1(n_9636),
.A2(n_8388),
.B1(n_8464),
.B2(n_8423),
.Y(n_11005)
);

AND2x2_ASAP7_75t_L g11006 ( 
.A(n_10360),
.B(n_9153),
.Y(n_11006)
);

AOI22xp33_ASAP7_75t_L g11007 ( 
.A1(n_9646),
.A2(n_8423),
.B1(n_8585),
.B2(n_8464),
.Y(n_11007)
);

AND2x4_ASAP7_75t_SL g11008 ( 
.A(n_9508),
.B(n_6965),
.Y(n_11008)
);

INVxp67_ASAP7_75t_L g11009 ( 
.A(n_10018),
.Y(n_11009)
);

AOI22xp33_ASAP7_75t_L g11010 ( 
.A1(n_9651),
.A2(n_8423),
.B1(n_8585),
.B2(n_8464),
.Y(n_11010)
);

AOI22xp33_ASAP7_75t_SL g11011 ( 
.A1(n_9650),
.A2(n_8763),
.B1(n_7353),
.B2(n_7342),
.Y(n_11011)
);

INVxp67_ASAP7_75t_SL g11012 ( 
.A(n_9825),
.Y(n_11012)
);

AOI22xp33_ASAP7_75t_L g11013 ( 
.A1(n_9653),
.A2(n_8585),
.B1(n_8639),
.B2(n_8637),
.Y(n_11013)
);

AOI22xp33_ASAP7_75t_L g11014 ( 
.A1(n_9653),
.A2(n_8585),
.B1(n_8639),
.B2(n_8637),
.Y(n_11014)
);

AOI22xp33_ASAP7_75t_L g11015 ( 
.A1(n_9663),
.A2(n_8637),
.B1(n_8740),
.B2(n_8639),
.Y(n_11015)
);

AND2x2_ASAP7_75t_L g11016 ( 
.A(n_10360),
.B(n_9153),
.Y(n_11016)
);

AOI22xp33_ASAP7_75t_L g11017 ( 
.A1(n_9663),
.A2(n_8637),
.B1(n_8740),
.B2(n_8639),
.Y(n_11017)
);

OAI22xp5_ASAP7_75t_L g11018 ( 
.A1(n_10214),
.A2(n_7915),
.B1(n_7334),
.B2(n_7362),
.Y(n_11018)
);

AOI22xp33_ASAP7_75t_L g11019 ( 
.A1(n_9665),
.A2(n_8740),
.B1(n_8791),
.B2(n_7681),
.Y(n_11019)
);

OAI22xp33_ASAP7_75t_L g11020 ( 
.A1(n_9850),
.A2(n_8218),
.B1(n_7870),
.B2(n_7825),
.Y(n_11020)
);

AOI22xp33_ASAP7_75t_L g11021 ( 
.A1(n_9665),
.A2(n_8740),
.B1(n_8791),
.B2(n_7681),
.Y(n_11021)
);

INVx1_ASAP7_75t_L g11022 ( 
.A(n_9641),
.Y(n_11022)
);

INVx1_ASAP7_75t_L g11023 ( 
.A(n_9645),
.Y(n_11023)
);

AOI22xp5_ASAP7_75t_L g11024 ( 
.A1(n_9982),
.A2(n_8122),
.B1(n_8132),
.B2(n_8799),
.Y(n_11024)
);

INVx1_ASAP7_75t_L g11025 ( 
.A(n_9648),
.Y(n_11025)
);

AOI221xp5_ASAP7_75t_L g11026 ( 
.A1(n_9666),
.A2(n_7210),
.B1(n_7209),
.B2(n_7183),
.C(n_8978),
.Y(n_11026)
);

OAI21xp5_ASAP7_75t_L g11027 ( 
.A1(n_10007),
.A2(n_8947),
.B(n_8928),
.Y(n_11027)
);

CKINVDCx20_ASAP7_75t_R g11028 ( 
.A(n_10090),
.Y(n_11028)
);

AOI22xp5_ASAP7_75t_L g11029 ( 
.A1(n_9650),
.A2(n_9662),
.B1(n_10165),
.B2(n_10150),
.Y(n_11029)
);

AOI22xp33_ASAP7_75t_L g11030 ( 
.A1(n_9667),
.A2(n_8791),
.B1(n_7681),
.B2(n_8090),
.Y(n_11030)
);

NAND2xp5_ASAP7_75t_L g11031 ( 
.A(n_10083),
.B(n_10096),
.Y(n_11031)
);

OAI22xp33_ASAP7_75t_L g11032 ( 
.A1(n_9627),
.A2(n_8218),
.B1(n_7870),
.B2(n_7825),
.Y(n_11032)
);

OR2x6_ASAP7_75t_L g11033 ( 
.A(n_9486),
.B(n_6647),
.Y(n_11033)
);

AOI21xp5_ASAP7_75t_L g11034 ( 
.A1(n_10185),
.A2(n_8680),
.B(n_7737),
.Y(n_11034)
);

INVx1_ASAP7_75t_L g11035 ( 
.A(n_9652),
.Y(n_11035)
);

AOI221xp5_ASAP7_75t_L g11036 ( 
.A1(n_9666),
.A2(n_7210),
.B1(n_7209),
.B2(n_7183),
.C(n_8978),
.Y(n_11036)
);

CKINVDCx20_ASAP7_75t_R g11037 ( 
.A(n_9507),
.Y(n_11037)
);

HB1xp67_ASAP7_75t_L g11038 ( 
.A(n_10098),
.Y(n_11038)
);

AOI22xp33_ASAP7_75t_L g11039 ( 
.A1(n_9667),
.A2(n_8791),
.B1(n_7681),
.B2(n_8090),
.Y(n_11039)
);

AOI22xp33_ASAP7_75t_L g11040 ( 
.A1(n_9678),
.A2(n_9683),
.B1(n_9684),
.B2(n_9681),
.Y(n_11040)
);

INVx2_ASAP7_75t_L g11041 ( 
.A(n_10224),
.Y(n_11041)
);

INVx1_ASAP7_75t_L g11042 ( 
.A(n_9654),
.Y(n_11042)
);

OAI22xp5_ASAP7_75t_L g11043 ( 
.A1(n_10214),
.A2(n_7915),
.B1(n_7334),
.B2(n_7362),
.Y(n_11043)
);

NAND2xp5_ASAP7_75t_L g11044 ( 
.A(n_10129),
.B(n_8300),
.Y(n_11044)
);

INVx1_ASAP7_75t_L g11045 ( 
.A(n_9655),
.Y(n_11045)
);

INVx1_ASAP7_75t_L g11046 ( 
.A(n_9657),
.Y(n_11046)
);

AOI22xp33_ASAP7_75t_L g11047 ( 
.A1(n_9678),
.A2(n_8045),
.B1(n_7881),
.B2(n_7784),
.Y(n_11047)
);

OAI22xp5_ASAP7_75t_L g11048 ( 
.A1(n_10214),
.A2(n_7334),
.B1(n_7362),
.B2(n_7161),
.Y(n_11048)
);

AOI221xp5_ASAP7_75t_L g11049 ( 
.A1(n_9714),
.A2(n_8989),
.B1(n_8997),
.B2(n_8981),
.C(n_8978),
.Y(n_11049)
);

NAND2xp5_ASAP7_75t_L g11050 ( 
.A(n_10153),
.B(n_9023),
.Y(n_11050)
);

OAI22xp5_ASAP7_75t_SL g11051 ( 
.A1(n_9525),
.A2(n_6649),
.B1(n_6499),
.B2(n_6561),
.Y(n_11051)
);

BUFx3_ASAP7_75t_L g11052 ( 
.A(n_9568),
.Y(n_11052)
);

BUFx5_ASAP7_75t_L g11053 ( 
.A(n_9625),
.Y(n_11053)
);

AOI22xp5_ASAP7_75t_L g11054 ( 
.A1(n_9662),
.A2(n_8122),
.B1(n_8132),
.B2(n_8806),
.Y(n_11054)
);

AOI21xp33_ASAP7_75t_L g11055 ( 
.A1(n_10212),
.A2(n_7220),
.B(n_7181),
.Y(n_11055)
);

OR2x6_ASAP7_75t_L g11056 ( 
.A(n_9591),
.B(n_6649),
.Y(n_11056)
);

AOI21xp5_ASAP7_75t_L g11057 ( 
.A1(n_10007),
.A2(n_8680),
.B(n_7737),
.Y(n_11057)
);

INVx1_ASAP7_75t_L g11058 ( 
.A(n_9671),
.Y(n_11058)
);

AND2x2_ASAP7_75t_L g11059 ( 
.A(n_10360),
.B(n_9153),
.Y(n_11059)
);

BUFx6f_ASAP7_75t_L g11060 ( 
.A(n_9508),
.Y(n_11060)
);

INVx1_ASAP7_75t_L g11061 ( 
.A(n_9679),
.Y(n_11061)
);

AO31x2_ASAP7_75t_L g11062 ( 
.A1(n_10358),
.A2(n_8710),
.A3(n_8658),
.B(n_8818),
.Y(n_11062)
);

AOI222xp33_ASAP7_75t_L g11063 ( 
.A1(n_9744),
.A2(n_9327),
.B1(n_8989),
.B2(n_9330),
.C1(n_8997),
.C2(n_8981),
.Y(n_11063)
);

INVx1_ASAP7_75t_SL g11064 ( 
.A(n_9466),
.Y(n_11064)
);

OAI21xp33_ASAP7_75t_L g11065 ( 
.A1(n_10165),
.A2(n_9419),
.B(n_9416),
.Y(n_11065)
);

INVx4_ASAP7_75t_L g11066 ( 
.A(n_10080),
.Y(n_11066)
);

HB1xp67_ASAP7_75t_L g11067 ( 
.A(n_10160),
.Y(n_11067)
);

AOI22xp33_ASAP7_75t_L g11068 ( 
.A1(n_9681),
.A2(n_8045),
.B1(n_7881),
.B2(n_7784),
.Y(n_11068)
);

NAND3xp33_ASAP7_75t_L g11069 ( 
.A(n_10178),
.B(n_9152),
.C(n_9077),
.Y(n_11069)
);

INVx1_ASAP7_75t_L g11070 ( 
.A(n_9687),
.Y(n_11070)
);

BUFx2_ASAP7_75t_L g11071 ( 
.A(n_9979),
.Y(n_11071)
);

AOI22xp33_ASAP7_75t_L g11072 ( 
.A1(n_9683),
.A2(n_7784),
.B1(n_8758),
.B2(n_8751),
.Y(n_11072)
);

AOI22xp33_ASAP7_75t_L g11073 ( 
.A1(n_9684),
.A2(n_7784),
.B1(n_8746),
.B2(n_8080),
.Y(n_11073)
);

AOI22xp33_ASAP7_75t_SL g11074 ( 
.A1(n_9744),
.A2(n_7353),
.B1(n_7342),
.B2(n_8775),
.Y(n_11074)
);

OAI22xp33_ASAP7_75t_L g11075 ( 
.A1(n_10223),
.A2(n_7870),
.B1(n_7825),
.B2(n_7914),
.Y(n_11075)
);

AOI22xp33_ASAP7_75t_SL g11076 ( 
.A1(n_10173),
.A2(n_7353),
.B1(n_7342),
.B2(n_8775),
.Y(n_11076)
);

BUFx2_ASAP7_75t_L g11077 ( 
.A(n_9508),
.Y(n_11077)
);

BUFx6f_ASAP7_75t_L g11078 ( 
.A(n_9555),
.Y(n_11078)
);

HB1xp67_ASAP7_75t_L g11079 ( 
.A(n_10181),
.Y(n_11079)
);

OAI221xp5_ASAP7_75t_L g11080 ( 
.A1(n_9697),
.A2(n_8837),
.B1(n_8869),
.B2(n_8749),
.C(n_8741),
.Y(n_11080)
);

AOI22xp33_ASAP7_75t_L g11081 ( 
.A1(n_9697),
.A2(n_7784),
.B1(n_8080),
.B2(n_8018),
.Y(n_11081)
);

INVx1_ASAP7_75t_L g11082 ( 
.A(n_9690),
.Y(n_11082)
);

AOI222xp33_ASAP7_75t_L g11083 ( 
.A1(n_9701),
.A2(n_9327),
.B1(n_8989),
.B2(n_9330),
.C1(n_8997),
.C2(n_8981),
.Y(n_11083)
);

AOI22xp33_ASAP7_75t_L g11084 ( 
.A1(n_9701),
.A2(n_7784),
.B1(n_8018),
.B2(n_7982),
.Y(n_11084)
);

AOI22xp33_ASAP7_75t_L g11085 ( 
.A1(n_9702),
.A2(n_7982),
.B1(n_7913),
.B2(n_8406),
.Y(n_11085)
);

OAI221xp5_ASAP7_75t_L g11086 ( 
.A1(n_9702),
.A2(n_8881),
.B1(n_8112),
.B2(n_8875),
.C(n_8855),
.Y(n_11086)
);

AOI221xp5_ASAP7_75t_SL g11087 ( 
.A1(n_10359),
.A2(n_7731),
.B1(n_7251),
.B2(n_7368),
.C(n_7307),
.Y(n_11087)
);

OAI211xp5_ASAP7_75t_L g11088 ( 
.A1(n_10363),
.A2(n_8710),
.B(n_8658),
.C(n_8775),
.Y(n_11088)
);

AND2x4_ASAP7_75t_L g11089 ( 
.A(n_9901),
.B(n_9032),
.Y(n_11089)
);

AOI22xp33_ASAP7_75t_L g11090 ( 
.A1(n_9706),
.A2(n_9719),
.B1(n_9725),
.B2(n_9711),
.Y(n_11090)
);

AOI22xp33_ASAP7_75t_L g11091 ( 
.A1(n_9706),
.A2(n_7913),
.B1(n_8421),
.B2(n_8406),
.Y(n_11091)
);

NOR2xp33_ASAP7_75t_L g11092 ( 
.A(n_9608),
.B(n_6223),
.Y(n_11092)
);

AOI22xp33_ASAP7_75t_L g11093 ( 
.A1(n_9711),
.A2(n_8421),
.B1(n_8494),
.B2(n_8406),
.Y(n_11093)
);

BUFx3_ASAP7_75t_L g11094 ( 
.A(n_9555),
.Y(n_11094)
);

AOI22xp33_ASAP7_75t_L g11095 ( 
.A1(n_9719),
.A2(n_8421),
.B1(n_8494),
.B2(n_8406),
.Y(n_11095)
);

AO21x2_ASAP7_75t_L g11096 ( 
.A1(n_9725),
.A2(n_8827),
.B(n_8824),
.Y(n_11096)
);

OAI22xp33_ASAP7_75t_L g11097 ( 
.A1(n_10223),
.A2(n_7870),
.B1(n_7825),
.B2(n_7914),
.Y(n_11097)
);

AOI22xp33_ASAP7_75t_L g11098 ( 
.A1(n_9468),
.A2(n_8421),
.B1(n_8494),
.B2(n_8406),
.Y(n_11098)
);

INVx2_ASAP7_75t_L g11099 ( 
.A(n_10412),
.Y(n_11099)
);

OAI22xp5_ASAP7_75t_L g11100 ( 
.A1(n_10223),
.A2(n_7334),
.B1(n_7362),
.B2(n_7161),
.Y(n_11100)
);

INVx2_ASAP7_75t_L g11101 ( 
.A(n_10412),
.Y(n_11101)
);

AOI22xp33_ASAP7_75t_L g11102 ( 
.A1(n_9468),
.A2(n_9470),
.B1(n_9488),
.B2(n_9479),
.Y(n_11102)
);

NAND3xp33_ASAP7_75t_L g11103 ( 
.A(n_10221),
.B(n_9167),
.C(n_9152),
.Y(n_11103)
);

AOI22xp33_ASAP7_75t_SL g11104 ( 
.A1(n_10173),
.A2(n_7353),
.B1(n_7342),
.B2(n_8775),
.Y(n_11104)
);

AOI22xp33_ASAP7_75t_L g11105 ( 
.A1(n_9470),
.A2(n_8421),
.B1(n_8494),
.B2(n_8406),
.Y(n_11105)
);

INVx1_ASAP7_75t_L g11106 ( 
.A(n_9693),
.Y(n_11106)
);

INVx1_ASAP7_75t_L g11107 ( 
.A(n_9694),
.Y(n_11107)
);

AOI22xp5_ASAP7_75t_L g11108 ( 
.A1(n_10220),
.A2(n_9619),
.B1(n_9488),
.B2(n_9491),
.Y(n_11108)
);

OAI22xp5_ASAP7_75t_L g11109 ( 
.A1(n_10241),
.A2(n_7334),
.B1(n_7362),
.B2(n_7161),
.Y(n_11109)
);

AOI22xp33_ASAP7_75t_L g11110 ( 
.A1(n_9479),
.A2(n_8494),
.B1(n_8518),
.B2(n_8421),
.Y(n_11110)
);

AOI22xp5_ASAP7_75t_L g11111 ( 
.A1(n_10220),
.A2(n_9619),
.B1(n_9501),
.B2(n_9503),
.Y(n_11111)
);

AOI22xp33_ASAP7_75t_L g11112 ( 
.A1(n_9491),
.A2(n_8518),
.B1(n_8556),
.B2(n_8494),
.Y(n_11112)
);

OA21x2_ASAP7_75t_L g11113 ( 
.A1(n_9443),
.A2(n_8832),
.B(n_8827),
.Y(n_11113)
);

NOR2x1_ASAP7_75t_L g11114 ( 
.A(n_10052),
.B(n_9032),
.Y(n_11114)
);

INVx2_ASAP7_75t_L g11115 ( 
.A(n_10365),
.Y(n_11115)
);

OAI211xp5_ASAP7_75t_L g11116 ( 
.A1(n_9551),
.A2(n_8710),
.B(n_8658),
.C(n_8857),
.Y(n_11116)
);

AOI33xp33_ASAP7_75t_L g11117 ( 
.A1(n_9766),
.A2(n_9773),
.A3(n_9551),
.B1(n_10146),
.B2(n_10135),
.B3(n_9619),
.Y(n_11117)
);

OAI22xp5_ASAP7_75t_L g11118 ( 
.A1(n_10241),
.A2(n_7429),
.B1(n_7596),
.B2(n_7161),
.Y(n_11118)
);

OAI22xp33_ASAP7_75t_L g11119 ( 
.A1(n_10241),
.A2(n_10258),
.B1(n_10281),
.B2(n_10248),
.Y(n_11119)
);

INVx1_ASAP7_75t_L g11120 ( 
.A(n_9695),
.Y(n_11120)
);

OAI211xp5_ASAP7_75t_L g11121 ( 
.A1(n_9825),
.A2(n_8934),
.B(n_8857),
.C(n_8945),
.Y(n_11121)
);

OR2x2_ASAP7_75t_L g11122 ( 
.A(n_9595),
.B(n_8192),
.Y(n_11122)
);

AOI22xp33_ASAP7_75t_SL g11123 ( 
.A1(n_10248),
.A2(n_7353),
.B1(n_7342),
.B2(n_8857),
.Y(n_11123)
);

OR2x2_ASAP7_75t_L g11124 ( 
.A(n_9595),
.B(n_7947),
.Y(n_11124)
);

AOI221xp5_ASAP7_75t_L g11125 ( 
.A1(n_9501),
.A2(n_9333),
.B1(n_9354),
.B2(n_9330),
.C(n_9327),
.Y(n_11125)
);

OAI211xp5_ASAP7_75t_L g11126 ( 
.A1(n_9825),
.A2(n_8934),
.B(n_8857),
.C(n_8945),
.Y(n_11126)
);

AND2x4_ASAP7_75t_L g11127 ( 
.A(n_10257),
.B(n_9032),
.Y(n_11127)
);

HB1xp67_ASAP7_75t_L g11128 ( 
.A(n_10245),
.Y(n_11128)
);

AOI22xp33_ASAP7_75t_L g11129 ( 
.A1(n_9503),
.A2(n_8556),
.B1(n_8605),
.B2(n_8518),
.Y(n_11129)
);

OAI221xp5_ASAP7_75t_L g11130 ( 
.A1(n_9504),
.A2(n_8879),
.B1(n_8810),
.B2(n_8912),
.C(n_8907),
.Y(n_11130)
);

AND2x2_ASAP7_75t_L g11131 ( 
.A(n_9766),
.B(n_9055),
.Y(n_11131)
);

INVx2_ASAP7_75t_L g11132 ( 
.A(n_10365),
.Y(n_11132)
);

OR2x2_ASAP7_75t_L g11133 ( 
.A(n_9631),
.B(n_7947),
.Y(n_11133)
);

INVx2_ASAP7_75t_L g11134 ( 
.A(n_10377),
.Y(n_11134)
);

OAI22xp5_ASAP7_75t_L g11135 ( 
.A1(n_10248),
.A2(n_7429),
.B1(n_7596),
.B2(n_7161),
.Y(n_11135)
);

AOI22xp33_ASAP7_75t_SL g11136 ( 
.A1(n_10258),
.A2(n_7353),
.B1(n_7342),
.B2(n_8934),
.Y(n_11136)
);

A2O1A1Ixp33_ASAP7_75t_L g11137 ( 
.A1(n_9942),
.A2(n_8921),
.B(n_7275),
.C(n_7238),
.Y(n_11137)
);

AOI221xp5_ASAP7_75t_L g11138 ( 
.A1(n_9504),
.A2(n_9361),
.B1(n_9381),
.B2(n_9354),
.C(n_9333),
.Y(n_11138)
);

OAI22xp33_ASAP7_75t_L g11139 ( 
.A1(n_10258),
.A2(n_8163),
.B1(n_8254),
.B2(n_7914),
.Y(n_11139)
);

BUFx3_ASAP7_75t_L g11140 ( 
.A(n_9555),
.Y(n_11140)
);

AOI22xp5_ASAP7_75t_L g11141 ( 
.A1(n_10281),
.A2(n_8019),
.B1(n_8224),
.B2(n_8209),
.Y(n_11141)
);

OAI22xp5_ASAP7_75t_L g11142 ( 
.A1(n_10281),
.A2(n_7596),
.B1(n_7655),
.B2(n_7429),
.Y(n_11142)
);

AND2x2_ASAP7_75t_L g11143 ( 
.A(n_9773),
.B(n_9055),
.Y(n_11143)
);

AOI22xp33_ASAP7_75t_L g11144 ( 
.A1(n_10380),
.A2(n_8556),
.B1(n_8605),
.B2(n_8518),
.Y(n_11144)
);

INVx1_ASAP7_75t_L g11145 ( 
.A(n_9698),
.Y(n_11145)
);

AOI22xp5_ASAP7_75t_L g11146 ( 
.A1(n_10319),
.A2(n_8019),
.B1(n_8224),
.B2(n_8209),
.Y(n_11146)
);

OAI211xp5_ASAP7_75t_L g11147 ( 
.A1(n_9825),
.A2(n_8934),
.B(n_9176),
.C(n_8945),
.Y(n_11147)
);

OAI211xp5_ASAP7_75t_SL g11148 ( 
.A1(n_10113),
.A2(n_7307),
.B(n_7368),
.C(n_7184),
.Y(n_11148)
);

AOI22xp33_ASAP7_75t_SL g11149 ( 
.A1(n_10319),
.A2(n_9176),
.B1(n_9294),
.B2(n_8945),
.Y(n_11149)
);

O2A1O1Ixp33_ASAP7_75t_L g11150 ( 
.A1(n_10249),
.A2(n_9419),
.B(n_9075),
.C(n_9096),
.Y(n_11150)
);

INVx1_ASAP7_75t_L g11151 ( 
.A(n_9700),
.Y(n_11151)
);

AOI221xp5_ASAP7_75t_L g11152 ( 
.A1(n_10380),
.A2(n_9361),
.B1(n_9381),
.B2(n_9354),
.C(n_9333),
.Y(n_11152)
);

OAI22xp5_ASAP7_75t_L g11153 ( 
.A1(n_10319),
.A2(n_10350),
.B1(n_10336),
.B2(n_9877),
.Y(n_11153)
);

BUFx3_ASAP7_75t_L g11154 ( 
.A(n_9555),
.Y(n_11154)
);

AND2x2_ASAP7_75t_L g11155 ( 
.A(n_9877),
.B(n_9055),
.Y(n_11155)
);

AND2x2_ASAP7_75t_L g11156 ( 
.A(n_9877),
.B(n_9059),
.Y(n_11156)
);

INVx2_ASAP7_75t_L g11157 ( 
.A(n_10377),
.Y(n_11157)
);

AOI22xp33_ASAP7_75t_SL g11158 ( 
.A1(n_10336),
.A2(n_9294),
.B1(n_9322),
.B2(n_9176),
.Y(n_11158)
);

INVx5_ASAP7_75t_L g11159 ( 
.A(n_9556),
.Y(n_11159)
);

INVx1_ASAP7_75t_L g11160 ( 
.A(n_9705),
.Y(n_11160)
);

OR2x2_ASAP7_75t_L g11161 ( 
.A(n_9631),
.B(n_7948),
.Y(n_11161)
);

INVxp67_ASAP7_75t_SL g11162 ( 
.A(n_9556),
.Y(n_11162)
);

AOI222xp33_ASAP7_75t_L g11163 ( 
.A1(n_10382),
.A2(n_9395),
.B1(n_9381),
.B2(n_9398),
.C1(n_9382),
.C2(n_9361),
.Y(n_11163)
);

AND2x4_ASAP7_75t_L g11164 ( 
.A(n_10257),
.B(n_9059),
.Y(n_11164)
);

AOI22xp5_ASAP7_75t_L g11165 ( 
.A1(n_10336),
.A2(n_8224),
.B1(n_8209),
.B2(n_7772),
.Y(n_11165)
);

BUFx2_ASAP7_75t_L g11166 ( 
.A(n_9556),
.Y(n_11166)
);

OAI21xp33_ASAP7_75t_L g11167 ( 
.A1(n_9792),
.A2(n_8868),
.B(n_7431),
.Y(n_11167)
);

OAI211xp5_ASAP7_75t_L g11168 ( 
.A1(n_10253),
.A2(n_10293),
.B(n_10332),
.C(n_10271),
.Y(n_11168)
);

INVx2_ASAP7_75t_L g11169 ( 
.A(n_9882),
.Y(n_11169)
);

OAI21x1_ASAP7_75t_L g11170 ( 
.A1(n_9443),
.A2(n_9379),
.B(n_9373),
.Y(n_11170)
);

INVx1_ASAP7_75t_L g11171 ( 
.A(n_9710),
.Y(n_11171)
);

OAI22xp33_ASAP7_75t_L g11172 ( 
.A1(n_10350),
.A2(n_8163),
.B1(n_8254),
.B2(n_7914),
.Y(n_11172)
);

INVx3_ASAP7_75t_L g11173 ( 
.A(n_9556),
.Y(n_11173)
);

AOI22xp33_ASAP7_75t_L g11174 ( 
.A1(n_10382),
.A2(n_8556),
.B1(n_8605),
.B2(n_8518),
.Y(n_11174)
);

AOI22xp5_ASAP7_75t_L g11175 ( 
.A1(n_10350),
.A2(n_8224),
.B1(n_8209),
.B2(n_7772),
.Y(n_11175)
);

OAI21xp33_ASAP7_75t_L g11176 ( 
.A1(n_9841),
.A2(n_8868),
.B(n_7431),
.Y(n_11176)
);

AND2x2_ASAP7_75t_L g11177 ( 
.A(n_9915),
.B(n_9059),
.Y(n_11177)
);

CKINVDCx5p33_ASAP7_75t_R g11178 ( 
.A(n_9640),
.Y(n_11178)
);

INVx2_ASAP7_75t_L g11179 ( 
.A(n_9882),
.Y(n_11179)
);

OR2x2_ASAP7_75t_L g11180 ( 
.A(n_9677),
.B(n_7948),
.Y(n_11180)
);

INVx2_ASAP7_75t_L g11181 ( 
.A(n_9884),
.Y(n_11181)
);

AND2x4_ASAP7_75t_L g11182 ( 
.A(n_10257),
.B(n_8929),
.Y(n_11182)
);

AOI22xp33_ASAP7_75t_L g11183 ( 
.A1(n_10388),
.A2(n_10409),
.B1(n_10410),
.B2(n_10400),
.Y(n_11183)
);

AOI22xp33_ASAP7_75t_L g11184 ( 
.A1(n_10388),
.A2(n_8556),
.B1(n_8605),
.B2(n_8518),
.Y(n_11184)
);

AOI22xp33_ASAP7_75t_L g11185 ( 
.A1(n_10400),
.A2(n_8605),
.B1(n_8649),
.B2(n_8556),
.Y(n_11185)
);

AOI22xp33_ASAP7_75t_L g11186 ( 
.A1(n_10409),
.A2(n_8649),
.B1(n_8661),
.B2(n_8605),
.Y(n_11186)
);

AOI21xp5_ASAP7_75t_L g11187 ( 
.A1(n_10135),
.A2(n_7405),
.B(n_9176),
.Y(n_11187)
);

OAI22xp5_ASAP7_75t_L g11188 ( 
.A1(n_9915),
.A2(n_9936),
.B1(n_9992),
.B2(n_9689),
.Y(n_11188)
);

NAND2xp5_ASAP7_75t_L g11189 ( 
.A(n_10273),
.B(n_9061),
.Y(n_11189)
);

AND2x2_ASAP7_75t_L g11190 ( 
.A(n_9915),
.B(n_8976),
.Y(n_11190)
);

OAI22xp5_ASAP7_75t_L g11191 ( 
.A1(n_9936),
.A2(n_7596),
.B1(n_7655),
.B2(n_7429),
.Y(n_11191)
);

INVx3_ASAP7_75t_L g11192 ( 
.A(n_9603),
.Y(n_11192)
);

BUFx3_ASAP7_75t_L g11193 ( 
.A(n_9603),
.Y(n_11193)
);

OAI21xp33_ASAP7_75t_SL g11194 ( 
.A1(n_9927),
.A2(n_10074),
.B(n_10022),
.Y(n_11194)
);

NAND2xp5_ASAP7_75t_L g11195 ( 
.A(n_10273),
.B(n_9111),
.Y(n_11195)
);

OAI22xp33_ASAP7_75t_L g11196 ( 
.A1(n_10410),
.A2(n_8254),
.B1(n_8163),
.B2(n_7200),
.Y(n_11196)
);

OAI22xp33_ASAP7_75t_L g11197 ( 
.A1(n_9746),
.A2(n_8254),
.B1(n_8163),
.B2(n_7200),
.Y(n_11197)
);

AOI211xp5_ASAP7_75t_L g11198 ( 
.A1(n_9447),
.A2(n_7238),
.B(n_7241),
.C(n_7483),
.Y(n_11198)
);

OAI22xp5_ASAP7_75t_L g11199 ( 
.A1(n_9936),
.A2(n_7596),
.B1(n_7655),
.B2(n_7429),
.Y(n_11199)
);

NOR2xp33_ASAP7_75t_L g11200 ( 
.A(n_9603),
.B(n_6867),
.Y(n_11200)
);

AOI22xp33_ASAP7_75t_L g11201 ( 
.A1(n_9746),
.A2(n_8661),
.B1(n_8679),
.B2(n_8649),
.Y(n_11201)
);

OAI221xp5_ASAP7_75t_L g11202 ( 
.A1(n_9750),
.A2(n_8912),
.B1(n_8907),
.B2(n_9322),
.C(n_9294),
.Y(n_11202)
);

AOI22xp33_ASAP7_75t_L g11203 ( 
.A1(n_9750),
.A2(n_8661),
.B1(n_8679),
.B2(n_8649),
.Y(n_11203)
);

INVx3_ASAP7_75t_L g11204 ( 
.A(n_9603),
.Y(n_11204)
);

OAI22xp5_ASAP7_75t_L g11205 ( 
.A1(n_9992),
.A2(n_7666),
.B1(n_7901),
.B2(n_7655),
.Y(n_11205)
);

OAI221xp5_ASAP7_75t_SL g11206 ( 
.A1(n_9884),
.A2(n_7826),
.B1(n_7801),
.B2(n_8283),
.C(n_8231),
.Y(n_11206)
);

OAI22xp5_ASAP7_75t_L g11207 ( 
.A1(n_9992),
.A2(n_7666),
.B1(n_7901),
.B2(n_7655),
.Y(n_11207)
);

AOI22xp33_ASAP7_75t_L g11208 ( 
.A1(n_9764),
.A2(n_8661),
.B1(n_8679),
.B2(n_8649),
.Y(n_11208)
);

OAI211xp5_ASAP7_75t_L g11209 ( 
.A1(n_9447),
.A2(n_9322),
.B(n_9341),
.C(n_9294),
.Y(n_11209)
);

AOI22xp33_ASAP7_75t_SL g11210 ( 
.A1(n_9764),
.A2(n_9341),
.B1(n_9363),
.B2(n_9322),
.Y(n_11210)
);

INVx1_ASAP7_75t_L g11211 ( 
.A(n_9712),
.Y(n_11211)
);

OAI22xp5_ASAP7_75t_L g11212 ( 
.A1(n_9677),
.A2(n_7901),
.B1(n_7666),
.B2(n_9038),
.Y(n_11212)
);

OAI221xp5_ASAP7_75t_L g11213 ( 
.A1(n_9767),
.A2(n_9782),
.B1(n_9783),
.B2(n_9776),
.C(n_9774),
.Y(n_11213)
);

INVx1_ASAP7_75t_L g11214 ( 
.A(n_9717),
.Y(n_11214)
);

CKINVDCx20_ASAP7_75t_R g11215 ( 
.A(n_10316),
.Y(n_11215)
);

AOI211xp5_ASAP7_75t_L g11216 ( 
.A1(n_9624),
.A2(n_7238),
.B(n_7241),
.C(n_7483),
.Y(n_11216)
);

AOI22xp33_ASAP7_75t_L g11217 ( 
.A1(n_9767),
.A2(n_8661),
.B1(n_8679),
.B2(n_8649),
.Y(n_11217)
);

INVx1_ASAP7_75t_L g11218 ( 
.A(n_9722),
.Y(n_11218)
);

OAI211xp5_ASAP7_75t_SL g11219 ( 
.A1(n_10113),
.A2(n_10122),
.B(n_10154),
.C(n_10121),
.Y(n_11219)
);

INVx1_ASAP7_75t_L g11220 ( 
.A(n_9726),
.Y(n_11220)
);

AOI22xp33_ASAP7_75t_SL g11221 ( 
.A1(n_9774),
.A2(n_9363),
.B1(n_9376),
.B2(n_9341),
.Y(n_11221)
);

A2O1A1Ixp33_ASAP7_75t_L g11222 ( 
.A1(n_10381),
.A2(n_8921),
.B(n_7959),
.C(n_7483),
.Y(n_11222)
);

AOI22xp33_ASAP7_75t_L g11223 ( 
.A1(n_9776),
.A2(n_8679),
.B1(n_8715),
.B2(n_8661),
.Y(n_11223)
);

AND2x2_ASAP7_75t_L g11224 ( 
.A(n_9927),
.B(n_8976),
.Y(n_11224)
);

OAI22xp5_ASAP7_75t_L g11225 ( 
.A1(n_9689),
.A2(n_7901),
.B1(n_7666),
.B2(n_9038),
.Y(n_11225)
);

BUFx6f_ASAP7_75t_L g11226 ( 
.A(n_9634),
.Y(n_11226)
);

HB1xp67_ASAP7_75t_L g11227 ( 
.A(n_9730),
.Y(n_11227)
);

AOI221xp5_ASAP7_75t_L g11228 ( 
.A1(n_9782),
.A2(n_9790),
.B1(n_9793),
.B2(n_9784),
.C(n_9783),
.Y(n_11228)
);

AOI22xp33_ASAP7_75t_L g11229 ( 
.A1(n_9784),
.A2(n_8715),
.B1(n_8717),
.B2(n_8679),
.Y(n_11229)
);

CKINVDCx5p33_ASAP7_75t_R g11230 ( 
.A(n_10324),
.Y(n_11230)
);

AND2x2_ASAP7_75t_L g11231 ( 
.A(n_10022),
.B(n_8976),
.Y(n_11231)
);

INVx1_ASAP7_75t_L g11232 ( 
.A(n_9734),
.Y(n_11232)
);

AOI21xp33_ASAP7_75t_L g11233 ( 
.A1(n_10212),
.A2(n_7220),
.B(n_7181),
.Y(n_11233)
);

INVx1_ASAP7_75t_L g11234 ( 
.A(n_11227),
.Y(n_11234)
);

AND2x2_ASAP7_75t_L g11235 ( 
.A(n_10437),
.B(n_9634),
.Y(n_11235)
);

INVx2_ASAP7_75t_L g11236 ( 
.A(n_10529),
.Y(n_11236)
);

OR2x2_ASAP7_75t_L g11237 ( 
.A(n_10428),
.B(n_9546),
.Y(n_11237)
);

INVx1_ASAP7_75t_L g11238 ( 
.A(n_10485),
.Y(n_11238)
);

INVx2_ASAP7_75t_L g11239 ( 
.A(n_10926),
.Y(n_11239)
);

AND2x4_ASAP7_75t_SL g11240 ( 
.A(n_10808),
.B(n_6965),
.Y(n_11240)
);

INVxp67_ASAP7_75t_SL g11241 ( 
.A(n_10544),
.Y(n_11241)
);

AND2x2_ASAP7_75t_L g11242 ( 
.A(n_11008),
.B(n_9634),
.Y(n_11242)
);

AND2x2_ASAP7_75t_L g11243 ( 
.A(n_10982),
.B(n_9634),
.Y(n_11243)
);

AND2x2_ASAP7_75t_L g11244 ( 
.A(n_10918),
.B(n_9686),
.Y(n_11244)
);

INVx2_ASAP7_75t_L g11245 ( 
.A(n_10950),
.Y(n_11245)
);

INVx1_ASAP7_75t_L g11246 ( 
.A(n_10502),
.Y(n_11246)
);

OR2x2_ASAP7_75t_L g11247 ( 
.A(n_10520),
.B(n_9546),
.Y(n_11247)
);

NAND2xp5_ASAP7_75t_L g11248 ( 
.A(n_10421),
.B(n_10570),
.Y(n_11248)
);

NAND2xp5_ASAP7_75t_L g11249 ( 
.A(n_10863),
.B(n_9686),
.Y(n_11249)
);

HB1xp67_ASAP7_75t_L g11250 ( 
.A(n_11009),
.Y(n_11250)
);

OR2x2_ASAP7_75t_L g11251 ( 
.A(n_10420),
.B(n_9617),
.Y(n_11251)
);

AND2x2_ASAP7_75t_L g11252 ( 
.A(n_10582),
.B(n_9686),
.Y(n_11252)
);

INVx2_ASAP7_75t_L g11253 ( 
.A(n_10972),
.Y(n_11253)
);

BUFx3_ASAP7_75t_L g11254 ( 
.A(n_10612),
.Y(n_11254)
);

INVx2_ASAP7_75t_L g11255 ( 
.A(n_10644),
.Y(n_11255)
);

INVxp67_ASAP7_75t_L g11256 ( 
.A(n_10739),
.Y(n_11256)
);

INVx1_ASAP7_75t_L g11257 ( 
.A(n_10433),
.Y(n_11257)
);

AND2x2_ASAP7_75t_L g11258 ( 
.A(n_10642),
.B(n_9686),
.Y(n_11258)
);

BUFx3_ASAP7_75t_L g11259 ( 
.A(n_10443),
.Y(n_11259)
);

INVxp67_ASAP7_75t_L g11260 ( 
.A(n_10531),
.Y(n_11260)
);

AND2x2_ASAP7_75t_L g11261 ( 
.A(n_10717),
.B(n_10649),
.Y(n_11261)
);

OR2x2_ASAP7_75t_L g11262 ( 
.A(n_10418),
.B(n_9617),
.Y(n_11262)
);

OR2x6_ASAP7_75t_L g11263 ( 
.A(n_10453),
.B(n_9878),
.Y(n_11263)
);

OR2x2_ASAP7_75t_L g11264 ( 
.A(n_10422),
.B(n_10466),
.Y(n_11264)
);

NOR2xp67_ASAP7_75t_L g11265 ( 
.A(n_10431),
.B(n_10146),
.Y(n_11265)
);

HB1xp67_ASAP7_75t_L g11266 ( 
.A(n_10790),
.Y(n_11266)
);

INVx2_ASAP7_75t_L g11267 ( 
.A(n_10543),
.Y(n_11267)
);

AND2x2_ASAP7_75t_L g11268 ( 
.A(n_10649),
.B(n_9664),
.Y(n_11268)
);

AND2x2_ASAP7_75t_L g11269 ( 
.A(n_10721),
.B(n_9675),
.Y(n_11269)
);

INVx2_ASAP7_75t_L g11270 ( 
.A(n_11052),
.Y(n_11270)
);

AND2x2_ASAP7_75t_L g11271 ( 
.A(n_10721),
.B(n_10766),
.Y(n_11271)
);

INVx1_ASAP7_75t_L g11272 ( 
.A(n_10438),
.Y(n_11272)
);

AND2x4_ASAP7_75t_L g11273 ( 
.A(n_10939),
.B(n_10807),
.Y(n_11273)
);

NOR2xp33_ASAP7_75t_L g11274 ( 
.A(n_10638),
.B(n_9691),
.Y(n_11274)
);

HB1xp67_ASAP7_75t_L g11275 ( 
.A(n_10815),
.Y(n_11275)
);

OR2x6_ASAP7_75t_L g11276 ( 
.A(n_10453),
.B(n_9878),
.Y(n_11276)
);

BUFx3_ASAP7_75t_L g11277 ( 
.A(n_10445),
.Y(n_11277)
);

AND2x2_ASAP7_75t_L g11278 ( 
.A(n_10766),
.B(n_9692),
.Y(n_11278)
);

NAND2xp5_ASAP7_75t_L g11279 ( 
.A(n_10490),
.B(n_10273),
.Y(n_11279)
);

INVx1_ASAP7_75t_L g11280 ( 
.A(n_10447),
.Y(n_11280)
);

INVx2_ASAP7_75t_L g11281 ( 
.A(n_11064),
.Y(n_11281)
);

AND2x2_ASAP7_75t_L g11282 ( 
.A(n_10770),
.B(n_9731),
.Y(n_11282)
);

INVx2_ASAP7_75t_L g11283 ( 
.A(n_11060),
.Y(n_11283)
);

INVx1_ASAP7_75t_SL g11284 ( 
.A(n_10639),
.Y(n_11284)
);

OR2x2_ASAP7_75t_L g11285 ( 
.A(n_10930),
.B(n_9789),
.Y(n_11285)
);

BUFx3_ASAP7_75t_L g11286 ( 
.A(n_11215),
.Y(n_11286)
);

HB1xp67_ASAP7_75t_L g11287 ( 
.A(n_10653),
.Y(n_11287)
);

INVx2_ASAP7_75t_L g11288 ( 
.A(n_11060),
.Y(n_11288)
);

BUFx2_ASAP7_75t_L g11289 ( 
.A(n_11028),
.Y(n_11289)
);

NAND3xp33_ASAP7_75t_L g11290 ( 
.A(n_10426),
.B(n_10126),
.C(n_10072),
.Y(n_11290)
);

AND2x4_ASAP7_75t_SL g11291 ( 
.A(n_10509),
.B(n_9493),
.Y(n_11291)
);

BUFx3_ASAP7_75t_L g11292 ( 
.A(n_10880),
.Y(n_11292)
);

INVx2_ASAP7_75t_SL g11293 ( 
.A(n_10628),
.Y(n_11293)
);

INVx1_ASAP7_75t_L g11294 ( 
.A(n_10462),
.Y(n_11294)
);

INVx1_ASAP7_75t_L g11295 ( 
.A(n_10468),
.Y(n_11295)
);

INVx2_ASAP7_75t_L g11296 ( 
.A(n_11060),
.Y(n_11296)
);

INVx5_ASAP7_75t_L g11297 ( 
.A(n_10491),
.Y(n_11297)
);

HB1xp67_ASAP7_75t_L g11298 ( 
.A(n_10788),
.Y(n_11298)
);

AND2x2_ASAP7_75t_L g11299 ( 
.A(n_10770),
.B(n_9765),
.Y(n_11299)
);

INVx1_ASAP7_75t_L g11300 ( 
.A(n_10470),
.Y(n_11300)
);

INVx2_ASAP7_75t_L g11301 ( 
.A(n_11078),
.Y(n_11301)
);

INVx3_ASAP7_75t_L g11302 ( 
.A(n_10780),
.Y(n_11302)
);

HB1xp67_ASAP7_75t_L g11303 ( 
.A(n_10414),
.Y(n_11303)
);

HB1xp67_ASAP7_75t_L g11304 ( 
.A(n_10641),
.Y(n_11304)
);

OR2x6_ASAP7_75t_L g11305 ( 
.A(n_10823),
.B(n_9878),
.Y(n_11305)
);

AND2x2_ASAP7_75t_L g11306 ( 
.A(n_10899),
.B(n_9791),
.Y(n_11306)
);

AND2x2_ASAP7_75t_L g11307 ( 
.A(n_10899),
.B(n_9808),
.Y(n_11307)
);

AND2x2_ASAP7_75t_L g11308 ( 
.A(n_11131),
.B(n_10052),
.Y(n_11308)
);

INVxp67_ASAP7_75t_L g11309 ( 
.A(n_10499),
.Y(n_11309)
);

OR2x2_ASAP7_75t_L g11310 ( 
.A(n_11031),
.B(n_9789),
.Y(n_11310)
);

INVx3_ASAP7_75t_L g11311 ( 
.A(n_10491),
.Y(n_11311)
);

AND2x2_ASAP7_75t_L g11312 ( 
.A(n_11143),
.B(n_9493),
.Y(n_11312)
);

INVx2_ASAP7_75t_L g11313 ( 
.A(n_11078),
.Y(n_11313)
);

INVx1_ASAP7_75t_L g11314 ( 
.A(n_10478),
.Y(n_11314)
);

AND2x4_ASAP7_75t_L g11315 ( 
.A(n_10807),
.B(n_9534),
.Y(n_11315)
);

AND2x2_ASAP7_75t_L g11316 ( 
.A(n_10524),
.B(n_9534),
.Y(n_11316)
);

INVx1_ASAP7_75t_L g11317 ( 
.A(n_10493),
.Y(n_11317)
);

INVx3_ASAP7_75t_L g11318 ( 
.A(n_10491),
.Y(n_11318)
);

INVx2_ASAP7_75t_SL g11319 ( 
.A(n_10628),
.Y(n_11319)
);

INVx1_ASAP7_75t_SL g11320 ( 
.A(n_10694),
.Y(n_11320)
);

BUFx3_ASAP7_75t_L g11321 ( 
.A(n_10509),
.Y(n_11321)
);

AND2x2_ASAP7_75t_L g11322 ( 
.A(n_10545),
.B(n_9820),
.Y(n_11322)
);

AND2x2_ASAP7_75t_L g11323 ( 
.A(n_10545),
.B(n_9820),
.Y(n_11323)
);

INVx2_ASAP7_75t_L g11324 ( 
.A(n_11078),
.Y(n_11324)
);

BUFx6f_ASAP7_75t_L g11325 ( 
.A(n_10509),
.Y(n_11325)
);

AND2x2_ASAP7_75t_L g11326 ( 
.A(n_10446),
.B(n_9835),
.Y(n_11326)
);

BUFx2_ASAP7_75t_L g11327 ( 
.A(n_10931),
.Y(n_11327)
);

BUFx3_ASAP7_75t_L g11328 ( 
.A(n_10546),
.Y(n_11328)
);

NAND2xp5_ASAP7_75t_L g11329 ( 
.A(n_10701),
.B(n_9835),
.Y(n_11329)
);

AND2x2_ASAP7_75t_L g11330 ( 
.A(n_10474),
.B(n_9852),
.Y(n_11330)
);

INVx1_ASAP7_75t_L g11331 ( 
.A(n_10504),
.Y(n_11331)
);

INVx2_ASAP7_75t_L g11332 ( 
.A(n_11226),
.Y(n_11332)
);

NAND2xp5_ASAP7_75t_L g11333 ( 
.A(n_10471),
.B(n_9852),
.Y(n_11333)
);

INVx1_ASAP7_75t_SL g11334 ( 
.A(n_10784),
.Y(n_11334)
);

INVx1_ASAP7_75t_L g11335 ( 
.A(n_10522),
.Y(n_11335)
);

AND2x2_ASAP7_75t_L g11336 ( 
.A(n_10540),
.B(n_9909),
.Y(n_11336)
);

HB1xp67_ASAP7_75t_L g11337 ( 
.A(n_10692),
.Y(n_11337)
);

AND2x2_ASAP7_75t_L g11338 ( 
.A(n_10832),
.B(n_9909),
.Y(n_11338)
);

INVx1_ASAP7_75t_L g11339 ( 
.A(n_10547),
.Y(n_11339)
);

INVx1_ASAP7_75t_L g11340 ( 
.A(n_10565),
.Y(n_11340)
);

HB1xp67_ASAP7_75t_L g11341 ( 
.A(n_11071),
.Y(n_11341)
);

AND2x2_ASAP7_75t_L g11342 ( 
.A(n_10465),
.B(n_9918),
.Y(n_11342)
);

AND2x2_ASAP7_75t_L g11343 ( 
.A(n_10569),
.B(n_9918),
.Y(n_11343)
);

BUFx2_ASAP7_75t_L g11344 ( 
.A(n_11037),
.Y(n_11344)
);

BUFx3_ASAP7_75t_L g11345 ( 
.A(n_10546),
.Y(n_11345)
);

INVx2_ASAP7_75t_L g11346 ( 
.A(n_11226),
.Y(n_11346)
);

AND2x2_ASAP7_75t_L g11347 ( 
.A(n_10571),
.B(n_9937),
.Y(n_11347)
);

AND2x2_ASAP7_75t_L g11348 ( 
.A(n_10618),
.B(n_9937),
.Y(n_11348)
);

HB1xp67_ASAP7_75t_L g11349 ( 
.A(n_10783),
.Y(n_11349)
);

AND2x2_ASAP7_75t_L g11350 ( 
.A(n_10625),
.B(n_9943),
.Y(n_11350)
);

INVx3_ASAP7_75t_SL g11351 ( 
.A(n_10687),
.Y(n_11351)
);

AND2x2_ASAP7_75t_L g11352 ( 
.A(n_10650),
.B(n_9943),
.Y(n_11352)
);

AND2x2_ASAP7_75t_L g11353 ( 
.A(n_10883),
.B(n_9972),
.Y(n_11353)
);

INVx2_ASAP7_75t_L g11354 ( 
.A(n_11226),
.Y(n_11354)
);

INVx2_ASAP7_75t_L g11355 ( 
.A(n_10572),
.Y(n_11355)
);

AND2x2_ASAP7_75t_L g11356 ( 
.A(n_10914),
.B(n_9972),
.Y(n_11356)
);

OR2x2_ASAP7_75t_L g11357 ( 
.A(n_10590),
.B(n_10023),
.Y(n_11357)
);

BUFx2_ASAP7_75t_L g11358 ( 
.A(n_10998),
.Y(n_11358)
);

NAND2xp5_ASAP7_75t_L g11359 ( 
.A(n_10854),
.B(n_10934),
.Y(n_11359)
);

AND2x2_ASAP7_75t_L g11360 ( 
.A(n_10945),
.B(n_10962),
.Y(n_11360)
);

AND2x2_ASAP7_75t_L g11361 ( 
.A(n_11006),
.B(n_10023),
.Y(n_11361)
);

INVx1_ASAP7_75t_L g11362 ( 
.A(n_10935),
.Y(n_11362)
);

AND2x2_ASAP7_75t_L g11363 ( 
.A(n_11016),
.B(n_10051),
.Y(n_11363)
);

INVx2_ASAP7_75t_L g11364 ( 
.A(n_10572),
.Y(n_11364)
);

AND2x2_ASAP7_75t_L g11365 ( 
.A(n_11059),
.B(n_10051),
.Y(n_11365)
);

INVx2_ASAP7_75t_L g11366 ( 
.A(n_10589),
.Y(n_11366)
);

INVx1_ASAP7_75t_L g11367 ( 
.A(n_11038),
.Y(n_11367)
);

OR2x2_ASAP7_75t_L g11368 ( 
.A(n_10631),
.B(n_9737),
.Y(n_11368)
);

NOR2xp33_ASAP7_75t_L g11369 ( 
.A(n_10546),
.B(n_10019),
.Y(n_11369)
);

INVx1_ASAP7_75t_L g11370 ( 
.A(n_11067),
.Y(n_11370)
);

AND2x2_ASAP7_75t_L g11371 ( 
.A(n_10560),
.B(n_8976),
.Y(n_11371)
);

BUFx2_ASAP7_75t_L g11372 ( 
.A(n_10441),
.Y(n_11372)
);

INVxp67_ASAP7_75t_SL g11373 ( 
.A(n_10497),
.Y(n_11373)
);

AND2x2_ASAP7_75t_L g11374 ( 
.A(n_10662),
.B(n_10668),
.Y(n_11374)
);

NOR2x1_ASAP7_75t_L g11375 ( 
.A(n_10627),
.B(n_10039),
.Y(n_11375)
);

INVx1_ASAP7_75t_L g11376 ( 
.A(n_11079),
.Y(n_11376)
);

INVx2_ASAP7_75t_L g11377 ( 
.A(n_10589),
.Y(n_11377)
);

INVx1_ASAP7_75t_L g11378 ( 
.A(n_11128),
.Y(n_11378)
);

INVx1_ASAP7_75t_L g11379 ( 
.A(n_10574),
.Y(n_11379)
);

INVx4_ASAP7_75t_SL g11380 ( 
.A(n_10913),
.Y(n_11380)
);

AND2x2_ASAP7_75t_L g11381 ( 
.A(n_10495),
.B(n_9030),
.Y(n_11381)
);

INVx2_ASAP7_75t_SL g11382 ( 
.A(n_11178),
.Y(n_11382)
);

INVx1_ASAP7_75t_L g11383 ( 
.A(n_10580),
.Y(n_11383)
);

INVx3_ASAP7_75t_L g11384 ( 
.A(n_10495),
.Y(n_11384)
);

INVx3_ASAP7_75t_L g11385 ( 
.A(n_10498),
.Y(n_11385)
);

AOI22xp33_ASAP7_75t_L g11386 ( 
.A1(n_10415),
.A2(n_9793),
.B1(n_9798),
.B2(n_9790),
.Y(n_11386)
);

INVx2_ASAP7_75t_L g11387 ( 
.A(n_11094),
.Y(n_11387)
);

OR2x2_ASAP7_75t_L g11388 ( 
.A(n_10779),
.B(n_9739),
.Y(n_11388)
);

INVx1_ASAP7_75t_L g11389 ( 
.A(n_10608),
.Y(n_11389)
);

INVx4_ASAP7_75t_L g11390 ( 
.A(n_10811),
.Y(n_11390)
);

OR2x2_ASAP7_75t_L g11391 ( 
.A(n_10924),
.B(n_9741),
.Y(n_11391)
);

OR2x2_ASAP7_75t_L g11392 ( 
.A(n_10953),
.B(n_9745),
.Y(n_11392)
);

OR2x2_ASAP7_75t_L g11393 ( 
.A(n_10961),
.B(n_9747),
.Y(n_11393)
);

AOI22xp33_ASAP7_75t_L g11394 ( 
.A1(n_10424),
.A2(n_9811),
.B1(n_9818),
.B2(n_9798),
.Y(n_11394)
);

HB1xp67_ASAP7_75t_L g11395 ( 
.A(n_10416),
.Y(n_11395)
);

OR2x2_ASAP7_75t_L g11396 ( 
.A(n_10430),
.B(n_9753),
.Y(n_11396)
);

OR2x2_ASAP7_75t_L g11397 ( 
.A(n_10969),
.B(n_9759),
.Y(n_11397)
);

AND2x2_ASAP7_75t_L g11398 ( 
.A(n_10498),
.B(n_9030),
.Y(n_11398)
);

AND2x2_ASAP7_75t_L g11399 ( 
.A(n_11155),
.B(n_9030),
.Y(n_11399)
);

AND2x2_ASAP7_75t_L g11400 ( 
.A(n_11156),
.B(n_11177),
.Y(n_11400)
);

INVx1_ASAP7_75t_L g11401 ( 
.A(n_10610),
.Y(n_11401)
);

AND2x2_ASAP7_75t_L g11402 ( 
.A(n_10716),
.B(n_10718),
.Y(n_11402)
);

INVx2_ASAP7_75t_L g11403 ( 
.A(n_11140),
.Y(n_11403)
);

INVx1_ASAP7_75t_L g11404 ( 
.A(n_10616),
.Y(n_11404)
);

INVx1_ASAP7_75t_L g11405 ( 
.A(n_10632),
.Y(n_11405)
);

INVx1_ASAP7_75t_L g11406 ( 
.A(n_10671),
.Y(n_11406)
);

INVxp67_ASAP7_75t_L g11407 ( 
.A(n_10796),
.Y(n_11407)
);

AO31x2_ASAP7_75t_L g11408 ( 
.A1(n_10555),
.A2(n_9890),
.A3(n_9898),
.B(n_9886),
.Y(n_11408)
);

INVx1_ASAP7_75t_L g11409 ( 
.A(n_10679),
.Y(n_11409)
);

AND2x2_ASAP7_75t_L g11410 ( 
.A(n_10723),
.B(n_9030),
.Y(n_11410)
);

AND2x2_ASAP7_75t_L g11411 ( 
.A(n_10731),
.B(n_9047),
.Y(n_11411)
);

INVx1_ASAP7_75t_L g11412 ( 
.A(n_10700),
.Y(n_11412)
);

AND2x4_ASAP7_75t_L g11413 ( 
.A(n_10419),
.B(n_8929),
.Y(n_11413)
);

AND2x2_ASAP7_75t_L g11414 ( 
.A(n_10733),
.B(n_9047),
.Y(n_11414)
);

HB1xp67_ASAP7_75t_L g11415 ( 
.A(n_11099),
.Y(n_11415)
);

INVx2_ASAP7_75t_L g11416 ( 
.A(n_11154),
.Y(n_11416)
);

INVx2_ASAP7_75t_L g11417 ( 
.A(n_11193),
.Y(n_11417)
);

INVx2_ASAP7_75t_L g11418 ( 
.A(n_10993),
.Y(n_11418)
);

INVx1_ASAP7_75t_L g11419 ( 
.A(n_10704),
.Y(n_11419)
);

AND2x2_ASAP7_75t_L g11420 ( 
.A(n_10748),
.B(n_9047),
.Y(n_11420)
);

AND2x2_ASAP7_75t_L g11421 ( 
.A(n_10799),
.B(n_9047),
.Y(n_11421)
);

INVx2_ASAP7_75t_SL g11422 ( 
.A(n_11230),
.Y(n_11422)
);

INVx2_ASAP7_75t_L g11423 ( 
.A(n_10993),
.Y(n_11423)
);

INVx2_ASAP7_75t_L g11424 ( 
.A(n_11173),
.Y(n_11424)
);

AND2x2_ASAP7_75t_L g11425 ( 
.A(n_10802),
.B(n_9199),
.Y(n_11425)
);

INVx2_ASAP7_75t_L g11426 ( 
.A(n_11173),
.Y(n_11426)
);

AND2x4_ASAP7_75t_L g11427 ( 
.A(n_10419),
.B(n_8929),
.Y(n_11427)
);

AND2x2_ASAP7_75t_L g11428 ( 
.A(n_10686),
.B(n_9199),
.Y(n_11428)
);

AND2x2_ASAP7_75t_L g11429 ( 
.A(n_10691),
.B(n_9199),
.Y(n_11429)
);

AND2x2_ASAP7_75t_L g11430 ( 
.A(n_10695),
.B(n_9199),
.Y(n_11430)
);

INVx1_ASAP7_75t_L g11431 ( 
.A(n_10730),
.Y(n_11431)
);

INVx2_ASAP7_75t_L g11432 ( 
.A(n_11192),
.Y(n_11432)
);

AND2x2_ASAP7_75t_L g11433 ( 
.A(n_10714),
.B(n_10019),
.Y(n_11433)
);

INVx2_ASAP7_75t_L g11434 ( 
.A(n_11192),
.Y(n_11434)
);

INVx2_ASAP7_75t_L g11435 ( 
.A(n_11204),
.Y(n_11435)
);

INVx2_ASAP7_75t_L g11436 ( 
.A(n_11204),
.Y(n_11436)
);

INVx1_ASAP7_75t_L g11437 ( 
.A(n_10735),
.Y(n_11437)
);

NAND2x1p5_ASAP7_75t_L g11438 ( 
.A(n_11159),
.B(n_8383),
.Y(n_11438)
);

AND2x2_ASAP7_75t_L g11439 ( 
.A(n_10627),
.B(n_10019),
.Y(n_11439)
);

INVx1_ASAP7_75t_L g11440 ( 
.A(n_10736),
.Y(n_11440)
);

INVx2_ASAP7_75t_L g11441 ( 
.A(n_11159),
.Y(n_11441)
);

AND2x4_ASAP7_75t_L g11442 ( 
.A(n_10720),
.B(n_8970),
.Y(n_11442)
);

BUFx2_ASAP7_75t_L g11443 ( 
.A(n_10659),
.Y(n_11443)
);

INVxp67_ASAP7_75t_SL g11444 ( 
.A(n_10512),
.Y(n_11444)
);

INVx2_ASAP7_75t_L g11445 ( 
.A(n_11159),
.Y(n_11445)
);

BUFx2_ASAP7_75t_L g11446 ( 
.A(n_10659),
.Y(n_11446)
);

INVx1_ASAP7_75t_L g11447 ( 
.A(n_10741),
.Y(n_11447)
);

AND2x4_ASAP7_75t_L g11448 ( 
.A(n_11182),
.B(n_8970),
.Y(n_11448)
);

AND2x2_ASAP7_75t_L g11449 ( 
.A(n_11224),
.B(n_11231),
.Y(n_11449)
);

INVx2_ASAP7_75t_L g11450 ( 
.A(n_11077),
.Y(n_11450)
);

AND2x2_ASAP7_75t_L g11451 ( 
.A(n_10827),
.B(n_8345),
.Y(n_11451)
);

OR2x2_ASAP7_75t_L g11452 ( 
.A(n_11002),
.B(n_9760),
.Y(n_11452)
);

INVx2_ASAP7_75t_L g11453 ( 
.A(n_11166),
.Y(n_11453)
);

INVx2_ASAP7_75t_L g11454 ( 
.A(n_11053),
.Y(n_11454)
);

BUFx3_ASAP7_75t_L g11455 ( 
.A(n_10436),
.Y(n_11455)
);

INVx1_ASAP7_75t_L g11456 ( 
.A(n_10775),
.Y(n_11456)
);

CKINVDCx20_ASAP7_75t_R g11457 ( 
.A(n_10481),
.Y(n_11457)
);

BUFx2_ASAP7_75t_L g11458 ( 
.A(n_10823),
.Y(n_11458)
);

AND2x2_ASAP7_75t_L g11459 ( 
.A(n_10830),
.B(n_8345),
.Y(n_11459)
);

INVxp67_ASAP7_75t_L g11460 ( 
.A(n_10959),
.Y(n_11460)
);

NAND2x1_ASAP7_75t_L g11461 ( 
.A(n_10551),
.B(n_9841),
.Y(n_11461)
);

AND2x2_ASAP7_75t_L g11462 ( 
.A(n_10831),
.B(n_8345),
.Y(n_11462)
);

INVxp67_ASAP7_75t_L g11463 ( 
.A(n_10577),
.Y(n_11463)
);

AND2x2_ASAP7_75t_L g11464 ( 
.A(n_11182),
.B(n_8345),
.Y(n_11464)
);

INVx1_ASAP7_75t_L g11465 ( 
.A(n_10792),
.Y(n_11465)
);

AND2x2_ASAP7_75t_L g11466 ( 
.A(n_11190),
.B(n_10074),
.Y(n_11466)
);

NAND2xp5_ASAP7_75t_L g11467 ( 
.A(n_11162),
.B(n_10794),
.Y(n_11467)
);

NOR2xp67_ASAP7_75t_L g11468 ( 
.A(n_10655),
.B(n_10243),
.Y(n_11468)
);

INVx1_ASAP7_75t_L g11469 ( 
.A(n_10805),
.Y(n_11469)
);

INVx1_ASAP7_75t_L g11470 ( 
.A(n_10819),
.Y(n_11470)
);

AND2x4_ASAP7_75t_L g11471 ( 
.A(n_11089),
.B(n_8970),
.Y(n_11471)
);

INVx2_ASAP7_75t_L g11472 ( 
.A(n_11053),
.Y(n_11472)
);

INVx2_ASAP7_75t_L g11473 ( 
.A(n_11053),
.Y(n_11473)
);

INVx1_ASAP7_75t_L g11474 ( 
.A(n_10826),
.Y(n_11474)
);

NOR2xp33_ASAP7_75t_L g11475 ( 
.A(n_10655),
.B(n_10956),
.Y(n_11475)
);

INVx3_ASAP7_75t_L g11476 ( 
.A(n_10481),
.Y(n_11476)
);

AND2x2_ASAP7_75t_L g11477 ( 
.A(n_10578),
.B(n_10072),
.Y(n_11477)
);

INVx1_ASAP7_75t_L g11478 ( 
.A(n_10843),
.Y(n_11478)
);

AND2x2_ASAP7_75t_L g11479 ( 
.A(n_10578),
.B(n_10072),
.Y(n_11479)
);

INVx4_ASAP7_75t_L g11480 ( 
.A(n_10643),
.Y(n_11480)
);

INVx5_ASAP7_75t_L g11481 ( 
.A(n_10577),
.Y(n_11481)
);

INVx2_ASAP7_75t_L g11482 ( 
.A(n_11053),
.Y(n_11482)
);

INVx2_ASAP7_75t_L g11483 ( 
.A(n_11053),
.Y(n_11483)
);

HB1xp67_ASAP7_75t_L g11484 ( 
.A(n_11101),
.Y(n_11484)
);

NOR2xp33_ASAP7_75t_L g11485 ( 
.A(n_10956),
.B(n_10995),
.Y(n_11485)
);

BUFx6f_ASAP7_75t_L g11486 ( 
.A(n_10577),
.Y(n_11486)
);

BUFx3_ASAP7_75t_L g11487 ( 
.A(n_10436),
.Y(n_11487)
);

HB1xp67_ASAP7_75t_L g11488 ( 
.A(n_11115),
.Y(n_11488)
);

INVx2_ASAP7_75t_L g11489 ( 
.A(n_11132),
.Y(n_11489)
);

NAND2xp5_ASAP7_75t_L g11490 ( 
.A(n_10816),
.B(n_10204),
.Y(n_11490)
);

BUFx6f_ASAP7_75t_L g11491 ( 
.A(n_10732),
.Y(n_11491)
);

OR2x2_ASAP7_75t_L g11492 ( 
.A(n_11050),
.B(n_9762),
.Y(n_11492)
);

AND2x2_ASAP7_75t_L g11493 ( 
.A(n_11127),
.B(n_10072),
.Y(n_11493)
);

INVx2_ASAP7_75t_L g11494 ( 
.A(n_11134),
.Y(n_11494)
);

INVx1_ASAP7_75t_L g11495 ( 
.A(n_10844),
.Y(n_11495)
);

HB1xp67_ASAP7_75t_L g11496 ( 
.A(n_11157),
.Y(n_11496)
);

AND2x2_ASAP7_75t_L g11497 ( 
.A(n_11127),
.B(n_10126),
.Y(n_11497)
);

AND2x2_ASAP7_75t_L g11498 ( 
.A(n_11164),
.B(n_10809),
.Y(n_11498)
);

AND2x2_ASAP7_75t_L g11499 ( 
.A(n_11164),
.B(n_10126),
.Y(n_11499)
);

INVx1_ASAP7_75t_L g11500 ( 
.A(n_10852),
.Y(n_11500)
);

BUFx2_ASAP7_75t_L g11501 ( 
.A(n_10877),
.Y(n_11501)
);

OR2x2_ASAP7_75t_L g11502 ( 
.A(n_11124),
.B(n_9772),
.Y(n_11502)
);

AND2x2_ASAP7_75t_L g11503 ( 
.A(n_10812),
.B(n_10126),
.Y(n_11503)
);

INVx1_ASAP7_75t_L g11504 ( 
.A(n_10853),
.Y(n_11504)
);

BUFx2_ASAP7_75t_L g11505 ( 
.A(n_10877),
.Y(n_11505)
);

INVx2_ASAP7_75t_R g11506 ( 
.A(n_10857),
.Y(n_11506)
);

AND2x2_ASAP7_75t_L g11507 ( 
.A(n_10988),
.B(n_10195),
.Y(n_11507)
);

OR2x2_ASAP7_75t_L g11508 ( 
.A(n_11133),
.B(n_9775),
.Y(n_11508)
);

INVx1_ASAP7_75t_L g11509 ( 
.A(n_10862),
.Y(n_11509)
);

AND2x2_ASAP7_75t_L g11510 ( 
.A(n_10988),
.B(n_10195),
.Y(n_11510)
);

OR2x2_ASAP7_75t_L g11511 ( 
.A(n_11161),
.B(n_9781),
.Y(n_11511)
);

HB1xp67_ASAP7_75t_L g11512 ( 
.A(n_10941),
.Y(n_11512)
);

INVx1_ASAP7_75t_L g11513 ( 
.A(n_10871),
.Y(n_11513)
);

AND2x2_ASAP7_75t_L g11514 ( 
.A(n_11033),
.B(n_10195),
.Y(n_11514)
);

HB1xp67_ASAP7_75t_L g11515 ( 
.A(n_11189),
.Y(n_11515)
);

AND2x2_ASAP7_75t_L g11516 ( 
.A(n_11033),
.B(n_10195),
.Y(n_11516)
);

AND2x2_ASAP7_75t_L g11517 ( 
.A(n_11056),
.B(n_11089),
.Y(n_11517)
);

AND2x2_ASAP7_75t_L g11518 ( 
.A(n_11056),
.B(n_10948),
.Y(n_11518)
);

AND2x2_ASAP7_75t_L g11519 ( 
.A(n_10948),
.B(n_10237),
.Y(n_11519)
);

AND2x2_ASAP7_75t_L g11520 ( 
.A(n_10955),
.B(n_10237),
.Y(n_11520)
);

AND2x2_ASAP7_75t_L g11521 ( 
.A(n_10955),
.B(n_10237),
.Y(n_11521)
);

INVx1_ASAP7_75t_L g11522 ( 
.A(n_10878),
.Y(n_11522)
);

INVx1_ASAP7_75t_L g11523 ( 
.A(n_10886),
.Y(n_11523)
);

INVx1_ASAP7_75t_L g11524 ( 
.A(n_10907),
.Y(n_11524)
);

BUFx2_ASAP7_75t_L g11525 ( 
.A(n_10436),
.Y(n_11525)
);

AND2x2_ASAP7_75t_L g11526 ( 
.A(n_10483),
.B(n_10237),
.Y(n_11526)
);

AND2x2_ASAP7_75t_L g11527 ( 
.A(n_10483),
.B(n_10275),
.Y(n_11527)
);

AND2x2_ASAP7_75t_L g11528 ( 
.A(n_10556),
.B(n_10275),
.Y(n_11528)
);

INVx2_ASAP7_75t_L g11529 ( 
.A(n_10439),
.Y(n_11529)
);

INVx2_ASAP7_75t_L g11530 ( 
.A(n_10439),
.Y(n_11530)
);

INVx1_ASAP7_75t_L g11531 ( 
.A(n_10922),
.Y(n_11531)
);

INVx1_ASAP7_75t_L g11532 ( 
.A(n_10940),
.Y(n_11532)
);

INVx1_ASAP7_75t_L g11533 ( 
.A(n_10952),
.Y(n_11533)
);

OAI22xp5_ASAP7_75t_L g11534 ( 
.A1(n_10463),
.A2(n_9038),
.B1(n_8096),
.B2(n_8181),
.Y(n_11534)
);

AND2x2_ASAP7_75t_L g11535 ( 
.A(n_10556),
.B(n_10275),
.Y(n_11535)
);

AND2x2_ASAP7_75t_L g11536 ( 
.A(n_10798),
.B(n_10275),
.Y(n_11536)
);

NAND2xp5_ASAP7_75t_L g11537 ( 
.A(n_10476),
.B(n_10204),
.Y(n_11537)
);

HB1xp67_ASAP7_75t_SL g11538 ( 
.A(n_10436),
.Y(n_11538)
);

AND2x4_ASAP7_75t_L g11539 ( 
.A(n_10734),
.B(n_10243),
.Y(n_11539)
);

INVx1_ASAP7_75t_L g11540 ( 
.A(n_10964),
.Y(n_11540)
);

HB1xp67_ASAP7_75t_L g11541 ( 
.A(n_11195),
.Y(n_11541)
);

AND2x2_ASAP7_75t_L g11542 ( 
.A(n_10798),
.B(n_10801),
.Y(n_11542)
);

INVx2_ASAP7_75t_L g11543 ( 
.A(n_11062),
.Y(n_11543)
);

AND2x2_ASAP7_75t_L g11544 ( 
.A(n_10801),
.B(n_10318),
.Y(n_11544)
);

INVx1_ASAP7_75t_L g11545 ( 
.A(n_10966),
.Y(n_11545)
);

INVx2_ASAP7_75t_L g11546 ( 
.A(n_11062),
.Y(n_11546)
);

NAND2xp5_ASAP7_75t_L g11547 ( 
.A(n_11012),
.B(n_10204),
.Y(n_11547)
);

INVx1_ASAP7_75t_L g11548 ( 
.A(n_10968),
.Y(n_11548)
);

INVx1_ASAP7_75t_L g11549 ( 
.A(n_10978),
.Y(n_11549)
);

AND2x2_ASAP7_75t_L g11550 ( 
.A(n_10566),
.B(n_10318),
.Y(n_11550)
);

CKINVDCx5p33_ASAP7_75t_R g11551 ( 
.A(n_10814),
.Y(n_11551)
);

BUFx2_ASAP7_75t_L g11552 ( 
.A(n_10436),
.Y(n_11552)
);

BUFx2_ASAP7_75t_L g11553 ( 
.A(n_11194),
.Y(n_11553)
);

INVx4_ASAP7_75t_L g11554 ( 
.A(n_10643),
.Y(n_11554)
);

INVx2_ASAP7_75t_L g11555 ( 
.A(n_11062),
.Y(n_11555)
);

INVx2_ASAP7_75t_L g11556 ( 
.A(n_10510),
.Y(n_11556)
);

HB1xp67_ASAP7_75t_L g11557 ( 
.A(n_10553),
.Y(n_11557)
);

INVx1_ASAP7_75t_SL g11558 ( 
.A(n_10881),
.Y(n_11558)
);

HB1xp67_ASAP7_75t_L g11559 ( 
.A(n_10564),
.Y(n_11559)
);

INVx3_ASAP7_75t_L g11560 ( 
.A(n_10732),
.Y(n_11560)
);

INVx1_ASAP7_75t_L g11561 ( 
.A(n_10981),
.Y(n_11561)
);

NAND2xp5_ASAP7_75t_L g11562 ( 
.A(n_10427),
.B(n_10413),
.Y(n_11562)
);

INVx1_ASAP7_75t_L g11563 ( 
.A(n_10986),
.Y(n_11563)
);

INVx2_ASAP7_75t_L g11564 ( 
.A(n_10535),
.Y(n_11564)
);

INVx1_ASAP7_75t_L g11565 ( 
.A(n_10991),
.Y(n_11565)
);

OR2x2_ASAP7_75t_L g11566 ( 
.A(n_11180),
.B(n_9787),
.Y(n_11566)
);

OR2x2_ASAP7_75t_L g11567 ( 
.A(n_10960),
.B(n_9799),
.Y(n_11567)
);

OAI22xp5_ASAP7_75t_L g11568 ( 
.A1(n_10442),
.A2(n_9038),
.B1(n_8096),
.B2(n_8181),
.Y(n_11568)
);

BUFx3_ASAP7_75t_L g11569 ( 
.A(n_10732),
.Y(n_11569)
);

NAND2xp5_ASAP7_75t_L g11570 ( 
.A(n_10666),
.B(n_10204),
.Y(n_11570)
);

INVx1_ASAP7_75t_L g11571 ( 
.A(n_11022),
.Y(n_11571)
);

BUFx6f_ASAP7_75t_L g11572 ( 
.A(n_10787),
.Y(n_11572)
);

INVx2_ASAP7_75t_L g11573 ( 
.A(n_10933),
.Y(n_11573)
);

OAI22xp5_ASAP7_75t_L g11574 ( 
.A1(n_10417),
.A2(n_8096),
.B1(n_8181),
.B2(n_7941),
.Y(n_11574)
);

INVx2_ASAP7_75t_L g11575 ( 
.A(n_10933),
.Y(n_11575)
);

AND2x2_ASAP7_75t_L g11576 ( 
.A(n_10566),
.B(n_10318),
.Y(n_11576)
);

AND2x4_ASAP7_75t_L g11577 ( 
.A(n_10751),
.B(n_10308),
.Y(n_11577)
);

AND2x2_ASAP7_75t_L g11578 ( 
.A(n_10861),
.B(n_10318),
.Y(n_11578)
);

INVx1_ASAP7_75t_L g11579 ( 
.A(n_11023),
.Y(n_11579)
);

BUFx2_ASAP7_75t_L g11580 ( 
.A(n_10787),
.Y(n_11580)
);

AND2x2_ASAP7_75t_L g11581 ( 
.A(n_10861),
.B(n_10406),
.Y(n_11581)
);

AND2x2_ASAP7_75t_L g11582 ( 
.A(n_11200),
.B(n_10406),
.Y(n_11582)
);

AND2x2_ASAP7_75t_L g11583 ( 
.A(n_10885),
.B(n_10406),
.Y(n_11583)
);

NAND2xp5_ASAP7_75t_L g11584 ( 
.A(n_11168),
.B(n_10204),
.Y(n_11584)
);

INVx1_ASAP7_75t_L g11585 ( 
.A(n_11025),
.Y(n_11585)
);

INVx2_ASAP7_75t_L g11586 ( 
.A(n_10933),
.Y(n_11586)
);

OR2x2_ASAP7_75t_L g11587 ( 
.A(n_10985),
.B(n_9801),
.Y(n_11587)
);

AND2x2_ASAP7_75t_L g11588 ( 
.A(n_10885),
.B(n_11029),
.Y(n_11588)
);

BUFx2_ASAP7_75t_L g11589 ( 
.A(n_10787),
.Y(n_11589)
);

AOI22xp33_ASAP7_75t_L g11590 ( 
.A1(n_10912),
.A2(n_9818),
.B1(n_9823),
.B2(n_9811),
.Y(n_11590)
);

CKINVDCx5p33_ASAP7_75t_R g11591 ( 
.A(n_11051),
.Y(n_11591)
);

INVx2_ASAP7_75t_L g11592 ( 
.A(n_10860),
.Y(n_11592)
);

NOR2x1p5_ASAP7_75t_L g11593 ( 
.A(n_11066),
.B(n_10995),
.Y(n_11593)
);

INVx1_ASAP7_75t_L g11594 ( 
.A(n_11035),
.Y(n_11594)
);

INVx1_ASAP7_75t_L g11595 ( 
.A(n_11042),
.Y(n_11595)
);

NAND2xp5_ASAP7_75t_L g11596 ( 
.A(n_10752),
.B(n_10308),
.Y(n_11596)
);

INVx1_ASAP7_75t_L g11597 ( 
.A(n_11045),
.Y(n_11597)
);

OR2x6_ASAP7_75t_L g11598 ( 
.A(n_10860),
.B(n_9878),
.Y(n_11598)
);

INVx1_ASAP7_75t_L g11599 ( 
.A(n_11046),
.Y(n_11599)
);

INVx2_ASAP7_75t_L g11600 ( 
.A(n_10860),
.Y(n_11600)
);

INVx1_ASAP7_75t_L g11601 ( 
.A(n_11058),
.Y(n_11601)
);

INVx1_ASAP7_75t_L g11602 ( 
.A(n_11061),
.Y(n_11602)
);

BUFx6f_ASAP7_75t_L g11603 ( 
.A(n_11066),
.Y(n_11603)
);

AND2x2_ASAP7_75t_L g11604 ( 
.A(n_11114),
.B(n_10406),
.Y(n_11604)
);

AND2x2_ASAP7_75t_L g11605 ( 
.A(n_10881),
.B(n_10321),
.Y(n_11605)
);

AOI22xp33_ASAP7_75t_L g11606 ( 
.A1(n_10912),
.A2(n_9829),
.B1(n_9830),
.B2(n_9823),
.Y(n_11606)
);

INVx2_ASAP7_75t_L g11607 ( 
.A(n_10963),
.Y(n_11607)
);

INVx2_ASAP7_75t_L g11608 ( 
.A(n_11041),
.Y(n_11608)
);

OR2x2_ASAP7_75t_L g11609 ( 
.A(n_11044),
.B(n_9805),
.Y(n_11609)
);

INVx2_ASAP7_75t_L g11610 ( 
.A(n_10594),
.Y(n_11610)
);

OR2x2_ASAP7_75t_L g11611 ( 
.A(n_10596),
.B(n_9809),
.Y(n_11611)
);

AND2x4_ASAP7_75t_L g11612 ( 
.A(n_10876),
.B(n_10321),
.Y(n_11612)
);

NAND2xp5_ASAP7_75t_L g11613 ( 
.A(n_10626),
.B(n_10459),
.Y(n_11613)
);

INVx1_ASAP7_75t_L g11614 ( 
.A(n_11070),
.Y(n_11614)
);

INVx1_ASAP7_75t_L g11615 ( 
.A(n_11082),
.Y(n_11615)
);

INVx1_ASAP7_75t_L g11616 ( 
.A(n_11106),
.Y(n_11616)
);

AND2x2_ASAP7_75t_L g11617 ( 
.A(n_10450),
.B(n_11092),
.Y(n_11617)
);

AND2x4_ASAP7_75t_SL g11618 ( 
.A(n_10908),
.B(n_8024),
.Y(n_11618)
);

AND2x2_ASAP7_75t_L g11619 ( 
.A(n_10900),
.B(n_10603),
.Y(n_11619)
);

AND2x2_ASAP7_75t_L g11620 ( 
.A(n_10630),
.B(n_10322),
.Y(n_11620)
);

AND2x2_ASAP7_75t_L g11621 ( 
.A(n_10636),
.B(n_10322),
.Y(n_11621)
);

NAND2xp5_ASAP7_75t_L g11622 ( 
.A(n_10584),
.B(n_10402),
.Y(n_11622)
);

AND2x2_ASAP7_75t_L g11623 ( 
.A(n_10647),
.B(n_10402),
.Y(n_11623)
);

INVx1_ASAP7_75t_L g11624 ( 
.A(n_11107),
.Y(n_11624)
);

AND2x2_ASAP7_75t_L g11625 ( 
.A(n_10665),
.B(n_10042),
.Y(n_11625)
);

INVx2_ASAP7_75t_L g11626 ( 
.A(n_10670),
.Y(n_11626)
);

AND2x2_ASAP7_75t_L g11627 ( 
.A(n_10673),
.B(n_10719),
.Y(n_11627)
);

INVx1_ASAP7_75t_L g11628 ( 
.A(n_11120),
.Y(n_11628)
);

OR2x2_ASAP7_75t_L g11629 ( 
.A(n_10606),
.B(n_9813),
.Y(n_11629)
);

AND2x2_ASAP7_75t_L g11630 ( 
.A(n_10722),
.B(n_10042),
.Y(n_11630)
);

AND2x2_ASAP7_75t_L g11631 ( 
.A(n_10738),
.B(n_10107),
.Y(n_11631)
);

AND2x2_ASAP7_75t_L g11632 ( 
.A(n_10858),
.B(n_10107),
.Y(n_11632)
);

INVx1_ASAP7_75t_L g11633 ( 
.A(n_11145),
.Y(n_11633)
);

INVx1_ASAP7_75t_L g11634 ( 
.A(n_11151),
.Y(n_11634)
);

AND2x2_ASAP7_75t_L g11635 ( 
.A(n_10897),
.B(n_10123),
.Y(n_11635)
);

AND2x2_ASAP7_75t_L g11636 ( 
.A(n_10909),
.B(n_10123),
.Y(n_11636)
);

HB1xp67_ASAP7_75t_L g11637 ( 
.A(n_10910),
.Y(n_11637)
);

INVx1_ASAP7_75t_L g11638 ( 
.A(n_11160),
.Y(n_11638)
);

INVx2_ASAP7_75t_SL g11639 ( 
.A(n_10803),
.Y(n_11639)
);

INVx2_ASAP7_75t_L g11640 ( 
.A(n_10947),
.Y(n_11640)
);

INVxp67_ASAP7_75t_SL g11641 ( 
.A(n_10839),
.Y(n_11641)
);

NOR2xp33_ASAP7_75t_L g11642 ( 
.A(n_10806),
.B(n_6867),
.Y(n_11642)
);

NAND2xp5_ASAP7_75t_L g11643 ( 
.A(n_10449),
.B(n_10425),
.Y(n_11643)
);

NAND2xp5_ASAP7_75t_L g11644 ( 
.A(n_10477),
.B(n_9001),
.Y(n_11644)
);

AND2x2_ASAP7_75t_L g11645 ( 
.A(n_11117),
.B(n_10134),
.Y(n_11645)
);

INVx1_ASAP7_75t_L g11646 ( 
.A(n_11171),
.Y(n_11646)
);

AOI22xp33_ASAP7_75t_L g11647 ( 
.A1(n_10477),
.A2(n_9830),
.B1(n_9834),
.B2(n_9829),
.Y(n_11647)
);

INVx2_ASAP7_75t_L g11648 ( 
.A(n_11122),
.Y(n_11648)
);

BUFx2_ASAP7_75t_L g11649 ( 
.A(n_10494),
.Y(n_11649)
);

AND2x2_ASAP7_75t_L g11650 ( 
.A(n_10689),
.B(n_10134),
.Y(n_11650)
);

AND2x2_ASAP7_75t_L g11651 ( 
.A(n_10624),
.B(n_8715),
.Y(n_11651)
);

AND2x2_ASAP7_75t_L g11652 ( 
.A(n_11001),
.B(n_8715),
.Y(n_11652)
);

INVx1_ASAP7_75t_L g11653 ( 
.A(n_11211),
.Y(n_11653)
);

BUFx3_ASAP7_75t_L g11654 ( 
.A(n_10652),
.Y(n_11654)
);

AOI22xp33_ASAP7_75t_L g11655 ( 
.A1(n_10473),
.A2(n_9836),
.B1(n_9843),
.B2(n_9834),
.Y(n_11655)
);

INVx2_ASAP7_75t_L g11656 ( 
.A(n_10440),
.Y(n_11656)
);

AND2x2_ASAP7_75t_L g11657 ( 
.A(n_11005),
.B(n_8715),
.Y(n_11657)
);

AND2x2_ASAP7_75t_L g11658 ( 
.A(n_11007),
.B(n_8715),
.Y(n_11658)
);

AND2x2_ASAP7_75t_L g11659 ( 
.A(n_11010),
.B(n_8717),
.Y(n_11659)
);

CKINVDCx14_ASAP7_75t_R g11660 ( 
.A(n_10765),
.Y(n_11660)
);

AND2x2_ASAP7_75t_L g11661 ( 
.A(n_11013),
.B(n_8717),
.Y(n_11661)
);

OAI22xp33_ASAP7_75t_L g11662 ( 
.A1(n_10586),
.A2(n_10423),
.B1(n_10711),
.B2(n_10432),
.Y(n_11662)
);

INVx1_ASAP7_75t_L g11663 ( 
.A(n_11214),
.Y(n_11663)
);

INVx1_ASAP7_75t_L g11664 ( 
.A(n_11218),
.Y(n_11664)
);

INVx1_ASAP7_75t_L g11665 ( 
.A(n_11220),
.Y(n_11665)
);

INVx2_ASAP7_75t_L g11666 ( 
.A(n_10444),
.Y(n_11666)
);

INVx3_ASAP7_75t_L g11667 ( 
.A(n_10448),
.Y(n_11667)
);

AND2x4_ASAP7_75t_SL g11668 ( 
.A(n_10987),
.B(n_8040),
.Y(n_11668)
);

OR2x2_ASAP7_75t_L g11669 ( 
.A(n_10506),
.B(n_9819),
.Y(n_11669)
);

BUFx3_ASAP7_75t_L g11670 ( 
.A(n_10777),
.Y(n_11670)
);

INVxp67_ASAP7_75t_L g11671 ( 
.A(n_10984),
.Y(n_11671)
);

INVx2_ASAP7_75t_SL g11672 ( 
.A(n_11188),
.Y(n_11672)
);

NAND2xp5_ASAP7_75t_L g11673 ( 
.A(n_10708),
.B(n_9001),
.Y(n_11673)
);

INVx3_ASAP7_75t_L g11674 ( 
.A(n_10448),
.Y(n_11674)
);

INVx2_ASAP7_75t_L g11675 ( 
.A(n_10761),
.Y(n_11675)
);

INVx2_ASAP7_75t_L g11676 ( 
.A(n_10761),
.Y(n_11676)
);

INVx2_ASAP7_75t_SL g11677 ( 
.A(n_10797),
.Y(n_11677)
);

INVxp67_ASAP7_75t_L g11678 ( 
.A(n_10685),
.Y(n_11678)
);

INVx1_ASAP7_75t_L g11679 ( 
.A(n_11232),
.Y(n_11679)
);

INVx2_ASAP7_75t_L g11680 ( 
.A(n_10448),
.Y(n_11680)
);

AND2x4_ASAP7_75t_L g11681 ( 
.A(n_10990),
.B(n_8383),
.Y(n_11681)
);

INVxp67_ASAP7_75t_L g11682 ( 
.A(n_10810),
.Y(n_11682)
);

INVx2_ASAP7_75t_L g11683 ( 
.A(n_11169),
.Y(n_11683)
);

INVx2_ASAP7_75t_SL g11684 ( 
.A(n_11153),
.Y(n_11684)
);

INVx2_ASAP7_75t_L g11685 ( 
.A(n_11179),
.Y(n_11685)
);

NAND2xp5_ASAP7_75t_L g11686 ( 
.A(n_10467),
.B(n_9007),
.Y(n_11686)
);

INVx1_ASAP7_75t_L g11687 ( 
.A(n_10769),
.Y(n_11687)
);

INVx1_ASAP7_75t_L g11688 ( 
.A(n_10769),
.Y(n_11688)
);

NOR2x1_ASAP7_75t_L g11689 ( 
.A(n_10469),
.B(n_10629),
.Y(n_11689)
);

AND2x2_ASAP7_75t_L g11690 ( 
.A(n_11014),
.B(n_8717),
.Y(n_11690)
);

INVx2_ASAP7_75t_L g11691 ( 
.A(n_11181),
.Y(n_11691)
);

INVx1_ASAP7_75t_L g11692 ( 
.A(n_10684),
.Y(n_11692)
);

BUFx3_ASAP7_75t_L g11693 ( 
.A(n_11069),
.Y(n_11693)
);

INVxp67_ASAP7_75t_R g11694 ( 
.A(n_10724),
.Y(n_11694)
);

INVx2_ASAP7_75t_L g11695 ( 
.A(n_10549),
.Y(n_11695)
);

INVx1_ASAP7_75t_L g11696 ( 
.A(n_10684),
.Y(n_11696)
);

INVxp67_ASAP7_75t_L g11697 ( 
.A(n_10585),
.Y(n_11697)
);

INVx2_ASAP7_75t_L g11698 ( 
.A(n_10549),
.Y(n_11698)
);

AND2x2_ASAP7_75t_L g11699 ( 
.A(n_11015),
.B(n_8717),
.Y(n_11699)
);

HB1xp67_ASAP7_75t_L g11700 ( 
.A(n_10837),
.Y(n_11700)
);

INVx1_ASAP7_75t_L g11701 ( 
.A(n_10576),
.Y(n_11701)
);

CKINVDCx5p33_ASAP7_75t_R g11702 ( 
.A(n_10728),
.Y(n_11702)
);

INVx1_ASAP7_75t_L g11703 ( 
.A(n_10576),
.Y(n_11703)
);

INVx1_ASAP7_75t_L g11704 ( 
.A(n_10895),
.Y(n_11704)
);

INVx2_ASAP7_75t_L g11705 ( 
.A(n_10518),
.Y(n_11705)
);

INVx2_ASAP7_75t_L g11706 ( 
.A(n_10592),
.Y(n_11706)
);

INVx1_ASAP7_75t_L g11707 ( 
.A(n_10818),
.Y(n_11707)
);

INVx1_ASAP7_75t_L g11708 ( 
.A(n_11213),
.Y(n_11708)
);

AND2x2_ASAP7_75t_L g11709 ( 
.A(n_11017),
.B(n_8717),
.Y(n_11709)
);

INVxp67_ASAP7_75t_L g11710 ( 
.A(n_11103),
.Y(n_11710)
);

AND2x2_ASAP7_75t_L g11711 ( 
.A(n_11087),
.B(n_9868),
.Y(n_11711)
);

AND2x2_ASAP7_75t_L g11712 ( 
.A(n_10911),
.B(n_9868),
.Y(n_11712)
);

INVx2_ASAP7_75t_L g11713 ( 
.A(n_10592),
.Y(n_11713)
);

AND2x2_ASAP7_75t_L g11714 ( 
.A(n_10515),
.B(n_9879),
.Y(n_11714)
);

NAND2xp5_ASAP7_75t_L g11715 ( 
.A(n_10460),
.B(n_9007),
.Y(n_11715)
);

AND2x2_ASAP7_75t_L g11716 ( 
.A(n_11108),
.B(n_9879),
.Y(n_11716)
);

NAND2xp5_ASAP7_75t_L g11717 ( 
.A(n_10605),
.B(n_9010),
.Y(n_11717)
);

AND2x2_ASAP7_75t_L g11718 ( 
.A(n_11111),
.B(n_9899),
.Y(n_11718)
);

NAND2xp5_ASAP7_75t_L g11719 ( 
.A(n_10429),
.B(n_9010),
.Y(n_11719)
);

INVx1_ASAP7_75t_L g11720 ( 
.A(n_10646),
.Y(n_11720)
);

INVx1_ASAP7_75t_L g11721 ( 
.A(n_10646),
.Y(n_11721)
);

AOI22xp33_ASAP7_75t_L g11722 ( 
.A1(n_10452),
.A2(n_9843),
.B1(n_9844),
.B2(n_9836),
.Y(n_11722)
);

INVx1_ASAP7_75t_L g11723 ( 
.A(n_10646),
.Y(n_11723)
);

OR2x2_ASAP7_75t_L g11724 ( 
.A(n_10579),
.B(n_10539),
.Y(n_11724)
);

INVx1_ASAP7_75t_L g11725 ( 
.A(n_10541),
.Y(n_11725)
);

INVx1_ASAP7_75t_L g11726 ( 
.A(n_10542),
.Y(n_11726)
);

INVx2_ASAP7_75t_L g11727 ( 
.A(n_10599),
.Y(n_11727)
);

AO21x2_ASAP7_75t_L g11728 ( 
.A1(n_10682),
.A2(n_10793),
.B(n_10710),
.Y(n_11728)
);

AND2x2_ASAP7_75t_L g11729 ( 
.A(n_11034),
.B(n_9899),
.Y(n_11729)
);

OAI22xp33_ASAP7_75t_L g11730 ( 
.A1(n_10754),
.A2(n_7666),
.B1(n_7901),
.B2(n_9844),
.Y(n_11730)
);

INVx2_ASAP7_75t_L g11731 ( 
.A(n_10599),
.Y(n_11731)
);

INVx2_ASAP7_75t_L g11732 ( 
.A(n_10435),
.Y(n_11732)
);

INVx2_ASAP7_75t_L g11733 ( 
.A(n_10702),
.Y(n_11733)
);

HB1xp67_ASAP7_75t_L g11734 ( 
.A(n_10703),
.Y(n_11734)
);

BUFx2_ASAP7_75t_L g11735 ( 
.A(n_10870),
.Y(n_11735)
);

AND2x2_ASAP7_75t_L g11736 ( 
.A(n_10615),
.B(n_9904),
.Y(n_11736)
);

INVx3_ASAP7_75t_SL g11737 ( 
.A(n_10527),
.Y(n_11737)
);

AND2x2_ASAP7_75t_L g11738 ( 
.A(n_10943),
.B(n_9904),
.Y(n_11738)
);

NAND2xp5_ASAP7_75t_L g11739 ( 
.A(n_10454),
.B(n_9824),
.Y(n_11739)
);

OR2x2_ASAP7_75t_L g11740 ( 
.A(n_10613),
.B(n_9826),
.Y(n_11740)
);

AND2x2_ASAP7_75t_L g11741 ( 
.A(n_10997),
.B(n_9910),
.Y(n_11741)
);

AND2x2_ASAP7_75t_L g11742 ( 
.A(n_10622),
.B(n_9910),
.Y(n_11742)
);

INVx1_ASAP7_75t_L g11743 ( 
.A(n_10658),
.Y(n_11743)
);

NAND2xp5_ASAP7_75t_L g11744 ( 
.A(n_10456),
.B(n_9828),
.Y(n_11744)
);

AND2x2_ASAP7_75t_L g11745 ( 
.A(n_10681),
.B(n_9940),
.Y(n_11745)
);

NAND2xp5_ASAP7_75t_L g11746 ( 
.A(n_10508),
.B(n_9831),
.Y(n_11746)
);

OR2x2_ASAP7_75t_L g11747 ( 
.A(n_10517),
.B(n_9842),
.Y(n_11747)
);

INVx1_ASAP7_75t_L g11748 ( 
.A(n_10658),
.Y(n_11748)
);

INVx2_ASAP7_75t_L g11749 ( 
.A(n_10702),
.Y(n_11749)
);

INVx1_ASAP7_75t_L g11750 ( 
.A(n_10677),
.Y(n_11750)
);

INVx1_ASAP7_75t_L g11751 ( 
.A(n_10677),
.Y(n_11751)
);

INVx1_ASAP7_75t_L g11752 ( 
.A(n_10920),
.Y(n_11752)
);

AND2x2_ASAP7_75t_L g11753 ( 
.A(n_11065),
.B(n_9940),
.Y(n_11753)
);

AND2x2_ASAP7_75t_L g11754 ( 
.A(n_11176),
.B(n_9990),
.Y(n_11754)
);

INVx1_ASAP7_75t_L g11755 ( 
.A(n_10920),
.Y(n_11755)
);

INVx1_ASAP7_75t_L g11756 ( 
.A(n_11150),
.Y(n_11756)
);

AND2x2_ASAP7_75t_L g11757 ( 
.A(n_11167),
.B(n_9990),
.Y(n_11757)
);

HB1xp67_ASAP7_75t_L g11758 ( 
.A(n_10795),
.Y(n_11758)
);

NAND2xp5_ASAP7_75t_L g11759 ( 
.A(n_10488),
.B(n_9848),
.Y(n_11759)
);

INVx1_ASAP7_75t_L g11760 ( 
.A(n_10709),
.Y(n_11760)
);

NAND2xp5_ASAP7_75t_L g11761 ( 
.A(n_10536),
.B(n_9855),
.Y(n_11761)
);

HB1xp67_ASAP7_75t_L g11762 ( 
.A(n_10609),
.Y(n_11762)
);

NAND2xp5_ASAP7_75t_L g11763 ( 
.A(n_10507),
.B(n_9856),
.Y(n_11763)
);

BUFx3_ASAP7_75t_L g11764 ( 
.A(n_10475),
.Y(n_11764)
);

AND2x2_ASAP7_75t_L g11765 ( 
.A(n_10654),
.B(n_9991),
.Y(n_11765)
);

OAI22xp33_ASAP7_75t_L g11766 ( 
.A1(n_11165),
.A2(n_9857),
.B1(n_9858),
.B2(n_9847),
.Y(n_11766)
);

AND2x2_ASAP7_75t_L g11767 ( 
.A(n_10656),
.B(n_9991),
.Y(n_11767)
);

AND2x2_ASAP7_75t_L g11768 ( 
.A(n_10753),
.B(n_10002),
.Y(n_11768)
);

HB1xp67_ASAP7_75t_L g11769 ( 
.A(n_10611),
.Y(n_11769)
);

AND2x2_ASAP7_75t_L g11770 ( 
.A(n_11098),
.B(n_10002),
.Y(n_11770)
);

OR2x2_ASAP7_75t_L g11771 ( 
.A(n_10588),
.B(n_9862),
.Y(n_11771)
);

AND2x2_ASAP7_75t_L g11772 ( 
.A(n_11105),
.B(n_10009),
.Y(n_11772)
);

INVx2_ASAP7_75t_L g11773 ( 
.A(n_10660),
.Y(n_11773)
);

INVx2_ASAP7_75t_L g11774 ( 
.A(n_10661),
.Y(n_11774)
);

NAND2xp5_ASAP7_75t_L g11775 ( 
.A(n_10464),
.B(n_9864),
.Y(n_11775)
);

INVx2_ASAP7_75t_L g11776 ( 
.A(n_11170),
.Y(n_11776)
);

INVx1_ASAP7_75t_L g11777 ( 
.A(n_10938),
.Y(n_11777)
);

OR2x2_ASAP7_75t_L g11778 ( 
.A(n_10800),
.B(n_9866),
.Y(n_11778)
);

BUFx2_ASAP7_75t_L g11779 ( 
.A(n_10866),
.Y(n_11779)
);

NAND2xp5_ASAP7_75t_L g11780 ( 
.A(n_10457),
.B(n_9867),
.Y(n_11780)
);

NAND2xp5_ASAP7_75t_L g11781 ( 
.A(n_10458),
.B(n_9869),
.Y(n_11781)
);

AND2x4_ASAP7_75t_L g11782 ( 
.A(n_10976),
.B(n_8383),
.Y(n_11782)
);

INVx2_ASAP7_75t_L g11783 ( 
.A(n_11113),
.Y(n_11783)
);

AND2x2_ASAP7_75t_L g11784 ( 
.A(n_11110),
.B(n_10009),
.Y(n_11784)
);

NAND2xp5_ASAP7_75t_L g11785 ( 
.A(n_10621),
.B(n_9870),
.Y(n_11785)
);

INVx1_ASAP7_75t_L g11786 ( 
.A(n_10938),
.Y(n_11786)
);

INVx2_ASAP7_75t_SL g11787 ( 
.A(n_10919),
.Y(n_11787)
);

HB1xp67_ASAP7_75t_L g11788 ( 
.A(n_10554),
.Y(n_11788)
);

INVx2_ASAP7_75t_L g11789 ( 
.A(n_11113),
.Y(n_11789)
);

AO21x2_ASAP7_75t_L g11790 ( 
.A1(n_10532),
.A2(n_9890),
.B(n_9886),
.Y(n_11790)
);

BUFx2_ASAP7_75t_L g11791 ( 
.A(n_10593),
.Y(n_11791)
);

AND2x2_ASAP7_75t_L g11792 ( 
.A(n_11112),
.B(n_10037),
.Y(n_11792)
);

BUFx3_ASAP7_75t_L g11793 ( 
.A(n_10974),
.Y(n_11793)
);

INVx1_ASAP7_75t_L g11794 ( 
.A(n_10755),
.Y(n_11794)
);

AND2x2_ASAP7_75t_L g11795 ( 
.A(n_11129),
.B(n_10037),
.Y(n_11795)
);

BUFx6f_ASAP7_75t_L g11796 ( 
.A(n_10896),
.Y(n_11796)
);

INVx2_ASAP7_75t_L g11797 ( 
.A(n_10841),
.Y(n_11797)
);

INVx2_ASAP7_75t_L g11798 ( 
.A(n_10847),
.Y(n_11798)
);

AND2x4_ASAP7_75t_L g11799 ( 
.A(n_10980),
.B(n_8383),
.Y(n_11799)
);

AND2x2_ASAP7_75t_L g11800 ( 
.A(n_11144),
.B(n_8373),
.Y(n_11800)
);

INVxp67_ASAP7_75t_SL g11801 ( 
.A(n_10633),
.Y(n_11801)
);

INVx2_ASAP7_75t_L g11802 ( 
.A(n_10764),
.Y(n_11802)
);

AND2x2_ASAP7_75t_L g11803 ( 
.A(n_11174),
.B(n_8373),
.Y(n_11803)
);

INVx2_ASAP7_75t_SL g11804 ( 
.A(n_10949),
.Y(n_11804)
);

INVx2_ASAP7_75t_L g11805 ( 
.A(n_10764),
.Y(n_11805)
);

AOI22xp33_ASAP7_75t_L g11806 ( 
.A1(n_10461),
.A2(n_10451),
.B1(n_10455),
.B2(n_10538),
.Y(n_11806)
);

AOI22xp33_ASAP7_75t_L g11807 ( 
.A1(n_10975),
.A2(n_10727),
.B1(n_10525),
.B2(n_10598),
.Y(n_11807)
);

INVx2_ASAP7_75t_L g11808 ( 
.A(n_11096),
.Y(n_11808)
);

INVx1_ASAP7_75t_L g11809 ( 
.A(n_11096),
.Y(n_11809)
);

AND2x2_ASAP7_75t_L g11810 ( 
.A(n_11184),
.B(n_8387),
.Y(n_11810)
);

AND2x2_ASAP7_75t_L g11811 ( 
.A(n_11185),
.B(n_8387),
.Y(n_11811)
);

NAND2xp5_ASAP7_75t_L g11812 ( 
.A(n_10472),
.B(n_9872),
.Y(n_11812)
);

INVx2_ASAP7_75t_L g11813 ( 
.A(n_10640),
.Y(n_11813)
);

INVx2_ASAP7_75t_L g11814 ( 
.A(n_10651),
.Y(n_11814)
);

INVx1_ASAP7_75t_L g11815 ( 
.A(n_10835),
.Y(n_11815)
);

INVx2_ASAP7_75t_SL g11816 ( 
.A(n_10951),
.Y(n_11816)
);

AND2x4_ASAP7_75t_L g11817 ( 
.A(n_11186),
.B(n_9152),
.Y(n_11817)
);

NAND2xp33_ASAP7_75t_SL g11818 ( 
.A(n_10480),
.B(n_6272),
.Y(n_11818)
);

INVx2_ASAP7_75t_L g11819 ( 
.A(n_10533),
.Y(n_11819)
);

AND2x2_ASAP7_75t_L g11820 ( 
.A(n_11201),
.B(n_8439),
.Y(n_11820)
);

INVx1_ASAP7_75t_L g11821 ( 
.A(n_10865),
.Y(n_11821)
);

NAND2x1_ASAP7_75t_L g11822 ( 
.A(n_10604),
.B(n_9281),
.Y(n_11822)
);

NOR2xp33_ASAP7_75t_L g11823 ( 
.A(n_10804),
.B(n_6867),
.Y(n_11823)
);

AND2x2_ASAP7_75t_L g11824 ( 
.A(n_11203),
.B(n_8439),
.Y(n_11824)
);

INVx1_ASAP7_75t_L g11825 ( 
.A(n_10888),
.Y(n_11825)
);

NAND2xp5_ASAP7_75t_L g11826 ( 
.A(n_10514),
.B(n_9876),
.Y(n_11826)
);

NAND2xp5_ASAP7_75t_L g11827 ( 
.A(n_10698),
.B(n_10905),
.Y(n_11827)
);

INVx1_ASAP7_75t_L g11828 ( 
.A(n_10890),
.Y(n_11828)
);

INVx2_ASAP7_75t_L g11829 ( 
.A(n_10915),
.Y(n_11829)
);

INVx1_ASAP7_75t_L g11830 ( 
.A(n_10999),
.Y(n_11830)
);

NAND2xp5_ASAP7_75t_L g11831 ( 
.A(n_10516),
.B(n_10942),
.Y(n_11831)
);

NAND2xp5_ASAP7_75t_L g11832 ( 
.A(n_10773),
.B(n_9881),
.Y(n_11832)
);

BUFx4f_ASAP7_75t_SL g11833 ( 
.A(n_10742),
.Y(n_11833)
);

HB1xp67_ASAP7_75t_L g11834 ( 
.A(n_10511),
.Y(n_11834)
);

INVx3_ASAP7_75t_L g11835 ( 
.A(n_10434),
.Y(n_11835)
);

INVx1_ASAP7_75t_L g11836 ( 
.A(n_11040),
.Y(n_11836)
);

AND2x2_ASAP7_75t_L g11837 ( 
.A(n_11208),
.B(n_8474),
.Y(n_11837)
);

AND2x2_ASAP7_75t_L g11838 ( 
.A(n_11217),
.B(n_8474),
.Y(n_11838)
);

AND2x2_ASAP7_75t_L g11839 ( 
.A(n_11223),
.B(n_8553),
.Y(n_11839)
);

INVx1_ASAP7_75t_L g11840 ( 
.A(n_11090),
.Y(n_11840)
);

BUFx2_ASAP7_75t_L g11841 ( 
.A(n_11119),
.Y(n_11841)
);

INVx1_ASAP7_75t_L g11842 ( 
.A(n_10567),
.Y(n_11842)
);

INVxp67_ASAP7_75t_L g11843 ( 
.A(n_10781),
.Y(n_11843)
);

AOI22xp33_ASAP7_75t_L g11844 ( 
.A1(n_10496),
.A2(n_10487),
.B1(n_10726),
.B2(n_10707),
.Y(n_11844)
);

INVx2_ASAP7_75t_L g11845 ( 
.A(n_11086),
.Y(n_11845)
);

INVx2_ASAP7_75t_L g11846 ( 
.A(n_11130),
.Y(n_11846)
);

INVx1_ASAP7_75t_L g11847 ( 
.A(n_10825),
.Y(n_11847)
);

OR2x2_ASAP7_75t_L g11848 ( 
.A(n_10848),
.B(n_10868),
.Y(n_11848)
);

INVx3_ASAP7_75t_L g11849 ( 
.A(n_10747),
.Y(n_11849)
);

INVx1_ASAP7_75t_L g11850 ( 
.A(n_10874),
.Y(n_11850)
);

INVx2_ASAP7_75t_L g11851 ( 
.A(n_11024),
.Y(n_11851)
);

INVx2_ASAP7_75t_L g11852 ( 
.A(n_10617),
.Y(n_11852)
);

INVx2_ASAP7_75t_L g11853 ( 
.A(n_10838),
.Y(n_11853)
);

OR2x2_ASAP7_75t_L g11854 ( 
.A(n_10901),
.B(n_9883),
.Y(n_11854)
);

INVx2_ASAP7_75t_L g11855 ( 
.A(n_10851),
.Y(n_11855)
);

AND2x2_ASAP7_75t_L g11856 ( 
.A(n_11229),
.B(n_8553),
.Y(n_11856)
);

NAND2x1_ASAP7_75t_L g11857 ( 
.A(n_10678),
.B(n_10813),
.Y(n_11857)
);

INVx3_ASAP7_75t_L g11858 ( 
.A(n_10743),
.Y(n_11858)
);

INVx2_ASAP7_75t_L g11859 ( 
.A(n_10923),
.Y(n_11859)
);

INVx1_ASAP7_75t_L g11860 ( 
.A(n_11102),
.Y(n_11860)
);

INVx1_ASAP7_75t_L g11861 ( 
.A(n_11183),
.Y(n_11861)
);

HB1xp67_ASAP7_75t_L g11862 ( 
.A(n_10521),
.Y(n_11862)
);

INVx2_ASAP7_75t_L g11863 ( 
.A(n_10925),
.Y(n_11863)
);

INVx1_ASAP7_75t_L g11864 ( 
.A(n_10791),
.Y(n_11864)
);

HB1xp67_ASAP7_75t_L g11865 ( 
.A(n_10558),
.Y(n_11865)
);

INVx1_ASAP7_75t_L g11866 ( 
.A(n_10904),
.Y(n_11866)
);

AND2x2_ASAP7_75t_L g11867 ( 
.A(n_10967),
.B(n_8624),
.Y(n_11867)
);

HB1xp67_ASAP7_75t_L g11868 ( 
.A(n_10559),
.Y(n_11868)
);

INVx2_ASAP7_75t_L g11869 ( 
.A(n_10927),
.Y(n_11869)
);

OR2x2_ASAP7_75t_L g11870 ( 
.A(n_10663),
.B(n_9887),
.Y(n_11870)
);

AND2x2_ASAP7_75t_L g11871 ( 
.A(n_10971),
.B(n_8624),
.Y(n_11871)
);

INVxp67_ASAP7_75t_L g11872 ( 
.A(n_10749),
.Y(n_11872)
);

INVx2_ASAP7_75t_L g11873 ( 
.A(n_11054),
.Y(n_11873)
);

INVx3_ASAP7_75t_L g11874 ( 
.A(n_10664),
.Y(n_11874)
);

AND2x2_ASAP7_75t_L g11875 ( 
.A(n_10977),
.B(n_9167),
.Y(n_11875)
);

INVx2_ASAP7_75t_L g11876 ( 
.A(n_10537),
.Y(n_11876)
);

INVx3_ASAP7_75t_L g11877 ( 
.A(n_10672),
.Y(n_11877)
);

AND2x2_ASAP7_75t_L g11878 ( 
.A(n_11093),
.B(n_9167),
.Y(n_11878)
);

INVx1_ASAP7_75t_L g11879 ( 
.A(n_11228),
.Y(n_11879)
);

INVx1_ASAP7_75t_L g11880 ( 
.A(n_10758),
.Y(n_11880)
);

INVx1_ASAP7_75t_L g11881 ( 
.A(n_11063),
.Y(n_11881)
);

INVx2_ASAP7_75t_L g11882 ( 
.A(n_10973),
.Y(n_11882)
);

OR2x2_ASAP7_75t_L g11883 ( 
.A(n_10829),
.B(n_9888),
.Y(n_11883)
);

BUFx3_ASAP7_75t_L g11884 ( 
.A(n_10822),
.Y(n_11884)
);

BUFx2_ASAP7_75t_L g11885 ( 
.A(n_10530),
.Y(n_11885)
);

INVx2_ASAP7_75t_L g11886 ( 
.A(n_11080),
.Y(n_11886)
);

HB1xp67_ASAP7_75t_L g11887 ( 
.A(n_10737),
.Y(n_11887)
);

AND2x2_ASAP7_75t_L g11888 ( 
.A(n_11095),
.B(n_9167),
.Y(n_11888)
);

HB1xp67_ASAP7_75t_L g11889 ( 
.A(n_10550),
.Y(n_11889)
);

INVx1_ASAP7_75t_L g11890 ( 
.A(n_10712),
.Y(n_11890)
);

INVx2_ASAP7_75t_L g11891 ( 
.A(n_11018),
.Y(n_11891)
);

INVx1_ASAP7_75t_L g11892 ( 
.A(n_10623),
.Y(n_11892)
);

INVx2_ASAP7_75t_L g11893 ( 
.A(n_11043),
.Y(n_11893)
);

AND2x4_ASAP7_75t_L g11894 ( 
.A(n_11057),
.B(n_9323),
.Y(n_11894)
);

INVx2_ASAP7_75t_L g11895 ( 
.A(n_10634),
.Y(n_11895)
);

INVx2_ASAP7_75t_L g11896 ( 
.A(n_10534),
.Y(n_11896)
);

INVx1_ASAP7_75t_L g11897 ( 
.A(n_10637),
.Y(n_11897)
);

INVx1_ASAP7_75t_L g11898 ( 
.A(n_10645),
.Y(n_11898)
);

INVx1_ASAP7_75t_L g11899 ( 
.A(n_10725),
.Y(n_11899)
);

OR2x2_ASAP7_75t_L g11900 ( 
.A(n_10489),
.B(n_9893),
.Y(n_11900)
);

AND2x2_ASAP7_75t_L g11901 ( 
.A(n_10864),
.B(n_9323),
.Y(n_11901)
);

INVx1_ASAP7_75t_L g11902 ( 
.A(n_10715),
.Y(n_11902)
);

INVx1_ASAP7_75t_L g11903 ( 
.A(n_10688),
.Y(n_11903)
);

INVx1_ASAP7_75t_L g11904 ( 
.A(n_10767),
.Y(n_11904)
);

INVx2_ASAP7_75t_L g11905 ( 
.A(n_10526),
.Y(n_11905)
);

INVx1_ASAP7_75t_L g11906 ( 
.A(n_10840),
.Y(n_11906)
);

NAND2xp5_ASAP7_75t_L g11907 ( 
.A(n_10785),
.B(n_9895),
.Y(n_11907)
);

AND2x2_ASAP7_75t_L g11908 ( 
.A(n_10884),
.B(n_9323),
.Y(n_11908)
);

NAND2x1p5_ASAP7_75t_L g11909 ( 
.A(n_10519),
.B(n_10039),
.Y(n_11909)
);

INVx2_ASAP7_75t_L g11910 ( 
.A(n_10859),
.Y(n_11910)
);

INVx2_ASAP7_75t_L g11911 ( 
.A(n_11212),
.Y(n_11911)
);

AND2x2_ASAP7_75t_L g11912 ( 
.A(n_10842),
.B(n_9323),
.Y(n_11912)
);

AND2x2_ASAP7_75t_L g11913 ( 
.A(n_11000),
.B(n_9375),
.Y(n_11913)
);

INVx2_ASAP7_75t_L g11914 ( 
.A(n_11225),
.Y(n_11914)
);

INVx1_ASAP7_75t_L g11915 ( 
.A(n_11004),
.Y(n_11915)
);

AOI22xp33_ASAP7_75t_SL g11916 ( 
.A1(n_10505),
.A2(n_9609),
.B1(n_9456),
.B2(n_9847),
.Y(n_11916)
);

BUFx3_ASAP7_75t_L g11917 ( 
.A(n_10979),
.Y(n_11917)
);

INVx1_ASAP7_75t_L g11918 ( 
.A(n_10937),
.Y(n_11918)
);

NOR2x1_ASAP7_75t_L g11919 ( 
.A(n_10600),
.B(n_10039),
.Y(n_11919)
);

AND2x2_ASAP7_75t_L g11920 ( 
.A(n_10591),
.B(n_9375),
.Y(n_11920)
);

HB1xp67_ASAP7_75t_L g11921 ( 
.A(n_10575),
.Y(n_11921)
);

AND2x2_ASAP7_75t_L g11922 ( 
.A(n_10581),
.B(n_9375),
.Y(n_11922)
);

INVx1_ASAP7_75t_L g11923 ( 
.A(n_10944),
.Y(n_11923)
);

INVx2_ASAP7_75t_SL g11924 ( 
.A(n_10563),
.Y(n_11924)
);

INVx1_ASAP7_75t_L g11925 ( 
.A(n_10561),
.Y(n_11925)
);

INVx1_ASAP7_75t_L g11926 ( 
.A(n_11083),
.Y(n_11926)
);

INVxp67_ASAP7_75t_SL g11927 ( 
.A(n_10746),
.Y(n_11927)
);

INVx2_ASAP7_75t_SL g11928 ( 
.A(n_10568),
.Y(n_11928)
);

AND2x2_ASAP7_75t_L g11929 ( 
.A(n_10916),
.B(n_9375),
.Y(n_11929)
);

INVx1_ASAP7_75t_L g11930 ( 
.A(n_11163),
.Y(n_11930)
);

BUFx6f_ASAP7_75t_L g11931 ( 
.A(n_10970),
.Y(n_11931)
);

INVx2_ASAP7_75t_L g11932 ( 
.A(n_11048),
.Y(n_11932)
);

INVx3_ASAP7_75t_L g11933 ( 
.A(n_10928),
.Y(n_11933)
);

AND2x4_ASAP7_75t_L g11934 ( 
.A(n_10696),
.B(n_9387),
.Y(n_11934)
);

NOR2x1_ASAP7_75t_SL g11935 ( 
.A(n_10479),
.B(n_9155),
.Y(n_11935)
);

AND2x4_ASAP7_75t_L g11936 ( 
.A(n_10889),
.B(n_9387),
.Y(n_11936)
);

BUFx3_ASAP7_75t_L g11937 ( 
.A(n_10932),
.Y(n_11937)
);

INVx1_ASAP7_75t_L g11938 ( 
.A(n_10557),
.Y(n_11938)
);

AND2x2_ASAP7_75t_L g11939 ( 
.A(n_11100),
.B(n_9387),
.Y(n_11939)
);

AND2x2_ASAP7_75t_L g11940 ( 
.A(n_11109),
.B(n_9387),
.Y(n_11940)
);

INVx1_ASAP7_75t_L g11941 ( 
.A(n_10683),
.Y(n_11941)
);

AND2x2_ASAP7_75t_L g11942 ( 
.A(n_11118),
.B(n_10128),
.Y(n_11942)
);

NAND2xp5_ASAP7_75t_L g11943 ( 
.A(n_10523),
.B(n_10484),
.Y(n_11943)
);

AND2x2_ASAP7_75t_L g11944 ( 
.A(n_11135),
.B(n_10128),
.Y(n_11944)
);

INVx2_ASAP7_75t_L g11945 ( 
.A(n_11142),
.Y(n_11945)
);

HB1xp67_ASAP7_75t_L g11946 ( 
.A(n_10501),
.Y(n_11946)
);

INVx2_ASAP7_75t_L g11947 ( 
.A(n_11202),
.Y(n_11947)
);

INVx1_ASAP7_75t_L g11948 ( 
.A(n_10965),
.Y(n_11948)
);

NAND2xp5_ASAP7_75t_L g11949 ( 
.A(n_10562),
.B(n_9897),
.Y(n_11949)
);

AND2x2_ASAP7_75t_L g11950 ( 
.A(n_10583),
.B(n_10128),
.Y(n_11950)
);

AND2x2_ASAP7_75t_L g11951 ( 
.A(n_10887),
.B(n_10270),
.Y(n_11951)
);

INVx2_ASAP7_75t_L g11952 ( 
.A(n_11205),
.Y(n_11952)
);

INVx1_ASAP7_75t_L g11953 ( 
.A(n_10983),
.Y(n_11953)
);

AND2x2_ASAP7_75t_L g11954 ( 
.A(n_10607),
.B(n_10270),
.Y(n_11954)
);

AND2x2_ASAP7_75t_L g11955 ( 
.A(n_10597),
.B(n_10270),
.Y(n_11955)
);

OR2x2_ASAP7_75t_L g11956 ( 
.A(n_11206),
.B(n_9900),
.Y(n_11956)
);

INVxp67_ASAP7_75t_SL g11957 ( 
.A(n_10921),
.Y(n_11957)
);

INVx2_ASAP7_75t_SL g11958 ( 
.A(n_11207),
.Y(n_11958)
);

INVx1_ASAP7_75t_L g11959 ( 
.A(n_10989),
.Y(n_11959)
);

BUFx2_ASAP7_75t_SL g11960 ( 
.A(n_10903),
.Y(n_11960)
);

AND2x2_ASAP7_75t_L g11961 ( 
.A(n_11019),
.B(n_9281),
.Y(n_11961)
);

BUFx6f_ASAP7_75t_L g11962 ( 
.A(n_10782),
.Y(n_11962)
);

BUFx6f_ASAP7_75t_L g11963 ( 
.A(n_10882),
.Y(n_11963)
);

OR2x2_ASAP7_75t_L g11964 ( 
.A(n_10486),
.B(n_9905),
.Y(n_11964)
);

OR2x2_ASAP7_75t_L g11965 ( 
.A(n_10879),
.B(n_9906),
.Y(n_11965)
);

INVx3_ASAP7_75t_L g11966 ( 
.A(n_10996),
.Y(n_11966)
);

INVx3_ASAP7_75t_L g11967 ( 
.A(n_11219),
.Y(n_11967)
);

BUFx2_ASAP7_75t_L g11968 ( 
.A(n_11027),
.Y(n_11968)
);

BUFx3_ASAP7_75t_L g11969 ( 
.A(n_11191),
.Y(n_11969)
);

AND2x2_ASAP7_75t_L g11970 ( 
.A(n_11021),
.B(n_9281),
.Y(n_11970)
);

OR2x2_ASAP7_75t_L g11971 ( 
.A(n_10482),
.B(n_9908),
.Y(n_11971)
);

INVx1_ASAP7_75t_L g11972 ( 
.A(n_10774),
.Y(n_11972)
);

AND2x2_ASAP7_75t_L g11973 ( 
.A(n_10573),
.B(n_9281),
.Y(n_11973)
);

INVxp67_ASAP7_75t_SL g11974 ( 
.A(n_10936),
.Y(n_11974)
);

AND2x4_ASAP7_75t_L g11975 ( 
.A(n_10992),
.B(n_8788),
.Y(n_11975)
);

NAND2x1_ASAP7_75t_L g11976 ( 
.A(n_10620),
.B(n_9295),
.Y(n_11976)
);

INVx2_ASAP7_75t_L g11977 ( 
.A(n_11199),
.Y(n_11977)
);

INVx1_ASAP7_75t_L g11978 ( 
.A(n_10954),
.Y(n_11978)
);

INVx5_ASAP7_75t_SL g11979 ( 
.A(n_11148),
.Y(n_11979)
);

HB1xp67_ASAP7_75t_L g11980 ( 
.A(n_11088),
.Y(n_11980)
);

AND2x2_ASAP7_75t_L g11981 ( 
.A(n_11011),
.B(n_9295),
.Y(n_11981)
);

NAND2xp5_ASAP7_75t_L g11982 ( 
.A(n_10693),
.B(n_10845),
.Y(n_11982)
);

INVx1_ASAP7_75t_L g11983 ( 
.A(n_10894),
.Y(n_11983)
);

INVx1_ASAP7_75t_L g11984 ( 
.A(n_10902),
.Y(n_11984)
);

INVx2_ASAP7_75t_L g11985 ( 
.A(n_11175),
.Y(n_11985)
);

HB1xp67_ASAP7_75t_L g11986 ( 
.A(n_10601),
.Y(n_11986)
);

BUFx3_ASAP7_75t_L g11987 ( 
.A(n_11141),
.Y(n_11987)
);

INVx1_ASAP7_75t_L g11988 ( 
.A(n_10906),
.Y(n_11988)
);

INVx2_ASAP7_75t_L g11989 ( 
.A(n_11146),
.Y(n_11989)
);

INVx2_ASAP7_75t_L g11990 ( 
.A(n_10898),
.Y(n_11990)
);

AND2x2_ASAP7_75t_L g11991 ( 
.A(n_11123),
.B(n_9295),
.Y(n_11991)
);

NAND2xp5_ASAP7_75t_L g11992 ( 
.A(n_10548),
.B(n_9911),
.Y(n_11992)
);

INVx1_ASAP7_75t_L g11993 ( 
.A(n_10929),
.Y(n_11993)
);

AND2x4_ASAP7_75t_L g11994 ( 
.A(n_11222),
.B(n_8788),
.Y(n_11994)
);

AND2x2_ASAP7_75t_L g11995 ( 
.A(n_11136),
.B(n_9295),
.Y(n_11995)
);

HB1xp67_ASAP7_75t_L g11996 ( 
.A(n_11116),
.Y(n_11996)
);

INVx1_ASAP7_75t_L g11997 ( 
.A(n_10768),
.Y(n_11997)
);

HB1xp67_ASAP7_75t_L g11998 ( 
.A(n_10821),
.Y(n_11998)
);

INVx2_ASAP7_75t_L g11999 ( 
.A(n_10817),
.Y(n_11999)
);

INVx2_ASAP7_75t_L g12000 ( 
.A(n_10676),
.Y(n_12000)
);

INVx1_ASAP7_75t_SL g12001 ( 
.A(n_11286),
.Y(n_12001)
);

INVx2_ASAP7_75t_L g12002 ( 
.A(n_11344),
.Y(n_12002)
);

INVx1_ASAP7_75t_L g12003 ( 
.A(n_11304),
.Y(n_12003)
);

INVx1_ASAP7_75t_L g12004 ( 
.A(n_11337),
.Y(n_12004)
);

INVx2_ASAP7_75t_L g12005 ( 
.A(n_11325),
.Y(n_12005)
);

INVx2_ASAP7_75t_L g12006 ( 
.A(n_11325),
.Y(n_12006)
);

NAND2xp5_ASAP7_75t_L g12007 ( 
.A(n_11241),
.B(n_11076),
.Y(n_12007)
);

INVx1_ASAP7_75t_L g12008 ( 
.A(n_11250),
.Y(n_12008)
);

HB1xp67_ASAP7_75t_L g12009 ( 
.A(n_11239),
.Y(n_12009)
);

INVx1_ASAP7_75t_SL g12010 ( 
.A(n_11240),
.Y(n_12010)
);

INVx1_ASAP7_75t_L g12011 ( 
.A(n_11238),
.Y(n_12011)
);

AND2x2_ASAP7_75t_L g12012 ( 
.A(n_11289),
.B(n_10102),
.Y(n_12012)
);

INVx2_ASAP7_75t_L g12013 ( 
.A(n_11325),
.Y(n_12013)
);

AND2x2_ASAP7_75t_L g12014 ( 
.A(n_11243),
.B(n_10102),
.Y(n_12014)
);

INVx1_ASAP7_75t_SL g12015 ( 
.A(n_11457),
.Y(n_12015)
);

AOI22xp33_ASAP7_75t_L g12016 ( 
.A1(n_11849),
.A2(n_10706),
.B1(n_10892),
.B2(n_10675),
.Y(n_12016)
);

HB1xp67_ASAP7_75t_L g12017 ( 
.A(n_11266),
.Y(n_12017)
);

INVx2_ASAP7_75t_L g12018 ( 
.A(n_11486),
.Y(n_12018)
);

INVx1_ASAP7_75t_L g12019 ( 
.A(n_11238),
.Y(n_12019)
);

NOR2xp33_ASAP7_75t_L g12020 ( 
.A(n_11259),
.B(n_10875),
.Y(n_12020)
);

AND2x2_ASAP7_75t_L g12021 ( 
.A(n_11261),
.B(n_10167),
.Y(n_12021)
);

NOR2xp67_ASAP7_75t_L g12022 ( 
.A(n_11302),
.B(n_10500),
.Y(n_12022)
);

NAND2xp5_ASAP7_75t_L g12023 ( 
.A(n_11281),
.B(n_11104),
.Y(n_12023)
);

INVx2_ASAP7_75t_L g12024 ( 
.A(n_11486),
.Y(n_12024)
);

NOR2x1_ASAP7_75t_L g12025 ( 
.A(n_11689),
.B(n_11121),
.Y(n_12025)
);

INVx1_ASAP7_75t_L g12026 ( 
.A(n_11667),
.Y(n_12026)
);

AND2x2_ASAP7_75t_L g12027 ( 
.A(n_11476),
.B(n_10167),
.Y(n_12027)
);

AND2x4_ASAP7_75t_L g12028 ( 
.A(n_11321),
.B(n_8921),
.Y(n_12028)
);

AOI22xp33_ASAP7_75t_SL g12029 ( 
.A1(n_11849),
.A2(n_11147),
.B1(n_11126),
.B2(n_11209),
.Y(n_12029)
);

AND2x2_ASAP7_75t_L g12030 ( 
.A(n_11476),
.B(n_9156),
.Y(n_12030)
);

NOR2xp33_ASAP7_75t_L g12031 ( 
.A(n_11351),
.B(n_6867),
.Y(n_12031)
);

NAND2xp5_ASAP7_75t_L g12032 ( 
.A(n_11349),
.B(n_10648),
.Y(n_12032)
);

INVx3_ASAP7_75t_L g12033 ( 
.A(n_11254),
.Y(n_12033)
);

AND2x2_ASAP7_75t_L g12034 ( 
.A(n_11444),
.B(n_9156),
.Y(n_12034)
);

INVx1_ASAP7_75t_L g12035 ( 
.A(n_11667),
.Y(n_12035)
);

HB1xp67_ASAP7_75t_L g12036 ( 
.A(n_11275),
.Y(n_12036)
);

OR2x2_ASAP7_75t_L g12037 ( 
.A(n_11267),
.B(n_11248),
.Y(n_12037)
);

INVx1_ASAP7_75t_L g12038 ( 
.A(n_11246),
.Y(n_12038)
);

NOR2xp33_ASAP7_75t_L g12039 ( 
.A(n_11382),
.B(n_6499),
.Y(n_12039)
);

INVx1_ASAP7_75t_L g12040 ( 
.A(n_11246),
.Y(n_12040)
);

NAND2xp5_ASAP7_75t_L g12041 ( 
.A(n_11256),
.B(n_10657),
.Y(n_12041)
);

OAI22xp5_ASAP7_75t_L g12042 ( 
.A1(n_11590),
.A2(n_10849),
.B1(n_10855),
.B2(n_10867),
.Y(n_12042)
);

AOI22xp33_ASAP7_75t_L g12043 ( 
.A1(n_11941),
.A2(n_10893),
.B1(n_10690),
.B2(n_10744),
.Y(n_12043)
);

INVxp67_ASAP7_75t_L g12044 ( 
.A(n_11327),
.Y(n_12044)
);

INVx2_ASAP7_75t_SL g12045 ( 
.A(n_11481),
.Y(n_12045)
);

INVx2_ASAP7_75t_L g12046 ( 
.A(n_11486),
.Y(n_12046)
);

INVxp67_ASAP7_75t_SL g12047 ( 
.A(n_11674),
.Y(n_12047)
);

AND2x2_ASAP7_75t_L g12048 ( 
.A(n_11358),
.B(n_9156),
.Y(n_12048)
);

AND2x2_ASAP7_75t_L g12049 ( 
.A(n_11374),
.B(n_9156),
.Y(n_12049)
);

INVx1_ASAP7_75t_L g12050 ( 
.A(n_11341),
.Y(n_12050)
);

NOR2xp33_ASAP7_75t_L g12051 ( 
.A(n_11302),
.B(n_6542),
.Y(n_12051)
);

NOR2xp33_ASAP7_75t_L g12052 ( 
.A(n_11481),
.B(n_11558),
.Y(n_12052)
);

INVx2_ASAP7_75t_L g12053 ( 
.A(n_11491),
.Y(n_12053)
);

INVx2_ASAP7_75t_L g12054 ( 
.A(n_11491),
.Y(n_12054)
);

AND2x2_ASAP7_75t_L g12055 ( 
.A(n_11271),
.B(n_9156),
.Y(n_12055)
);

INVx1_ASAP7_75t_L g12056 ( 
.A(n_11287),
.Y(n_12056)
);

INVx3_ASAP7_75t_L g12057 ( 
.A(n_11277),
.Y(n_12057)
);

NAND2xp5_ASAP7_75t_L g12058 ( 
.A(n_11927),
.B(n_11972),
.Y(n_12058)
);

INVx1_ASAP7_75t_L g12059 ( 
.A(n_11298),
.Y(n_12059)
);

INVx1_ASAP7_75t_L g12060 ( 
.A(n_11674),
.Y(n_12060)
);

AND2x2_ASAP7_75t_L g12061 ( 
.A(n_11252),
.B(n_9156),
.Y(n_12061)
);

INVx1_ASAP7_75t_L g12062 ( 
.A(n_11687),
.Y(n_12062)
);

AND2x2_ASAP7_75t_L g12063 ( 
.A(n_11258),
.B(n_9186),
.Y(n_12063)
);

INVx2_ASAP7_75t_L g12064 ( 
.A(n_11491),
.Y(n_12064)
);

AND2x4_ASAP7_75t_L g12065 ( 
.A(n_11328),
.B(n_8868),
.Y(n_12065)
);

AND2x2_ASAP7_75t_L g12066 ( 
.A(n_11273),
.B(n_9186),
.Y(n_12066)
);

AND2x2_ASAP7_75t_L g12067 ( 
.A(n_11273),
.B(n_9186),
.Y(n_12067)
);

INVx1_ASAP7_75t_L g12068 ( 
.A(n_11687),
.Y(n_12068)
);

AND2x4_ASAP7_75t_L g12069 ( 
.A(n_11345),
.B(n_9186),
.Y(n_12069)
);

INVx2_ASAP7_75t_L g12070 ( 
.A(n_11572),
.Y(n_12070)
);

HB1xp67_ASAP7_75t_L g12071 ( 
.A(n_11236),
.Y(n_12071)
);

INVx3_ASAP7_75t_L g12072 ( 
.A(n_11572),
.Y(n_12072)
);

AND2x2_ASAP7_75t_L g12073 ( 
.A(n_11402),
.B(n_9186),
.Y(n_12073)
);

INVx3_ASAP7_75t_L g12074 ( 
.A(n_11572),
.Y(n_12074)
);

BUFx3_ASAP7_75t_L g12075 ( 
.A(n_11292),
.Y(n_12075)
);

AND2x2_ASAP7_75t_L g12076 ( 
.A(n_11274),
.B(n_9186),
.Y(n_12076)
);

AND2x2_ASAP7_75t_L g12077 ( 
.A(n_11694),
.B(n_9389),
.Y(n_12077)
);

OR2x2_ASAP7_75t_L g12078 ( 
.A(n_11648),
.B(n_9912),
.Y(n_12078)
);

INVxp67_ASAP7_75t_SL g12079 ( 
.A(n_11407),
.Y(n_12079)
);

INVx1_ASAP7_75t_L g12080 ( 
.A(n_11688),
.Y(n_12080)
);

INVx1_ASAP7_75t_L g12081 ( 
.A(n_11688),
.Y(n_12081)
);

INVx1_ASAP7_75t_L g12082 ( 
.A(n_11743),
.Y(n_12082)
);

INVx2_ASAP7_75t_L g12083 ( 
.A(n_11422),
.Y(n_12083)
);

AND2x2_ASAP7_75t_L g12084 ( 
.A(n_11373),
.B(n_9389),
.Y(n_12084)
);

INVx1_ASAP7_75t_L g12085 ( 
.A(n_11743),
.Y(n_12085)
);

AND2x2_ASAP7_75t_L g12086 ( 
.A(n_11498),
.B(n_9389),
.Y(n_12086)
);

AND2x2_ASAP7_75t_L g12087 ( 
.A(n_11372),
.B(n_11235),
.Y(n_12087)
);

NAND2x1p5_ASAP7_75t_L g12088 ( 
.A(n_11297),
.B(n_8788),
.Y(n_12088)
);

INVx1_ASAP7_75t_L g12089 ( 
.A(n_11748),
.Y(n_12089)
);

INVx2_ASAP7_75t_L g12090 ( 
.A(n_11569),
.Y(n_12090)
);

INVx1_ASAP7_75t_L g12091 ( 
.A(n_11748),
.Y(n_12091)
);

AND2x2_ASAP7_75t_L g12092 ( 
.A(n_11291),
.B(n_9389),
.Y(n_12092)
);

AND2x2_ASAP7_75t_L g12093 ( 
.A(n_11583),
.B(n_9389),
.Y(n_12093)
);

AOI22xp33_ASAP7_75t_L g12094 ( 
.A1(n_11941),
.A2(n_10891),
.B1(n_10873),
.B2(n_10713),
.Y(n_12094)
);

AND2x2_ASAP7_75t_L g12095 ( 
.A(n_11428),
.B(n_9389),
.Y(n_12095)
);

INVx1_ASAP7_75t_L g12096 ( 
.A(n_11750),
.Y(n_12096)
);

AND2x2_ASAP7_75t_L g12097 ( 
.A(n_11429),
.B(n_9432),
.Y(n_12097)
);

HB1xp67_ASAP7_75t_L g12098 ( 
.A(n_11255),
.Y(n_12098)
);

AND2x2_ASAP7_75t_L g12099 ( 
.A(n_11430),
.B(n_9432),
.Y(n_12099)
);

OAI221xp5_ASAP7_75t_SL g12100 ( 
.A1(n_11606),
.A2(n_10619),
.B1(n_10614),
.B2(n_10872),
.C(n_10869),
.Y(n_12100)
);

AND2x2_ASAP7_75t_L g12101 ( 
.A(n_11268),
.B(n_9432),
.Y(n_12101)
);

BUFx2_ASAP7_75t_SL g12102 ( 
.A(n_11481),
.Y(n_12102)
);

INVx2_ASAP7_75t_L g12103 ( 
.A(n_11560),
.Y(n_12103)
);

INVx1_ASAP7_75t_SL g12104 ( 
.A(n_11380),
.Y(n_12104)
);

BUFx3_ASAP7_75t_L g12105 ( 
.A(n_11580),
.Y(n_12105)
);

AND2x2_ASAP7_75t_L g12106 ( 
.A(n_11269),
.B(n_11278),
.Y(n_12106)
);

AND2x2_ASAP7_75t_L g12107 ( 
.A(n_11282),
.B(n_9432),
.Y(n_12107)
);

INVx1_ASAP7_75t_L g12108 ( 
.A(n_11750),
.Y(n_12108)
);

AND2x2_ASAP7_75t_L g12109 ( 
.A(n_11299),
.B(n_9432),
.Y(n_12109)
);

INVx1_ASAP7_75t_L g12110 ( 
.A(n_11751),
.Y(n_12110)
);

INVx1_ASAP7_75t_L g12111 ( 
.A(n_11751),
.Y(n_12111)
);

INVx1_ASAP7_75t_L g12112 ( 
.A(n_11695),
.Y(n_12112)
);

AND2x2_ASAP7_75t_L g12113 ( 
.A(n_11306),
.B(n_9432),
.Y(n_12113)
);

OR2x2_ASAP7_75t_L g12114 ( 
.A(n_11359),
.B(n_9913),
.Y(n_12114)
);

INVx1_ASAP7_75t_L g12115 ( 
.A(n_11698),
.Y(n_12115)
);

INVx1_ASAP7_75t_L g12116 ( 
.A(n_11362),
.Y(n_12116)
);

INVx2_ASAP7_75t_L g12117 ( 
.A(n_11560),
.Y(n_12117)
);

INVx4_ASAP7_75t_L g12118 ( 
.A(n_11380),
.Y(n_12118)
);

AND2x2_ASAP7_75t_L g12119 ( 
.A(n_11307),
.B(n_9434),
.Y(n_12119)
);

INVx2_ASAP7_75t_L g12120 ( 
.A(n_11589),
.Y(n_12120)
);

INVx2_ASAP7_75t_L g12121 ( 
.A(n_11297),
.Y(n_12121)
);

AND2x2_ASAP7_75t_L g12122 ( 
.A(n_11244),
.B(n_9434),
.Y(n_12122)
);

OR2x2_ASAP7_75t_L g12123 ( 
.A(n_11704),
.B(n_9917),
.Y(n_12123)
);

INVx2_ASAP7_75t_L g12124 ( 
.A(n_11297),
.Y(n_12124)
);

INVx2_ASAP7_75t_L g12125 ( 
.A(n_11311),
.Y(n_12125)
);

AND2x4_ASAP7_75t_SL g12126 ( 
.A(n_11390),
.B(n_8040),
.Y(n_12126)
);

INVx1_ASAP7_75t_L g12127 ( 
.A(n_11367),
.Y(n_12127)
);

AOI22xp33_ASAP7_75t_L g12128 ( 
.A1(n_11899),
.A2(n_10705),
.B1(n_10697),
.B2(n_10745),
.Y(n_12128)
);

NOR2xp33_ASAP7_75t_L g12129 ( 
.A(n_11480),
.B(n_6771),
.Y(n_12129)
);

AND2x4_ASAP7_75t_L g12130 ( 
.A(n_11315),
.B(n_9434),
.Y(n_12130)
);

HB1xp67_ASAP7_75t_L g12131 ( 
.A(n_11760),
.Y(n_12131)
);

AOI22xp33_ASAP7_75t_L g12132 ( 
.A1(n_11899),
.A2(n_10763),
.B1(n_10528),
.B2(n_10503),
.Y(n_12132)
);

INVx1_ASAP7_75t_L g12133 ( 
.A(n_11370),
.Y(n_12133)
);

NAND2xp5_ASAP7_75t_L g12134 ( 
.A(n_11972),
.B(n_10669),
.Y(n_12134)
);

INVx1_ASAP7_75t_L g12135 ( 
.A(n_11376),
.Y(n_12135)
);

AND2x2_ASAP7_75t_L g12136 ( 
.A(n_11360),
.B(n_9434),
.Y(n_12136)
);

INVx1_ASAP7_75t_L g12137 ( 
.A(n_11378),
.Y(n_12137)
);

AND2x2_ASAP7_75t_L g12138 ( 
.A(n_11242),
.B(n_9434),
.Y(n_12138)
);

INVx1_ASAP7_75t_L g12139 ( 
.A(n_11303),
.Y(n_12139)
);

INVx1_ASAP7_75t_L g12140 ( 
.A(n_11704),
.Y(n_12140)
);

INVx1_ASAP7_75t_L g12141 ( 
.A(n_11257),
.Y(n_12141)
);

NAND2xp5_ASAP7_75t_L g12142 ( 
.A(n_11847),
.B(n_11187),
.Y(n_12142)
);

OR2x2_ASAP7_75t_L g12143 ( 
.A(n_11724),
.B(n_9920),
.Y(n_12143)
);

AND2x4_ASAP7_75t_L g12144 ( 
.A(n_11315),
.B(n_9434),
.Y(n_12144)
);

AND2x2_ASAP7_75t_L g12145 ( 
.A(n_11493),
.B(n_9042),
.Y(n_12145)
);

AND2x4_ASAP7_75t_L g12146 ( 
.A(n_11245),
.B(n_8788),
.Y(n_12146)
);

INVx1_ASAP7_75t_L g12147 ( 
.A(n_11257),
.Y(n_12147)
);

AND2x2_ASAP7_75t_L g12148 ( 
.A(n_11497),
.B(n_9042),
.Y(n_12148)
);

AND2x2_ASAP7_75t_L g12149 ( 
.A(n_11499),
.B(n_9050),
.Y(n_12149)
);

INVxp67_ASAP7_75t_SL g12150 ( 
.A(n_11265),
.Y(n_12150)
);

INVx1_ASAP7_75t_L g12151 ( 
.A(n_11272),
.Y(n_12151)
);

OAI222xp33_ASAP7_75t_L g12152 ( 
.A1(n_11827),
.A2(n_11074),
.B1(n_10635),
.B2(n_10595),
.C1(n_11221),
.C2(n_11210),
.Y(n_12152)
);

INVx1_ASAP7_75t_L g12153 ( 
.A(n_11272),
.Y(n_12153)
);

INVx1_ASAP7_75t_L g12154 ( 
.A(n_11280),
.Y(n_12154)
);

AND2x2_ASAP7_75t_L g12155 ( 
.A(n_11400),
.B(n_9050),
.Y(n_12155)
);

INVx1_ASAP7_75t_L g12156 ( 
.A(n_11280),
.Y(n_12156)
);

AOI22xp33_ASAP7_75t_L g12157 ( 
.A1(n_11892),
.A2(n_10680),
.B1(n_10492),
.B2(n_10602),
.Y(n_12157)
);

INVx3_ASAP7_75t_L g12158 ( 
.A(n_11390),
.Y(n_12158)
);

INVx2_ASAP7_75t_L g12159 ( 
.A(n_11311),
.Y(n_12159)
);

INVx1_ASAP7_75t_L g12160 ( 
.A(n_11294),
.Y(n_12160)
);

NAND2xp5_ASAP7_75t_L g12161 ( 
.A(n_11847),
.B(n_10946),
.Y(n_12161)
);

HB1xp67_ASAP7_75t_L g12162 ( 
.A(n_11253),
.Y(n_12162)
);

INVx2_ASAP7_75t_L g12163 ( 
.A(n_11318),
.Y(n_12163)
);

AND2x2_ASAP7_75t_L g12164 ( 
.A(n_11316),
.B(n_9105),
.Y(n_12164)
);

INVx1_ASAP7_75t_L g12165 ( 
.A(n_11294),
.Y(n_12165)
);

BUFx2_ASAP7_75t_L g12166 ( 
.A(n_11263),
.Y(n_12166)
);

INVx1_ASAP7_75t_L g12167 ( 
.A(n_11295),
.Y(n_12167)
);

INVx1_ASAP7_75t_L g12168 ( 
.A(n_11295),
.Y(n_12168)
);

INVx1_ASAP7_75t_L g12169 ( 
.A(n_11300),
.Y(n_12169)
);

AND2x2_ASAP7_75t_L g12170 ( 
.A(n_11526),
.B(n_9105),
.Y(n_12170)
);

OR2x2_ASAP7_75t_SL g12171 ( 
.A(n_11831),
.B(n_9341),
.Y(n_12171)
);

INVx3_ASAP7_75t_L g12172 ( 
.A(n_11480),
.Y(n_12172)
);

OAI22xp5_ASAP7_75t_L g12173 ( 
.A1(n_11979),
.A2(n_11647),
.B1(n_11735),
.B2(n_11801),
.Y(n_12173)
);

INVx2_ASAP7_75t_L g12174 ( 
.A(n_11318),
.Y(n_12174)
);

INVx3_ASAP7_75t_L g12175 ( 
.A(n_11554),
.Y(n_12175)
);

AND2x2_ASAP7_75t_L g12176 ( 
.A(n_11527),
.B(n_9131),
.Y(n_12176)
);

INVx2_ASAP7_75t_L g12177 ( 
.A(n_11384),
.Y(n_12177)
);

INVx2_ASAP7_75t_L g12178 ( 
.A(n_11384),
.Y(n_12178)
);

OAI221xp5_ASAP7_75t_L g12179 ( 
.A1(n_11807),
.A2(n_10856),
.B1(n_10957),
.B2(n_10958),
.C(n_10917),
.Y(n_12179)
);

OR2x2_ASAP7_75t_L g12180 ( 
.A(n_11725),
.B(n_9924),
.Y(n_12180)
);

INVx1_ASAP7_75t_L g12181 ( 
.A(n_11300),
.Y(n_12181)
);

AND2x2_ASAP7_75t_L g12182 ( 
.A(n_11528),
.B(n_9131),
.Y(n_12182)
);

OR2x2_ASAP7_75t_L g12183 ( 
.A(n_11725),
.B(n_9929),
.Y(n_12183)
);

INVx1_ASAP7_75t_L g12184 ( 
.A(n_11314),
.Y(n_12184)
);

NAND2xp5_ASAP7_75t_L g12185 ( 
.A(n_11726),
.B(n_9931),
.Y(n_12185)
);

INVx1_ASAP7_75t_L g12186 ( 
.A(n_11314),
.Y(n_12186)
);

NOR2xp33_ASAP7_75t_L g12187 ( 
.A(n_11554),
.B(n_6771),
.Y(n_12187)
);

NAND2xp5_ASAP7_75t_L g12188 ( 
.A(n_11726),
.B(n_9933),
.Y(n_12188)
);

AND2x2_ASAP7_75t_L g12189 ( 
.A(n_11535),
.B(n_9151),
.Y(n_12189)
);

INVx1_ASAP7_75t_L g12190 ( 
.A(n_11317),
.Y(n_12190)
);

AND2x2_ASAP7_75t_L g12191 ( 
.A(n_11433),
.B(n_9151),
.Y(n_12191)
);

INVx2_ASAP7_75t_L g12192 ( 
.A(n_11385),
.Y(n_12192)
);

NAND3xp33_ASAP7_75t_L g12193 ( 
.A(n_11978),
.B(n_11198),
.C(n_11216),
.Y(n_12193)
);

AND2x2_ASAP7_75t_L g12194 ( 
.A(n_11714),
.B(n_9160),
.Y(n_12194)
);

INVx2_ASAP7_75t_L g12195 ( 
.A(n_11385),
.Y(n_12195)
);

OAI22xp5_ASAP7_75t_L g12196 ( 
.A1(n_11979),
.A2(n_11158),
.B1(n_11149),
.B2(n_10587),
.Y(n_12196)
);

AOI22xp33_ASAP7_75t_L g12197 ( 
.A1(n_11892),
.A2(n_10789),
.B1(n_11068),
.B2(n_11047),
.Y(n_12197)
);

NAND2xp5_ASAP7_75t_L g12198 ( 
.A(n_11978),
.B(n_9935),
.Y(n_12198)
);

OAI22xp5_ASAP7_75t_L g12199 ( 
.A1(n_11562),
.A2(n_10513),
.B1(n_11137),
.B2(n_10776),
.Y(n_12199)
);

AND2x2_ASAP7_75t_L g12200 ( 
.A(n_11617),
.B(n_11449),
.Y(n_12200)
);

INVx1_ASAP7_75t_L g12201 ( 
.A(n_11317),
.Y(n_12201)
);

INVx1_ASAP7_75t_L g12202 ( 
.A(n_11331),
.Y(n_12202)
);

INVx1_ASAP7_75t_L g12203 ( 
.A(n_11331),
.Y(n_12203)
);

INVx1_ASAP7_75t_L g12204 ( 
.A(n_11335),
.Y(n_12204)
);

AOI22xp33_ASAP7_75t_L g12205 ( 
.A1(n_11897),
.A2(n_10786),
.B1(n_11073),
.B2(n_11091),
.Y(n_12205)
);

AND2x2_ASAP7_75t_L g12206 ( 
.A(n_11425),
.B(n_9160),
.Y(n_12206)
);

INVx3_ASAP7_75t_L g12207 ( 
.A(n_11603),
.Y(n_12207)
);

AND2x2_ASAP7_75t_L g12208 ( 
.A(n_11598),
.B(n_9165),
.Y(n_12208)
);

OR2x2_ASAP7_75t_L g12209 ( 
.A(n_11669),
.B(n_11264),
.Y(n_12209)
);

INVx1_ASAP7_75t_L g12210 ( 
.A(n_11335),
.Y(n_12210)
);

NAND2xp5_ASAP7_75t_L g12211 ( 
.A(n_11488),
.B(n_9939),
.Y(n_12211)
);

NAND2xp5_ASAP7_75t_L g12212 ( 
.A(n_11496),
.B(n_9947),
.Y(n_12212)
);

INVx1_ASAP7_75t_L g12213 ( 
.A(n_11339),
.Y(n_12213)
);

INVx2_ASAP7_75t_L g12214 ( 
.A(n_11443),
.Y(n_12214)
);

INVx2_ASAP7_75t_L g12215 ( 
.A(n_11446),
.Y(n_12215)
);

INVx2_ASAP7_75t_L g12216 ( 
.A(n_11270),
.Y(n_12216)
);

OR2x2_ASAP7_75t_SL g12217 ( 
.A(n_11734),
.B(n_9363),
.Y(n_12217)
);

INVx1_ASAP7_75t_L g12218 ( 
.A(n_11339),
.Y(n_12218)
);

AND2x2_ASAP7_75t_L g12219 ( 
.A(n_11598),
.B(n_9165),
.Y(n_12219)
);

OR2x2_ASAP7_75t_L g12220 ( 
.A(n_11948),
.B(n_9952),
.Y(n_12220)
);

HB1xp67_ASAP7_75t_L g12221 ( 
.A(n_11309),
.Y(n_12221)
);

INVx1_ASAP7_75t_L g12222 ( 
.A(n_11340),
.Y(n_12222)
);

INVx1_ASAP7_75t_L g12223 ( 
.A(n_11340),
.Y(n_12223)
);

NAND2x1_ASAP7_75t_L g12224 ( 
.A(n_11975),
.B(n_10113),
.Y(n_12224)
);

INVx1_ASAP7_75t_L g12225 ( 
.A(n_11389),
.Y(n_12225)
);

AND2x2_ASAP7_75t_L g12226 ( 
.A(n_11841),
.B(n_9207),
.Y(n_12226)
);

BUFx2_ASAP7_75t_L g12227 ( 
.A(n_11263),
.Y(n_12227)
);

OAI22xp5_ASAP7_75t_L g12228 ( 
.A1(n_11553),
.A2(n_10552),
.B1(n_10850),
.B2(n_11081),
.Y(n_12228)
);

INVx1_ASAP7_75t_L g12229 ( 
.A(n_11389),
.Y(n_12229)
);

AND2x2_ASAP7_75t_L g12230 ( 
.A(n_11519),
.B(n_9207),
.Y(n_12230)
);

INVx2_ASAP7_75t_L g12231 ( 
.A(n_11355),
.Y(n_12231)
);

AND2x4_ASAP7_75t_L g12232 ( 
.A(n_11413),
.B(n_6779),
.Y(n_12232)
);

NAND2xp5_ASAP7_75t_L g12233 ( 
.A(n_11627),
.B(n_9956),
.Y(n_12233)
);

NOR2x1_ASAP7_75t_L g12234 ( 
.A(n_11593),
.B(n_8860),
.Y(n_12234)
);

NAND2xp5_ASAP7_75t_L g12235 ( 
.A(n_11998),
.B(n_9961),
.Y(n_12235)
);

INVx1_ASAP7_75t_L g12236 ( 
.A(n_11401),
.Y(n_12236)
);

NAND2xp5_ASAP7_75t_L g12237 ( 
.A(n_11887),
.B(n_9963),
.Y(n_12237)
);

NAND2xp5_ASAP7_75t_SL g12238 ( 
.A(n_11975),
.B(n_10674),
.Y(n_12238)
);

NAND2xp5_ASAP7_75t_L g12239 ( 
.A(n_11515),
.B(n_11541),
.Y(n_12239)
);

INVx1_ASAP7_75t_L g12240 ( 
.A(n_11401),
.Y(n_12240)
);

NAND2xp5_ASAP7_75t_SL g12241 ( 
.A(n_11933),
.B(n_11936),
.Y(n_12241)
);

INVx2_ASAP7_75t_SL g12242 ( 
.A(n_11603),
.Y(n_12242)
);

AND2x4_ASAP7_75t_L g12243 ( 
.A(n_11413),
.B(n_6779),
.Y(n_12243)
);

AND2x2_ASAP7_75t_L g12244 ( 
.A(n_11520),
.B(n_9214),
.Y(n_12244)
);

AND2x2_ASAP7_75t_L g12245 ( 
.A(n_11521),
.B(n_9214),
.Y(n_12245)
);

HB1xp67_ASAP7_75t_L g12246 ( 
.A(n_11260),
.Y(n_12246)
);

INVx1_ASAP7_75t_L g12247 ( 
.A(n_11404),
.Y(n_12247)
);

AND2x4_ASAP7_75t_L g12248 ( 
.A(n_11427),
.B(n_6272),
.Y(n_12248)
);

INVxp67_ASAP7_75t_SL g12249 ( 
.A(n_11701),
.Y(n_12249)
);

HB1xp67_ASAP7_75t_L g12250 ( 
.A(n_11249),
.Y(n_12250)
);

NAND2xp5_ASAP7_75t_L g12251 ( 
.A(n_11557),
.B(n_9967),
.Y(n_12251)
);

AND2x2_ASAP7_75t_L g12252 ( 
.A(n_11276),
.B(n_9217),
.Y(n_12252)
);

NOR2xp67_ASAP7_75t_L g12253 ( 
.A(n_11460),
.B(n_9125),
.Y(n_12253)
);

INVx1_ASAP7_75t_L g12254 ( 
.A(n_11404),
.Y(n_12254)
);

NAND2xp5_ASAP7_75t_L g12255 ( 
.A(n_11559),
.B(n_11637),
.Y(n_12255)
);

INVxp33_ASAP7_75t_SL g12256 ( 
.A(n_11551),
.Y(n_12256)
);

AND2x2_ASAP7_75t_L g12257 ( 
.A(n_11276),
.B(n_9217),
.Y(n_12257)
);

AND2x2_ASAP7_75t_L g12258 ( 
.A(n_11477),
.B(n_9222),
.Y(n_12258)
);

INVx1_ASAP7_75t_L g12259 ( 
.A(n_11405),
.Y(n_12259)
);

INVx2_ASAP7_75t_SL g12260 ( 
.A(n_11603),
.Y(n_12260)
);

INVx1_ASAP7_75t_L g12261 ( 
.A(n_11405),
.Y(n_12261)
);

AOI22xp33_ASAP7_75t_L g12262 ( 
.A1(n_11897),
.A2(n_11085),
.B1(n_11003),
.B2(n_9858),
.Y(n_12262)
);

INVx3_ASAP7_75t_L g12263 ( 
.A(n_11539),
.Y(n_12263)
);

NOR2xp67_ASAP7_75t_L g12264 ( 
.A(n_11463),
.B(n_9128),
.Y(n_12264)
);

INVx3_ASAP7_75t_SL g12265 ( 
.A(n_11334),
.Y(n_12265)
);

INVx1_ASAP7_75t_L g12266 ( 
.A(n_11406),
.Y(n_12266)
);

INVx1_ASAP7_75t_L g12267 ( 
.A(n_11406),
.Y(n_12267)
);

NAND2xp5_ASAP7_75t_L g12268 ( 
.A(n_11395),
.B(n_9974),
.Y(n_12268)
);

NAND2x1_ASAP7_75t_L g12269 ( 
.A(n_11936),
.B(n_10121),
.Y(n_12269)
);

AND2x2_ASAP7_75t_L g12270 ( 
.A(n_11479),
.B(n_9222),
.Y(n_12270)
);

CKINVDCx14_ASAP7_75t_R g12271 ( 
.A(n_11660),
.Y(n_12271)
);

INVx1_ASAP7_75t_L g12272 ( 
.A(n_11431),
.Y(n_12272)
);

AND2x2_ASAP7_75t_L g12273 ( 
.A(n_11464),
.B(n_9240),
.Y(n_12273)
);

OR2x2_ASAP7_75t_L g12274 ( 
.A(n_11948),
.B(n_9977),
.Y(n_12274)
);

INVx2_ASAP7_75t_L g12275 ( 
.A(n_11364),
.Y(n_12275)
);

INVx1_ASAP7_75t_L g12276 ( 
.A(n_11431),
.Y(n_12276)
);

AND2x2_ASAP7_75t_L g12277 ( 
.A(n_11588),
.B(n_11330),
.Y(n_12277)
);

INVx2_ASAP7_75t_L g12278 ( 
.A(n_11366),
.Y(n_12278)
);

INVx1_ASAP7_75t_L g12279 ( 
.A(n_11437),
.Y(n_12279)
);

INVx2_ASAP7_75t_L g12280 ( 
.A(n_11377),
.Y(n_12280)
);

INVx1_ASAP7_75t_L g12281 ( 
.A(n_11437),
.Y(n_12281)
);

AND2x2_ASAP7_75t_L g12282 ( 
.A(n_11336),
.B(n_9240),
.Y(n_12282)
);

INVx2_ASAP7_75t_SL g12283 ( 
.A(n_11605),
.Y(n_12283)
);

INVx1_ASAP7_75t_L g12284 ( 
.A(n_11440),
.Y(n_12284)
);

NAND2xp5_ASAP7_75t_L g12285 ( 
.A(n_11415),
.B(n_9980),
.Y(n_12285)
);

HB1xp67_ASAP7_75t_L g12286 ( 
.A(n_11573),
.Y(n_12286)
);

AND2x2_ASAP7_75t_L g12287 ( 
.A(n_11312),
.B(n_9304),
.Y(n_12287)
);

INVx2_ASAP7_75t_L g12288 ( 
.A(n_11575),
.Y(n_12288)
);

AND2x2_ASAP7_75t_L g12289 ( 
.A(n_11550),
.B(n_9304),
.Y(n_12289)
);

NAND2xp5_ASAP7_75t_L g12290 ( 
.A(n_11484),
.B(n_9983),
.Y(n_12290)
);

INVx2_ASAP7_75t_L g12291 ( 
.A(n_11586),
.Y(n_12291)
);

INVx1_ASAP7_75t_L g12292 ( 
.A(n_11440),
.Y(n_12292)
);

AND2x4_ASAP7_75t_L g12293 ( 
.A(n_11427),
.B(n_6353),
.Y(n_12293)
);

AND2x2_ASAP7_75t_L g12294 ( 
.A(n_11576),
.B(n_9396),
.Y(n_12294)
);

AND2x4_ASAP7_75t_L g12295 ( 
.A(n_11448),
.B(n_6353),
.Y(n_12295)
);

INVx2_ASAP7_75t_L g12296 ( 
.A(n_11592),
.Y(n_12296)
);

HB1xp67_ASAP7_75t_L g12297 ( 
.A(n_11600),
.Y(n_12297)
);

AND2x2_ASAP7_75t_L g12298 ( 
.A(n_11578),
.B(n_9396),
.Y(n_12298)
);

HB1xp67_ASAP7_75t_L g12299 ( 
.A(n_11450),
.Y(n_12299)
);

INVx1_ASAP7_75t_L g12300 ( 
.A(n_11701),
.Y(n_12300)
);

NAND2xp5_ASAP7_75t_L g12301 ( 
.A(n_11512),
.B(n_11902),
.Y(n_12301)
);

INVx2_ASAP7_75t_SL g12302 ( 
.A(n_11448),
.Y(n_12302)
);

INVx1_ASAP7_75t_L g12303 ( 
.A(n_11703),
.Y(n_12303)
);

INVx2_ASAP7_75t_SL g12304 ( 
.A(n_11503),
.Y(n_12304)
);

INVx1_ASAP7_75t_L g12305 ( 
.A(n_11703),
.Y(n_12305)
);

NAND2xp5_ASAP7_75t_L g12306 ( 
.A(n_11902),
.B(n_9985),
.Y(n_12306)
);

INVxp67_ASAP7_75t_SL g12307 ( 
.A(n_11279),
.Y(n_12307)
);

AND2x4_ASAP7_75t_L g12308 ( 
.A(n_11471),
.B(n_7077),
.Y(n_12308)
);

AND2x2_ASAP7_75t_L g12309 ( 
.A(n_11581),
.B(n_9397),
.Y(n_12309)
);

NAND2xp5_ASAP7_75t_L g12310 ( 
.A(n_11903),
.B(n_9988),
.Y(n_12310)
);

INVxp67_ASAP7_75t_SL g12311 ( 
.A(n_11680),
.Y(n_12311)
);

INVx1_ASAP7_75t_L g12312 ( 
.A(n_11752),
.Y(n_12312)
);

INVx1_ASAP7_75t_L g12313 ( 
.A(n_11752),
.Y(n_12313)
);

INVx2_ASAP7_75t_SL g12314 ( 
.A(n_11471),
.Y(n_12314)
);

NAND2xp5_ASAP7_75t_L g12315 ( 
.A(n_11903),
.B(n_9994),
.Y(n_12315)
);

INVx1_ASAP7_75t_L g12316 ( 
.A(n_11447),
.Y(n_12316)
);

INVx2_ASAP7_75t_L g12317 ( 
.A(n_11322),
.Y(n_12317)
);

AND2x2_ASAP7_75t_L g12318 ( 
.A(n_11343),
.B(n_9397),
.Y(n_12318)
);

INVxp67_ASAP7_75t_L g12319 ( 
.A(n_11538),
.Y(n_12319)
);

HB1xp67_ASAP7_75t_L g12320 ( 
.A(n_11453),
.Y(n_12320)
);

CKINVDCx5p33_ASAP7_75t_R g12321 ( 
.A(n_11320),
.Y(n_12321)
);

INVx2_ASAP7_75t_L g12322 ( 
.A(n_11323),
.Y(n_12322)
);

OR2x2_ASAP7_75t_L g12323 ( 
.A(n_11953),
.B(n_9996),
.Y(n_12323)
);

INVx2_ASAP7_75t_L g12324 ( 
.A(n_11612),
.Y(n_12324)
);

INVx2_ASAP7_75t_L g12325 ( 
.A(n_11612),
.Y(n_12325)
);

INVx1_ASAP7_75t_L g12326 ( 
.A(n_11447),
.Y(n_12326)
);

AND2x2_ASAP7_75t_L g12327 ( 
.A(n_11347),
.B(n_9411),
.Y(n_12327)
);

AOI22xp33_ASAP7_75t_L g12328 ( 
.A1(n_11898),
.A2(n_9857),
.B1(n_11072),
.B2(n_10771),
.Y(n_12328)
);

AND2x2_ASAP7_75t_L g12329 ( 
.A(n_11348),
.B(n_9411),
.Y(n_12329)
);

NAND2xp5_ASAP7_75t_L g12330 ( 
.A(n_11489),
.B(n_9998),
.Y(n_12330)
);

INVxp67_ASAP7_75t_SL g12331 ( 
.A(n_11468),
.Y(n_12331)
);

AND2x2_ASAP7_75t_L g12332 ( 
.A(n_11350),
.B(n_8860),
.Y(n_12332)
);

INVx3_ASAP7_75t_L g12333 ( 
.A(n_11539),
.Y(n_12333)
);

INVx2_ASAP7_75t_L g12334 ( 
.A(n_11796),
.Y(n_12334)
);

NAND2xp5_ASAP7_75t_L g12335 ( 
.A(n_11494),
.B(n_9999),
.Y(n_12335)
);

OR2x2_ASAP7_75t_L g12336 ( 
.A(n_11953),
.B(n_10001),
.Y(n_12336)
);

NAND2xp5_ASAP7_75t_L g12337 ( 
.A(n_11644),
.B(n_10003),
.Y(n_12337)
);

AND2x2_ASAP7_75t_L g12338 ( 
.A(n_11352),
.B(n_9091),
.Y(n_12338)
);

INVx2_ASAP7_75t_L g12339 ( 
.A(n_11796),
.Y(n_12339)
);

AND2x2_ASAP7_75t_L g12340 ( 
.A(n_11308),
.B(n_11451),
.Y(n_12340)
);

AND2x2_ASAP7_75t_L g12341 ( 
.A(n_11459),
.B(n_9091),
.Y(n_12341)
);

NAND2xp5_ASAP7_75t_L g12342 ( 
.A(n_11607),
.B(n_10005),
.Y(n_12342)
);

AND2x2_ASAP7_75t_L g12343 ( 
.A(n_11462),
.B(n_11342),
.Y(n_12343)
);

NAND2xp5_ASAP7_75t_L g12344 ( 
.A(n_11608),
.B(n_11671),
.Y(n_12344)
);

BUFx8_ASAP7_75t_SL g12345 ( 
.A(n_11525),
.Y(n_12345)
);

BUFx6f_ASAP7_75t_L g12346 ( 
.A(n_11455),
.Y(n_12346)
);

INVxp67_ASAP7_75t_SL g12347 ( 
.A(n_11980),
.Y(n_12347)
);

INVx1_ASAP7_75t_L g12348 ( 
.A(n_11456),
.Y(n_12348)
);

INVx2_ASAP7_75t_L g12349 ( 
.A(n_11796),
.Y(n_12349)
);

INVx1_ASAP7_75t_SL g12350 ( 
.A(n_11284),
.Y(n_12350)
);

OR2x2_ASAP7_75t_L g12351 ( 
.A(n_11959),
.B(n_10006),
.Y(n_12351)
);

HB1xp67_ASAP7_75t_L g12352 ( 
.A(n_11619),
.Y(n_12352)
);

OR2x2_ASAP7_75t_L g12353 ( 
.A(n_11959),
.B(n_10011),
.Y(n_12353)
);

BUFx2_ASAP7_75t_L g12354 ( 
.A(n_11670),
.Y(n_12354)
);

AND2x4_ASAP7_75t_L g12355 ( 
.A(n_11517),
.B(n_7077),
.Y(n_12355)
);

AND2x2_ASAP7_75t_L g12356 ( 
.A(n_11466),
.B(n_9162),
.Y(n_12356)
);

INVx1_ASAP7_75t_L g12357 ( 
.A(n_11456),
.Y(n_12357)
);

BUFx3_ASAP7_75t_L g12358 ( 
.A(n_11458),
.Y(n_12358)
);

INVx2_ASAP7_75t_L g12359 ( 
.A(n_11733),
.Y(n_12359)
);

AO22x1_ASAP7_75t_L g12360 ( 
.A1(n_11641),
.A2(n_4175),
.B1(n_4226),
.B2(n_4164),
.Y(n_12360)
);

BUFx2_ASAP7_75t_L g12361 ( 
.A(n_11833),
.Y(n_12361)
);

INVx1_ASAP7_75t_L g12362 ( 
.A(n_11465),
.Y(n_12362)
);

INVx1_ASAP7_75t_L g12363 ( 
.A(n_11465),
.Y(n_12363)
);

INVx2_ASAP7_75t_SL g12364 ( 
.A(n_11604),
.Y(n_12364)
);

AND2x2_ASAP7_75t_L g12365 ( 
.A(n_11371),
.B(n_9162),
.Y(n_12365)
);

AND2x2_ASAP7_75t_L g12366 ( 
.A(n_11353),
.B(n_11356),
.Y(n_12366)
);

NOR2xp67_ASAP7_75t_L g12367 ( 
.A(n_11290),
.B(n_9188),
.Y(n_12367)
);

AND2x2_ASAP7_75t_L g12368 ( 
.A(n_11361),
.B(n_11363),
.Y(n_12368)
);

AND2x2_ASAP7_75t_L g12369 ( 
.A(n_11365),
.B(n_9212),
.Y(n_12369)
);

AND2x2_ASAP7_75t_L g12370 ( 
.A(n_11326),
.B(n_9212),
.Y(n_12370)
);

INVx1_ASAP7_75t_L g12371 ( 
.A(n_11469),
.Y(n_12371)
);

CKINVDCx20_ASAP7_75t_R g12372 ( 
.A(n_11591),
.Y(n_12372)
);

AND2x2_ASAP7_75t_L g12373 ( 
.A(n_11410),
.B(n_8786),
.Y(n_12373)
);

INVx2_ASAP7_75t_L g12374 ( 
.A(n_11749),
.Y(n_12374)
);

INVx1_ASAP7_75t_L g12375 ( 
.A(n_11469),
.Y(n_12375)
);

AND2x2_ASAP7_75t_SL g12376 ( 
.A(n_11643),
.B(n_7951),
.Y(n_12376)
);

INVx2_ASAP7_75t_L g12377 ( 
.A(n_11283),
.Y(n_12377)
);

AND2x2_ASAP7_75t_L g12378 ( 
.A(n_11411),
.B(n_11414),
.Y(n_12378)
);

HB1xp67_ASAP7_75t_L g12379 ( 
.A(n_11237),
.Y(n_12379)
);

INVx1_ASAP7_75t_SL g12380 ( 
.A(n_11518),
.Y(n_12380)
);

OAI22xp5_ASAP7_75t_L g12381 ( 
.A1(n_11857),
.A2(n_7941),
.B1(n_8181),
.B2(n_8096),
.Y(n_12381)
);

INVx1_ASAP7_75t_L g12382 ( 
.A(n_11470),
.Y(n_12382)
);

AND2x2_ASAP7_75t_L g12383 ( 
.A(n_11420),
.B(n_8786),
.Y(n_12383)
);

NAND2xp5_ASAP7_75t_L g12384 ( 
.A(n_11906),
.B(n_10014),
.Y(n_12384)
);

INVx2_ASAP7_75t_L g12385 ( 
.A(n_11288),
.Y(n_12385)
);

NOR2x1_ASAP7_75t_L g12386 ( 
.A(n_11487),
.B(n_10846),
.Y(n_12386)
);

INVx1_ASAP7_75t_L g12387 ( 
.A(n_11470),
.Y(n_12387)
);

AND2x2_ASAP7_75t_L g12388 ( 
.A(n_11421),
.B(n_8829),
.Y(n_12388)
);

AND3x2_ASAP7_75t_L g12389 ( 
.A(n_11552),
.B(n_8039),
.C(n_9898),
.Y(n_12389)
);

INVx1_ASAP7_75t_L g12390 ( 
.A(n_11474),
.Y(n_12390)
);

INVx3_ASAP7_75t_L g12391 ( 
.A(n_11577),
.Y(n_12391)
);

HB1xp67_ASAP7_75t_L g12392 ( 
.A(n_11247),
.Y(n_12392)
);

AND2x2_ASAP7_75t_L g12393 ( 
.A(n_11338),
.B(n_8829),
.Y(n_12393)
);

AND2x2_ASAP7_75t_L g12394 ( 
.A(n_11399),
.B(n_8713),
.Y(n_12394)
);

INVx3_ASAP7_75t_L g12395 ( 
.A(n_11577),
.Y(n_12395)
);

AND2x2_ASAP7_75t_L g12396 ( 
.A(n_11439),
.B(n_8713),
.Y(n_12396)
);

INVx1_ASAP7_75t_L g12397 ( 
.A(n_11474),
.Y(n_12397)
);

AOI22xp33_ASAP7_75t_L g12398 ( 
.A1(n_11898),
.A2(n_11084),
.B1(n_11030),
.B2(n_11039),
.Y(n_12398)
);

INVx2_ASAP7_75t_L g12399 ( 
.A(n_11296),
.Y(n_12399)
);

AND2x4_ASAP7_75t_L g12400 ( 
.A(n_11542),
.B(n_8357),
.Y(n_12400)
);

AOI22xp5_ASAP7_75t_L g12401 ( 
.A1(n_11960),
.A2(n_10667),
.B1(n_10699),
.B2(n_11020),
.Y(n_12401)
);

INVx1_ASAP7_75t_L g12402 ( 
.A(n_11478),
.Y(n_12402)
);

INVxp67_ASAP7_75t_SL g12403 ( 
.A(n_11996),
.Y(n_12403)
);

AND2x2_ASAP7_75t_L g12404 ( 
.A(n_11507),
.B(n_11510),
.Y(n_12404)
);

AOI22xp33_ASAP7_75t_L g12405 ( 
.A1(n_11987),
.A2(n_10834),
.B1(n_11233),
.B2(n_11055),
.Y(n_12405)
);

BUFx6f_ASAP7_75t_L g12406 ( 
.A(n_11441),
.Y(n_12406)
);

NOR2x1_ASAP7_75t_SL g12407 ( 
.A(n_11305),
.B(n_11963),
.Y(n_12407)
);

AOI22xp33_ASAP7_75t_L g12408 ( 
.A1(n_11880),
.A2(n_10778),
.B1(n_10182),
.B2(n_10189),
.Y(n_12408)
);

AND2x2_ASAP7_75t_L g12409 ( 
.A(n_11514),
.B(n_8739),
.Y(n_12409)
);

NAND3xp33_ASAP7_75t_L g12410 ( 
.A(n_11707),
.B(n_11036),
.C(n_11026),
.Y(n_12410)
);

OR2x2_ASAP7_75t_L g12411 ( 
.A(n_11391),
.B(n_10017),
.Y(n_12411)
);

INVx1_ASAP7_75t_L g12412 ( 
.A(n_11478),
.Y(n_12412)
);

OAI21xp5_ASAP7_75t_L g12413 ( 
.A1(n_11943),
.A2(n_9659),
.B(n_9624),
.Y(n_12413)
);

INVx1_ASAP7_75t_L g12414 ( 
.A(n_11500),
.Y(n_12414)
);

NAND2xp5_ASAP7_75t_L g12415 ( 
.A(n_11906),
.B(n_10020),
.Y(n_12415)
);

INVx1_ASAP7_75t_L g12416 ( 
.A(n_11500),
.Y(n_12416)
);

NAND2xp5_ASAP7_75t_L g12417 ( 
.A(n_11610),
.B(n_10021),
.Y(n_12417)
);

INVx2_ASAP7_75t_L g12418 ( 
.A(n_11301),
.Y(n_12418)
);

NAND2x1p5_ASAP7_75t_L g12419 ( 
.A(n_11375),
.B(n_7795),
.Y(n_12419)
);

INVx1_ASAP7_75t_L g12420 ( 
.A(n_11504),
.Y(n_12420)
);

NAND2xp5_ASAP7_75t_L g12421 ( 
.A(n_11626),
.B(n_10028),
.Y(n_12421)
);

INVx2_ASAP7_75t_L g12422 ( 
.A(n_11313),
.Y(n_12422)
);

AND2x4_ASAP7_75t_L g12423 ( 
.A(n_11293),
.B(n_8357),
.Y(n_12423)
);

INVx1_ASAP7_75t_L g12424 ( 
.A(n_11504),
.Y(n_12424)
);

OR2x2_ASAP7_75t_L g12425 ( 
.A(n_11392),
.B(n_10036),
.Y(n_12425)
);

AOI22xp33_ASAP7_75t_SL g12426 ( 
.A1(n_11997),
.A2(n_9609),
.B1(n_9456),
.B2(n_10038),
.Y(n_12426)
);

INVx1_ASAP7_75t_L g12427 ( 
.A(n_11509),
.Y(n_12427)
);

AND2x2_ASAP7_75t_L g12428 ( 
.A(n_11516),
.B(n_8739),
.Y(n_12428)
);

HB1xp67_ASAP7_75t_L g12429 ( 
.A(n_11672),
.Y(n_12429)
);

AND2x4_ASAP7_75t_SL g12430 ( 
.A(n_11305),
.B(n_6876),
.Y(n_12430)
);

NOR2xp33_ASAP7_75t_L g12431 ( 
.A(n_11501),
.B(n_6899),
.Y(n_12431)
);

AND2x2_ASAP7_75t_L g12432 ( 
.A(n_11536),
.B(n_8742),
.Y(n_12432)
);

INVx1_ASAP7_75t_L g12433 ( 
.A(n_11509),
.Y(n_12433)
);

AND2x2_ASAP7_75t_L g12434 ( 
.A(n_11544),
.B(n_11625),
.Y(n_12434)
);

INVx1_ASAP7_75t_L g12435 ( 
.A(n_11522),
.Y(n_12435)
);

BUFx2_ASAP7_75t_L g12436 ( 
.A(n_11702),
.Y(n_12436)
);

AND2x2_ASAP7_75t_L g12437 ( 
.A(n_11630),
.B(n_11631),
.Y(n_12437)
);

INVx2_ASAP7_75t_L g12438 ( 
.A(n_11324),
.Y(n_12438)
);

INVx1_ASAP7_75t_L g12439 ( 
.A(n_11522),
.Y(n_12439)
);

AND2x4_ASAP7_75t_SL g12440 ( 
.A(n_11369),
.B(n_6896),
.Y(n_12440)
);

OR2x2_ASAP7_75t_L g12441 ( 
.A(n_11393),
.B(n_10044),
.Y(n_12441)
);

OR2x2_ASAP7_75t_L g12442 ( 
.A(n_11397),
.B(n_10047),
.Y(n_12442)
);

AND2x2_ASAP7_75t_L g12443 ( 
.A(n_11632),
.B(n_8742),
.Y(n_12443)
);

INVx1_ASAP7_75t_L g12444 ( 
.A(n_11523),
.Y(n_12444)
);

INVx4_ASAP7_75t_L g12445 ( 
.A(n_11505),
.Y(n_12445)
);

AND2x2_ASAP7_75t_L g12446 ( 
.A(n_11635),
.B(n_11636),
.Y(n_12446)
);

BUFx2_ASAP7_75t_L g12447 ( 
.A(n_11793),
.Y(n_12447)
);

INVx1_ASAP7_75t_L g12448 ( 
.A(n_11523),
.Y(n_12448)
);

AND2x2_ASAP7_75t_L g12449 ( 
.A(n_11582),
.B(n_11716),
.Y(n_12449)
);

BUFx2_ASAP7_75t_L g12450 ( 
.A(n_11779),
.Y(n_12450)
);

INVx1_ASAP7_75t_L g12451 ( 
.A(n_11524),
.Y(n_12451)
);

AND2x4_ASAP7_75t_L g12452 ( 
.A(n_11319),
.B(n_8458),
.Y(n_12452)
);

INVxp67_ASAP7_75t_SL g12453 ( 
.A(n_11329),
.Y(n_12453)
);

OR2x2_ASAP7_75t_L g12454 ( 
.A(n_11452),
.B(n_10050),
.Y(n_12454)
);

NAND2xp5_ASAP7_75t_L g12455 ( 
.A(n_11640),
.B(n_10055),
.Y(n_12455)
);

INVx2_ASAP7_75t_L g12456 ( 
.A(n_11332),
.Y(n_12456)
);

INVx3_ASAP7_75t_L g12457 ( 
.A(n_11438),
.Y(n_12457)
);

INVx1_ASAP7_75t_L g12458 ( 
.A(n_11524),
.Y(n_12458)
);

INVx1_ASAP7_75t_L g12459 ( 
.A(n_11531),
.Y(n_12459)
);

AND2x2_ASAP7_75t_L g12460 ( 
.A(n_11718),
.B(n_8458),
.Y(n_12460)
);

AND2x4_ASAP7_75t_SL g12461 ( 
.A(n_11387),
.B(n_6899),
.Y(n_12461)
);

INVx1_ASAP7_75t_L g12462 ( 
.A(n_11531),
.Y(n_12462)
);

AND2x4_ASAP7_75t_L g12463 ( 
.A(n_11403),
.B(n_8485),
.Y(n_12463)
);

BUFx2_ASAP7_75t_L g12464 ( 
.A(n_11442),
.Y(n_12464)
);

AOI22xp33_ASAP7_75t_SL g12465 ( 
.A1(n_11997),
.A2(n_9609),
.B1(n_9456),
.B2(n_10038),
.Y(n_12465)
);

INVx1_ASAP7_75t_L g12466 ( 
.A(n_11532),
.Y(n_12466)
);

OR2x2_ASAP7_75t_L g12467 ( 
.A(n_11567),
.B(n_10058),
.Y(n_12467)
);

INVx1_ASAP7_75t_L g12468 ( 
.A(n_11532),
.Y(n_12468)
);

INVx2_ASAP7_75t_L g12469 ( 
.A(n_11346),
.Y(n_12469)
);

AND2x2_ASAP7_75t_L g12470 ( 
.A(n_11738),
.B(n_8485),
.Y(n_12470)
);

AND2x2_ASAP7_75t_L g12471 ( 
.A(n_11381),
.B(n_8523),
.Y(n_12471)
);

AND2x2_ASAP7_75t_L g12472 ( 
.A(n_11398),
.B(n_8523),
.Y(n_12472)
);

AND2x2_ASAP7_75t_L g12473 ( 
.A(n_11729),
.B(n_8529),
.Y(n_12473)
);

INVx2_ASAP7_75t_SL g12474 ( 
.A(n_11442),
.Y(n_12474)
);

INVx1_ASAP7_75t_L g12475 ( 
.A(n_11533),
.Y(n_12475)
);

BUFx2_ASAP7_75t_L g12476 ( 
.A(n_11654),
.Y(n_12476)
);

BUFx2_ASAP7_75t_SL g12477 ( 
.A(n_11445),
.Y(n_12477)
);

NAND2xp5_ASAP7_75t_L g12478 ( 
.A(n_11707),
.B(n_10066),
.Y(n_12478)
);

INVx1_ASAP7_75t_L g12479 ( 
.A(n_11533),
.Y(n_12479)
);

AND2x2_ASAP7_75t_L g12480 ( 
.A(n_11650),
.B(n_8529),
.Y(n_12480)
);

INVx1_ASAP7_75t_L g12481 ( 
.A(n_11540),
.Y(n_12481)
);

OR2x2_ASAP7_75t_L g12482 ( 
.A(n_11587),
.B(n_10077),
.Y(n_12482)
);

INVx1_ASAP7_75t_L g12483 ( 
.A(n_11540),
.Y(n_12483)
);

INVx1_ASAP7_75t_L g12484 ( 
.A(n_11545),
.Y(n_12484)
);

INVx1_ASAP7_75t_L g12485 ( 
.A(n_11545),
.Y(n_12485)
);

INVxp67_ASAP7_75t_SL g12486 ( 
.A(n_11678),
.Y(n_12486)
);

INVx1_ASAP7_75t_L g12487 ( 
.A(n_11548),
.Y(n_12487)
);

INVx3_ASAP7_75t_L g12488 ( 
.A(n_11782),
.Y(n_12488)
);

AND2x2_ASAP7_75t_L g12489 ( 
.A(n_11765),
.B(n_8559),
.Y(n_12489)
);

INVxp67_ASAP7_75t_SL g12490 ( 
.A(n_11931),
.Y(n_12490)
);

NAND2xp5_ASAP7_75t_L g12491 ( 
.A(n_11845),
.B(n_11556),
.Y(n_12491)
);

INVx1_ASAP7_75t_L g12492 ( 
.A(n_11548),
.Y(n_12492)
);

INVx1_ASAP7_75t_L g12493 ( 
.A(n_11549),
.Y(n_12493)
);

INVx1_ASAP7_75t_L g12494 ( 
.A(n_11549),
.Y(n_12494)
);

NAND2xp5_ASAP7_75t_L g12495 ( 
.A(n_11564),
.B(n_10079),
.Y(n_12495)
);

INVx2_ASAP7_75t_L g12496 ( 
.A(n_11354),
.Y(n_12496)
);

NOR2xp33_ASAP7_75t_L g12497 ( 
.A(n_11475),
.B(n_11485),
.Y(n_12497)
);

OR2x2_ASAP7_75t_L g12498 ( 
.A(n_11609),
.B(n_10086),
.Y(n_12498)
);

OR2x2_ASAP7_75t_L g12499 ( 
.A(n_11502),
.B(n_10088),
.Y(n_12499)
);

AND2x2_ASAP7_75t_L g12500 ( 
.A(n_11767),
.B(n_8559),
.Y(n_12500)
);

AND2x2_ASAP7_75t_L g12501 ( 
.A(n_11736),
.B(n_8584),
.Y(n_12501)
);

AND2x4_ASAP7_75t_SL g12502 ( 
.A(n_11416),
.B(n_11417),
.Y(n_12502)
);

AND2x2_ASAP7_75t_L g12503 ( 
.A(n_11753),
.B(n_8584),
.Y(n_12503)
);

BUFx8_ASAP7_75t_SL g12504 ( 
.A(n_11649),
.Y(n_12504)
);

INVx1_ASAP7_75t_L g12505 ( 
.A(n_11561),
.Y(n_12505)
);

INVx1_ASAP7_75t_L g12506 ( 
.A(n_11561),
.Y(n_12506)
);

INVx1_ASAP7_75t_L g12507 ( 
.A(n_11563),
.Y(n_12507)
);

AND2x2_ASAP7_75t_L g12508 ( 
.A(n_11954),
.B(n_8600),
.Y(n_12508)
);

OR2x2_ASAP7_75t_L g12509 ( 
.A(n_11508),
.B(n_10089),
.Y(n_12509)
);

INVx2_ASAP7_75t_L g12510 ( 
.A(n_11677),
.Y(n_12510)
);

INVx1_ASAP7_75t_L g12511 ( 
.A(n_11563),
.Y(n_12511)
);

BUFx3_ASAP7_75t_L g12512 ( 
.A(n_11684),
.Y(n_12512)
);

INVx1_ASAP7_75t_L g12513 ( 
.A(n_11565),
.Y(n_12513)
);

AND2x4_ASAP7_75t_L g12514 ( 
.A(n_11639),
.B(n_8600),
.Y(n_12514)
);

INVx1_ASAP7_75t_L g12515 ( 
.A(n_11565),
.Y(n_12515)
);

NAND2xp5_ASAP7_75t_L g12516 ( 
.A(n_11788),
.B(n_10093),
.Y(n_12516)
);

INVx2_ASAP7_75t_SL g12517 ( 
.A(n_11262),
.Y(n_12517)
);

AND2x2_ASAP7_75t_L g12518 ( 
.A(n_11754),
.B(n_8622),
.Y(n_12518)
);

INVx4_ASAP7_75t_L g12519 ( 
.A(n_11454),
.Y(n_12519)
);

INVx1_ASAP7_75t_SL g12520 ( 
.A(n_11885),
.Y(n_12520)
);

OR2x2_ASAP7_75t_L g12521 ( 
.A(n_11511),
.B(n_10094),
.Y(n_12521)
);

AND2x2_ASAP7_75t_L g12522 ( 
.A(n_11757),
.B(n_8622),
.Y(n_12522)
);

AND2x2_ASAP7_75t_L g12523 ( 
.A(n_11768),
.B(n_8636),
.Y(n_12523)
);

INVx2_ASAP7_75t_L g12524 ( 
.A(n_11418),
.Y(n_12524)
);

NAND2xp5_ASAP7_75t_L g12525 ( 
.A(n_11868),
.B(n_10095),
.Y(n_12525)
);

INVx2_ASAP7_75t_L g12526 ( 
.A(n_11423),
.Y(n_12526)
);

AND2x2_ASAP7_75t_L g12527 ( 
.A(n_11741),
.B(n_8636),
.Y(n_12527)
);

AOI222xp33_ASAP7_75t_L g12528 ( 
.A1(n_11806),
.A2(n_10757),
.B1(n_10760),
.B2(n_10762),
.C1(n_10750),
.C2(n_10740),
.Y(n_12528)
);

INVx2_ASAP7_75t_L g12529 ( 
.A(n_11424),
.Y(n_12529)
);

AND2x2_ASAP7_75t_L g12530 ( 
.A(n_11742),
.B(n_8691),
.Y(n_12530)
);

INVx6_ASAP7_75t_L g12531 ( 
.A(n_11251),
.Y(n_12531)
);

INVx2_ASAP7_75t_L g12532 ( 
.A(n_11426),
.Y(n_12532)
);

AND2x2_ASAP7_75t_L g12533 ( 
.A(n_11745),
.B(n_8691),
.Y(n_12533)
);

INVx1_ASAP7_75t_L g12534 ( 
.A(n_11571),
.Y(n_12534)
);

OR2x2_ASAP7_75t_L g12535 ( 
.A(n_11566),
.B(n_10097),
.Y(n_12535)
);

OR2x2_ASAP7_75t_L g12536 ( 
.A(n_11611),
.B(n_10101),
.Y(n_12536)
);

NAND2xp5_ASAP7_75t_L g12537 ( 
.A(n_11234),
.B(n_10104),
.Y(n_12537)
);

AND2x4_ASAP7_75t_L g12538 ( 
.A(n_11234),
.B(n_8703),
.Y(n_12538)
);

OR2x2_ASAP7_75t_L g12539 ( 
.A(n_11629),
.B(n_11673),
.Y(n_12539)
);

OR2x2_ASAP7_75t_L g12540 ( 
.A(n_11368),
.B(n_10105),
.Y(n_12540)
);

AOI22xp33_ASAP7_75t_L g12541 ( 
.A1(n_11880),
.A2(n_10187),
.B1(n_10189),
.B2(n_10182),
.Y(n_12541)
);

AND2x2_ASAP7_75t_L g12542 ( 
.A(n_11645),
.B(n_8703),
.Y(n_12542)
);

AND2x2_ASAP7_75t_L g12543 ( 
.A(n_11712),
.B(n_7184),
.Y(n_12543)
);

AND2x2_ASAP7_75t_L g12544 ( 
.A(n_11620),
.B(n_7517),
.Y(n_12544)
);

AND2x2_ASAP7_75t_L g12545 ( 
.A(n_11621),
.B(n_7517),
.Y(n_12545)
);

AND2x4_ASAP7_75t_L g12546 ( 
.A(n_11623),
.B(n_6905),
.Y(n_12546)
);

OR2x2_ASAP7_75t_L g12547 ( 
.A(n_11388),
.B(n_10106),
.Y(n_12547)
);

AND2x4_ASAP7_75t_SL g12548 ( 
.A(n_11823),
.B(n_6905),
.Y(n_12548)
);

BUFx2_ASAP7_75t_L g12549 ( 
.A(n_11682),
.Y(n_12549)
);

NAND2xp5_ASAP7_75t_L g12550 ( 
.A(n_11865),
.B(n_10110),
.Y(n_12550)
);

OR2x2_ASAP7_75t_L g12551 ( 
.A(n_11622),
.B(n_11761),
.Y(n_12551)
);

NAND2xp5_ASAP7_75t_L g12552 ( 
.A(n_11759),
.B(n_10112),
.Y(n_12552)
);

INVx1_ASAP7_75t_L g12553 ( 
.A(n_11571),
.Y(n_12553)
);

NAND2xp5_ASAP7_75t_L g12554 ( 
.A(n_12000),
.B(n_10115),
.Y(n_12554)
);

AND2x2_ASAP7_75t_L g12555 ( 
.A(n_11867),
.B(n_7518),
.Y(n_12555)
);

INVx1_ASAP7_75t_L g12556 ( 
.A(n_11579),
.Y(n_12556)
);

HB1xp67_ASAP7_75t_L g12557 ( 
.A(n_11467),
.Y(n_12557)
);

INVxp67_ASAP7_75t_L g12558 ( 
.A(n_11946),
.Y(n_12558)
);

AND2x4_ASAP7_75t_SL g12559 ( 
.A(n_11642),
.B(n_7033),
.Y(n_12559)
);

OR2x2_ASAP7_75t_L g12560 ( 
.A(n_11715),
.B(n_10119),
.Y(n_12560)
);

AND2x2_ASAP7_75t_L g12561 ( 
.A(n_11871),
.B(n_7518),
.Y(n_12561)
);

INVx1_ASAP7_75t_L g12562 ( 
.A(n_11579),
.Y(n_12562)
);

INVxp33_ASAP7_75t_SL g12563 ( 
.A(n_11758),
.Y(n_12563)
);

BUFx2_ASAP7_75t_L g12564 ( 
.A(n_11909),
.Y(n_12564)
);

INVx1_ASAP7_75t_L g12565 ( 
.A(n_11585),
.Y(n_12565)
);

HB1xp67_ASAP7_75t_L g12566 ( 
.A(n_11814),
.Y(n_12566)
);

INVx2_ASAP7_75t_SL g12567 ( 
.A(n_11651),
.Y(n_12567)
);

AND2x2_ASAP7_75t_L g12568 ( 
.A(n_11901),
.B(n_11668),
.Y(n_12568)
);

INVx2_ASAP7_75t_L g12569 ( 
.A(n_11432),
.Y(n_12569)
);

NAND2xp5_ASAP7_75t_L g12570 ( 
.A(n_11762),
.B(n_10125),
.Y(n_12570)
);

NAND2xp5_ASAP7_75t_L g12571 ( 
.A(n_11769),
.B(n_10130),
.Y(n_12571)
);

INVx2_ASAP7_75t_L g12572 ( 
.A(n_11434),
.Y(n_12572)
);

AND2x2_ASAP7_75t_L g12573 ( 
.A(n_11804),
.B(n_7610),
.Y(n_12573)
);

INVx2_ASAP7_75t_L g12574 ( 
.A(n_11435),
.Y(n_12574)
);

AND2x2_ASAP7_75t_L g12575 ( 
.A(n_11816),
.B(n_7610),
.Y(n_12575)
);

OR2x2_ASAP7_75t_L g12576 ( 
.A(n_11883),
.B(n_10138),
.Y(n_12576)
);

AOI22xp33_ASAP7_75t_L g12577 ( 
.A1(n_11937),
.A2(n_10192),
.B1(n_10209),
.B2(n_10187),
.Y(n_12577)
);

INVx2_ASAP7_75t_L g12578 ( 
.A(n_11436),
.Y(n_12578)
);

BUFx6f_ASAP7_75t_L g12579 ( 
.A(n_11529),
.Y(n_12579)
);

OAI22xp5_ASAP7_75t_L g12580 ( 
.A1(n_11613),
.A2(n_7941),
.B1(n_8181),
.B2(n_8096),
.Y(n_12580)
);

AND2x2_ASAP7_75t_L g12581 ( 
.A(n_11711),
.B(n_7642),
.Y(n_12581)
);

INVx1_ASAP7_75t_L g12582 ( 
.A(n_11585),
.Y(n_12582)
);

INVx1_ASAP7_75t_L g12583 ( 
.A(n_11594),
.Y(n_12583)
);

BUFx2_ASAP7_75t_L g12584 ( 
.A(n_11933),
.Y(n_12584)
);

AND2x2_ASAP7_75t_L g12585 ( 
.A(n_11800),
.B(n_7642),
.Y(n_12585)
);

INVx1_ASAP7_75t_L g12586 ( 
.A(n_11594),
.Y(n_12586)
);

INVx2_ASAP7_75t_L g12587 ( 
.A(n_11357),
.Y(n_12587)
);

INVx2_ASAP7_75t_L g12588 ( 
.A(n_11310),
.Y(n_12588)
);

AND2x2_ASAP7_75t_L g12589 ( 
.A(n_11803),
.B(n_7676),
.Y(n_12589)
);

HB1xp67_ASAP7_75t_L g12590 ( 
.A(n_11819),
.Y(n_12590)
);

INVx1_ASAP7_75t_L g12591 ( 
.A(n_11595),
.Y(n_12591)
);

AND2x2_ASAP7_75t_L g12592 ( 
.A(n_11810),
.B(n_7676),
.Y(n_12592)
);

INVx2_ASAP7_75t_SL g12593 ( 
.A(n_11782),
.Y(n_12593)
);

INVx2_ASAP7_75t_L g12594 ( 
.A(n_11285),
.Y(n_12594)
);

INVxp67_ASAP7_75t_L g12595 ( 
.A(n_11834),
.Y(n_12595)
);

OR2x2_ASAP7_75t_L g12596 ( 
.A(n_11492),
.B(n_11965),
.Y(n_12596)
);

AOI22xp33_ASAP7_75t_L g12597 ( 
.A1(n_11986),
.A2(n_10209),
.B1(n_10215),
.B2(n_10192),
.Y(n_12597)
);

AND2x2_ASAP7_75t_L g12598 ( 
.A(n_11811),
.B(n_7696),
.Y(n_12598)
);

INVx1_ASAP7_75t_L g12599 ( 
.A(n_11595),
.Y(n_12599)
);

NAND2xp5_ASAP7_75t_L g12600 ( 
.A(n_11683),
.B(n_10140),
.Y(n_12600)
);

INVx1_ASAP7_75t_L g12601 ( 
.A(n_11597),
.Y(n_12601)
);

INVx2_ASAP7_75t_L g12602 ( 
.A(n_11790),
.Y(n_12602)
);

NAND2xp5_ASAP7_75t_L g12603 ( 
.A(n_11685),
.B(n_10148),
.Y(n_12603)
);

INVxp67_ASAP7_75t_L g12604 ( 
.A(n_11862),
.Y(n_12604)
);

INVx1_ASAP7_75t_L g12605 ( 
.A(n_11597),
.Y(n_12605)
);

AOI22xp33_ASAP7_75t_L g12606 ( 
.A1(n_11985),
.A2(n_10218),
.B1(n_10231),
.B2(n_10215),
.Y(n_12606)
);

INVx2_ASAP7_75t_L g12607 ( 
.A(n_11790),
.Y(n_12607)
);

INVx2_ASAP7_75t_L g12608 ( 
.A(n_11472),
.Y(n_12608)
);

NOR2xp33_ASAP7_75t_L g12609 ( 
.A(n_11537),
.B(n_7033),
.Y(n_12609)
);

INVx1_ASAP7_75t_L g12610 ( 
.A(n_11599),
.Y(n_12610)
);

INVx2_ASAP7_75t_L g12611 ( 
.A(n_11473),
.Y(n_12611)
);

INVx1_ASAP7_75t_L g12612 ( 
.A(n_11599),
.Y(n_12612)
);

INVx2_ASAP7_75t_L g12613 ( 
.A(n_11482),
.Y(n_12613)
);

AND2x4_ASAP7_75t_L g12614 ( 
.A(n_11799),
.B(n_7074),
.Y(n_12614)
);

INVx2_ASAP7_75t_L g12615 ( 
.A(n_11483),
.Y(n_12615)
);

INVx3_ASAP7_75t_L g12616 ( 
.A(n_11799),
.Y(n_12616)
);

INVx2_ASAP7_75t_L g12617 ( 
.A(n_11652),
.Y(n_12617)
);

NAND2xp5_ASAP7_75t_L g12618 ( 
.A(n_11691),
.B(n_10149),
.Y(n_12618)
);

AND2x2_ASAP7_75t_L g12619 ( 
.A(n_11820),
.B(n_7696),
.Y(n_12619)
);

INVx2_ASAP7_75t_L g12620 ( 
.A(n_11657),
.Y(n_12620)
);

INVxp67_ASAP7_75t_L g12621 ( 
.A(n_11957),
.Y(n_12621)
);

AND2x2_ASAP7_75t_L g12622 ( 
.A(n_11824),
.B(n_7727),
.Y(n_12622)
);

INVx1_ASAP7_75t_L g12623 ( 
.A(n_11601),
.Y(n_12623)
);

INVxp33_ASAP7_75t_L g12624 ( 
.A(n_11976),
.Y(n_12624)
);

NAND2xp5_ASAP7_75t_L g12625 ( 
.A(n_11697),
.B(n_10151),
.Y(n_12625)
);

INVx1_ASAP7_75t_L g12626 ( 
.A(n_11601),
.Y(n_12626)
);

INVxp67_ASAP7_75t_SL g12627 ( 
.A(n_11931),
.Y(n_12627)
);

OR2x2_ASAP7_75t_L g12628 ( 
.A(n_11785),
.B(n_10152),
.Y(n_12628)
);

OR2x2_ASAP7_75t_L g12629 ( 
.A(n_11717),
.B(n_10155),
.Y(n_12629)
);

INVx2_ASAP7_75t_L g12630 ( 
.A(n_11658),
.Y(n_12630)
);

INVx2_ASAP7_75t_L g12631 ( 
.A(n_11659),
.Y(n_12631)
);

INVx1_ASAP7_75t_L g12632 ( 
.A(n_11755),
.Y(n_12632)
);

INVx1_ASAP7_75t_L g12633 ( 
.A(n_11755),
.Y(n_12633)
);

INVx1_ASAP7_75t_L g12634 ( 
.A(n_11777),
.Y(n_12634)
);

INVx2_ASAP7_75t_L g12635 ( 
.A(n_11661),
.Y(n_12635)
);

NOR2xp33_ASAP7_75t_L g12636 ( 
.A(n_11843),
.B(n_7074),
.Y(n_12636)
);

INVx1_ASAP7_75t_L g12637 ( 
.A(n_11777),
.Y(n_12637)
);

NAND2xp5_ASAP7_75t_L g12638 ( 
.A(n_11910),
.B(n_10163),
.Y(n_12638)
);

AND2x2_ASAP7_75t_L g12639 ( 
.A(n_11837),
.B(n_7727),
.Y(n_12639)
);

INVxp67_ASAP7_75t_SL g12640 ( 
.A(n_11931),
.Y(n_12640)
);

INVx1_ASAP7_75t_L g12641 ( 
.A(n_11602),
.Y(n_12641)
);

INVx1_ASAP7_75t_L g12642 ( 
.A(n_11602),
.Y(n_12642)
);

AND2x2_ASAP7_75t_L g12643 ( 
.A(n_11838),
.B(n_9155),
.Y(n_12643)
);

AND2x2_ASAP7_75t_L g12644 ( 
.A(n_11839),
.B(n_9231),
.Y(n_12644)
);

NOR2x1p5_ASAP7_75t_L g12645 ( 
.A(n_11461),
.B(n_9231),
.Y(n_12645)
);

NAND2xp5_ASAP7_75t_L g12646 ( 
.A(n_11853),
.B(n_10168),
.Y(n_12646)
);

INVx1_ASAP7_75t_L g12647 ( 
.A(n_11614),
.Y(n_12647)
);

INVx1_ASAP7_75t_L g12648 ( 
.A(n_11614),
.Y(n_12648)
);

AND2x4_ASAP7_75t_L g12649 ( 
.A(n_11935),
.B(n_6941),
.Y(n_12649)
);

INVx1_ASAP7_75t_L g12650 ( 
.A(n_11615),
.Y(n_12650)
);

INVxp67_ASAP7_75t_L g12651 ( 
.A(n_11700),
.Y(n_12651)
);

INVx1_ASAP7_75t_L g12652 ( 
.A(n_11615),
.Y(n_12652)
);

INVx1_ASAP7_75t_L g12653 ( 
.A(n_11616),
.Y(n_12653)
);

AND2x2_ASAP7_75t_L g12654 ( 
.A(n_11856),
.B(n_8289),
.Y(n_12654)
);

AND2x2_ASAP7_75t_L g12655 ( 
.A(n_12015),
.B(n_11859),
.Y(n_12655)
);

AND2x2_ASAP7_75t_L g12656 ( 
.A(n_12265),
.B(n_11863),
.Y(n_12656)
);

INVx2_ASAP7_75t_L g12657 ( 
.A(n_12057),
.Y(n_12657)
);

AND2x2_ASAP7_75t_L g12658 ( 
.A(n_12057),
.B(n_11869),
.Y(n_12658)
);

NAND2xp5_ASAP7_75t_L g12659 ( 
.A(n_12001),
.B(n_11921),
.Y(n_12659)
);

AND2x2_ASAP7_75t_L g12660 ( 
.A(n_12447),
.B(n_11618),
.Y(n_12660)
);

AND2x4_ASAP7_75t_SL g12661 ( 
.A(n_12118),
.B(n_11681),
.Y(n_12661)
);

INVx1_ASAP7_75t_L g12662 ( 
.A(n_12009),
.Y(n_12662)
);

BUFx6f_ASAP7_75t_L g12663 ( 
.A(n_12118),
.Y(n_12663)
);

INVx2_ASAP7_75t_L g12664 ( 
.A(n_12075),
.Y(n_12664)
);

INVx3_ASAP7_75t_L g12665 ( 
.A(n_12232),
.Y(n_12665)
);

NAND2x1p5_ASAP7_75t_SL g12666 ( 
.A(n_12242),
.B(n_11787),
.Y(n_12666)
);

INVx2_ASAP7_75t_L g12667 ( 
.A(n_12354),
.Y(n_12667)
);

NOR2xp33_ASAP7_75t_L g12668 ( 
.A(n_12271),
.B(n_11884),
.Y(n_12668)
);

BUFx3_ASAP7_75t_L g12669 ( 
.A(n_12033),
.Y(n_12669)
);

INVx2_ASAP7_75t_L g12670 ( 
.A(n_12033),
.Y(n_12670)
);

INVxp67_ASAP7_75t_SL g12671 ( 
.A(n_12504),
.Y(n_12671)
);

AND2x2_ASAP7_75t_L g12672 ( 
.A(n_12077),
.B(n_11756),
.Y(n_12672)
);

INVx2_ASAP7_75t_L g12673 ( 
.A(n_12602),
.Y(n_12673)
);

INVx1_ASAP7_75t_L g12674 ( 
.A(n_12221),
.Y(n_12674)
);

BUFx3_ASAP7_75t_L g12675 ( 
.A(n_12345),
.Y(n_12675)
);

AND2x2_ASAP7_75t_L g12676 ( 
.A(n_12104),
.B(n_11912),
.Y(n_12676)
);

AOI221xp5_ASAP7_75t_L g12677 ( 
.A1(n_12152),
.A2(n_11662),
.B1(n_11766),
.B2(n_11982),
.C(n_11386),
.Y(n_12677)
);

INVx1_ASAP7_75t_L g12678 ( 
.A(n_12026),
.Y(n_12678)
);

AND2x2_ASAP7_75t_L g12679 ( 
.A(n_12226),
.B(n_11872),
.Y(n_12679)
);

INVx1_ASAP7_75t_L g12680 ( 
.A(n_12026),
.Y(n_12680)
);

HB1xp67_ASAP7_75t_L g12681 ( 
.A(n_12429),
.Y(n_12681)
);

AND2x2_ASAP7_75t_L g12682 ( 
.A(n_12340),
.B(n_11882),
.Y(n_12682)
);

AOI22xp33_ASAP7_75t_L g12683 ( 
.A1(n_12016),
.A2(n_11794),
.B1(n_11915),
.B2(n_11989),
.Y(n_12683)
);

AND2x2_ASAP7_75t_L g12684 ( 
.A(n_12437),
.B(n_12446),
.Y(n_12684)
);

NAND2xp5_ASAP7_75t_L g12685 ( 
.A(n_12520),
.B(n_11886),
.Y(n_12685)
);

AND2x2_ASAP7_75t_L g12686 ( 
.A(n_12476),
.B(n_11693),
.Y(n_12686)
);

INVx1_ASAP7_75t_L g12687 ( 
.A(n_12035),
.Y(n_12687)
);

OAI21xp5_ASAP7_75t_SL g12688 ( 
.A1(n_12025),
.A2(n_11570),
.B(n_11791),
.Y(n_12688)
);

INVx1_ASAP7_75t_L g12689 ( 
.A(n_12035),
.Y(n_12689)
);

INVx2_ASAP7_75t_L g12690 ( 
.A(n_12607),
.Y(n_12690)
);

HB1xp67_ASAP7_75t_L g12691 ( 
.A(n_12512),
.Y(n_12691)
);

NAND2xp5_ASAP7_75t_L g12692 ( 
.A(n_12563),
.B(n_11764),
.Y(n_12692)
);

AND2x2_ASAP7_75t_L g12693 ( 
.A(n_12449),
.B(n_11770),
.Y(n_12693)
);

INVx3_ASAP7_75t_L g12694 ( 
.A(n_12232),
.Y(n_12694)
);

AND2x2_ASAP7_75t_L g12695 ( 
.A(n_12010),
.B(n_11772),
.Y(n_12695)
);

HB1xp67_ASAP7_75t_L g12696 ( 
.A(n_12253),
.Y(n_12696)
);

BUFx6f_ASAP7_75t_L g12697 ( 
.A(n_12321),
.Y(n_12697)
);

INVx4_ASAP7_75t_L g12698 ( 
.A(n_12158),
.Y(n_12698)
);

OR2x2_ASAP7_75t_L g12699 ( 
.A(n_12549),
.B(n_11900),
.Y(n_12699)
);

INVx2_ASAP7_75t_L g12700 ( 
.A(n_12436),
.Y(n_12700)
);

INVx3_ASAP7_75t_L g12701 ( 
.A(n_12243),
.Y(n_12701)
);

INVx5_ASAP7_75t_SL g12702 ( 
.A(n_12346),
.Y(n_12702)
);

INVx2_ASAP7_75t_L g12703 ( 
.A(n_12263),
.Y(n_12703)
);

HB1xp67_ASAP7_75t_L g12704 ( 
.A(n_12264),
.Y(n_12704)
);

BUFx2_ASAP7_75t_L g12705 ( 
.A(n_12249),
.Y(n_12705)
);

INVx2_ASAP7_75t_L g12706 ( 
.A(n_12263),
.Y(n_12706)
);

AND2x2_ASAP7_75t_L g12707 ( 
.A(n_12243),
.B(n_11784),
.Y(n_12707)
);

INVx2_ASAP7_75t_L g12708 ( 
.A(n_12333),
.Y(n_12708)
);

INVx1_ASAP7_75t_L g12709 ( 
.A(n_12017),
.Y(n_12709)
);

AO21x2_ASAP7_75t_L g12710 ( 
.A1(n_12058),
.A2(n_11530),
.B(n_11786),
.Y(n_12710)
);

BUFx2_ASAP7_75t_L g12711 ( 
.A(n_12490),
.Y(n_12711)
);

INVx2_ASAP7_75t_L g12712 ( 
.A(n_12333),
.Y(n_12712)
);

NAND2xp5_ASAP7_75t_L g12713 ( 
.A(n_12350),
.B(n_11889),
.Y(n_12713)
);

OR2x2_ASAP7_75t_L g12714 ( 
.A(n_12595),
.B(n_11396),
.Y(n_12714)
);

AND2x2_ASAP7_75t_L g12715 ( 
.A(n_12200),
.B(n_11792),
.Y(n_12715)
);

BUFx2_ASAP7_75t_L g12716 ( 
.A(n_12627),
.Y(n_12716)
);

AND2x2_ASAP7_75t_L g12717 ( 
.A(n_12366),
.B(n_11795),
.Y(n_12717)
);

NAND2xp5_ASAP7_75t_L g12718 ( 
.A(n_12453),
.B(n_11746),
.Y(n_12718)
);

INVx1_ASAP7_75t_L g12719 ( 
.A(n_12036),
.Y(n_12719)
);

BUFx2_ASAP7_75t_L g12720 ( 
.A(n_12640),
.Y(n_12720)
);

OR2x2_ASAP7_75t_L g12721 ( 
.A(n_12604),
.B(n_12596),
.Y(n_12721)
);

AND2x2_ASAP7_75t_L g12722 ( 
.A(n_12368),
.B(n_11891),
.Y(n_12722)
);

AND2x4_ASAP7_75t_L g12723 ( 
.A(n_12546),
.B(n_11681),
.Y(n_12723)
);

AND2x2_ASAP7_75t_L g12724 ( 
.A(n_12087),
.B(n_11893),
.Y(n_12724)
);

INVxp67_ASAP7_75t_SL g12725 ( 
.A(n_12352),
.Y(n_12725)
);

AND2x2_ASAP7_75t_L g12726 ( 
.A(n_12361),
.B(n_11875),
.Y(n_12726)
);

INVx1_ASAP7_75t_L g12727 ( 
.A(n_12047),
.Y(n_12727)
);

INVx2_ASAP7_75t_L g12728 ( 
.A(n_12391),
.Y(n_12728)
);

OR2x6_ASAP7_75t_L g12729 ( 
.A(n_12102),
.B(n_11547),
.Y(n_12729)
);

INVx1_ASAP7_75t_L g12730 ( 
.A(n_12246),
.Y(n_12730)
);

AND2x2_ASAP7_75t_L g12731 ( 
.A(n_12106),
.B(n_11974),
.Y(n_12731)
);

BUFx2_ASAP7_75t_L g12732 ( 
.A(n_12372),
.Y(n_12732)
);

AND2x2_ASAP7_75t_L g12733 ( 
.A(n_12343),
.B(n_11710),
.Y(n_12733)
);

AND2x2_ASAP7_75t_L g12734 ( 
.A(n_12546),
.B(n_11951),
.Y(n_12734)
);

AOI22xp33_ASAP7_75t_L g12735 ( 
.A1(n_12551),
.A2(n_11794),
.B1(n_11915),
.B2(n_11983),
.Y(n_12735)
);

HB1xp67_ASAP7_75t_L g12736 ( 
.A(n_12044),
.Y(n_12736)
);

INVx1_ASAP7_75t_L g12737 ( 
.A(n_12071),
.Y(n_12737)
);

HB1xp67_ASAP7_75t_L g12738 ( 
.A(n_12358),
.Y(n_12738)
);

INVx2_ASAP7_75t_L g12739 ( 
.A(n_12391),
.Y(n_12739)
);

AND2x2_ASAP7_75t_L g12740 ( 
.A(n_12502),
.B(n_11690),
.Y(n_12740)
);

AND2x2_ASAP7_75t_L g12741 ( 
.A(n_12308),
.B(n_11699),
.Y(n_12741)
);

OR2x2_ASAP7_75t_L g12742 ( 
.A(n_12486),
.B(n_11780),
.Y(n_12742)
);

AOI221xp5_ASAP7_75t_L g12743 ( 
.A1(n_12100),
.A2(n_11925),
.B1(n_11938),
.B2(n_11844),
.C(n_11907),
.Y(n_12743)
);

INVx2_ASAP7_75t_L g12744 ( 
.A(n_12395),
.Y(n_12744)
);

AND2x2_ASAP7_75t_L g12745 ( 
.A(n_12308),
.B(n_11709),
.Y(n_12745)
);

INVx4_ASAP7_75t_L g12746 ( 
.A(n_12158),
.Y(n_12746)
);

NAND2x1p5_ASAP7_75t_L g12747 ( 
.A(n_12072),
.B(n_11963),
.Y(n_12747)
);

BUFx3_ASAP7_75t_L g12748 ( 
.A(n_12461),
.Y(n_12748)
);

OR2x2_ASAP7_75t_L g12749 ( 
.A(n_12209),
.B(n_11781),
.Y(n_12749)
);

INVx1_ASAP7_75t_L g12750 ( 
.A(n_12098),
.Y(n_12750)
);

BUFx6f_ASAP7_75t_L g12751 ( 
.A(n_12406),
.Y(n_12751)
);

INVxp67_ASAP7_75t_L g12752 ( 
.A(n_12431),
.Y(n_12752)
);

AND2x2_ASAP7_75t_L g12753 ( 
.A(n_12277),
.B(n_11506),
.Y(n_12753)
);

AND2x2_ASAP7_75t_L g12754 ( 
.A(n_12248),
.B(n_11950),
.Y(n_12754)
);

INVx2_ASAP7_75t_L g12755 ( 
.A(n_12395),
.Y(n_12755)
);

INVx2_ASAP7_75t_L g12756 ( 
.A(n_12445),
.Y(n_12756)
);

INVx1_ASAP7_75t_L g12757 ( 
.A(n_12579),
.Y(n_12757)
);

OR2x2_ASAP7_75t_L g12758 ( 
.A(n_12403),
.B(n_11812),
.Y(n_12758)
);

INVx1_ASAP7_75t_L g12759 ( 
.A(n_12579),
.Y(n_12759)
);

AND2x2_ASAP7_75t_L g12760 ( 
.A(n_12248),
.B(n_12293),
.Y(n_12760)
);

AND2x2_ASAP7_75t_L g12761 ( 
.A(n_12293),
.B(n_11967),
.Y(n_12761)
);

INVx1_ASAP7_75t_L g12762 ( 
.A(n_12579),
.Y(n_12762)
);

AND2x2_ASAP7_75t_L g12763 ( 
.A(n_12355),
.B(n_11967),
.Y(n_12763)
);

INVx1_ASAP7_75t_L g12764 ( 
.A(n_12002),
.Y(n_12764)
);

AND2x2_ASAP7_75t_L g12765 ( 
.A(n_12355),
.B(n_11969),
.Y(n_12765)
);

INVx1_ASAP7_75t_L g12766 ( 
.A(n_12079),
.Y(n_12766)
);

NOR2x1_ASAP7_75t_L g12767 ( 
.A(n_12102),
.B(n_11584),
.Y(n_12767)
);

NAND2xp5_ASAP7_75t_L g12768 ( 
.A(n_12307),
.B(n_11686),
.Y(n_12768)
);

INVx3_ASAP7_75t_L g12769 ( 
.A(n_12295),
.Y(n_12769)
);

INVx1_ASAP7_75t_L g12770 ( 
.A(n_12060),
.Y(n_12770)
);

INVx5_ASAP7_75t_SL g12771 ( 
.A(n_12346),
.Y(n_12771)
);

INVx3_ASAP7_75t_L g12772 ( 
.A(n_12295),
.Y(n_12772)
);

INVx1_ASAP7_75t_L g12773 ( 
.A(n_12312),
.Y(n_12773)
);

INVx1_ASAP7_75t_L g12774 ( 
.A(n_12312),
.Y(n_12774)
);

INVx3_ASAP7_75t_L g12775 ( 
.A(n_12105),
.Y(n_12775)
);

HB1xp67_ASAP7_75t_L g12776 ( 
.A(n_12450),
.Y(n_12776)
);

OR2x2_ASAP7_75t_L g12777 ( 
.A(n_12347),
.B(n_11719),
.Y(n_12777)
);

INVx1_ASAP7_75t_L g12778 ( 
.A(n_12313),
.Y(n_12778)
);

HB1xp67_ASAP7_75t_L g12779 ( 
.A(n_12162),
.Y(n_12779)
);

NAND2xp5_ASAP7_75t_L g12780 ( 
.A(n_12445),
.B(n_11956),
.Y(n_12780)
);

INVx2_ASAP7_75t_L g12781 ( 
.A(n_12464),
.Y(n_12781)
);

AO21x2_ASAP7_75t_L g12782 ( 
.A1(n_12300),
.A2(n_11786),
.B(n_11728),
.Y(n_12782)
);

INVx2_ASAP7_75t_L g12783 ( 
.A(n_12072),
.Y(n_12783)
);

INVx2_ASAP7_75t_L g12784 ( 
.A(n_12074),
.Y(n_12784)
);

INVx1_ASAP7_75t_L g12785 ( 
.A(n_12313),
.Y(n_12785)
);

INVx3_ASAP7_75t_L g12786 ( 
.A(n_12130),
.Y(n_12786)
);

AND2x4_ASAP7_75t_L g12787 ( 
.A(n_12407),
.B(n_11379),
.Y(n_12787)
);

AND2x4_ASAP7_75t_L g12788 ( 
.A(n_12407),
.B(n_11383),
.Y(n_12788)
);

OR2x2_ASAP7_75t_L g12789 ( 
.A(n_12539),
.B(n_11739),
.Y(n_12789)
);

HB1xp67_ASAP7_75t_L g12790 ( 
.A(n_12299),
.Y(n_12790)
);

AO21x2_ASAP7_75t_L g12791 ( 
.A1(n_12300),
.A2(n_11728),
.B(n_11696),
.Y(n_12791)
);

OR2x2_ASAP7_75t_L g12792 ( 
.A(n_12558),
.B(n_11744),
.Y(n_12792)
);

INVx3_ASAP7_75t_L g12793 ( 
.A(n_12130),
.Y(n_12793)
);

NOR2xp33_ASAP7_75t_L g12794 ( 
.A(n_12256),
.B(n_11966),
.Y(n_12794)
);

INVx3_ASAP7_75t_L g12795 ( 
.A(n_12144),
.Y(n_12795)
);

AND2x2_ASAP7_75t_L g12796 ( 
.A(n_12434),
.B(n_11966),
.Y(n_12796)
);

AND2x2_ASAP7_75t_L g12797 ( 
.A(n_12126),
.B(n_11981),
.Y(n_12797)
);

INVx2_ASAP7_75t_L g12798 ( 
.A(n_12074),
.Y(n_12798)
);

INVx4_ASAP7_75t_L g12799 ( 
.A(n_12207),
.Y(n_12799)
);

INVx1_ASAP7_75t_L g12800 ( 
.A(n_12632),
.Y(n_12800)
);

AND2x2_ASAP7_75t_L g12801 ( 
.A(n_12164),
.B(n_11911),
.Y(n_12801)
);

AO21x2_ASAP7_75t_L g12802 ( 
.A1(n_12303),
.A2(n_12305),
.B(n_12241),
.Y(n_12802)
);

OR2x2_ASAP7_75t_L g12803 ( 
.A(n_12301),
.B(n_11964),
.Y(n_12803)
);

INVx1_ASAP7_75t_L g12804 ( 
.A(n_12632),
.Y(n_12804)
);

INVx2_ASAP7_75t_SL g12805 ( 
.A(n_12531),
.Y(n_12805)
);

INVx3_ASAP7_75t_L g12806 ( 
.A(n_12144),
.Y(n_12806)
);

OR2x2_ASAP7_75t_L g12807 ( 
.A(n_12239),
.B(n_11826),
.Y(n_12807)
);

AND2x2_ASAP7_75t_L g12808 ( 
.A(n_12489),
.B(n_11914),
.Y(n_12808)
);

O2A1O1Ixp33_ASAP7_75t_L g12809 ( 
.A1(n_12651),
.A2(n_12621),
.B(n_12131),
.C(n_12173),
.Y(n_12809)
);

INVx2_ASAP7_75t_L g12810 ( 
.A(n_12531),
.Y(n_12810)
);

INVx2_ASAP7_75t_L g12811 ( 
.A(n_12207),
.Y(n_12811)
);

INVx2_ASAP7_75t_L g12812 ( 
.A(n_12406),
.Y(n_12812)
);

INVx2_ASAP7_75t_L g12813 ( 
.A(n_12406),
.Y(n_12813)
);

INVx3_ASAP7_75t_L g12814 ( 
.A(n_12614),
.Y(n_12814)
);

INVx1_ASAP7_75t_L g12815 ( 
.A(n_12633),
.Y(n_12815)
);

INVx1_ASAP7_75t_L g12816 ( 
.A(n_12633),
.Y(n_12816)
);

HB1xp67_ASAP7_75t_L g12817 ( 
.A(n_12320),
.Y(n_12817)
);

HB1xp67_ASAP7_75t_L g12818 ( 
.A(n_12324),
.Y(n_12818)
);

INVx1_ASAP7_75t_L g12819 ( 
.A(n_12634),
.Y(n_12819)
);

AND2x2_ASAP7_75t_L g12820 ( 
.A(n_12500),
.B(n_11973),
.Y(n_12820)
);

INVx2_ASAP7_75t_L g12821 ( 
.A(n_12510),
.Y(n_12821)
);

OR2x2_ASAP7_75t_L g12822 ( 
.A(n_12255),
.B(n_11775),
.Y(n_12822)
);

INVx1_ASAP7_75t_L g12823 ( 
.A(n_12634),
.Y(n_12823)
);

AND2x2_ASAP7_75t_L g12824 ( 
.A(n_12287),
.B(n_11908),
.Y(n_12824)
);

INVx1_ASAP7_75t_L g12825 ( 
.A(n_12637),
.Y(n_12825)
);

OR2x6_ASAP7_75t_L g12826 ( 
.A(n_12083),
.B(n_11879),
.Y(n_12826)
);

INVx2_ASAP7_75t_L g12827 ( 
.A(n_12302),
.Y(n_12827)
);

INVx2_ASAP7_75t_L g12828 ( 
.A(n_12314),
.Y(n_12828)
);

HB1xp67_ASAP7_75t_L g12829 ( 
.A(n_12325),
.Y(n_12829)
);

AND2x2_ASAP7_75t_L g12830 ( 
.A(n_12021),
.B(n_11991),
.Y(n_12830)
);

INVx2_ASAP7_75t_L g12831 ( 
.A(n_12514),
.Y(n_12831)
);

INVx1_ASAP7_75t_L g12832 ( 
.A(n_12637),
.Y(n_12832)
);

OR2x2_ASAP7_75t_L g12833 ( 
.A(n_12139),
.B(n_11832),
.Y(n_12833)
);

AOI21xp5_ASAP7_75t_SL g12834 ( 
.A1(n_12150),
.A2(n_11963),
.B(n_11934),
.Y(n_12834)
);

HB1xp67_ASAP7_75t_L g12835 ( 
.A(n_12214),
.Y(n_12835)
);

INVx1_ASAP7_75t_L g12836 ( 
.A(n_12311),
.Y(n_12836)
);

NAND2xp5_ASAP7_75t_L g12837 ( 
.A(n_12557),
.B(n_12517),
.Y(n_12837)
);

INVx1_ASAP7_75t_L g12838 ( 
.A(n_12082),
.Y(n_12838)
);

INVx1_ASAP7_75t_L g12839 ( 
.A(n_12085),
.Y(n_12839)
);

AND2x2_ASAP7_75t_L g12840 ( 
.A(n_12012),
.B(n_12378),
.Y(n_12840)
);

AND2x2_ASAP7_75t_L g12841 ( 
.A(n_12194),
.B(n_11995),
.Y(n_12841)
);

AND2x2_ASAP7_75t_L g12842 ( 
.A(n_12544),
.B(n_11932),
.Y(n_12842)
);

BUFx2_ASAP7_75t_L g12843 ( 
.A(n_12303),
.Y(n_12843)
);

INVx1_ASAP7_75t_L g12844 ( 
.A(n_12089),
.Y(n_12844)
);

INVx2_ASAP7_75t_L g12845 ( 
.A(n_12514),
.Y(n_12845)
);

NAND2x1_ASAP7_75t_SL g12846 ( 
.A(n_12379),
.B(n_11919),
.Y(n_12846)
);

HB1xp67_ASAP7_75t_L g12847 ( 
.A(n_12215),
.Y(n_12847)
);

INVx1_ASAP7_75t_L g12848 ( 
.A(n_12091),
.Y(n_12848)
);

INVx4_ASAP7_75t_L g12849 ( 
.A(n_12172),
.Y(n_12849)
);

AND2x2_ASAP7_75t_L g12850 ( 
.A(n_12545),
.B(n_11945),
.Y(n_12850)
);

AND2x4_ASAP7_75t_L g12851 ( 
.A(n_12614),
.B(n_12304),
.Y(n_12851)
);

INVx1_ASAP7_75t_L g12852 ( 
.A(n_12096),
.Y(n_12852)
);

INVx1_ASAP7_75t_L g12853 ( 
.A(n_12108),
.Y(n_12853)
);

AND2x2_ASAP7_75t_L g12854 ( 
.A(n_12086),
.B(n_11977),
.Y(n_12854)
);

AND2x2_ASAP7_75t_L g12855 ( 
.A(n_12191),
.B(n_11958),
.Y(n_12855)
);

INVx1_ASAP7_75t_L g12856 ( 
.A(n_12110),
.Y(n_12856)
);

AND2x2_ASAP7_75t_L g12857 ( 
.A(n_12573),
.B(n_11952),
.Y(n_12857)
);

NAND2xp5_ASAP7_75t_L g12858 ( 
.A(n_12392),
.B(n_11855),
.Y(n_12858)
);

INVxp67_ASAP7_75t_SL g12859 ( 
.A(n_12022),
.Y(n_12859)
);

INVxp67_ASAP7_75t_SL g12860 ( 
.A(n_12636),
.Y(n_12860)
);

INVx1_ASAP7_75t_L g12861 ( 
.A(n_12111),
.Y(n_12861)
);

HB1xp67_ASAP7_75t_L g12862 ( 
.A(n_12367),
.Y(n_12862)
);

INVx2_ASAP7_75t_L g12863 ( 
.A(n_12155),
.Y(n_12863)
);

INVx4_ASAP7_75t_L g12864 ( 
.A(n_12172),
.Y(n_12864)
);

INVx1_ASAP7_75t_L g12865 ( 
.A(n_12305),
.Y(n_12865)
);

INVx2_ASAP7_75t_L g12866 ( 
.A(n_12045),
.Y(n_12866)
);

AND2x2_ASAP7_75t_L g12867 ( 
.A(n_12575),
.B(n_11920),
.Y(n_12867)
);

AND2x2_ASAP7_75t_L g12868 ( 
.A(n_12380),
.B(n_11878),
.Y(n_12868)
);

INVx1_ASAP7_75t_L g12869 ( 
.A(n_12050),
.Y(n_12869)
);

INVx1_ASAP7_75t_L g12870 ( 
.A(n_12062),
.Y(n_12870)
);

OR2x2_ASAP7_75t_L g12871 ( 
.A(n_12037),
.B(n_11990),
.Y(n_12871)
);

INVx2_ASAP7_75t_L g12872 ( 
.A(n_12488),
.Y(n_12872)
);

AND2x2_ASAP7_75t_L g12873 ( 
.A(n_12073),
.B(n_11888),
.Y(n_12873)
);

INVx1_ASAP7_75t_L g12874 ( 
.A(n_12068),
.Y(n_12874)
);

BUFx2_ASAP7_75t_L g12875 ( 
.A(n_12584),
.Y(n_12875)
);

INVx2_ASAP7_75t_L g12876 ( 
.A(n_12488),
.Y(n_12876)
);

BUFx2_ASAP7_75t_L g12877 ( 
.A(n_12331),
.Y(n_12877)
);

OR2x2_ASAP7_75t_L g12878 ( 
.A(n_12143),
.B(n_11596),
.Y(n_12878)
);

INVx1_ASAP7_75t_L g12879 ( 
.A(n_12080),
.Y(n_12879)
);

NAND3xp33_ASAP7_75t_L g12880 ( 
.A(n_12029),
.B(n_11923),
.C(n_11918),
.Y(n_12880)
);

INVx2_ASAP7_75t_L g12881 ( 
.A(n_12616),
.Y(n_12881)
);

OR2x2_ASAP7_75t_L g12882 ( 
.A(n_12525),
.B(n_11333),
.Y(n_12882)
);

INVx2_ASAP7_75t_L g12883 ( 
.A(n_12616),
.Y(n_12883)
);

AND2x2_ASAP7_75t_L g12884 ( 
.A(n_12084),
.B(n_11737),
.Y(n_12884)
);

AND2x2_ASAP7_75t_L g12885 ( 
.A(n_12049),
.B(n_11961),
.Y(n_12885)
);

NOR2xp33_ASAP7_75t_L g12886 ( 
.A(n_12175),
.B(n_11490),
.Y(n_12886)
);

NOR2xp33_ASAP7_75t_L g12887 ( 
.A(n_12175),
.B(n_11924),
.Y(n_12887)
);

HB1xp67_ASAP7_75t_L g12888 ( 
.A(n_12286),
.Y(n_12888)
);

INVx1_ASAP7_75t_L g12889 ( 
.A(n_12081),
.Y(n_12889)
);

AND2x4_ASAP7_75t_L g12890 ( 
.A(n_12474),
.B(n_11409),
.Y(n_12890)
);

INVx1_ASAP7_75t_L g12891 ( 
.A(n_12008),
.Y(n_12891)
);

BUFx2_ASAP7_75t_L g12892 ( 
.A(n_12171),
.Y(n_12892)
);

INVx1_ASAP7_75t_L g12893 ( 
.A(n_12003),
.Y(n_12893)
);

HB1xp67_ASAP7_75t_L g12894 ( 
.A(n_12297),
.Y(n_12894)
);

OR2x2_ASAP7_75t_L g12895 ( 
.A(n_12550),
.B(n_12516),
.Y(n_12895)
);

INVx2_ASAP7_75t_L g12896 ( 
.A(n_12443),
.Y(n_12896)
);

HB1xp67_ASAP7_75t_L g12897 ( 
.A(n_12250),
.Y(n_12897)
);

OR2x2_ASAP7_75t_L g12898 ( 
.A(n_12570),
.B(n_11992),
.Y(n_12898)
);

INVx2_ASAP7_75t_L g12899 ( 
.A(n_12393),
.Y(n_12899)
);

BUFx3_ASAP7_75t_L g12900 ( 
.A(n_12166),
.Y(n_12900)
);

HB1xp67_ASAP7_75t_L g12901 ( 
.A(n_12120),
.Y(n_12901)
);

INVx2_ASAP7_75t_L g12902 ( 
.A(n_12282),
.Y(n_12902)
);

AND2x2_ASAP7_75t_L g12903 ( 
.A(n_12404),
.B(n_12470),
.Y(n_12903)
);

AND2x2_ASAP7_75t_L g12904 ( 
.A(n_12568),
.B(n_11970),
.Y(n_12904)
);

INVx2_ASAP7_75t_L g12905 ( 
.A(n_12318),
.Y(n_12905)
);

AND2x2_ASAP7_75t_L g12906 ( 
.A(n_12227),
.B(n_11922),
.Y(n_12906)
);

BUFx3_ASAP7_75t_L g12907 ( 
.A(n_12048),
.Y(n_12907)
);

AND2x4_ASAP7_75t_L g12908 ( 
.A(n_12283),
.B(n_11412),
.Y(n_12908)
);

BUFx2_ASAP7_75t_L g12909 ( 
.A(n_12564),
.Y(n_12909)
);

BUFx3_ASAP7_75t_L g12910 ( 
.A(n_12076),
.Y(n_12910)
);

AND2x2_ASAP7_75t_L g12911 ( 
.A(n_12460),
.B(n_11934),
.Y(n_12911)
);

INVx1_ASAP7_75t_L g12912 ( 
.A(n_12004),
.Y(n_12912)
);

AND2x2_ASAP7_75t_L g12913 ( 
.A(n_12136),
.B(n_11929),
.Y(n_12913)
);

NAND2xp5_ASAP7_75t_L g12914 ( 
.A(n_12588),
.B(n_11419),
.Y(n_12914)
);

BUFx2_ASAP7_75t_L g12915 ( 
.A(n_12007),
.Y(n_12915)
);

INVx1_ASAP7_75t_L g12916 ( 
.A(n_12566),
.Y(n_12916)
);

INVx2_ASAP7_75t_L g12917 ( 
.A(n_12327),
.Y(n_12917)
);

NAND3xp33_ASAP7_75t_L g12918 ( 
.A(n_12410),
.B(n_12528),
.C(n_12193),
.Y(n_12918)
);

AND2x2_ASAP7_75t_L g12919 ( 
.A(n_12101),
.B(n_11913),
.Y(n_12919)
);

INVx1_ASAP7_75t_L g12920 ( 
.A(n_12590),
.Y(n_12920)
);

INVx2_ASAP7_75t_L g12921 ( 
.A(n_12329),
.Y(n_12921)
);

INVx1_ASAP7_75t_L g12922 ( 
.A(n_12112),
.Y(n_12922)
);

HB1xp67_ASAP7_75t_L g12923 ( 
.A(n_12103),
.Y(n_12923)
);

INVx1_ASAP7_75t_L g12924 ( 
.A(n_12115),
.Y(n_12924)
);

INVx2_ASAP7_75t_L g12925 ( 
.A(n_12346),
.Y(n_12925)
);

NOR2xp33_ASAP7_75t_L g12926 ( 
.A(n_12360),
.B(n_11928),
.Y(n_12926)
);

AND2x2_ASAP7_75t_L g12927 ( 
.A(n_12107),
.B(n_11955),
.Y(n_12927)
);

INVx2_ASAP7_75t_L g12928 ( 
.A(n_12480),
.Y(n_12928)
);

BUFx3_ASAP7_75t_L g12929 ( 
.A(n_12364),
.Y(n_12929)
);

INVx1_ASAP7_75t_L g12930 ( 
.A(n_12056),
.Y(n_12930)
);

INVx2_ASAP7_75t_L g12931 ( 
.A(n_12034),
.Y(n_12931)
);

INVx4_ASAP7_75t_L g12932 ( 
.A(n_12260),
.Y(n_12932)
);

INVx1_ASAP7_75t_L g12933 ( 
.A(n_12059),
.Y(n_12933)
);

HB1xp67_ASAP7_75t_L g12934 ( 
.A(n_12117),
.Y(n_12934)
);

INVx3_ASAP7_75t_L g12935 ( 
.A(n_12649),
.Y(n_12935)
);

INVx2_ASAP7_75t_L g12936 ( 
.A(n_12069),
.Y(n_12936)
);

AND2x2_ASAP7_75t_L g12937 ( 
.A(n_12109),
.B(n_11894),
.Y(n_12937)
);

AND2x2_ASAP7_75t_L g12938 ( 
.A(n_12113),
.B(n_11894),
.Y(n_12938)
);

OR2x2_ASAP7_75t_L g12939 ( 
.A(n_12571),
.B(n_11949),
.Y(n_12939)
);

INVx1_ASAP7_75t_L g12940 ( 
.A(n_12467),
.Y(n_12940)
);

AND2x2_ASAP7_75t_L g12941 ( 
.A(n_12119),
.B(n_11817),
.Y(n_12941)
);

AND2x4_ASAP7_75t_L g12942 ( 
.A(n_12649),
.B(n_11495),
.Y(n_12942)
);

AND2x2_ASAP7_75t_L g12943 ( 
.A(n_12430),
.B(n_11817),
.Y(n_12943)
);

AND2x2_ASAP7_75t_L g12944 ( 
.A(n_12473),
.B(n_11942),
.Y(n_12944)
);

BUFx2_ASAP7_75t_SL g12945 ( 
.A(n_12121),
.Y(n_12945)
);

INVx2_ASAP7_75t_L g12946 ( 
.A(n_12069),
.Y(n_12946)
);

INVx2_ASAP7_75t_L g12947 ( 
.A(n_12373),
.Y(n_12947)
);

BUFx2_ASAP7_75t_L g12948 ( 
.A(n_12142),
.Y(n_12948)
);

INVx2_ASAP7_75t_L g12949 ( 
.A(n_12383),
.Y(n_12949)
);

AND2x4_ASAP7_75t_L g12950 ( 
.A(n_12317),
.B(n_11513),
.Y(n_12950)
);

INVx1_ASAP7_75t_L g12951 ( 
.A(n_12482),
.Y(n_12951)
);

AND2x2_ASAP7_75t_L g12952 ( 
.A(n_12014),
.B(n_11944),
.Y(n_12952)
);

OR2x2_ASAP7_75t_L g12953 ( 
.A(n_12576),
.B(n_11624),
.Y(n_12953)
);

INVx2_ASAP7_75t_L g12954 ( 
.A(n_12388),
.Y(n_12954)
);

HB1xp67_ASAP7_75t_L g12955 ( 
.A(n_12177),
.Y(n_12955)
);

INVx2_ASAP7_75t_SL g12956 ( 
.A(n_12548),
.Y(n_12956)
);

INVx1_ASAP7_75t_L g12957 ( 
.A(n_12498),
.Y(n_12957)
);

NOR2xp33_ASAP7_75t_L g12958 ( 
.A(n_12360),
.B(n_11917),
.Y(n_12958)
);

HB1xp67_ASAP7_75t_L g12959 ( 
.A(n_12178),
.Y(n_12959)
);

BUFx2_ASAP7_75t_L g12960 ( 
.A(n_12030),
.Y(n_12960)
);

INVx1_ASAP7_75t_L g12961 ( 
.A(n_12411),
.Y(n_12961)
);

AND2x2_ASAP7_75t_L g12962 ( 
.A(n_12027),
.B(n_11939),
.Y(n_12962)
);

BUFx2_ASAP7_75t_L g12963 ( 
.A(n_12146),
.Y(n_12963)
);

INVx1_ASAP7_75t_L g12964 ( 
.A(n_12425),
.Y(n_12964)
);

NAND2xp5_ASAP7_75t_L g12965 ( 
.A(n_12594),
.B(n_11628),
.Y(n_12965)
);

HB1xp67_ASAP7_75t_L g12966 ( 
.A(n_12192),
.Y(n_12966)
);

INVx2_ASAP7_75t_SL g12967 ( 
.A(n_12559),
.Y(n_12967)
);

OR2x2_ASAP7_75t_L g12968 ( 
.A(n_12344),
.B(n_12629),
.Y(n_12968)
);

INVx3_ASAP7_75t_L g12969 ( 
.A(n_12065),
.Y(n_12969)
);

INVx2_ASAP7_75t_L g12970 ( 
.A(n_12206),
.Y(n_12970)
);

AND2x2_ASAP7_75t_L g12971 ( 
.A(n_12370),
.B(n_11940),
.Y(n_12971)
);

INVx2_ASAP7_75t_L g12972 ( 
.A(n_12005),
.Y(n_12972)
);

OAI33xp33_ASAP7_75t_L g12973 ( 
.A1(n_12199),
.A2(n_11938),
.A3(n_11925),
.B1(n_11918),
.B2(n_11923),
.B3(n_11879),
.Y(n_12973)
);

INVx3_ASAP7_75t_L g12974 ( 
.A(n_12065),
.Y(n_12974)
);

INVx1_ASAP7_75t_L g12975 ( 
.A(n_12441),
.Y(n_12975)
);

HB1xp67_ASAP7_75t_L g12976 ( 
.A(n_12195),
.Y(n_12976)
);

BUFx3_ASAP7_75t_L g12977 ( 
.A(n_12052),
.Y(n_12977)
);

INVx1_ASAP7_75t_L g12978 ( 
.A(n_12442),
.Y(n_12978)
);

AND2x4_ASAP7_75t_L g12979 ( 
.A(n_12322),
.B(n_11633),
.Y(n_12979)
);

AND2x4_ASAP7_75t_L g12980 ( 
.A(n_12440),
.B(n_11634),
.Y(n_12980)
);

HB1xp67_ASAP7_75t_L g12981 ( 
.A(n_12006),
.Y(n_12981)
);

INVx2_ASAP7_75t_L g12982 ( 
.A(n_12013),
.Y(n_12982)
);

HB1xp67_ASAP7_75t_L g12983 ( 
.A(n_12018),
.Y(n_12983)
);

HB1xp67_ASAP7_75t_L g12984 ( 
.A(n_12024),
.Y(n_12984)
);

INVx2_ASAP7_75t_L g12985 ( 
.A(n_12046),
.Y(n_12985)
);

INVx1_ASAP7_75t_L g12986 ( 
.A(n_12454),
.Y(n_12986)
);

INVx2_ASAP7_75t_L g12987 ( 
.A(n_12053),
.Y(n_12987)
);

NAND2xp5_ASAP7_75t_L g12988 ( 
.A(n_12587),
.B(n_11638),
.Y(n_12988)
);

AND2x2_ASAP7_75t_L g12989 ( 
.A(n_12092),
.B(n_11732),
.Y(n_12989)
);

INVx1_ASAP7_75t_L g12990 ( 
.A(n_12540),
.Y(n_12990)
);

INVx1_ASAP7_75t_L g12991 ( 
.A(n_12547),
.Y(n_12991)
);

INVx1_ASAP7_75t_L g12992 ( 
.A(n_12499),
.Y(n_12992)
);

INVx2_ASAP7_75t_L g12993 ( 
.A(n_12054),
.Y(n_12993)
);

BUFx2_ASAP7_75t_L g12994 ( 
.A(n_12146),
.Y(n_12994)
);

NAND2xp5_ASAP7_75t_L g12995 ( 
.A(n_12216),
.B(n_11663),
.Y(n_12995)
);

AND2x2_ASAP7_75t_L g12996 ( 
.A(n_12138),
.B(n_11664),
.Y(n_12996)
);

AND2x2_ASAP7_75t_L g12997 ( 
.A(n_12061),
.B(n_11665),
.Y(n_12997)
);

INVx1_ASAP7_75t_L g12998 ( 
.A(n_12509),
.Y(n_12998)
);

INVx1_ASAP7_75t_L g12999 ( 
.A(n_12521),
.Y(n_12999)
);

AND2x2_ASAP7_75t_L g13000 ( 
.A(n_12063),
.B(n_11968),
.Y(n_13000)
);

INVx2_ASAP7_75t_L g13001 ( 
.A(n_12064),
.Y(n_13001)
);

INVx2_ASAP7_75t_L g13002 ( 
.A(n_12070),
.Y(n_13002)
);

INVx2_ASAP7_75t_SL g13003 ( 
.A(n_12028),
.Y(n_13003)
);

HB1xp67_ASAP7_75t_L g13004 ( 
.A(n_12090),
.Y(n_13004)
);

OAI31xp33_ASAP7_75t_SL g13005 ( 
.A1(n_12196),
.A2(n_11568),
.A3(n_11534),
.B(n_11730),
.Y(n_13005)
);

NAND2xp5_ASAP7_75t_L g13006 ( 
.A(n_12538),
.B(n_11896),
.Y(n_13006)
);

INVx1_ASAP7_75t_L g13007 ( 
.A(n_12535),
.Y(n_13007)
);

NAND2xp5_ASAP7_75t_L g13008 ( 
.A(n_12538),
.B(n_11616),
.Y(n_13008)
);

AND2x2_ASAP7_75t_L g13009 ( 
.A(n_12581),
.B(n_11705),
.Y(n_13009)
);

INVx2_ASAP7_75t_L g13010 ( 
.A(n_12394),
.Y(n_13010)
);

INVx1_ASAP7_75t_L g13011 ( 
.A(n_12180),
.Y(n_13011)
);

INVx2_ASAP7_75t_L g13012 ( 
.A(n_12258),
.Y(n_13012)
);

INVx2_ASAP7_75t_L g13013 ( 
.A(n_12270),
.Y(n_13013)
);

NAND2xp5_ASAP7_75t_L g13014 ( 
.A(n_12231),
.B(n_12275),
.Y(n_13014)
);

OR2x2_ASAP7_75t_L g13015 ( 
.A(n_12237),
.B(n_11763),
.Y(n_13015)
);

INVx3_ASAP7_75t_L g13016 ( 
.A(n_12028),
.Y(n_13016)
);

INVxp67_ASAP7_75t_L g13017 ( 
.A(n_12051),
.Y(n_13017)
);

AND2x2_ASAP7_75t_L g13018 ( 
.A(n_12508),
.B(n_11822),
.Y(n_13018)
);

NOR2xp33_ASAP7_75t_L g13019 ( 
.A(n_12319),
.B(n_11646),
.Y(n_13019)
);

INVx2_ASAP7_75t_L g13020 ( 
.A(n_12463),
.Y(n_13020)
);

AND2x2_ASAP7_75t_L g13021 ( 
.A(n_12122),
.B(n_11646),
.Y(n_13021)
);

NAND2xp5_ASAP7_75t_L g13022 ( 
.A(n_12278),
.B(n_11653),
.Y(n_13022)
);

INVx1_ASAP7_75t_L g13023 ( 
.A(n_12183),
.Y(n_13023)
);

INVx1_ASAP7_75t_L g13024 ( 
.A(n_12235),
.Y(n_13024)
);

AND2x2_ASAP7_75t_L g13025 ( 
.A(n_12055),
.B(n_12093),
.Y(n_13025)
);

INVx1_ASAP7_75t_L g13026 ( 
.A(n_12198),
.Y(n_13026)
);

INVx3_ASAP7_75t_L g13027 ( 
.A(n_12463),
.Y(n_13027)
);

OR2x2_ASAP7_75t_L g13028 ( 
.A(n_12625),
.B(n_11740),
.Y(n_13028)
);

OR2x2_ASAP7_75t_L g13029 ( 
.A(n_12560),
.B(n_12233),
.Y(n_13029)
);

BUFx3_ASAP7_75t_L g13030 ( 
.A(n_12031),
.Y(n_13030)
);

AND2x2_ASAP7_75t_L g13031 ( 
.A(n_12654),
.B(n_12208),
.Y(n_13031)
);

INVx1_ASAP7_75t_L g13032 ( 
.A(n_12140),
.Y(n_13032)
);

INVxp67_ASAP7_75t_SL g13033 ( 
.A(n_12039),
.Y(n_13033)
);

AND2x2_ASAP7_75t_L g13034 ( 
.A(n_12219),
.B(n_11653),
.Y(n_13034)
);

HB1xp67_ASAP7_75t_L g13035 ( 
.A(n_12125),
.Y(n_13035)
);

INVx2_ASAP7_75t_L g13036 ( 
.A(n_12273),
.Y(n_13036)
);

AND2x2_ASAP7_75t_L g13037 ( 
.A(n_12396),
.B(n_11679),
.Y(n_13037)
);

BUFx6f_ASAP7_75t_L g13038 ( 
.A(n_12124),
.Y(n_13038)
);

NOR2xp67_ASAP7_75t_L g13039 ( 
.A(n_12593),
.B(n_11773),
.Y(n_13039)
);

INVx1_ASAP7_75t_L g13040 ( 
.A(n_12123),
.Y(n_13040)
);

AND2x2_ASAP7_75t_L g13041 ( 
.A(n_12555),
.B(n_11679),
.Y(n_13041)
);

INVx1_ASAP7_75t_L g13042 ( 
.A(n_12211),
.Y(n_13042)
);

AND2x2_ASAP7_75t_L g13043 ( 
.A(n_12561),
.B(n_11797),
.Y(n_13043)
);

INVx1_ASAP7_75t_L g13044 ( 
.A(n_12212),
.Y(n_13044)
);

AOI22xp33_ASAP7_75t_L g13045 ( 
.A1(n_12134),
.A2(n_11983),
.B1(n_11988),
.B2(n_11984),
.Y(n_13045)
);

AND2x2_ASAP7_75t_L g13046 ( 
.A(n_12543),
.B(n_11798),
.Y(n_13046)
);

INVx1_ASAP7_75t_L g13047 ( 
.A(n_12078),
.Y(n_13047)
);

AND2x2_ASAP7_75t_L g13048 ( 
.A(n_12542),
.B(n_11776),
.Y(n_13048)
);

OR2x2_ASAP7_75t_L g13049 ( 
.A(n_12536),
.B(n_11747),
.Y(n_13049)
);

AND2x2_ASAP7_75t_L g13050 ( 
.A(n_12095),
.B(n_11813),
.Y(n_13050)
);

HB1xp67_ASAP7_75t_L g13051 ( 
.A(n_12159),
.Y(n_13051)
);

AND2x4_ASAP7_75t_L g13052 ( 
.A(n_12280),
.B(n_11656),
.Y(n_13052)
);

OAI221xp5_ASAP7_75t_L g13053 ( 
.A1(n_12179),
.A2(n_11394),
.B1(n_11655),
.B2(n_11916),
.C(n_11722),
.Y(n_13053)
);

INVx1_ASAP7_75t_L g13054 ( 
.A(n_12141),
.Y(n_13054)
);

AND2x2_ASAP7_75t_L g13055 ( 
.A(n_12097),
.B(n_11774),
.Y(n_13055)
);

OR2x6_ASAP7_75t_L g13056 ( 
.A(n_12477),
.B(n_12288),
.Y(n_13056)
);

INVx1_ASAP7_75t_L g13057 ( 
.A(n_12147),
.Y(n_13057)
);

HB1xp67_ASAP7_75t_L g13058 ( 
.A(n_12163),
.Y(n_13058)
);

INVxp67_ASAP7_75t_SL g13059 ( 
.A(n_12088),
.Y(n_13059)
);

NOR2xp67_ASAP7_75t_L g13060 ( 
.A(n_12457),
.B(n_11994),
.Y(n_13060)
);

INVx1_ASAP7_75t_L g13061 ( 
.A(n_12151),
.Y(n_13061)
);

INVx2_ASAP7_75t_L g13062 ( 
.A(n_12230),
.Y(n_13062)
);

HB1xp67_ASAP7_75t_L g13063 ( 
.A(n_12174),
.Y(n_13063)
);

INVx2_ASAP7_75t_L g13064 ( 
.A(n_12244),
.Y(n_13064)
);

INVx2_ASAP7_75t_L g13065 ( 
.A(n_12245),
.Y(n_13065)
);

INVx2_ASAP7_75t_L g13066 ( 
.A(n_12289),
.Y(n_13066)
);

NAND2x1p5_ASAP7_75t_L g13067 ( 
.A(n_12234),
.B(n_7987),
.Y(n_13067)
);

INVx1_ASAP7_75t_L g13068 ( 
.A(n_12153),
.Y(n_13068)
);

AND2x2_ASAP7_75t_L g13069 ( 
.A(n_12099),
.B(n_11994),
.Y(n_13069)
);

OR2x6_ASAP7_75t_L g13070 ( 
.A(n_12477),
.B(n_11815),
.Y(n_13070)
);

INVx1_ASAP7_75t_L g13071 ( 
.A(n_12154),
.Y(n_13071)
);

AND2x2_ASAP7_75t_L g13072 ( 
.A(n_12332),
.B(n_11574),
.Y(n_13072)
);

INVx2_ASAP7_75t_L g13073 ( 
.A(n_12294),
.Y(n_13073)
);

HB1xp67_ASAP7_75t_L g13074 ( 
.A(n_12617),
.Y(n_13074)
);

OR2x2_ASAP7_75t_L g13075 ( 
.A(n_12032),
.B(n_11971),
.Y(n_13075)
);

INVxp67_ASAP7_75t_L g13076 ( 
.A(n_12129),
.Y(n_13076)
);

AOI22xp33_ASAP7_75t_L g13077 ( 
.A1(n_12094),
.A2(n_11988),
.B1(n_11984),
.B2(n_11993),
.Y(n_13077)
);

INVx1_ASAP7_75t_L g13078 ( 
.A(n_12156),
.Y(n_13078)
);

INVx2_ASAP7_75t_L g13079 ( 
.A(n_12298),
.Y(n_13079)
);

AO21x2_ASAP7_75t_L g13080 ( 
.A1(n_12023),
.A2(n_11696),
.B(n_11692),
.Y(n_13080)
);

OR2x2_ASAP7_75t_L g13081 ( 
.A(n_12554),
.B(n_11771),
.Y(n_13081)
);

INVx1_ASAP7_75t_L g13082 ( 
.A(n_12160),
.Y(n_13082)
);

NAND2xp5_ASAP7_75t_L g13083 ( 
.A(n_12020),
.B(n_11890),
.Y(n_13083)
);

INVx2_ASAP7_75t_L g13084 ( 
.A(n_12309),
.Y(n_13084)
);

OR2x2_ASAP7_75t_L g13085 ( 
.A(n_12220),
.B(n_11778),
.Y(n_13085)
);

AND2x2_ASAP7_75t_L g13086 ( 
.A(n_12338),
.B(n_11675),
.Y(n_13086)
);

AND2x2_ASAP7_75t_L g13087 ( 
.A(n_12252),
.B(n_12257),
.Y(n_13087)
);

INVx2_ASAP7_75t_SL g13088 ( 
.A(n_12645),
.Y(n_13088)
);

AND2x2_ASAP7_75t_L g13089 ( 
.A(n_12585),
.B(n_11676),
.Y(n_13089)
);

BUFx2_ASAP7_75t_L g13090 ( 
.A(n_12457),
.Y(n_13090)
);

AOI22xp33_ASAP7_75t_L g13091 ( 
.A1(n_12043),
.A2(n_11993),
.B1(n_11881),
.B2(n_11890),
.Y(n_13091)
);

INVx2_ASAP7_75t_L g13092 ( 
.A(n_12145),
.Y(n_13092)
);

HB1xp67_ASAP7_75t_L g13093 ( 
.A(n_12620),
.Y(n_13093)
);

INVx1_ASAP7_75t_L g13094 ( 
.A(n_12165),
.Y(n_13094)
);

INVx3_ASAP7_75t_L g13095 ( 
.A(n_12400),
.Y(n_13095)
);

INVx1_ASAP7_75t_L g13096 ( 
.A(n_12167),
.Y(n_13096)
);

AND2x2_ASAP7_75t_L g13097 ( 
.A(n_12589),
.B(n_11947),
.Y(n_13097)
);

INVx1_ASAP7_75t_L g13098 ( 
.A(n_12168),
.Y(n_13098)
);

HB1xp67_ASAP7_75t_L g13099 ( 
.A(n_12630),
.Y(n_13099)
);

INVx1_ASAP7_75t_L g13100 ( 
.A(n_12169),
.Y(n_13100)
);

AND2x2_ASAP7_75t_L g13101 ( 
.A(n_12592),
.B(n_11543),
.Y(n_13101)
);

AOI22xp5_ASAP7_75t_L g13102 ( 
.A1(n_12042),
.A2(n_11842),
.B1(n_11852),
.B2(n_11876),
.Y(n_13102)
);

AND2x2_ASAP7_75t_L g13103 ( 
.A(n_12598),
.B(n_11546),
.Y(n_13103)
);

AND2x2_ASAP7_75t_L g13104 ( 
.A(n_12619),
.B(n_11555),
.Y(n_13104)
);

INVx1_ASAP7_75t_L g13105 ( 
.A(n_12181),
.Y(n_13105)
);

AND2x2_ASAP7_75t_L g13106 ( 
.A(n_12622),
.B(n_12639),
.Y(n_13106)
);

INVx1_ASAP7_75t_L g13107 ( 
.A(n_12184),
.Y(n_13107)
);

INVx2_ASAP7_75t_L g13108 ( 
.A(n_12148),
.Y(n_13108)
);

AO21x2_ASAP7_75t_L g13109 ( 
.A1(n_12161),
.A2(n_11692),
.B(n_11706),
.Y(n_13109)
);

AND2x2_ASAP7_75t_L g13110 ( 
.A(n_12369),
.B(n_11846),
.Y(n_13110)
);

AND2x2_ASAP7_75t_L g13111 ( 
.A(n_12631),
.B(n_6941),
.Y(n_13111)
);

NAND2xp5_ASAP7_75t_L g13112 ( 
.A(n_12291),
.B(n_11842),
.Y(n_13112)
);

AND2x2_ASAP7_75t_L g13113 ( 
.A(n_12635),
.B(n_6960),
.Y(n_13113)
);

INVx5_ASAP7_75t_L g13114 ( 
.A(n_12519),
.Y(n_13114)
);

OR2x2_ASAP7_75t_L g13115 ( 
.A(n_12274),
.B(n_12323),
.Y(n_13115)
);

INVx2_ASAP7_75t_L g13116 ( 
.A(n_12149),
.Y(n_13116)
);

AND2x4_ASAP7_75t_L g13117 ( 
.A(n_12296),
.B(n_11666),
.Y(n_13117)
);

INVx2_ASAP7_75t_L g13118 ( 
.A(n_12170),
.Y(n_13118)
);

AND2x2_ASAP7_75t_L g13119 ( 
.A(n_12643),
.B(n_6960),
.Y(n_13119)
);

BUFx2_ASAP7_75t_L g13120 ( 
.A(n_12011),
.Y(n_13120)
);

OR2x2_ASAP7_75t_L g13121 ( 
.A(n_12336),
.B(n_11854),
.Y(n_13121)
);

INVx1_ASAP7_75t_L g13122 ( 
.A(n_12186),
.Y(n_13122)
);

AND2x2_ASAP7_75t_L g13123 ( 
.A(n_12644),
.B(n_6971),
.Y(n_13123)
);

AND2x2_ASAP7_75t_L g13124 ( 
.A(n_12530),
.B(n_6971),
.Y(n_13124)
);

HB1xp67_ASAP7_75t_L g13125 ( 
.A(n_12334),
.Y(n_13125)
);

INVx2_ASAP7_75t_L g13126 ( 
.A(n_12176),
.Y(n_13126)
);

HB1xp67_ASAP7_75t_L g13127 ( 
.A(n_12339),
.Y(n_13127)
);

NAND2xp5_ASAP7_75t_L g13128 ( 
.A(n_12377),
.B(n_11408),
.Y(n_13128)
);

INVx1_ASAP7_75t_L g13129 ( 
.A(n_12190),
.Y(n_13129)
);

OR2x2_ASAP7_75t_L g13130 ( 
.A(n_12351),
.B(n_11870),
.Y(n_13130)
);

INVx2_ASAP7_75t_L g13131 ( 
.A(n_12182),
.Y(n_13131)
);

NAND2xp5_ASAP7_75t_L g13132 ( 
.A(n_12385),
.B(n_11408),
.Y(n_13132)
);

INVx3_ASAP7_75t_L g13133 ( 
.A(n_12400),
.Y(n_13133)
);

BUFx2_ASAP7_75t_L g13134 ( 
.A(n_12019),
.Y(n_13134)
);

AND2x2_ASAP7_75t_L g13135 ( 
.A(n_12533),
.B(n_7004),
.Y(n_13135)
);

AND2x2_ASAP7_75t_L g13136 ( 
.A(n_12527),
.B(n_7004),
.Y(n_13136)
);

INVx2_ASAP7_75t_L g13137 ( 
.A(n_12189),
.Y(n_13137)
);

AND2x2_ASAP7_75t_L g13138 ( 
.A(n_12409),
.B(n_11962),
.Y(n_13138)
);

INVx3_ASAP7_75t_L g13139 ( 
.A(n_12423),
.Y(n_13139)
);

AND2x2_ASAP7_75t_L g13140 ( 
.A(n_12428),
.B(n_11962),
.Y(n_13140)
);

NAND2xp5_ASAP7_75t_L g13141 ( 
.A(n_12399),
.B(n_11408),
.Y(n_13141)
);

AO21x2_ASAP7_75t_L g13142 ( 
.A1(n_12349),
.A2(n_12413),
.B(n_12310),
.Y(n_13142)
);

INVx2_ASAP7_75t_L g13143 ( 
.A(n_12217),
.Y(n_13143)
);

AND2x2_ASAP7_75t_L g13144 ( 
.A(n_12501),
.B(n_11962),
.Y(n_13144)
);

INVx2_ASAP7_75t_L g13145 ( 
.A(n_12432),
.Y(n_13145)
);

AND2x2_ASAP7_75t_L g13146 ( 
.A(n_12365),
.B(n_8289),
.Y(n_13146)
);

HB1xp67_ASAP7_75t_L g13147 ( 
.A(n_12524),
.Y(n_13147)
);

INVx3_ASAP7_75t_L g13148 ( 
.A(n_12423),
.Y(n_13148)
);

INVx1_ASAP7_75t_L g13149 ( 
.A(n_12201),
.Y(n_13149)
);

INVx1_ASAP7_75t_L g13150 ( 
.A(n_12202),
.Y(n_13150)
);

AND2x2_ASAP7_75t_L g13151 ( 
.A(n_12066),
.B(n_9243),
.Y(n_13151)
);

INVx1_ASAP7_75t_L g13152 ( 
.A(n_12203),
.Y(n_13152)
);

BUFx2_ASAP7_75t_L g13153 ( 
.A(n_12038),
.Y(n_13153)
);

OAI21xp5_ASAP7_75t_SL g13154 ( 
.A1(n_12419),
.A2(n_11861),
.B(n_11860),
.Y(n_13154)
);

OR2x2_ASAP7_75t_L g13155 ( 
.A(n_12353),
.B(n_11835),
.Y(n_13155)
);

AND2x2_ASAP7_75t_L g13156 ( 
.A(n_12067),
.B(n_9246),
.Y(n_13156)
);

AND2x2_ASAP7_75t_L g13157 ( 
.A(n_12356),
.B(n_9284),
.Y(n_13157)
);

NOR2xp33_ASAP7_75t_L g13158 ( 
.A(n_12187),
.B(n_11818),
.Y(n_13158)
);

INVx2_ASAP7_75t_SL g13159 ( 
.A(n_12341),
.Y(n_13159)
);

AND2x2_ASAP7_75t_L g13160 ( 
.A(n_12503),
.B(n_9320),
.Y(n_13160)
);

AND2x2_ASAP7_75t_L g13161 ( 
.A(n_12518),
.B(n_9339),
.Y(n_13161)
);

OR2x2_ASAP7_75t_L g13162 ( 
.A(n_12337),
.B(n_11835),
.Y(n_13162)
);

AOI221xp5_ASAP7_75t_L g13163 ( 
.A1(n_12405),
.A2(n_11904),
.B1(n_11905),
.B2(n_11881),
.C(n_11828),
.Y(n_13163)
);

AND2x2_ASAP7_75t_L g13164 ( 
.A(n_12522),
.B(n_9351),
.Y(n_13164)
);

INVx1_ASAP7_75t_SL g13165 ( 
.A(n_12376),
.Y(n_13165)
);

NAND2xp5_ASAP7_75t_L g13166 ( 
.A(n_12418),
.B(n_11858),
.Y(n_13166)
);

BUFx3_ASAP7_75t_L g13167 ( 
.A(n_12497),
.Y(n_13167)
);

INVx2_ASAP7_75t_L g13168 ( 
.A(n_12471),
.Y(n_13168)
);

AND2x2_ASAP7_75t_L g13169 ( 
.A(n_12523),
.B(n_9358),
.Y(n_13169)
);

INVx2_ASAP7_75t_L g13170 ( 
.A(n_12472),
.Y(n_13170)
);

AND2x2_ASAP7_75t_L g13171 ( 
.A(n_12567),
.B(n_9374),
.Y(n_13171)
);

BUFx6f_ASAP7_75t_L g13172 ( 
.A(n_12422),
.Y(n_13172)
);

AND2x2_ASAP7_75t_L g13173 ( 
.A(n_12609),
.B(n_9392),
.Y(n_13173)
);

INVx2_ASAP7_75t_L g13174 ( 
.A(n_12452),
.Y(n_13174)
);

AND2x2_ASAP7_75t_L g13175 ( 
.A(n_12452),
.B(n_10177),
.Y(n_13175)
);

INVx1_ASAP7_75t_L g13176 ( 
.A(n_12204),
.Y(n_13176)
);

OR2x2_ASAP7_75t_L g13177 ( 
.A(n_12552),
.B(n_11848),
.Y(n_13177)
);

INVx1_ASAP7_75t_L g13178 ( 
.A(n_12210),
.Y(n_13178)
);

BUFx4f_ASAP7_75t_L g13179 ( 
.A(n_12438),
.Y(n_13179)
);

INVx1_ASAP7_75t_L g13180 ( 
.A(n_12213),
.Y(n_13180)
);

AND2x2_ASAP7_75t_L g13181 ( 
.A(n_12456),
.B(n_10196),
.Y(n_13181)
);

INVx3_ASAP7_75t_L g13182 ( 
.A(n_12469),
.Y(n_13182)
);

INVx1_ASAP7_75t_L g13183 ( 
.A(n_12218),
.Y(n_13183)
);

NAND2xp5_ASAP7_75t_L g13184 ( 
.A(n_12496),
.B(n_11858),
.Y(n_13184)
);

INVx1_ASAP7_75t_SL g13185 ( 
.A(n_12041),
.Y(n_13185)
);

INVx2_ASAP7_75t_L g13186 ( 
.A(n_12519),
.Y(n_13186)
);

INVx1_ASAP7_75t_L g13187 ( 
.A(n_12222),
.Y(n_13187)
);

INVx2_ASAP7_75t_L g13188 ( 
.A(n_12224),
.Y(n_13188)
);

INVx1_ASAP7_75t_L g13189 ( 
.A(n_12223),
.Y(n_13189)
);

AND2x2_ASAP7_75t_L g13190 ( 
.A(n_12526),
.B(n_10197),
.Y(n_13190)
);

AND2x2_ASAP7_75t_L g13191 ( 
.A(n_12529),
.B(n_10200),
.Y(n_13191)
);

AND2x2_ASAP7_75t_L g13192 ( 
.A(n_12532),
.B(n_10201),
.Y(n_13192)
);

INVxp67_ASAP7_75t_SL g13193 ( 
.A(n_12624),
.Y(n_13193)
);

AND2x2_ASAP7_75t_L g13194 ( 
.A(n_12569),
.B(n_10205),
.Y(n_13194)
);

BUFx2_ASAP7_75t_L g13195 ( 
.A(n_12040),
.Y(n_13195)
);

INVx1_ASAP7_75t_L g13196 ( 
.A(n_12225),
.Y(n_13196)
);

OR2x2_ASAP7_75t_L g13197 ( 
.A(n_12384),
.B(n_12415),
.Y(n_13197)
);

INVx1_ASAP7_75t_L g13198 ( 
.A(n_12229),
.Y(n_13198)
);

INVx4_ASAP7_75t_L g13199 ( 
.A(n_12572),
.Y(n_13199)
);

BUFx2_ASAP7_75t_L g13200 ( 
.A(n_12306),
.Y(n_13200)
);

INVx1_ASAP7_75t_L g13201 ( 
.A(n_12236),
.Y(n_13201)
);

INVx2_ASAP7_75t_L g13202 ( 
.A(n_12224),
.Y(n_13202)
);

INVxp67_ASAP7_75t_SL g13203 ( 
.A(n_12638),
.Y(n_13203)
);

AND2x4_ASAP7_75t_L g13204 ( 
.A(n_12574),
.B(n_11713),
.Y(n_13204)
);

BUFx2_ASAP7_75t_L g13205 ( 
.A(n_12315),
.Y(n_13205)
);

AND2x2_ASAP7_75t_L g13206 ( 
.A(n_12578),
.B(n_10206),
.Y(n_13206)
);

NAND2xp5_ASAP7_75t_L g13207 ( 
.A(n_12478),
.B(n_11874),
.Y(n_13207)
);

NAND2xp5_ASAP7_75t_L g13208 ( 
.A(n_12116),
.B(n_11874),
.Y(n_13208)
);

INVxp67_ASAP7_75t_SL g13209 ( 
.A(n_12386),
.Y(n_13209)
);

INVx1_ASAP7_75t_L g13210 ( 
.A(n_12240),
.Y(n_13210)
);

OR2x2_ASAP7_75t_L g13211 ( 
.A(n_12628),
.B(n_11821),
.Y(n_13211)
);

AND2x2_ASAP7_75t_L g13212 ( 
.A(n_12127),
.B(n_10210),
.Y(n_13212)
);

NAND2xp5_ASAP7_75t_L g13213 ( 
.A(n_12133),
.B(n_11877),
.Y(n_13213)
);

HB1xp67_ASAP7_75t_L g13214 ( 
.A(n_12135),
.Y(n_13214)
);

OR2x2_ASAP7_75t_L g13215 ( 
.A(n_12137),
.B(n_11825),
.Y(n_13215)
);

INVx2_ASAP7_75t_L g13216 ( 
.A(n_12608),
.Y(n_13216)
);

HB1xp67_ASAP7_75t_L g13217 ( 
.A(n_12611),
.Y(n_13217)
);

NAND2x1p5_ASAP7_75t_L g13218 ( 
.A(n_12269),
.B(n_7987),
.Y(n_13218)
);

NOR2xp67_ASAP7_75t_L g13219 ( 
.A(n_12381),
.B(n_11727),
.Y(n_13219)
);

AND2x2_ASAP7_75t_L g13220 ( 
.A(n_12613),
.B(n_10213),
.Y(n_13220)
);

INVx2_ASAP7_75t_L g13221 ( 
.A(n_12615),
.Y(n_13221)
);

INVx1_ASAP7_75t_L g13222 ( 
.A(n_12247),
.Y(n_13222)
);

INVx1_ASAP7_75t_L g13223 ( 
.A(n_12254),
.Y(n_13223)
);

HB1xp67_ASAP7_75t_L g13224 ( 
.A(n_12646),
.Y(n_13224)
);

BUFx6f_ASAP7_75t_L g13225 ( 
.A(n_12491),
.Y(n_13225)
);

INVx2_ASAP7_75t_L g13226 ( 
.A(n_12114),
.Y(n_13226)
);

INVx2_ASAP7_75t_L g13227 ( 
.A(n_12732),
.Y(n_13227)
);

AND2x2_ASAP7_75t_L g13228 ( 
.A(n_12732),
.B(n_12671),
.Y(n_13228)
);

AND2x4_ASAP7_75t_L g13229 ( 
.A(n_12669),
.B(n_12259),
.Y(n_13229)
);

INVx1_ASAP7_75t_L g13230 ( 
.A(n_12779),
.Y(n_13230)
);

INVx1_ASAP7_75t_L g13231 ( 
.A(n_12790),
.Y(n_13231)
);

INVx1_ASAP7_75t_L g13232 ( 
.A(n_12817),
.Y(n_13232)
);

OR2x2_ASAP7_75t_L g13233 ( 
.A(n_12713),
.B(n_12251),
.Y(n_13233)
);

INVx2_ASAP7_75t_L g13234 ( 
.A(n_12697),
.Y(n_13234)
);

HB1xp67_ASAP7_75t_L g13235 ( 
.A(n_12802),
.Y(n_13235)
);

INVx1_ASAP7_75t_L g13236 ( 
.A(n_12711),
.Y(n_13236)
);

AND2x2_ASAP7_75t_L g13237 ( 
.A(n_12697),
.B(n_12268),
.Y(n_13237)
);

AND2x2_ASAP7_75t_L g13238 ( 
.A(n_12684),
.B(n_12285),
.Y(n_13238)
);

AND2x2_ASAP7_75t_L g13239 ( 
.A(n_12903),
.B(n_12290),
.Y(n_13239)
);

AND2x4_ASAP7_75t_L g13240 ( 
.A(n_12675),
.B(n_12261),
.Y(n_13240)
);

INVx2_ASAP7_75t_L g13241 ( 
.A(n_12751),
.Y(n_13241)
);

HB1xp67_ASAP7_75t_L g13242 ( 
.A(n_13056),
.Y(n_13242)
);

INVx1_ASAP7_75t_L g13243 ( 
.A(n_12711),
.Y(n_13243)
);

NOR2xp33_ASAP7_75t_L g13244 ( 
.A(n_13165),
.B(n_12330),
.Y(n_13244)
);

NAND2xp5_ASAP7_75t_L g13245 ( 
.A(n_12948),
.B(n_12185),
.Y(n_13245)
);

HB1xp67_ASAP7_75t_L g13246 ( 
.A(n_13056),
.Y(n_13246)
);

AND2x2_ASAP7_75t_L g13247 ( 
.A(n_12731),
.B(n_12188),
.Y(n_13247)
);

AND2x2_ASAP7_75t_L g13248 ( 
.A(n_12753),
.B(n_12266),
.Y(n_13248)
);

INVx1_ASAP7_75t_L g13249 ( 
.A(n_12716),
.Y(n_13249)
);

AND2x2_ASAP7_75t_L g13250 ( 
.A(n_12693),
.B(n_12267),
.Y(n_13250)
);

AND2x2_ASAP7_75t_SL g13251 ( 
.A(n_12915),
.B(n_11860),
.Y(n_13251)
);

AND2x2_ASAP7_75t_L g13252 ( 
.A(n_12724),
.B(n_12272),
.Y(n_13252)
);

OR2x2_ASAP7_75t_L g13253 ( 
.A(n_12721),
.B(n_12335),
.Y(n_13253)
);

INVx1_ASAP7_75t_L g13254 ( 
.A(n_12716),
.Y(n_13254)
);

AND2x2_ASAP7_75t_L g13255 ( 
.A(n_12796),
.B(n_12276),
.Y(n_13255)
);

OR2x2_ASAP7_75t_L g13256 ( 
.A(n_12659),
.B(n_12342),
.Y(n_13256)
);

INVx2_ASAP7_75t_L g13257 ( 
.A(n_12751),
.Y(n_13257)
);

INVx1_ASAP7_75t_L g13258 ( 
.A(n_12720),
.Y(n_13258)
);

OR2x2_ASAP7_75t_L g13259 ( 
.A(n_12699),
.B(n_12417),
.Y(n_13259)
);

NAND2x1_ASAP7_75t_SL g13260 ( 
.A(n_12691),
.B(n_11731),
.Y(n_13260)
);

INVx2_ASAP7_75t_L g13261 ( 
.A(n_12702),
.Y(n_13261)
);

NAND2xp5_ASAP7_75t_L g13262 ( 
.A(n_12948),
.B(n_12421),
.Y(n_13262)
);

AND2x4_ASAP7_75t_SL g13263 ( 
.A(n_12765),
.B(n_12279),
.Y(n_13263)
);

AND2x2_ASAP7_75t_L g13264 ( 
.A(n_12656),
.B(n_12281),
.Y(n_13264)
);

BUFx2_ASAP7_75t_L g13265 ( 
.A(n_12846),
.Y(n_13265)
);

INVx2_ASAP7_75t_L g13266 ( 
.A(n_12702),
.Y(n_13266)
);

HB1xp67_ASAP7_75t_L g13267 ( 
.A(n_12705),
.Y(n_13267)
);

OA211x2_ASAP7_75t_L g13268 ( 
.A1(n_12668),
.A2(n_12958),
.B(n_12794),
.C(n_12926),
.Y(n_13268)
);

AND2x2_ASAP7_75t_L g13269 ( 
.A(n_12715),
.B(n_12284),
.Y(n_13269)
);

INVx1_ASAP7_75t_L g13270 ( 
.A(n_12720),
.Y(n_13270)
);

AND2x4_ASAP7_75t_L g13271 ( 
.A(n_12805),
.B(n_12292),
.Y(n_13271)
);

INVx1_ASAP7_75t_L g13272 ( 
.A(n_12888),
.Y(n_13272)
);

INVx1_ASAP7_75t_L g13273 ( 
.A(n_12894),
.Y(n_13273)
);

INVx2_ASAP7_75t_L g13274 ( 
.A(n_12771),
.Y(n_13274)
);

NAND2xp5_ASAP7_75t_L g13275 ( 
.A(n_13209),
.B(n_12455),
.Y(n_13275)
);

INVx1_ASAP7_75t_L g13276 ( 
.A(n_12681),
.Y(n_13276)
);

AND2x2_ASAP7_75t_L g13277 ( 
.A(n_12682),
.B(n_12316),
.Y(n_13277)
);

AND2x2_ASAP7_75t_L g13278 ( 
.A(n_12717),
.B(n_12326),
.Y(n_13278)
);

INVx2_ASAP7_75t_L g13279 ( 
.A(n_12771),
.Y(n_13279)
);

HB1xp67_ASAP7_75t_L g13280 ( 
.A(n_12705),
.Y(n_13280)
);

NAND2xp5_ASAP7_75t_L g13281 ( 
.A(n_12738),
.B(n_12495),
.Y(n_13281)
);

AND2x2_ASAP7_75t_L g13282 ( 
.A(n_12722),
.B(n_12348),
.Y(n_13282)
);

INVxp67_ASAP7_75t_SL g13283 ( 
.A(n_12846),
.Y(n_13283)
);

AND2x2_ASAP7_75t_L g13284 ( 
.A(n_12840),
.B(n_12357),
.Y(n_13284)
);

AND2x2_ASAP7_75t_L g13285 ( 
.A(n_12686),
.B(n_12362),
.Y(n_13285)
);

AND2x2_ASAP7_75t_L g13286 ( 
.A(n_13106),
.B(n_12363),
.Y(n_13286)
);

OR2x2_ASAP7_75t_L g13287 ( 
.A(n_12776),
.B(n_12600),
.Y(n_13287)
);

NOR3xp33_ASAP7_75t_L g13288 ( 
.A(n_12880),
.B(n_12238),
.C(n_12228),
.Y(n_13288)
);

INVx1_ASAP7_75t_L g13289 ( 
.A(n_12843),
.Y(n_13289)
);

NAND2xp5_ASAP7_75t_L g13290 ( 
.A(n_12679),
.B(n_12371),
.Y(n_13290)
);

INVx3_ASAP7_75t_L g13291 ( 
.A(n_12663),
.Y(n_13291)
);

AND2x2_ASAP7_75t_L g13292 ( 
.A(n_12655),
.B(n_12375),
.Y(n_13292)
);

AND2x2_ASAP7_75t_L g13293 ( 
.A(n_12658),
.B(n_12740),
.Y(n_13293)
);

AND2x2_ASAP7_75t_L g13294 ( 
.A(n_13136),
.B(n_12855),
.Y(n_13294)
);

INVx2_ASAP7_75t_L g13295 ( 
.A(n_12663),
.Y(n_13295)
);

OR2x2_ASAP7_75t_L g13296 ( 
.A(n_13115),
.B(n_12758),
.Y(n_13296)
);

AND2x2_ASAP7_75t_L g13297 ( 
.A(n_12695),
.B(n_13124),
.Y(n_13297)
);

NAND2xp5_ASAP7_75t_L g13298 ( 
.A(n_12875),
.B(n_12382),
.Y(n_13298)
);

NAND2xp5_ASAP7_75t_L g13299 ( 
.A(n_12875),
.B(n_12387),
.Y(n_13299)
);

INVx2_ASAP7_75t_L g13300 ( 
.A(n_12900),
.Y(n_13300)
);

INVx2_ASAP7_75t_L g13301 ( 
.A(n_12747),
.Y(n_13301)
);

NAND2xp5_ASAP7_75t_L g13302 ( 
.A(n_13200),
.B(n_12390),
.Y(n_13302)
);

NOR2xp33_ASAP7_75t_L g13303 ( 
.A(n_13167),
.B(n_12603),
.Y(n_13303)
);

AND2x2_ASAP7_75t_L g13304 ( 
.A(n_13135),
.B(n_12397),
.Y(n_13304)
);

INVx1_ASAP7_75t_L g13305 ( 
.A(n_12843),
.Y(n_13305)
);

INVx1_ASAP7_75t_L g13306 ( 
.A(n_12835),
.Y(n_13306)
);

AND2x2_ASAP7_75t_L g13307 ( 
.A(n_12763),
.B(n_13138),
.Y(n_13307)
);

INVx2_ASAP7_75t_L g13308 ( 
.A(n_13114),
.Y(n_13308)
);

INVx1_ASAP7_75t_L g13309 ( 
.A(n_12847),
.Y(n_13309)
);

INVx1_ASAP7_75t_L g13310 ( 
.A(n_12897),
.Y(n_13310)
);

AND2x2_ASAP7_75t_L g13311 ( 
.A(n_13140),
.B(n_12402),
.Y(n_13311)
);

NAND2xp5_ASAP7_75t_L g13312 ( 
.A(n_13200),
.B(n_12412),
.Y(n_13312)
);

AND2x2_ASAP7_75t_L g13313 ( 
.A(n_12734),
.B(n_12414),
.Y(n_13313)
);

NAND2xp5_ASAP7_75t_L g13314 ( 
.A(n_13205),
.B(n_13027),
.Y(n_13314)
);

OR2x2_ASAP7_75t_L g13315 ( 
.A(n_12742),
.B(n_12618),
.Y(n_13315)
);

AND2x2_ASAP7_75t_L g13316 ( 
.A(n_12808),
.B(n_12416),
.Y(n_13316)
);

OR2x2_ASAP7_75t_L g13317 ( 
.A(n_12725),
.B(n_12537),
.Y(n_13317)
);

NAND2xp5_ASAP7_75t_L g13318 ( 
.A(n_13205),
.B(n_12420),
.Y(n_13318)
);

INVx1_ASAP7_75t_L g13319 ( 
.A(n_12736),
.Y(n_13319)
);

AND2x2_ASAP7_75t_L g13320 ( 
.A(n_12733),
.B(n_12424),
.Y(n_13320)
);

OR2x2_ASAP7_75t_L g13321 ( 
.A(n_12662),
.B(n_12427),
.Y(n_13321)
);

AND2x2_ASAP7_75t_L g13322 ( 
.A(n_12801),
.B(n_12433),
.Y(n_13322)
);

HB1xp67_ASAP7_75t_L g13323 ( 
.A(n_13070),
.Y(n_13323)
);

INVx1_ASAP7_75t_L g13324 ( 
.A(n_12818),
.Y(n_13324)
);

AND2x2_ASAP7_75t_L g13325 ( 
.A(n_13144),
.B(n_12435),
.Y(n_13325)
);

INVx1_ASAP7_75t_L g13326 ( 
.A(n_12829),
.Y(n_13326)
);

AND2x4_ASAP7_75t_L g13327 ( 
.A(n_12748),
.B(n_12439),
.Y(n_13327)
);

INVx1_ASAP7_75t_L g13328 ( 
.A(n_13147),
.Y(n_13328)
);

AND2x2_ASAP7_75t_L g13329 ( 
.A(n_13000),
.B(n_12444),
.Y(n_13329)
);

INVx1_ASAP7_75t_L g13330 ( 
.A(n_13074),
.Y(n_13330)
);

INVx1_ASAP7_75t_L g13331 ( 
.A(n_13093),
.Y(n_13331)
);

AND2x4_ASAP7_75t_SL g13332 ( 
.A(n_12664),
.B(n_12448),
.Y(n_13332)
);

HB1xp67_ASAP7_75t_L g13333 ( 
.A(n_13070),
.Y(n_13333)
);

AND2x2_ASAP7_75t_L g13334 ( 
.A(n_13018),
.B(n_12451),
.Y(n_13334)
);

AND2x4_ASAP7_75t_L g13335 ( 
.A(n_12810),
.B(n_12458),
.Y(n_13335)
);

INVx1_ASAP7_75t_SL g13336 ( 
.A(n_12909),
.Y(n_13336)
);

INVx2_ASAP7_75t_L g13337 ( 
.A(n_13114),
.Y(n_13337)
);

NAND2xp5_ASAP7_75t_L g13338 ( 
.A(n_13037),
.B(n_12459),
.Y(n_13338)
);

AND2x4_ASAP7_75t_L g13339 ( 
.A(n_12851),
.B(n_12462),
.Y(n_13339)
);

INVx1_ASAP7_75t_L g13340 ( 
.A(n_13099),
.Y(n_13340)
);

NOR2xp67_ASAP7_75t_L g13341 ( 
.A(n_12775),
.B(n_12704),
.Y(n_13341)
);

OR2x2_ASAP7_75t_L g13342 ( 
.A(n_12968),
.B(n_12466),
.Y(n_13342)
);

INVx2_ASAP7_75t_L g13343 ( 
.A(n_13114),
.Y(n_13343)
);

AND2x4_ASAP7_75t_L g13344 ( 
.A(n_12851),
.B(n_12468),
.Y(n_13344)
);

OR2x2_ASAP7_75t_L g13345 ( 
.A(n_12768),
.B(n_12475),
.Y(n_13345)
);

INVxp67_ASAP7_75t_SL g13346 ( 
.A(n_12692),
.Y(n_13346)
);

AND2x2_ASAP7_75t_L g13347 ( 
.A(n_12761),
.B(n_12479),
.Y(n_13347)
);

OR2x2_ASAP7_75t_L g13348 ( 
.A(n_12737),
.B(n_12481),
.Y(n_13348)
);

INVxp67_ASAP7_75t_L g13349 ( 
.A(n_12945),
.Y(n_13349)
);

NAND2xp5_ASAP7_75t_SL g13350 ( 
.A(n_13172),
.B(n_12426),
.Y(n_13350)
);

INVx1_ASAP7_75t_L g13351 ( 
.A(n_12901),
.Y(n_13351)
);

NAND2xp5_ASAP7_75t_L g13352 ( 
.A(n_12877),
.B(n_12483),
.Y(n_13352)
);

NOR2xp33_ASAP7_75t_SL g13353 ( 
.A(n_12660),
.B(n_12887),
.Y(n_13353)
);

AND2x2_ASAP7_75t_L g13354 ( 
.A(n_12904),
.B(n_12484),
.Y(n_13354)
);

AND2x2_ASAP7_75t_L g13355 ( 
.A(n_12854),
.B(n_12485),
.Y(n_13355)
);

AND2x2_ASAP7_75t_L g13356 ( 
.A(n_12707),
.B(n_12487),
.Y(n_13356)
);

AND2x2_ASAP7_75t_L g13357 ( 
.A(n_12842),
.B(n_12492),
.Y(n_13357)
);

NAND2xp5_ASAP7_75t_L g13358 ( 
.A(n_12877),
.B(n_13041),
.Y(n_13358)
);

AND2x2_ASAP7_75t_L g13359 ( 
.A(n_12850),
.B(n_12493),
.Y(n_13359)
);

OR2x2_ASAP7_75t_L g13360 ( 
.A(n_12750),
.B(n_12494),
.Y(n_13360)
);

INVxp67_ASAP7_75t_SL g13361 ( 
.A(n_12696),
.Y(n_13361)
);

INVx1_ASAP7_75t_L g13362 ( 
.A(n_13120),
.Y(n_13362)
);

NAND2xp5_ASAP7_75t_L g13363 ( 
.A(n_12909),
.B(n_12505),
.Y(n_13363)
);

INVx1_ASAP7_75t_L g13364 ( 
.A(n_13120),
.Y(n_13364)
);

INVx2_ASAP7_75t_L g13365 ( 
.A(n_12960),
.Y(n_13365)
);

INVx2_ASAP7_75t_L g13366 ( 
.A(n_12960),
.Y(n_13366)
);

NAND2xp5_ASAP7_75t_L g13367 ( 
.A(n_13203),
.B(n_12506),
.Y(n_13367)
);

NAND2x1p5_ASAP7_75t_L g13368 ( 
.A(n_13179),
.B(n_12269),
.Y(n_13368)
);

INVx2_ASAP7_75t_L g13369 ( 
.A(n_13225),
.Y(n_13369)
);

HB1xp67_ASAP7_75t_L g13370 ( 
.A(n_12892),
.Y(n_13370)
);

AND2x4_ASAP7_75t_L g13371 ( 
.A(n_12929),
.B(n_12507),
.Y(n_13371)
);

INVx1_ASAP7_75t_L g13372 ( 
.A(n_13134),
.Y(n_13372)
);

INVx1_ASAP7_75t_L g13373 ( 
.A(n_13134),
.Y(n_13373)
);

OR2x2_ASAP7_75t_L g13374 ( 
.A(n_12714),
.B(n_12511),
.Y(n_13374)
);

AND2x4_ASAP7_75t_SL g13375 ( 
.A(n_13119),
.B(n_12513),
.Y(n_13375)
);

AND2x2_ASAP7_75t_L g13376 ( 
.A(n_12670),
.B(n_12515),
.Y(n_13376)
);

INVx1_ASAP7_75t_L g13377 ( 
.A(n_13153),
.Y(n_13377)
);

INVx1_ASAP7_75t_L g13378 ( 
.A(n_13153),
.Y(n_13378)
);

HB1xp67_ASAP7_75t_L g13379 ( 
.A(n_12892),
.Y(n_13379)
);

HB1xp67_ASAP7_75t_L g13380 ( 
.A(n_12710),
.Y(n_13380)
);

AND2x2_ASAP7_75t_L g13381 ( 
.A(n_13111),
.B(n_12534),
.Y(n_13381)
);

OR2x2_ASAP7_75t_L g13382 ( 
.A(n_12777),
.B(n_12553),
.Y(n_13382)
);

INVx1_ASAP7_75t_L g13383 ( 
.A(n_13195),
.Y(n_13383)
);

AND2x2_ASAP7_75t_L g13384 ( 
.A(n_13113),
.B(n_12556),
.Y(n_13384)
);

OAI21xp5_ASAP7_75t_SL g13385 ( 
.A1(n_13005),
.A2(n_12389),
.B(n_12465),
.Y(n_13385)
);

HB1xp67_ASAP7_75t_L g13386 ( 
.A(n_13039),
.Y(n_13386)
);

AND2x2_ASAP7_75t_L g13387 ( 
.A(n_12911),
.B(n_12562),
.Y(n_13387)
);

INVx1_ASAP7_75t_L g13388 ( 
.A(n_13195),
.Y(n_13388)
);

NAND2xp5_ASAP7_75t_L g13389 ( 
.A(n_13021),
.B(n_12565),
.Y(n_13389)
);

INVx1_ASAP7_75t_L g13390 ( 
.A(n_12791),
.Y(n_13390)
);

INVx1_ASAP7_75t_L g13391 ( 
.A(n_12782),
.Y(n_13391)
);

AND2x2_ASAP7_75t_L g13392 ( 
.A(n_13095),
.B(n_12582),
.Y(n_13392)
);

INVx2_ASAP7_75t_L g13393 ( 
.A(n_13225),
.Y(n_13393)
);

INVx1_ASAP7_75t_L g13394 ( 
.A(n_13004),
.Y(n_13394)
);

NAND2xp5_ASAP7_75t_L g13395 ( 
.A(n_13199),
.B(n_12583),
.Y(n_13395)
);

AND2x2_ASAP7_75t_L g13396 ( 
.A(n_13133),
.B(n_12586),
.Y(n_13396)
);

OR2x2_ASAP7_75t_L g13397 ( 
.A(n_12789),
.B(n_12591),
.Y(n_13397)
);

OR2x2_ASAP7_75t_L g13398 ( 
.A(n_13049),
.B(n_13085),
.Y(n_13398)
);

OR2x2_ASAP7_75t_L g13399 ( 
.A(n_13121),
.B(n_12599),
.Y(n_13399)
);

OR2x2_ASAP7_75t_L g13400 ( 
.A(n_13130),
.B(n_12601),
.Y(n_13400)
);

AND2x2_ASAP7_75t_L g13401 ( 
.A(n_13139),
.B(n_12605),
.Y(n_13401)
);

AND2x2_ASAP7_75t_L g13402 ( 
.A(n_13148),
.B(n_12610),
.Y(n_13402)
);

AND2x2_ASAP7_75t_L g13403 ( 
.A(n_12820),
.B(n_12612),
.Y(n_13403)
);

INVx2_ASAP7_75t_L g13404 ( 
.A(n_13090),
.Y(n_13404)
);

AND2x2_ASAP7_75t_L g13405 ( 
.A(n_13031),
.B(n_12623),
.Y(n_13405)
);

HB1xp67_ASAP7_75t_L g13406 ( 
.A(n_13090),
.Y(n_13406)
);

AND2x2_ASAP7_75t_L g13407 ( 
.A(n_12841),
.B(n_12626),
.Y(n_13407)
);

AND2x2_ASAP7_75t_L g13408 ( 
.A(n_12830),
.B(n_12641),
.Y(n_13408)
);

AND2x2_ASAP7_75t_L g13409 ( 
.A(n_12760),
.B(n_12642),
.Y(n_13409)
);

NAND2xp5_ASAP7_75t_L g13410 ( 
.A(n_13199),
.B(n_12647),
.Y(n_13410)
);

NOR2xp67_ASAP7_75t_L g13411 ( 
.A(n_12935),
.B(n_12648),
.Y(n_13411)
);

OR2x2_ASAP7_75t_L g13412 ( 
.A(n_12781),
.B(n_12650),
.Y(n_13412)
);

INVx1_ASAP7_75t_L g13413 ( 
.A(n_13155),
.Y(n_13413)
);

NAND2xp5_ASAP7_75t_L g13414 ( 
.A(n_13185),
.B(n_12652),
.Y(n_13414)
);

OR2x2_ASAP7_75t_L g13415 ( 
.A(n_12792),
.B(n_12653),
.Y(n_13415)
);

OR2x2_ASAP7_75t_L g13416 ( 
.A(n_13197),
.B(n_11830),
.Y(n_13416)
);

INVx1_ASAP7_75t_L g13417 ( 
.A(n_12953),
.Y(n_13417)
);

NAND2xp5_ASAP7_75t_L g13418 ( 
.A(n_13172),
.B(n_11836),
.Y(n_13418)
);

AND2x2_ASAP7_75t_L g13419 ( 
.A(n_12726),
.B(n_12580),
.Y(n_13419)
);

INVx1_ASAP7_75t_L g13420 ( 
.A(n_13224),
.Y(n_13420)
);

INVx1_ASAP7_75t_L g13421 ( 
.A(n_13217),
.Y(n_13421)
);

INVx1_ASAP7_75t_L g13422 ( 
.A(n_12837),
.Y(n_13422)
);

AND2x2_ASAP7_75t_L g13423 ( 
.A(n_13123),
.B(n_11999),
.Y(n_13423)
);

INVx4_ASAP7_75t_L g13424 ( 
.A(n_13038),
.Y(n_13424)
);

INVx2_ASAP7_75t_L g13425 ( 
.A(n_12787),
.Y(n_13425)
);

INVx1_ASAP7_75t_L g13426 ( 
.A(n_12709),
.Y(n_13426)
);

INVx2_ASAP7_75t_L g13427 ( 
.A(n_12787),
.Y(n_13427)
);

OR2x2_ASAP7_75t_L g13428 ( 
.A(n_12915),
.B(n_11840),
.Y(n_13428)
);

HB1xp67_ASAP7_75t_L g13429 ( 
.A(n_12756),
.Y(n_13429)
);

OAI21xp5_ASAP7_75t_SL g13430 ( 
.A1(n_13154),
.A2(n_12132),
.B(n_12128),
.Y(n_13430)
);

INVx1_ASAP7_75t_L g13431 ( 
.A(n_12719),
.Y(n_13431)
);

NAND2xp5_ASAP7_75t_L g13432 ( 
.A(n_12812),
.B(n_12157),
.Y(n_13432)
);

HB1xp67_ASAP7_75t_L g13433 ( 
.A(n_12857),
.Y(n_13433)
);

AND2x2_ASAP7_75t_L g13434 ( 
.A(n_12952),
.B(n_10216),
.Y(n_13434)
);

AND2x2_ASAP7_75t_L g13435 ( 
.A(n_13025),
.B(n_10222),
.Y(n_13435)
);

INVx4_ASAP7_75t_L g13436 ( 
.A(n_13038),
.Y(n_13436)
);

INVx2_ASAP7_75t_L g13437 ( 
.A(n_12788),
.Y(n_13437)
);

INVx1_ASAP7_75t_L g13438 ( 
.A(n_13125),
.Y(n_13438)
);

INVx1_ASAP7_75t_L g13439 ( 
.A(n_13127),
.Y(n_13439)
);

AND2x2_ASAP7_75t_L g13440 ( 
.A(n_12741),
.B(n_10225),
.Y(n_13440)
);

AND2x2_ASAP7_75t_L g13441 ( 
.A(n_12745),
.B(n_10227),
.Y(n_13441)
);

AND2x2_ASAP7_75t_L g13442 ( 
.A(n_12944),
.B(n_10228),
.Y(n_13442)
);

OR2x2_ASAP7_75t_L g13443 ( 
.A(n_12667),
.B(n_11861),
.Y(n_13443)
);

AND2x2_ASAP7_75t_L g13444 ( 
.A(n_12969),
.B(n_10230),
.Y(n_13444)
);

OAI21xp5_ASAP7_75t_L g13445 ( 
.A1(n_12918),
.A2(n_11789),
.B(n_11783),
.Y(n_13445)
);

INVx1_ASAP7_75t_L g13446 ( 
.A(n_12923),
.Y(n_13446)
);

OR2x2_ASAP7_75t_L g13447 ( 
.A(n_12749),
.B(n_12895),
.Y(n_13447)
);

AND2x4_ASAP7_75t_L g13448 ( 
.A(n_12788),
.B(n_12359),
.Y(n_13448)
);

NAND2xp5_ASAP7_75t_L g13449 ( 
.A(n_12813),
.B(n_11708),
.Y(n_13449)
);

NOR2xp67_ASAP7_75t_SL g13450 ( 
.A(n_12977),
.B(n_4175),
.Y(n_13450)
);

NAND2xp5_ASAP7_75t_L g13451 ( 
.A(n_13182),
.B(n_11708),
.Y(n_13451)
);

AND2x2_ASAP7_75t_L g13452 ( 
.A(n_12974),
.B(n_10233),
.Y(n_13452)
);

OR2x2_ASAP7_75t_L g13453 ( 
.A(n_13081),
.B(n_11873),
.Y(n_13453)
);

NAND2xp5_ASAP7_75t_L g13454 ( 
.A(n_12890),
.B(n_11877),
.Y(n_13454)
);

INVx2_ASAP7_75t_L g13455 ( 
.A(n_12666),
.Y(n_13455)
);

NAND2xp5_ASAP7_75t_L g13456 ( 
.A(n_12890),
.B(n_11850),
.Y(n_13456)
);

INVx2_ASAP7_75t_L g13457 ( 
.A(n_12910),
.Y(n_13457)
);

AND2x2_ASAP7_75t_L g13458 ( 
.A(n_12868),
.B(n_10236),
.Y(n_13458)
);

AND2x4_ASAP7_75t_L g13459 ( 
.A(n_12657),
.B(n_12723),
.Y(n_13459)
);

INVx1_ASAP7_75t_L g13460 ( 
.A(n_12934),
.Y(n_13460)
);

AND2x2_ASAP7_75t_L g13461 ( 
.A(n_13089),
.B(n_10238),
.Y(n_13461)
);

INVx1_ASAP7_75t_L g13462 ( 
.A(n_13035),
.Y(n_13462)
);

AND2x2_ASAP7_75t_L g13463 ( 
.A(n_12937),
.B(n_10239),
.Y(n_13463)
);

INVx1_ASAP7_75t_L g13464 ( 
.A(n_13051),
.Y(n_13464)
);

NOR2x1_ASAP7_75t_L g13465 ( 
.A(n_12834),
.B(n_12374),
.Y(n_13465)
);

AND2x4_ASAP7_75t_L g13466 ( 
.A(n_12723),
.B(n_12703),
.Y(n_13466)
);

INVx1_ASAP7_75t_L g13467 ( 
.A(n_13058),
.Y(n_13467)
);

INVx1_ASAP7_75t_L g13468 ( 
.A(n_13063),
.Y(n_13468)
);

INVx2_ASAP7_75t_L g13469 ( 
.A(n_13016),
.Y(n_13469)
);

INVx1_ASAP7_75t_L g13470 ( 
.A(n_12955),
.Y(n_13470)
);

INVx2_ASAP7_75t_L g13471 ( 
.A(n_12963),
.Y(n_13471)
);

AND2x4_ASAP7_75t_L g13472 ( 
.A(n_12706),
.B(n_11851),
.Y(n_13472)
);

NAND2xp5_ASAP7_75t_L g13473 ( 
.A(n_12908),
.B(n_11850),
.Y(n_13473)
);

AND2x4_ASAP7_75t_L g13474 ( 
.A(n_12708),
.B(n_11829),
.Y(n_13474)
);

OR2x2_ASAP7_75t_L g13475 ( 
.A(n_13015),
.B(n_11864),
.Y(n_13475)
);

AND2x2_ASAP7_75t_L g13476 ( 
.A(n_12938),
.B(n_10240),
.Y(n_13476)
);

INVx1_ASAP7_75t_L g13477 ( 
.A(n_12959),
.Y(n_13477)
);

AND2x2_ASAP7_75t_L g13478 ( 
.A(n_12797),
.B(n_12884),
.Y(n_13478)
);

INVx2_ASAP7_75t_L g13479 ( 
.A(n_12963),
.Y(n_13479)
);

NAND3xp33_ASAP7_75t_L g13480 ( 
.A(n_12688),
.B(n_11904),
.C(n_12262),
.Y(n_13480)
);

INVx2_ASAP7_75t_L g13481 ( 
.A(n_12994),
.Y(n_13481)
);

INVx1_ASAP7_75t_L g13482 ( 
.A(n_12966),
.Y(n_13482)
);

BUFx2_ASAP7_75t_SL g13483 ( 
.A(n_12700),
.Y(n_13483)
);

HB1xp67_ASAP7_75t_L g13484 ( 
.A(n_12994),
.Y(n_13484)
);

OR2x6_ASAP7_75t_L g13485 ( 
.A(n_12945),
.B(n_8545),
.Y(n_13485)
);

INVx2_ASAP7_75t_L g13486 ( 
.A(n_12826),
.Y(n_13486)
);

AND2x4_ASAP7_75t_L g13487 ( 
.A(n_13003),
.B(n_4226),
.Y(n_13487)
);

NAND2xp5_ASAP7_75t_L g13488 ( 
.A(n_12908),
.B(n_11864),
.Y(n_13488)
);

INVx1_ASAP7_75t_L g13489 ( 
.A(n_12976),
.Y(n_13489)
);

INVx1_ASAP7_75t_L g13490 ( 
.A(n_12981),
.Y(n_13490)
);

AND2x2_ASAP7_75t_L g13491 ( 
.A(n_12906),
.B(n_10246),
.Y(n_13491)
);

INVx1_ASAP7_75t_L g13492 ( 
.A(n_12983),
.Y(n_13492)
);

AND2x2_ASAP7_75t_L g13493 ( 
.A(n_12769),
.B(n_10247),
.Y(n_13493)
);

HB1xp67_ASAP7_75t_L g13494 ( 
.A(n_12862),
.Y(n_13494)
);

OAI22xp5_ASAP7_75t_L g13495 ( 
.A1(n_13053),
.A2(n_12401),
.B1(n_12328),
.B2(n_12398),
.Y(n_13495)
);

AND2x2_ASAP7_75t_L g13496 ( 
.A(n_12772),
.B(n_10259),
.Y(n_13496)
);

INVx2_ASAP7_75t_L g13497 ( 
.A(n_12826),
.Y(n_13497)
);

NAND2xp5_ASAP7_75t_L g13498 ( 
.A(n_12928),
.B(n_11866),
.Y(n_13498)
);

NAND2xp5_ASAP7_75t_L g13499 ( 
.A(n_13034),
.B(n_11866),
.Y(n_13499)
);

INVx1_ASAP7_75t_L g13500 ( 
.A(n_12984),
.Y(n_13500)
);

INVx1_ASAP7_75t_L g13501 ( 
.A(n_12859),
.Y(n_13501)
);

AND2x4_ASAP7_75t_L g13502 ( 
.A(n_12712),
.B(n_11802),
.Y(n_13502)
);

AND2x2_ASAP7_75t_L g13503 ( 
.A(n_12885),
.B(n_10260),
.Y(n_13503)
);

AND2x2_ASAP7_75t_L g13504 ( 
.A(n_12665),
.B(n_10266),
.Y(n_13504)
);

AND2x4_ASAP7_75t_SL g13505 ( 
.A(n_12694),
.B(n_12701),
.Y(n_13505)
);

INVx1_ASAP7_75t_L g13506 ( 
.A(n_13214),
.Y(n_13506)
);

HB1xp67_ASAP7_75t_L g13507 ( 
.A(n_12728),
.Y(n_13507)
);

OR2x2_ASAP7_75t_L g13508 ( 
.A(n_12807),
.B(n_11895),
.Y(n_13508)
);

AND2x2_ASAP7_75t_L g13509 ( 
.A(n_13087),
.B(n_10267),
.Y(n_13509)
);

INVx1_ASAP7_75t_L g13510 ( 
.A(n_12764),
.Y(n_13510)
);

INVx2_ASAP7_75t_L g13511 ( 
.A(n_12907),
.Y(n_13511)
);

INVxp67_ASAP7_75t_L g13512 ( 
.A(n_12676),
.Y(n_13512)
);

INVxp67_ASAP7_75t_SL g13513 ( 
.A(n_12685),
.Y(n_13513)
);

NAND2xp5_ASAP7_75t_L g13514 ( 
.A(n_13145),
.B(n_12205),
.Y(n_13514)
);

INVx1_ASAP7_75t_L g13515 ( 
.A(n_12916),
.Y(n_13515)
);

AND2x2_ASAP7_75t_L g13516 ( 
.A(n_13069),
.B(n_10269),
.Y(n_13516)
);

INVx1_ASAP7_75t_L g13517 ( 
.A(n_12920),
.Y(n_13517)
);

AND2x2_ASAP7_75t_L g13518 ( 
.A(n_12672),
.B(n_10274),
.Y(n_13518)
);

INVx1_ASAP7_75t_L g13519 ( 
.A(n_13029),
.Y(n_13519)
);

INVx1_ASAP7_75t_L g13520 ( 
.A(n_13028),
.Y(n_13520)
);

INVx1_ASAP7_75t_L g13521 ( 
.A(n_12674),
.Y(n_13521)
);

NAND2xp5_ASAP7_75t_L g13522 ( 
.A(n_13117),
.B(n_11805),
.Y(n_13522)
);

NAND2xp5_ASAP7_75t_L g13523 ( 
.A(n_13117),
.B(n_12597),
.Y(n_13523)
);

AND2x2_ASAP7_75t_L g13524 ( 
.A(n_12824),
.B(n_10277),
.Y(n_13524)
);

INVx2_ASAP7_75t_L g13525 ( 
.A(n_12799),
.Y(n_13525)
);

AND2x2_ASAP7_75t_L g13526 ( 
.A(n_12867),
.B(n_10279),
.Y(n_13526)
);

BUFx2_ASAP7_75t_L g13527 ( 
.A(n_13142),
.Y(n_13527)
);

INVx1_ASAP7_75t_L g13528 ( 
.A(n_12730),
.Y(n_13528)
);

INVx1_ASAP7_75t_L g13529 ( 
.A(n_12773),
.Y(n_13529)
);

INVx1_ASAP7_75t_L g13530 ( 
.A(n_12774),
.Y(n_13530)
);

NAND2x1p5_ASAP7_75t_L g13531 ( 
.A(n_12932),
.B(n_7987),
.Y(n_13531)
);

INVx3_ASAP7_75t_L g13532 ( 
.A(n_12932),
.Y(n_13532)
);

AND2x2_ASAP7_75t_L g13533 ( 
.A(n_12941),
.B(n_10283),
.Y(n_13533)
);

INVx1_ASAP7_75t_L g13534 ( 
.A(n_12778),
.Y(n_13534)
);

INVx1_ASAP7_75t_L g13535 ( 
.A(n_12785),
.Y(n_13535)
);

AND2x2_ASAP7_75t_L g13536 ( 
.A(n_12831),
.B(n_10288),
.Y(n_13536)
);

NAND2xp5_ASAP7_75t_L g13537 ( 
.A(n_12970),
.B(n_12606),
.Y(n_13537)
);

AND2x2_ASAP7_75t_L g13538 ( 
.A(n_12845),
.B(n_10290),
.Y(n_13538)
);

NOR2x1_ASAP7_75t_L g13539 ( 
.A(n_12799),
.B(n_11809),
.Y(n_13539)
);

INVxp67_ASAP7_75t_L g13540 ( 
.A(n_12767),
.Y(n_13540)
);

OR2x2_ASAP7_75t_L g13541 ( 
.A(n_12766),
.B(n_10295),
.Y(n_13541)
);

NAND2xp5_ASAP7_75t_L g13542 ( 
.A(n_13024),
.B(n_12197),
.Y(n_13542)
);

NAND2xp5_ASAP7_75t_L g13543 ( 
.A(n_13024),
.B(n_12577),
.Y(n_13543)
);

AND2x2_ASAP7_75t_L g13544 ( 
.A(n_12927),
.B(n_10300),
.Y(n_13544)
);

NAND2xp5_ASAP7_75t_L g13545 ( 
.A(n_13012),
.B(n_12408),
.Y(n_13545)
);

AND2x2_ASAP7_75t_L g13546 ( 
.A(n_13174),
.B(n_10303),
.Y(n_13546)
);

INVx2_ASAP7_75t_L g13547 ( 
.A(n_12729),
.Y(n_13547)
);

INVx2_ASAP7_75t_L g13548 ( 
.A(n_12729),
.Y(n_13548)
);

INVx1_ASAP7_75t_L g13549 ( 
.A(n_12800),
.Y(n_13549)
);

AND2x2_ASAP7_75t_L g13550 ( 
.A(n_13020),
.B(n_10304),
.Y(n_13550)
);

INVx1_ASAP7_75t_L g13551 ( 
.A(n_12804),
.Y(n_13551)
);

AND2x2_ASAP7_75t_L g13552 ( 
.A(n_12943),
.B(n_10306),
.Y(n_13552)
);

AND2x2_ASAP7_75t_L g13553 ( 
.A(n_12814),
.B(n_10307),
.Y(n_13553)
);

AND2x2_ASAP7_75t_L g13554 ( 
.A(n_12919),
.B(n_10310),
.Y(n_13554)
);

NAND2x1_ASAP7_75t_SL g13555 ( 
.A(n_12980),
.B(n_10121),
.Y(n_13555)
);

AND2x2_ASAP7_75t_L g13556 ( 
.A(n_12913),
.B(n_10312),
.Y(n_13556)
);

INVx1_ASAP7_75t_L g13557 ( 
.A(n_12815),
.Y(n_13557)
);

INVx1_ASAP7_75t_L g13558 ( 
.A(n_12816),
.Y(n_13558)
);

AND2x2_ASAP7_75t_L g13559 ( 
.A(n_13013),
.B(n_10315),
.Y(n_13559)
);

AND2x2_ASAP7_75t_L g13560 ( 
.A(n_13062),
.B(n_10328),
.Y(n_13560)
);

OR2x6_ASAP7_75t_L g13561 ( 
.A(n_12739),
.B(n_8545),
.Y(n_13561)
);

INVx2_ASAP7_75t_SL g13562 ( 
.A(n_12661),
.Y(n_13562)
);

OAI32xp33_ASAP7_75t_L g13563 ( 
.A1(n_13143),
.A2(n_11926),
.A3(n_11930),
.B1(n_10158),
.B2(n_10171),
.Y(n_13563)
);

OR2x2_ASAP7_75t_L g13564 ( 
.A(n_13226),
.B(n_10334),
.Y(n_13564)
);

INVxp67_ASAP7_75t_SL g13565 ( 
.A(n_12780),
.Y(n_13565)
);

INVx1_ASAP7_75t_L g13566 ( 
.A(n_12819),
.Y(n_13566)
);

AND2x2_ASAP7_75t_L g13567 ( 
.A(n_13064),
.B(n_10335),
.Y(n_13567)
);

NAND2xp5_ASAP7_75t_L g13568 ( 
.A(n_13065),
.B(n_11926),
.Y(n_13568)
);

INVx1_ASAP7_75t_L g13569 ( 
.A(n_12823),
.Y(n_13569)
);

AND2x2_ASAP7_75t_L g13570 ( 
.A(n_13066),
.B(n_10345),
.Y(n_13570)
);

AND2x2_ASAP7_75t_L g13571 ( 
.A(n_13073),
.B(n_10347),
.Y(n_13571)
);

HB1xp67_ASAP7_75t_L g13572 ( 
.A(n_12744),
.Y(n_13572)
);

INVx1_ASAP7_75t_L g13573 ( 
.A(n_12825),
.Y(n_13573)
);

AND2x2_ASAP7_75t_L g13574 ( 
.A(n_13079),
.B(n_10348),
.Y(n_13574)
);

INVx1_ASAP7_75t_L g13575 ( 
.A(n_12832),
.Y(n_13575)
);

INVx2_ASAP7_75t_SL g13576 ( 
.A(n_12755),
.Y(n_13576)
);

INVx4_ASAP7_75t_L g13577 ( 
.A(n_12698),
.Y(n_13577)
);

INVx1_ASAP7_75t_L g13578 ( 
.A(n_12865),
.Y(n_13578)
);

INVx1_ASAP7_75t_L g13579 ( 
.A(n_12727),
.Y(n_13579)
);

INVx1_ASAP7_75t_L g13580 ( 
.A(n_13204),
.Y(n_13580)
);

AND2x2_ASAP7_75t_L g13581 ( 
.A(n_13084),
.B(n_10349),
.Y(n_13581)
);

OR2x2_ASAP7_75t_L g13582 ( 
.A(n_13177),
.B(n_10351),
.Y(n_13582)
);

INVx1_ASAP7_75t_L g13583 ( 
.A(n_13204),
.Y(n_13583)
);

NAND2x1p5_ASAP7_75t_L g13584 ( 
.A(n_12698),
.B(n_7996),
.Y(n_13584)
);

INVx2_ASAP7_75t_L g13585 ( 
.A(n_12746),
.Y(n_13585)
);

AND2x2_ASAP7_75t_L g13586 ( 
.A(n_13092),
.B(n_13108),
.Y(n_13586)
);

OR2x2_ASAP7_75t_L g13587 ( 
.A(n_12878),
.B(n_13047),
.Y(n_13587)
);

INVx1_ASAP7_75t_L g13588 ( 
.A(n_13011),
.Y(n_13588)
);

NAND2xp5_ASAP7_75t_L g13589 ( 
.A(n_13116),
.B(n_11930),
.Y(n_13589)
);

AND2x4_ASAP7_75t_L g13590 ( 
.A(n_12872),
.B(n_10355),
.Y(n_13590)
);

NAND2x1p5_ASAP7_75t_L g13591 ( 
.A(n_12746),
.B(n_7996),
.Y(n_13591)
);

INVx1_ASAP7_75t_L g13592 ( 
.A(n_13023),
.Y(n_13592)
);

OR2x2_ASAP7_75t_L g13593 ( 
.A(n_12939),
.B(n_10356),
.Y(n_13593)
);

NAND2xp5_ASAP7_75t_L g13594 ( 
.A(n_13118),
.B(n_12541),
.Y(n_13594)
);

AND2x4_ASAP7_75t_L g13595 ( 
.A(n_12827),
.B(n_7996),
.Y(n_13595)
);

NAND2xp5_ASAP7_75t_L g13596 ( 
.A(n_13126),
.B(n_9914),
.Y(n_13596)
);

NOR2xp33_ASAP7_75t_L g13597 ( 
.A(n_12849),
.B(n_7843),
.Y(n_13597)
);

NOR2xp33_ASAP7_75t_SL g13598 ( 
.A(n_13193),
.B(n_12752),
.Y(n_13598)
);

OR2x2_ASAP7_75t_L g13599 ( 
.A(n_12821),
.B(n_10361),
.Y(n_13599)
);

INVx1_ASAP7_75t_L g13600 ( 
.A(n_13040),
.Y(n_13600)
);

OR2x2_ASAP7_75t_L g13601 ( 
.A(n_12822),
.B(n_10364),
.Y(n_13601)
);

NAND2xp5_ASAP7_75t_L g13602 ( 
.A(n_13131),
.B(n_9914),
.Y(n_13602)
);

INVx2_ASAP7_75t_L g13603 ( 
.A(n_12980),
.Y(n_13603)
);

AND2x2_ASAP7_75t_L g13604 ( 
.A(n_13137),
.B(n_10372),
.Y(n_13604)
);

AND2x2_ASAP7_75t_L g13605 ( 
.A(n_12996),
.B(n_10373),
.Y(n_13605)
);

INVx2_ASAP7_75t_L g13606 ( 
.A(n_12876),
.Y(n_13606)
);

AND2x2_ASAP7_75t_L g13607 ( 
.A(n_12997),
.B(n_10374),
.Y(n_13607)
);

AND2x2_ASAP7_75t_L g13608 ( 
.A(n_12828),
.B(n_13009),
.Y(n_13608)
);

INVx2_ASAP7_75t_L g13609 ( 
.A(n_12881),
.Y(n_13609)
);

AND2x2_ASAP7_75t_L g13610 ( 
.A(n_12754),
.B(n_10379),
.Y(n_13610)
);

AND2x2_ASAP7_75t_L g13611 ( 
.A(n_12962),
.B(n_10389),
.Y(n_13611)
);

OR2x2_ASAP7_75t_L g13612 ( 
.A(n_12833),
.B(n_10397),
.Y(n_13612)
);

NAND2xp5_ASAP7_75t_L g13613 ( 
.A(n_12899),
.B(n_9916),
.Y(n_13613)
);

AND2x2_ASAP7_75t_L g13614 ( 
.A(n_12873),
.B(n_10399),
.Y(n_13614)
);

INVx1_ASAP7_75t_L g13615 ( 
.A(n_12836),
.Y(n_13615)
);

NAND2xp5_ASAP7_75t_L g13616 ( 
.A(n_12896),
.B(n_9916),
.Y(n_13616)
);

OR2x2_ASAP7_75t_L g13617 ( 
.A(n_12940),
.B(n_10401),
.Y(n_13617)
);

AND2x2_ASAP7_75t_L g13618 ( 
.A(n_12863),
.B(n_7180),
.Y(n_13618)
);

INVx1_ASAP7_75t_L g13619 ( 
.A(n_13022),
.Y(n_13619)
);

AND2x2_ASAP7_75t_L g13620 ( 
.A(n_13036),
.B(n_7203),
.Y(n_13620)
);

NAND2xp5_ASAP7_75t_L g13621 ( 
.A(n_12950),
.B(n_9922),
.Y(n_13621)
);

AND2x4_ASAP7_75t_L g13622 ( 
.A(n_13168),
.B(n_7996),
.Y(n_13622)
);

INVx2_ASAP7_75t_L g13623 ( 
.A(n_12883),
.Y(n_13623)
);

INVx1_ASAP7_75t_L g13624 ( 
.A(n_12673),
.Y(n_13624)
);

INVx1_ASAP7_75t_L g13625 ( 
.A(n_12690),
.Y(n_13625)
);

INVx3_ASAP7_75t_L g13626 ( 
.A(n_12849),
.Y(n_13626)
);

NAND2x1p5_ASAP7_75t_L g13627 ( 
.A(n_12864),
.B(n_7859),
.Y(n_13627)
);

NAND3xp33_ASAP7_75t_L g13628 ( 
.A(n_12743),
.B(n_11721),
.C(n_11720),
.Y(n_13628)
);

NAND3xp33_ASAP7_75t_L g13629 ( 
.A(n_12677),
.B(n_11721),
.C(n_11720),
.Y(n_13629)
);

AND2x2_ASAP7_75t_L g13630 ( 
.A(n_12902),
.B(n_7291),
.Y(n_13630)
);

OR2x6_ASAP7_75t_L g13631 ( 
.A(n_12809),
.B(n_11808),
.Y(n_13631)
);

INVxp67_ASAP7_75t_L g13632 ( 
.A(n_12886),
.Y(n_13632)
);

AND2x4_ASAP7_75t_L g13633 ( 
.A(n_13170),
.B(n_12905),
.Y(n_13633)
);

AND2x2_ASAP7_75t_L g13634 ( 
.A(n_12917),
.B(n_7766),
.Y(n_13634)
);

INVx2_ASAP7_75t_SL g13635 ( 
.A(n_12942),
.Y(n_13635)
);

AND2x2_ASAP7_75t_L g13636 ( 
.A(n_12921),
.B(n_7766),
.Y(n_13636)
);

INVx1_ASAP7_75t_L g13637 ( 
.A(n_13181),
.Y(n_13637)
);

HB1xp67_ASAP7_75t_L g13638 ( 
.A(n_13043),
.Y(n_13638)
);

NAND3xp33_ASAP7_75t_L g13639 ( 
.A(n_13083),
.B(n_11723),
.C(n_9930),
.Y(n_13639)
);

AND2x2_ASAP7_75t_L g13640 ( 
.A(n_13048),
.B(n_7766),
.Y(n_13640)
);

INVx1_ASAP7_75t_L g13641 ( 
.A(n_13008),
.Y(n_13641)
);

NAND2xp5_ASAP7_75t_L g13642 ( 
.A(n_12950),
.B(n_9922),
.Y(n_13642)
);

NAND2xp5_ASAP7_75t_L g13643 ( 
.A(n_12979),
.B(n_9930),
.Y(n_13643)
);

NOR2xp33_ASAP7_75t_L g13644 ( 
.A(n_12864),
.B(n_7859),
.Y(n_13644)
);

AND2x2_ASAP7_75t_L g13645 ( 
.A(n_12947),
.B(n_7818),
.Y(n_13645)
);

INVx2_ASAP7_75t_SL g13646 ( 
.A(n_12942),
.Y(n_13646)
);

HB1xp67_ASAP7_75t_L g13647 ( 
.A(n_12866),
.Y(n_13647)
);

AND2x4_ASAP7_75t_L g13648 ( 
.A(n_12949),
.B(n_12954),
.Y(n_13648)
);

INVx1_ASAP7_75t_L g13649 ( 
.A(n_13220),
.Y(n_13649)
);

NAND2x1_ASAP7_75t_L g13650 ( 
.A(n_12786),
.B(n_10122),
.Y(n_13650)
);

AND2x2_ASAP7_75t_L g13651 ( 
.A(n_13010),
.B(n_13055),
.Y(n_13651)
);

OR2x2_ASAP7_75t_L g13652 ( 
.A(n_12951),
.B(n_12957),
.Y(n_13652)
);

INVx1_ASAP7_75t_L g13653 ( 
.A(n_12979),
.Y(n_13653)
);

INVx2_ASAP7_75t_L g13654 ( 
.A(n_13188),
.Y(n_13654)
);

OR2x2_ASAP7_75t_L g13655 ( 
.A(n_12898),
.B(n_8284),
.Y(n_13655)
);

NAND3xp33_ASAP7_75t_L g13656 ( 
.A(n_13163),
.B(n_11723),
.C(n_10729),
.Y(n_13656)
);

OR2x2_ASAP7_75t_L g13657 ( 
.A(n_12961),
.B(n_8284),
.Y(n_13657)
);

OAI221xp5_ASAP7_75t_SL g13658 ( 
.A1(n_12803),
.A2(n_10158),
.B1(n_10171),
.B2(n_10154),
.C(n_10122),
.Y(n_13658)
);

AOI22xp33_ASAP7_75t_SL g13659 ( 
.A1(n_13075),
.A2(n_10211),
.B1(n_10038),
.B2(n_10158),
.Y(n_13659)
);

NOR2xp33_ASAP7_75t_L g13660 ( 
.A(n_12925),
.B(n_8285),
.Y(n_13660)
);

INVx1_ASAP7_75t_L g13661 ( 
.A(n_13190),
.Y(n_13661)
);

INVx1_ASAP7_75t_L g13662 ( 
.A(n_13191),
.Y(n_13662)
);

INVx1_ASAP7_75t_L g13663 ( 
.A(n_13192),
.Y(n_13663)
);

INVx1_ASAP7_75t_L g13664 ( 
.A(n_13194),
.Y(n_13664)
);

NAND2xp5_ASAP7_75t_L g13665 ( 
.A(n_13097),
.B(n_9944),
.Y(n_13665)
);

HB1xp67_ASAP7_75t_L g13666 ( 
.A(n_13128),
.Y(n_13666)
);

OR2x2_ASAP7_75t_L g13667 ( 
.A(n_12964),
.B(n_8285),
.Y(n_13667)
);

AND2x6_ASAP7_75t_SL g13668 ( 
.A(n_12718),
.B(n_6829),
.Y(n_13668)
);

NAND2xp5_ASAP7_75t_L g13669 ( 
.A(n_13052),
.B(n_9944),
.Y(n_13669)
);

OR2x2_ASAP7_75t_L g13670 ( 
.A(n_12975),
.B(n_8105),
.Y(n_13670)
);

INVx1_ASAP7_75t_L g13671 ( 
.A(n_13206),
.Y(n_13671)
);

NAND2xp5_ASAP7_75t_L g13672 ( 
.A(n_13052),
.B(n_9945),
.Y(n_13672)
);

AND2x2_ASAP7_75t_L g13673 ( 
.A(n_12860),
.B(n_7818),
.Y(n_13673)
);

AND2x2_ASAP7_75t_L g13674 ( 
.A(n_13033),
.B(n_7818),
.Y(n_13674)
);

INVxp67_ASAP7_75t_SL g13675 ( 
.A(n_13132),
.Y(n_13675)
);

NAND2xp5_ASAP7_75t_L g13676 ( 
.A(n_13026),
.B(n_9945),
.Y(n_13676)
);

OR2x2_ASAP7_75t_L g13677 ( 
.A(n_12978),
.B(n_8105),
.Y(n_13677)
);

BUFx2_ASAP7_75t_L g13678 ( 
.A(n_13141),
.Y(n_13678)
);

BUFx2_ASAP7_75t_L g13679 ( 
.A(n_13202),
.Y(n_13679)
);

AOI22xp33_ASAP7_75t_L g13680 ( 
.A1(n_12973),
.A2(n_10231),
.B1(n_10242),
.B2(n_10218),
.Y(n_13680)
);

INVx1_ASAP7_75t_L g13681 ( 
.A(n_12678),
.Y(n_13681)
);

INVx1_ASAP7_75t_L g13682 ( 
.A(n_12680),
.Y(n_13682)
);

HB1xp67_ASAP7_75t_L g13683 ( 
.A(n_12811),
.Y(n_13683)
);

AND2x2_ASAP7_75t_L g13684 ( 
.A(n_13160),
.B(n_7833),
.Y(n_13684)
);

INVx2_ASAP7_75t_L g13685 ( 
.A(n_12793),
.Y(n_13685)
);

NAND2xp5_ASAP7_75t_L g13686 ( 
.A(n_13026),
.B(n_13175),
.Y(n_13686)
);

INVx1_ASAP7_75t_L g13687 ( 
.A(n_12687),
.Y(n_13687)
);

INVx1_ASAP7_75t_L g13688 ( 
.A(n_12689),
.Y(n_13688)
);

AND2x2_ASAP7_75t_L g13689 ( 
.A(n_13161),
.B(n_7833),
.Y(n_13689)
);

AND2x2_ASAP7_75t_SL g13690 ( 
.A(n_12871),
.B(n_7951),
.Y(n_13690)
);

AND2x2_ASAP7_75t_L g13691 ( 
.A(n_13164),
.B(n_7833),
.Y(n_13691)
);

INVx1_ASAP7_75t_L g13692 ( 
.A(n_12988),
.Y(n_13692)
);

AND2x2_ASAP7_75t_L g13693 ( 
.A(n_13169),
.B(n_7882),
.Y(n_13693)
);

OR2x2_ASAP7_75t_L g13694 ( 
.A(n_12986),
.B(n_8111),
.Y(n_13694)
);

AND2x2_ASAP7_75t_L g13695 ( 
.A(n_12971),
.B(n_7882),
.Y(n_13695)
);

BUFx2_ASAP7_75t_SL g13696 ( 
.A(n_12783),
.Y(n_13696)
);

AND2x4_ASAP7_75t_L g13697 ( 
.A(n_12956),
.B(n_10056),
.Y(n_13697)
);

INVx2_ASAP7_75t_L g13698 ( 
.A(n_12795),
.Y(n_13698)
);

OR2x2_ASAP7_75t_L g13699 ( 
.A(n_12990),
.B(n_8111),
.Y(n_13699)
);

AND2x2_ASAP7_75t_L g13700 ( 
.A(n_13050),
.B(n_13086),
.Y(n_13700)
);

INVx1_ASAP7_75t_L g13701 ( 
.A(n_12914),
.Y(n_13701)
);

AND2x2_ASAP7_75t_L g13702 ( 
.A(n_12931),
.B(n_7882),
.Y(n_13702)
);

NAND2xp5_ASAP7_75t_L g13703 ( 
.A(n_12991),
.B(n_9951),
.Y(n_13703)
);

INVx1_ASAP7_75t_L g13704 ( 
.A(n_12965),
.Y(n_13704)
);

NAND2xp5_ASAP7_75t_L g13705 ( 
.A(n_12992),
.B(n_12998),
.Y(n_13705)
);

INVx1_ASAP7_75t_L g13706 ( 
.A(n_13014),
.Y(n_13706)
);

AND2x2_ASAP7_75t_L g13707 ( 
.A(n_12967),
.B(n_7926),
.Y(n_13707)
);

OAI21xp33_ASAP7_75t_L g13708 ( 
.A1(n_13006),
.A2(n_10251),
.B(n_10250),
.Y(n_13708)
);

HB1xp67_ASAP7_75t_L g13709 ( 
.A(n_13219),
.Y(n_13709)
);

AND2x4_ASAP7_75t_SL g13710 ( 
.A(n_13088),
.B(n_7926),
.Y(n_13710)
);

INVx1_ASAP7_75t_L g13711 ( 
.A(n_12995),
.Y(n_13711)
);

INVx1_ASAP7_75t_L g13712 ( 
.A(n_13212),
.Y(n_13712)
);

NAND2xp5_ASAP7_75t_L g13713 ( 
.A(n_12999),
.B(n_9951),
.Y(n_13713)
);

INVx1_ASAP7_75t_L g13714 ( 
.A(n_13007),
.Y(n_13714)
);

NAND2xp5_ASAP7_75t_L g13715 ( 
.A(n_13101),
.B(n_9957),
.Y(n_13715)
);

AND2x4_ASAP7_75t_L g13716 ( 
.A(n_12784),
.B(n_10056),
.Y(n_13716)
);

HB1xp67_ASAP7_75t_L g13717 ( 
.A(n_12798),
.Y(n_13717)
);

BUFx2_ASAP7_75t_L g13718 ( 
.A(n_12806),
.Y(n_13718)
);

INVx1_ASAP7_75t_L g13719 ( 
.A(n_13208),
.Y(n_13719)
);

OR2x2_ASAP7_75t_L g13720 ( 
.A(n_12858),
.B(n_8116),
.Y(n_13720)
);

NAND3xp33_ASAP7_75t_L g13721 ( 
.A(n_13045),
.B(n_10994),
.C(n_9958),
.Y(n_13721)
);

OR2x2_ASAP7_75t_L g13722 ( 
.A(n_13215),
.B(n_8116),
.Y(n_13722)
);

HB1xp67_ASAP7_75t_L g13723 ( 
.A(n_13103),
.Y(n_13723)
);

INVx2_ASAP7_75t_L g13724 ( 
.A(n_13218),
.Y(n_13724)
);

INVx1_ASAP7_75t_L g13725 ( 
.A(n_13213),
.Y(n_13725)
);

HB1xp67_ASAP7_75t_L g13726 ( 
.A(n_13104),
.Y(n_13726)
);

INVx1_ASAP7_75t_L g13727 ( 
.A(n_13068),
.Y(n_13727)
);

INVx1_ASAP7_75t_L g13728 ( 
.A(n_13068),
.Y(n_13728)
);

OR2x2_ASAP7_75t_L g13729 ( 
.A(n_13162),
.B(n_8118),
.Y(n_13729)
);

AND2x2_ASAP7_75t_L g13730 ( 
.A(n_13046),
.B(n_7926),
.Y(n_13730)
);

NAND2xp5_ASAP7_75t_L g13731 ( 
.A(n_13186),
.B(n_9957),
.Y(n_13731)
);

AND2x2_ASAP7_75t_L g13732 ( 
.A(n_13159),
.B(n_7935),
.Y(n_13732)
);

NAND2xp5_ASAP7_75t_L g13733 ( 
.A(n_13171),
.B(n_9958),
.Y(n_13733)
);

OR2x6_ASAP7_75t_L g13734 ( 
.A(n_12972),
.B(n_8797),
.Y(n_13734)
);

AND2x2_ASAP7_75t_L g13735 ( 
.A(n_13146),
.B(n_7935),
.Y(n_13735)
);

INVx1_ASAP7_75t_L g13736 ( 
.A(n_13129),
.Y(n_13736)
);

NAND2xp5_ASAP7_75t_L g13737 ( 
.A(n_13216),
.B(n_9959),
.Y(n_13737)
);

INVx1_ASAP7_75t_L g13738 ( 
.A(n_13129),
.Y(n_13738)
);

AND2x2_ASAP7_75t_L g13739 ( 
.A(n_12989),
.B(n_7935),
.Y(n_13739)
);

HB1xp67_ASAP7_75t_L g13740 ( 
.A(n_12936),
.Y(n_13740)
);

AND2x2_ASAP7_75t_SL g13741 ( 
.A(n_13211),
.B(n_10820),
.Y(n_13741)
);

OR2x2_ASAP7_75t_L g13742 ( 
.A(n_13207),
.B(n_8118),
.Y(n_13742)
);

AND2x2_ASAP7_75t_L g13743 ( 
.A(n_13110),
.B(n_7950),
.Y(n_13743)
);

INVx2_ASAP7_75t_L g13744 ( 
.A(n_12946),
.Y(n_13744)
);

NAND2xp5_ASAP7_75t_L g13745 ( 
.A(n_13221),
.B(n_9959),
.Y(n_13745)
);

INVx2_ASAP7_75t_L g13746 ( 
.A(n_13228),
.Y(n_13746)
);

AOI22xp33_ASAP7_75t_L g13747 ( 
.A1(n_13480),
.A2(n_13077),
.B1(n_13091),
.B2(n_12683),
.Y(n_13747)
);

HB1xp67_ASAP7_75t_L g13748 ( 
.A(n_13433),
.Y(n_13748)
);

INVx1_ASAP7_75t_L g13749 ( 
.A(n_13406),
.Y(n_13749)
);

INVx1_ASAP7_75t_L g13750 ( 
.A(n_13484),
.Y(n_13750)
);

OR2x2_ASAP7_75t_L g13751 ( 
.A(n_13336),
.B(n_13166),
.Y(n_13751)
);

INVx2_ASAP7_75t_SL g13752 ( 
.A(n_13505),
.Y(n_13752)
);

AND2x2_ASAP7_75t_L g13753 ( 
.A(n_13307),
.B(n_13173),
.Y(n_13753)
);

INVx1_ASAP7_75t_L g13754 ( 
.A(n_13380),
.Y(n_13754)
);

HB1xp67_ASAP7_75t_L g13755 ( 
.A(n_13527),
.Y(n_13755)
);

INVx1_ASAP7_75t_L g13756 ( 
.A(n_13527),
.Y(n_13756)
);

AND2x2_ASAP7_75t_L g13757 ( 
.A(n_13293),
.B(n_13158),
.Y(n_13757)
);

AND2x2_ASAP7_75t_L g13758 ( 
.A(n_13700),
.B(n_13017),
.Y(n_13758)
);

INVx1_ASAP7_75t_L g13759 ( 
.A(n_13235),
.Y(n_13759)
);

AND2x2_ASAP7_75t_L g13760 ( 
.A(n_13297),
.B(n_13030),
.Y(n_13760)
);

HB1xp67_ASAP7_75t_L g13761 ( 
.A(n_13265),
.Y(n_13761)
);

AND2x2_ASAP7_75t_L g13762 ( 
.A(n_13294),
.B(n_13059),
.Y(n_13762)
);

NAND2xp5_ASAP7_75t_L g13763 ( 
.A(n_13251),
.B(n_12757),
.Y(n_13763)
);

OR2x2_ASAP7_75t_L g13764 ( 
.A(n_13447),
.B(n_13184),
.Y(n_13764)
);

INVx1_ASAP7_75t_L g13765 ( 
.A(n_13267),
.Y(n_13765)
);

OR2x2_ASAP7_75t_L g13766 ( 
.A(n_13398),
.B(n_12882),
.Y(n_13766)
);

INVx1_ASAP7_75t_L g13767 ( 
.A(n_13280),
.Y(n_13767)
);

NAND2xp5_ASAP7_75t_L g13768 ( 
.A(n_13355),
.B(n_12759),
.Y(n_13768)
);

AND2x2_ASAP7_75t_L g13769 ( 
.A(n_13478),
.B(n_12982),
.Y(n_13769)
);

HB1xp67_ASAP7_75t_L g13770 ( 
.A(n_13265),
.Y(n_13770)
);

AND2x2_ASAP7_75t_L g13771 ( 
.A(n_13354),
.B(n_12985),
.Y(n_13771)
);

HB1xp67_ASAP7_75t_L g13772 ( 
.A(n_13638),
.Y(n_13772)
);

AND2x2_ASAP7_75t_L g13773 ( 
.A(n_13408),
.B(n_12987),
.Y(n_13773)
);

NAND2xp5_ASAP7_75t_L g13774 ( 
.A(n_13277),
.B(n_12762),
.Y(n_13774)
);

INVx2_ASAP7_75t_L g13775 ( 
.A(n_13555),
.Y(n_13775)
);

AND2x2_ASAP7_75t_L g13776 ( 
.A(n_13282),
.B(n_13316),
.Y(n_13776)
);

AND2x2_ASAP7_75t_L g13777 ( 
.A(n_13322),
.B(n_13357),
.Y(n_13777)
);

NAND2xp5_ASAP7_75t_L g13778 ( 
.A(n_13359),
.B(n_12993),
.Y(n_13778)
);

AND2x2_ASAP7_75t_L g13779 ( 
.A(n_13247),
.B(n_13001),
.Y(n_13779)
);

AND2x2_ASAP7_75t_L g13780 ( 
.A(n_13252),
.B(n_13002),
.Y(n_13780)
);

AND2x2_ASAP7_75t_L g13781 ( 
.A(n_13292),
.B(n_13157),
.Y(n_13781)
);

INVx1_ASAP7_75t_L g13782 ( 
.A(n_13723),
.Y(n_13782)
);

BUFx3_ASAP7_75t_L g13783 ( 
.A(n_13466),
.Y(n_13783)
);

INVx1_ASAP7_75t_L g13784 ( 
.A(n_13726),
.Y(n_13784)
);

NAND2xp5_ASAP7_75t_L g13785 ( 
.A(n_13407),
.B(n_13019),
.Y(n_13785)
);

INVx1_ASAP7_75t_L g13786 ( 
.A(n_13718),
.Y(n_13786)
);

INVx1_ASAP7_75t_L g13787 ( 
.A(n_13718),
.Y(n_13787)
);

OR2x2_ASAP7_75t_L g13788 ( 
.A(n_13296),
.B(n_13365),
.Y(n_13788)
);

AND2x2_ASAP7_75t_L g13789 ( 
.A(n_13403),
.B(n_13076),
.Y(n_13789)
);

AND2x2_ASAP7_75t_L g13790 ( 
.A(n_13227),
.B(n_13072),
.Y(n_13790)
);

OR2x2_ASAP7_75t_L g13791 ( 
.A(n_13366),
.B(n_12869),
.Y(n_13791)
);

INVx2_ASAP7_75t_L g13792 ( 
.A(n_13424),
.Y(n_13792)
);

AND2x2_ASAP7_75t_L g13793 ( 
.A(n_13651),
.B(n_13151),
.Y(n_13793)
);

AND2x2_ASAP7_75t_L g13794 ( 
.A(n_13250),
.B(n_13156),
.Y(n_13794)
);

OR2x2_ASAP7_75t_L g13795 ( 
.A(n_13358),
.B(n_13471),
.Y(n_13795)
);

INVx2_ASAP7_75t_L g13796 ( 
.A(n_13436),
.Y(n_13796)
);

INVx2_ASAP7_75t_SL g13797 ( 
.A(n_13263),
.Y(n_13797)
);

OR2x2_ASAP7_75t_L g13798 ( 
.A(n_13479),
.B(n_12891),
.Y(n_13798)
);

INVx1_ASAP7_75t_L g13799 ( 
.A(n_13507),
.Y(n_13799)
);

AND2x4_ASAP7_75t_L g13800 ( 
.A(n_13459),
.B(n_12930),
.Y(n_13800)
);

INVx1_ASAP7_75t_SL g13801 ( 
.A(n_13260),
.Y(n_13801)
);

NAND2xp5_ASAP7_75t_L g13802 ( 
.A(n_13405),
.B(n_13269),
.Y(n_13802)
);

AND2x2_ASAP7_75t_L g13803 ( 
.A(n_13278),
.B(n_13042),
.Y(n_13803)
);

INVx1_ASAP7_75t_L g13804 ( 
.A(n_13572),
.Y(n_13804)
);

AND2x2_ASAP7_75t_L g13805 ( 
.A(n_13284),
.B(n_13044),
.Y(n_13805)
);

OR2x2_ASAP7_75t_L g13806 ( 
.A(n_13481),
.B(n_12933),
.Y(n_13806)
);

NAND2xp5_ASAP7_75t_L g13807 ( 
.A(n_13329),
.B(n_13112),
.Y(n_13807)
);

BUFx2_ASAP7_75t_L g13808 ( 
.A(n_13283),
.Y(n_13808)
);

INVx1_ASAP7_75t_L g13809 ( 
.A(n_13404),
.Y(n_13809)
);

AND2x2_ASAP7_75t_L g13810 ( 
.A(n_13313),
.B(n_13060),
.Y(n_13810)
);

AND2x2_ASAP7_75t_L g13811 ( 
.A(n_13459),
.B(n_12893),
.Y(n_13811)
);

INVx2_ASAP7_75t_L g13812 ( 
.A(n_13466),
.Y(n_13812)
);

AND2x2_ASAP7_75t_L g13813 ( 
.A(n_13286),
.B(n_12912),
.Y(n_13813)
);

NOR2x1_ASAP7_75t_L g13814 ( 
.A(n_13631),
.B(n_12838),
.Y(n_13814)
);

NAND2xp5_ASAP7_75t_L g13815 ( 
.A(n_13635),
.B(n_13032),
.Y(n_13815)
);

INVx1_ASAP7_75t_L g13816 ( 
.A(n_13740),
.Y(n_13816)
);

INVx1_ASAP7_75t_L g13817 ( 
.A(n_13453),
.Y(n_13817)
);

OR2x2_ASAP7_75t_L g13818 ( 
.A(n_13587),
.B(n_13397),
.Y(n_13818)
);

NAND2xp5_ASAP7_75t_L g13819 ( 
.A(n_13646),
.B(n_13054),
.Y(n_13819)
);

NAND5xp2_ASAP7_75t_L g13820 ( 
.A(n_13385),
.B(n_13353),
.C(n_13598),
.D(n_13288),
.E(n_13368),
.Y(n_13820)
);

NAND2xp5_ASAP7_75t_L g13821 ( 
.A(n_13320),
.B(n_13057),
.Y(n_13821)
);

AND2x2_ASAP7_75t_L g13822 ( 
.A(n_13674),
.B(n_13673),
.Y(n_13822)
);

OR2x6_ASAP7_75t_L g13823 ( 
.A(n_13483),
.B(n_12922),
.Y(n_13823)
);

AND2x2_ASAP7_75t_L g13824 ( 
.A(n_13608),
.B(n_13311),
.Y(n_13824)
);

AND2x2_ASAP7_75t_L g13825 ( 
.A(n_13325),
.B(n_13067),
.Y(n_13825)
);

INVx2_ASAP7_75t_L g13826 ( 
.A(n_13743),
.Y(n_13826)
);

OR2x2_ASAP7_75t_L g13827 ( 
.A(n_13314),
.B(n_12839),
.Y(n_13827)
);

INVx1_ASAP7_75t_L g13828 ( 
.A(n_13647),
.Y(n_13828)
);

OR2x2_ASAP7_75t_L g13829 ( 
.A(n_13259),
.B(n_12844),
.Y(n_13829)
);

INVx1_ASAP7_75t_L g13830 ( 
.A(n_13391),
.Y(n_13830)
);

AND2x2_ASAP7_75t_L g13831 ( 
.A(n_13264),
.B(n_12770),
.Y(n_13831)
);

AND2x2_ASAP7_75t_L g13832 ( 
.A(n_13238),
.B(n_13356),
.Y(n_13832)
);

INVxp67_ASAP7_75t_SL g13833 ( 
.A(n_13370),
.Y(n_13833)
);

AND2x4_ASAP7_75t_L g13834 ( 
.A(n_13562),
.B(n_13061),
.Y(n_13834)
);

NOR2xp33_ASAP7_75t_L g13835 ( 
.A(n_13540),
.B(n_13071),
.Y(n_13835)
);

AND2x2_ASAP7_75t_L g13836 ( 
.A(n_13239),
.B(n_12848),
.Y(n_13836)
);

AND2x2_ASAP7_75t_L g13837 ( 
.A(n_13387),
.B(n_12852),
.Y(n_13837)
);

INVx1_ASAP7_75t_L g13838 ( 
.A(n_13494),
.Y(n_13838)
);

AND2x2_ASAP7_75t_L g13839 ( 
.A(n_13334),
.B(n_12853),
.Y(n_13839)
);

AND2x2_ASAP7_75t_L g13840 ( 
.A(n_13603),
.B(n_12856),
.Y(n_13840)
);

AND2x2_ASAP7_75t_L g13841 ( 
.A(n_13285),
.B(n_12861),
.Y(n_13841)
);

OR2x2_ASAP7_75t_L g13842 ( 
.A(n_13324),
.B(n_13078),
.Y(n_13842)
);

INVx2_ASAP7_75t_L g13843 ( 
.A(n_13472),
.Y(n_13843)
);

AND2x4_ASAP7_75t_L g13844 ( 
.A(n_13341),
.B(n_13082),
.Y(n_13844)
);

AND2x2_ASAP7_75t_L g13845 ( 
.A(n_13375),
.B(n_13094),
.Y(n_13845)
);

NAND2xp5_ASAP7_75t_L g13846 ( 
.A(n_13255),
.B(n_13339),
.Y(n_13846)
);

AND2x2_ASAP7_75t_L g13847 ( 
.A(n_13237),
.B(n_13096),
.Y(n_13847)
);

INVx1_ASAP7_75t_L g13848 ( 
.A(n_13361),
.Y(n_13848)
);

INVx1_ASAP7_75t_L g13849 ( 
.A(n_13683),
.Y(n_13849)
);

INVx1_ASAP7_75t_L g13850 ( 
.A(n_13717),
.Y(n_13850)
);

AND2x2_ASAP7_75t_L g13851 ( 
.A(n_13409),
.B(n_13098),
.Y(n_13851)
);

NAND2xp5_ASAP7_75t_L g13852 ( 
.A(n_13344),
.B(n_13100),
.Y(n_13852)
);

AND2x2_ASAP7_75t_L g13853 ( 
.A(n_13300),
.B(n_13105),
.Y(n_13853)
);

AND2x4_ASAP7_75t_L g13854 ( 
.A(n_13487),
.B(n_13107),
.Y(n_13854)
);

AND2x2_ASAP7_75t_L g13855 ( 
.A(n_13261),
.B(n_13122),
.Y(n_13855)
);

AND2x2_ASAP7_75t_L g13856 ( 
.A(n_13266),
.B(n_13149),
.Y(n_13856)
);

NOR3xp33_ASAP7_75t_SL g13857 ( 
.A(n_13350),
.B(n_13303),
.C(n_13244),
.Y(n_13857)
);

INVxp67_ASAP7_75t_SL g13858 ( 
.A(n_13379),
.Y(n_13858)
);

BUFx3_ASAP7_75t_L g13859 ( 
.A(n_13240),
.Y(n_13859)
);

NAND2xp5_ASAP7_75t_L g13860 ( 
.A(n_13347),
.B(n_13150),
.Y(n_13860)
);

AND2x2_ASAP7_75t_L g13861 ( 
.A(n_13274),
.B(n_13152),
.Y(n_13861)
);

INVx1_ASAP7_75t_L g13862 ( 
.A(n_13679),
.Y(n_13862)
);

INVx2_ASAP7_75t_L g13863 ( 
.A(n_13472),
.Y(n_13863)
);

NAND2xp5_ASAP7_75t_L g13864 ( 
.A(n_13242),
.B(n_13176),
.Y(n_13864)
);

INVx1_ASAP7_75t_L g13865 ( 
.A(n_13679),
.Y(n_13865)
);

INVx1_ASAP7_75t_L g13866 ( 
.A(n_13289),
.Y(n_13866)
);

OR2x2_ASAP7_75t_L g13867 ( 
.A(n_13326),
.B(n_13178),
.Y(n_13867)
);

INVx1_ASAP7_75t_L g13868 ( 
.A(n_13305),
.Y(n_13868)
);

HB1xp67_ASAP7_75t_L g13869 ( 
.A(n_13386),
.Y(n_13869)
);

INVx1_ASAP7_75t_L g13870 ( 
.A(n_13363),
.Y(n_13870)
);

INVx1_ASAP7_75t_L g13871 ( 
.A(n_13390),
.Y(n_13871)
);

AND2x2_ASAP7_75t_L g13872 ( 
.A(n_13279),
.B(n_13180),
.Y(n_13872)
);

AND2x2_ASAP7_75t_L g13873 ( 
.A(n_13455),
.B(n_13183),
.Y(n_13873)
);

OR2x2_ASAP7_75t_L g13874 ( 
.A(n_13501),
.B(n_13187),
.Y(n_13874)
);

INVx1_ASAP7_75t_L g13875 ( 
.A(n_13342),
.Y(n_13875)
);

NAND2xp5_ASAP7_75t_L g13876 ( 
.A(n_13246),
.B(n_13189),
.Y(n_13876)
);

NAND2xp5_ASAP7_75t_L g13877 ( 
.A(n_13332),
.B(n_13196),
.Y(n_13877)
);

NAND2xp5_ASAP7_75t_L g13878 ( 
.A(n_13434),
.B(n_13198),
.Y(n_13878)
);

BUFx3_ASAP7_75t_L g13879 ( 
.A(n_13240),
.Y(n_13879)
);

AND2x2_ASAP7_75t_SL g13880 ( 
.A(n_13428),
.B(n_12735),
.Y(n_13880)
);

INVx2_ASAP7_75t_L g13881 ( 
.A(n_13448),
.Y(n_13881)
);

NAND2xp5_ASAP7_75t_L g13882 ( 
.A(n_13323),
.B(n_13201),
.Y(n_13882)
);

NAND2xp5_ASAP7_75t_L g13883 ( 
.A(n_13333),
.B(n_13448),
.Y(n_13883)
);

NAND3xp33_ASAP7_75t_L g13884 ( 
.A(n_13430),
.B(n_12924),
.C(n_13102),
.Y(n_13884)
);

NOR2xp33_ASAP7_75t_L g13885 ( 
.A(n_13532),
.B(n_13222),
.Y(n_13885)
);

AOI22xp33_ASAP7_75t_L g13886 ( 
.A1(n_13656),
.A2(n_13109),
.B1(n_13080),
.B2(n_12870),
.Y(n_13886)
);

INVx2_ASAP7_75t_L g13887 ( 
.A(n_13425),
.Y(n_13887)
);

NAND3xp33_ASAP7_75t_L g13888 ( 
.A(n_13709),
.B(n_13223),
.C(n_13210),
.Y(n_13888)
);

AND2x2_ASAP7_75t_L g13889 ( 
.A(n_13586),
.B(n_13210),
.Y(n_13889)
);

INVx2_ASAP7_75t_L g13890 ( 
.A(n_13427),
.Y(n_13890)
);

INVx3_ASAP7_75t_L g13891 ( 
.A(n_13271),
.Y(n_13891)
);

NAND2xp5_ASAP7_75t_L g13892 ( 
.A(n_13513),
.B(n_12874),
.Y(n_13892)
);

AND2x2_ASAP7_75t_L g13893 ( 
.A(n_13707),
.B(n_12879),
.Y(n_13893)
);

AND2x2_ASAP7_75t_L g13894 ( 
.A(n_13457),
.B(n_12889),
.Y(n_13894)
);

AND2x2_ASAP7_75t_L g13895 ( 
.A(n_13419),
.B(n_7950),
.Y(n_13895)
);

OR2x2_ASAP7_75t_L g13896 ( 
.A(n_13394),
.B(n_13653),
.Y(n_13896)
);

AND2x2_ASAP7_75t_L g13897 ( 
.A(n_13248),
.B(n_7950),
.Y(n_13897)
);

AND2x2_ASAP7_75t_L g13898 ( 
.A(n_13511),
.B(n_7990),
.Y(n_13898)
);

HB1xp67_ASAP7_75t_L g13899 ( 
.A(n_13411),
.Y(n_13899)
);

INVx1_ASAP7_75t_L g13900 ( 
.A(n_13580),
.Y(n_13900)
);

AND2x4_ASAP7_75t_L g13901 ( 
.A(n_13633),
.B(n_7941),
.Y(n_13901)
);

AND2x2_ASAP7_75t_L g13902 ( 
.A(n_13648),
.B(n_7990),
.Y(n_13902)
);

INVx2_ASAP7_75t_L g13903 ( 
.A(n_13437),
.Y(n_13903)
);

AND2x2_ASAP7_75t_L g13904 ( 
.A(n_13512),
.B(n_7990),
.Y(n_13904)
);

NAND2xp5_ASAP7_75t_L g13905 ( 
.A(n_13518),
.B(n_9960),
.Y(n_13905)
);

AND2x2_ASAP7_75t_L g13906 ( 
.A(n_13327),
.B(n_8028),
.Y(n_13906)
);

INVx1_ASAP7_75t_L g13907 ( 
.A(n_13583),
.Y(n_13907)
);

NAND2xp5_ASAP7_75t_L g13908 ( 
.A(n_13544),
.B(n_9960),
.Y(n_13908)
);

INVx2_ASAP7_75t_L g13909 ( 
.A(n_13508),
.Y(n_13909)
);

AND2x2_ASAP7_75t_L g13910 ( 
.A(n_13304),
.B(n_8028),
.Y(n_13910)
);

NAND2x1_ASAP7_75t_SL g13911 ( 
.A(n_13423),
.B(n_10154),
.Y(n_13911)
);

AND2x2_ASAP7_75t_L g13912 ( 
.A(n_13234),
.B(n_8028),
.Y(n_13912)
);

AND2x2_ASAP7_75t_L g13913 ( 
.A(n_13450),
.B(n_8083),
.Y(n_13913)
);

INVx2_ASAP7_75t_L g13914 ( 
.A(n_13640),
.Y(n_13914)
);

NAND2xp5_ASAP7_75t_L g13915 ( 
.A(n_13503),
.B(n_9962),
.Y(n_13915)
);

INVx2_ASAP7_75t_L g13916 ( 
.A(n_13695),
.Y(n_13916)
);

NAND2xp5_ASAP7_75t_L g13917 ( 
.A(n_13519),
.B(n_13229),
.Y(n_13917)
);

OR2x2_ASAP7_75t_L g13918 ( 
.A(n_13306),
.B(n_10250),
.Y(n_13918)
);

BUFx2_ASAP7_75t_L g13919 ( 
.A(n_13631),
.Y(n_13919)
);

AND2x2_ASAP7_75t_L g13920 ( 
.A(n_13469),
.B(n_8083),
.Y(n_13920)
);

INVx1_ASAP7_75t_L g13921 ( 
.A(n_13362),
.Y(n_13921)
);

INVx3_ASAP7_75t_L g13922 ( 
.A(n_13271),
.Y(n_13922)
);

INVx1_ASAP7_75t_L g13923 ( 
.A(n_13364),
.Y(n_13923)
);

INVx1_ASAP7_75t_L g13924 ( 
.A(n_13372),
.Y(n_13924)
);

HB1xp67_ASAP7_75t_L g13925 ( 
.A(n_13349),
.Y(n_13925)
);

AND2x2_ASAP7_75t_L g13926 ( 
.A(n_13381),
.B(n_8083),
.Y(n_13926)
);

INVx1_ASAP7_75t_L g13927 ( 
.A(n_13373),
.Y(n_13927)
);

NOR2xp33_ASAP7_75t_L g13928 ( 
.A(n_13291),
.B(n_9962),
.Y(n_13928)
);

OR2x2_ASAP7_75t_L g13929 ( 
.A(n_13309),
.B(n_10251),
.Y(n_13929)
);

INVx2_ASAP7_75t_L g13930 ( 
.A(n_13730),
.Y(n_13930)
);

NAND2x1_ASAP7_75t_L g13931 ( 
.A(n_13485),
.B(n_10171),
.Y(n_13931)
);

OR2x2_ASAP7_75t_L g13932 ( 
.A(n_13351),
.B(n_10254),
.Y(n_13932)
);

AND2x2_ASAP7_75t_L g13933 ( 
.A(n_13384),
.B(n_8124),
.Y(n_13933)
);

NOR2xp33_ASAP7_75t_L g13934 ( 
.A(n_13632),
.B(n_9964),
.Y(n_13934)
);

AND2x2_ASAP7_75t_L g13935 ( 
.A(n_13547),
.B(n_8124),
.Y(n_13935)
);

HB1xp67_ASAP7_75t_L g13936 ( 
.A(n_13377),
.Y(n_13936)
);

INVx2_ASAP7_75t_L g13937 ( 
.A(n_13739),
.Y(n_13937)
);

INVx1_ASAP7_75t_L g13938 ( 
.A(n_13378),
.Y(n_13938)
);

INVx2_ASAP7_75t_L g13939 ( 
.A(n_13399),
.Y(n_13939)
);

AND2x2_ASAP7_75t_L g13940 ( 
.A(n_13548),
.B(n_8124),
.Y(n_13940)
);

AND2x4_ASAP7_75t_L g13941 ( 
.A(n_13229),
.B(n_10183),
.Y(n_13941)
);

AND2x4_ASAP7_75t_SL g13942 ( 
.A(n_13485),
.B(n_10254),
.Y(n_13942)
);

AND2x2_ASAP7_75t_L g13943 ( 
.A(n_13732),
.B(n_8144),
.Y(n_13943)
);

OAI21xp5_ASAP7_75t_L g13944 ( 
.A1(n_13445),
.A2(n_9659),
.B(n_9742),
.Y(n_13944)
);

INVx1_ASAP7_75t_L g13945 ( 
.A(n_13383),
.Y(n_13945)
);

AND2x4_ASAP7_75t_SL g13946 ( 
.A(n_13371),
.B(n_10255),
.Y(n_13946)
);

OR2x2_ASAP7_75t_L g13947 ( 
.A(n_13317),
.B(n_10255),
.Y(n_13947)
);

OR2x2_ASAP7_75t_L g13948 ( 
.A(n_13438),
.B(n_13439),
.Y(n_13948)
);

OR2x2_ASAP7_75t_L g13949 ( 
.A(n_13490),
.B(n_10262),
.Y(n_13949)
);

NAND2xp5_ASAP7_75t_L g13950 ( 
.A(n_13442),
.B(n_9964),
.Y(n_13950)
);

AND2x2_ASAP7_75t_L g13951 ( 
.A(n_13565),
.B(n_8144),
.Y(n_13951)
);

INVx2_ASAP7_75t_SL g13952 ( 
.A(n_13392),
.Y(n_13952)
);

BUFx2_ASAP7_75t_L g13953 ( 
.A(n_13465),
.Y(n_13953)
);

INVxp67_ASAP7_75t_L g13954 ( 
.A(n_13696),
.Y(n_13954)
);

BUFx2_ASAP7_75t_L g13955 ( 
.A(n_13388),
.Y(n_13955)
);

INVx1_ASAP7_75t_L g13956 ( 
.A(n_13236),
.Y(n_13956)
);

INVx1_ASAP7_75t_L g13957 ( 
.A(n_13243),
.Y(n_13957)
);

NAND2xp5_ASAP7_75t_L g13958 ( 
.A(n_13520),
.B(n_9965),
.Y(n_13958)
);

INVx1_ASAP7_75t_SL g13959 ( 
.A(n_13416),
.Y(n_13959)
);

NOR2xp33_ASAP7_75t_L g13960 ( 
.A(n_13577),
.B(n_9965),
.Y(n_13960)
);

AOI22xp5_ASAP7_75t_L g13961 ( 
.A1(n_13495),
.A2(n_11032),
.B1(n_10759),
.B2(n_10756),
.Y(n_13961)
);

AND2x2_ASAP7_75t_L g13962 ( 
.A(n_13533),
.B(n_8144),
.Y(n_13962)
);

NAND2x1p5_ASAP7_75t_L g13963 ( 
.A(n_13301),
.B(n_6790),
.Y(n_13963)
);

INVx1_ASAP7_75t_L g13964 ( 
.A(n_13249),
.Y(n_13964)
);

NAND2xp5_ASAP7_75t_L g13965 ( 
.A(n_13712),
.B(n_9968),
.Y(n_13965)
);

INVx1_ASAP7_75t_L g13966 ( 
.A(n_13254),
.Y(n_13966)
);

NAND2xp5_ASAP7_75t_L g13967 ( 
.A(n_13637),
.B(n_9968),
.Y(n_13967)
);

AND2x2_ASAP7_75t_L g13968 ( 
.A(n_13516),
.B(n_8149),
.Y(n_13968)
);

OR2x2_ASAP7_75t_L g13969 ( 
.A(n_13492),
.B(n_10262),
.Y(n_13969)
);

NAND2xp5_ASAP7_75t_L g13970 ( 
.A(n_13649),
.B(n_9973),
.Y(n_13970)
);

AND2x2_ASAP7_75t_L g13971 ( 
.A(n_13685),
.B(n_8149),
.Y(n_13971)
);

OR2x2_ASAP7_75t_L g13972 ( 
.A(n_13500),
.B(n_10268),
.Y(n_13972)
);

INVx2_ASAP7_75t_L g13973 ( 
.A(n_13400),
.Y(n_13973)
);

NAND2xp5_ASAP7_75t_L g13974 ( 
.A(n_13661),
.B(n_9973),
.Y(n_13974)
);

NOR2x1_ASAP7_75t_L g13975 ( 
.A(n_13258),
.B(n_10183),
.Y(n_13975)
);

INVx2_ASAP7_75t_SL g13976 ( 
.A(n_13396),
.Y(n_13976)
);

AND2x2_ASAP7_75t_L g13977 ( 
.A(n_13698),
.B(n_8149),
.Y(n_13977)
);

AND2x2_ASAP7_75t_L g13978 ( 
.A(n_13346),
.B(n_8179),
.Y(n_13978)
);

AND2x2_ASAP7_75t_L g13979 ( 
.A(n_13611),
.B(n_13634),
.Y(n_13979)
);

NAND2x1p5_ASAP7_75t_L g13980 ( 
.A(n_13369),
.B(n_6790),
.Y(n_13980)
);

NAND2xp5_ASAP7_75t_L g13981 ( 
.A(n_13662),
.B(n_13663),
.Y(n_13981)
);

AND2x2_ASAP7_75t_L g13982 ( 
.A(n_13636),
.B(n_8179),
.Y(n_13982)
);

AND2x2_ASAP7_75t_L g13983 ( 
.A(n_13645),
.B(n_8179),
.Y(n_13983)
);

NAND2xp5_ASAP7_75t_L g13984 ( 
.A(n_13664),
.B(n_9981),
.Y(n_13984)
);

BUFx2_ASAP7_75t_L g13985 ( 
.A(n_13678),
.Y(n_13985)
);

HB1xp67_ASAP7_75t_L g13986 ( 
.A(n_13270),
.Y(n_13986)
);

NAND2xp5_ASAP7_75t_L g13987 ( 
.A(n_13671),
.B(n_9981),
.Y(n_13987)
);

INVx2_ASAP7_75t_L g13988 ( 
.A(n_13486),
.Y(n_13988)
);

INVx2_ASAP7_75t_L g13989 ( 
.A(n_13497),
.Y(n_13989)
);

AND2x2_ASAP7_75t_L g13990 ( 
.A(n_13524),
.B(n_8233),
.Y(n_13990)
);

NOR2x1_ASAP7_75t_L g13991 ( 
.A(n_13626),
.B(n_10183),
.Y(n_13991)
);

AND2x2_ASAP7_75t_L g13992 ( 
.A(n_13561),
.B(n_8233),
.Y(n_13992)
);

AND2x2_ASAP7_75t_L g13993 ( 
.A(n_13561),
.B(n_8233),
.Y(n_13993)
);

INVx1_ASAP7_75t_L g13994 ( 
.A(n_13429),
.Y(n_13994)
);

NAND2xp5_ASAP7_75t_L g13995 ( 
.A(n_13554),
.B(n_9986),
.Y(n_13995)
);

AND2x2_ASAP7_75t_L g13996 ( 
.A(n_13556),
.B(n_8265),
.Y(n_13996)
);

INVx1_ASAP7_75t_SL g13997 ( 
.A(n_13415),
.Y(n_13997)
);

AND2x2_ASAP7_75t_L g13998 ( 
.A(n_13463),
.B(n_8265),
.Y(n_13998)
);

INVx1_ASAP7_75t_L g13999 ( 
.A(n_13315),
.Y(n_13999)
);

AND2x4_ASAP7_75t_SL g14000 ( 
.A(n_13393),
.B(n_13335),
.Y(n_14000)
);

AND2x2_ASAP7_75t_L g14001 ( 
.A(n_13476),
.B(n_8265),
.Y(n_14001)
);

AND2x4_ASAP7_75t_L g14002 ( 
.A(n_13576),
.B(n_10184),
.Y(n_14002)
);

INVx2_ASAP7_75t_L g14003 ( 
.A(n_13531),
.Y(n_14003)
);

OR2x2_ASAP7_75t_L g14004 ( 
.A(n_13245),
.B(n_13330),
.Y(n_14004)
);

NOR3xp33_ASAP7_75t_SL g14005 ( 
.A(n_13275),
.B(n_11097),
.C(n_11075),
.Y(n_14005)
);

INVx1_ASAP7_75t_SL g14006 ( 
.A(n_13443),
.Y(n_14006)
);

AND2x2_ASAP7_75t_L g14007 ( 
.A(n_13526),
.B(n_13491),
.Y(n_14007)
);

INVx2_ASAP7_75t_SL g14008 ( 
.A(n_13401),
.Y(n_14008)
);

OR2x2_ASAP7_75t_L g14009 ( 
.A(n_13331),
.B(n_10268),
.Y(n_14009)
);

INVx6_ASAP7_75t_L g14010 ( 
.A(n_13595),
.Y(n_14010)
);

NAND2xp5_ASAP7_75t_L g14011 ( 
.A(n_13605),
.B(n_9986),
.Y(n_14011)
);

OR2x2_ASAP7_75t_L g14012 ( 
.A(n_13340),
.B(n_10276),
.Y(n_14012)
);

AND2x2_ASAP7_75t_L g14013 ( 
.A(n_13614),
.B(n_10276),
.Y(n_14013)
);

INVx1_ASAP7_75t_L g14014 ( 
.A(n_13389),
.Y(n_14014)
);

NAND2xp5_ASAP7_75t_L g14015 ( 
.A(n_13607),
.B(n_9997),
.Y(n_14015)
);

INVx2_ASAP7_75t_L g14016 ( 
.A(n_13627),
.Y(n_14016)
);

AND2x4_ASAP7_75t_L g14017 ( 
.A(n_13446),
.B(n_10184),
.Y(n_14017)
);

INVx6_ASAP7_75t_L g14018 ( 
.A(n_13652),
.Y(n_14018)
);

NAND2xp5_ASAP7_75t_L g14019 ( 
.A(n_13435),
.B(n_9997),
.Y(n_14019)
);

NAND2xp5_ASAP7_75t_L g14020 ( 
.A(n_13458),
.B(n_10008),
.Y(n_14020)
);

NAND2xp5_ASAP7_75t_L g14021 ( 
.A(n_13461),
.B(n_10008),
.Y(n_14021)
);

AND2x2_ASAP7_75t_L g14022 ( 
.A(n_13710),
.B(n_10291),
.Y(n_14022)
);

AND2x2_ASAP7_75t_L g14023 ( 
.A(n_13413),
.B(n_10291),
.Y(n_14023)
);

AND2x4_ASAP7_75t_L g14024 ( 
.A(n_13460),
.B(n_10184),
.Y(n_14024)
);

INVx1_ASAP7_75t_L g14025 ( 
.A(n_13382),
.Y(n_14025)
);

INVx3_ASAP7_75t_L g14026 ( 
.A(n_13474),
.Y(n_14026)
);

INVx1_ASAP7_75t_L g14027 ( 
.A(n_13352),
.Y(n_14027)
);

OR2x2_ASAP7_75t_L g14028 ( 
.A(n_13290),
.B(n_10294),
.Y(n_14028)
);

INVx1_ASAP7_75t_L g14029 ( 
.A(n_13262),
.Y(n_14029)
);

NAND2xp5_ASAP7_75t_L g14030 ( 
.A(n_13610),
.B(n_10013),
.Y(n_14030)
);

AND3x1_ASAP7_75t_L g14031 ( 
.A(n_13597),
.B(n_10297),
.C(n_10294),
.Y(n_14031)
);

NOR2xp67_ASAP7_75t_SL g14032 ( 
.A(n_13319),
.B(n_7195),
.Y(n_14032)
);

NAND2xp5_ASAP7_75t_L g14033 ( 
.A(n_13376),
.B(n_10013),
.Y(n_14033)
);

INVx1_ASAP7_75t_L g14034 ( 
.A(n_13338),
.Y(n_14034)
);

INVx3_ASAP7_75t_L g14035 ( 
.A(n_13474),
.Y(n_14035)
);

HB1xp67_ASAP7_75t_L g14036 ( 
.A(n_13462),
.Y(n_14036)
);

INVx1_ASAP7_75t_L g14037 ( 
.A(n_13475),
.Y(n_14037)
);

AND2x2_ASAP7_75t_L g14038 ( 
.A(n_13552),
.B(n_10297),
.Y(n_14038)
);

AND2x2_ASAP7_75t_L g14039 ( 
.A(n_13440),
.B(n_10302),
.Y(n_14039)
);

AND2x2_ASAP7_75t_L g14040 ( 
.A(n_13441),
.B(n_10302),
.Y(n_14040)
);

INVx3_ASAP7_75t_L g14041 ( 
.A(n_13650),
.Y(n_14041)
);

NAND2xp5_ASAP7_75t_L g14042 ( 
.A(n_13417),
.B(n_10015),
.Y(n_14042)
);

AND2x2_ASAP7_75t_L g14043 ( 
.A(n_13702),
.B(n_10311),
.Y(n_14043)
);

OR2x2_ASAP7_75t_L g14044 ( 
.A(n_13464),
.B(n_10311),
.Y(n_14044)
);

AND2x2_ASAP7_75t_L g14045 ( 
.A(n_13402),
.B(n_10314),
.Y(n_14045)
);

INVx4_ASAP7_75t_L g14046 ( 
.A(n_13295),
.Y(n_14046)
);

AND2x2_ASAP7_75t_L g14047 ( 
.A(n_13618),
.B(n_10314),
.Y(n_14047)
);

AND2x2_ASAP7_75t_L g14048 ( 
.A(n_13620),
.B(n_10325),
.Y(n_14048)
);

AND2x2_ASAP7_75t_L g14049 ( 
.A(n_13630),
.B(n_10325),
.Y(n_14049)
);

OR2x2_ASAP7_75t_L g14050 ( 
.A(n_13467),
.B(n_13468),
.Y(n_14050)
);

INVx1_ASAP7_75t_L g14051 ( 
.A(n_13298),
.Y(n_14051)
);

AND2x4_ASAP7_75t_SL g14052 ( 
.A(n_13606),
.B(n_10329),
.Y(n_14052)
);

OR2x2_ASAP7_75t_L g14053 ( 
.A(n_13470),
.B(n_13477),
.Y(n_14053)
);

AOI22xp33_ASAP7_75t_L g14054 ( 
.A1(n_13542),
.A2(n_10242),
.B1(n_10211),
.B2(n_11125),
.Y(n_14054)
);

AND2x2_ASAP7_75t_L g14055 ( 
.A(n_13482),
.B(n_10329),
.Y(n_14055)
);

INVx3_ASAP7_75t_L g14056 ( 
.A(n_13584),
.Y(n_14056)
);

INVx1_ASAP7_75t_L g14057 ( 
.A(n_13299),
.Y(n_14057)
);

NAND2xp5_ASAP7_75t_L g14058 ( 
.A(n_13509),
.B(n_10015),
.Y(n_14058)
);

INVx1_ASAP7_75t_L g14059 ( 
.A(n_13302),
.Y(n_14059)
);

INVx1_ASAP7_75t_L g14060 ( 
.A(n_13312),
.Y(n_14060)
);

BUFx2_ASAP7_75t_L g14061 ( 
.A(n_13678),
.Y(n_14061)
);

NAND2xp5_ASAP7_75t_SL g14062 ( 
.A(n_13489),
.B(n_11139),
.Y(n_14062)
);

OR2x2_ASAP7_75t_L g14063 ( 
.A(n_13253),
.B(n_10330),
.Y(n_14063)
);

INVx2_ASAP7_75t_L g14064 ( 
.A(n_13735),
.Y(n_14064)
);

INVx1_ASAP7_75t_L g14065 ( 
.A(n_13318),
.Y(n_14065)
);

HB1xp67_ASAP7_75t_L g14066 ( 
.A(n_13502),
.Y(n_14066)
);

NOR2xp33_ASAP7_75t_R g14067 ( 
.A(n_13276),
.B(n_9423),
.Y(n_14067)
);

INVx2_ASAP7_75t_L g14068 ( 
.A(n_13591),
.Y(n_14068)
);

NOR2xp33_ASAP7_75t_L g14069 ( 
.A(n_13525),
.B(n_10024),
.Y(n_14069)
);

AND2x2_ASAP7_75t_L g14070 ( 
.A(n_13622),
.B(n_10330),
.Y(n_14070)
);

INVx2_ASAP7_75t_SL g14071 ( 
.A(n_13412),
.Y(n_14071)
);

AND2x2_ASAP7_75t_L g14072 ( 
.A(n_13328),
.B(n_10331),
.Y(n_14072)
);

NAND2xp5_ASAP7_75t_L g14073 ( 
.A(n_13421),
.B(n_10024),
.Y(n_14073)
);

INVx1_ASAP7_75t_SL g14074 ( 
.A(n_13287),
.Y(n_14074)
);

AND2x2_ASAP7_75t_L g14075 ( 
.A(n_13609),
.B(n_10331),
.Y(n_14075)
);

INVx2_ASAP7_75t_L g14076 ( 
.A(n_13601),
.Y(n_14076)
);

NAND2xp5_ASAP7_75t_L g14077 ( 
.A(n_13623),
.B(n_13619),
.Y(n_14077)
);

INVx2_ASAP7_75t_L g14078 ( 
.A(n_13374),
.Y(n_14078)
);

AND2x2_ASAP7_75t_L g14079 ( 
.A(n_13684),
.B(n_10337),
.Y(n_14079)
);

INVx1_ASAP7_75t_L g14080 ( 
.A(n_13414),
.Y(n_14080)
);

INVx1_ASAP7_75t_L g14081 ( 
.A(n_13456),
.Y(n_14081)
);

NAND2xp5_ASAP7_75t_L g14082 ( 
.A(n_13692),
.B(n_10025),
.Y(n_14082)
);

AND2x2_ASAP7_75t_L g14083 ( 
.A(n_13689),
.B(n_10337),
.Y(n_14083)
);

INVx3_ASAP7_75t_L g14084 ( 
.A(n_13744),
.Y(n_14084)
);

INVx2_ASAP7_75t_L g14085 ( 
.A(n_13593),
.Y(n_14085)
);

INVx1_ASAP7_75t_L g14086 ( 
.A(n_13256),
.Y(n_14086)
);

INVx1_ASAP7_75t_L g14087 ( 
.A(n_13686),
.Y(n_14087)
);

AND2x4_ASAP7_75t_L g14088 ( 
.A(n_13241),
.B(n_7941),
.Y(n_14088)
);

INVx2_ASAP7_75t_L g14089 ( 
.A(n_13655),
.Y(n_14089)
);

HB1xp67_ASAP7_75t_L g14090 ( 
.A(n_13502),
.Y(n_14090)
);

OR2x2_ASAP7_75t_L g14091 ( 
.A(n_13233),
.B(n_10338),
.Y(n_14091)
);

INVx1_ASAP7_75t_L g14092 ( 
.A(n_13418),
.Y(n_14092)
);

NAND2xp5_ASAP7_75t_L g14093 ( 
.A(n_13701),
.B(n_10025),
.Y(n_14093)
);

INVx1_ASAP7_75t_L g14094 ( 
.A(n_13473),
.Y(n_14094)
);

AND2x2_ASAP7_75t_L g14095 ( 
.A(n_13691),
.B(n_10338),
.Y(n_14095)
);

NAND2xp5_ASAP7_75t_L g14096 ( 
.A(n_13704),
.B(n_10030),
.Y(n_14096)
);

AND2x2_ASAP7_75t_L g14097 ( 
.A(n_13693),
.B(n_10340),
.Y(n_14097)
);

AND2x2_ASAP7_75t_L g14098 ( 
.A(n_13257),
.B(n_10340),
.Y(n_14098)
);

HB1xp67_ASAP7_75t_L g14099 ( 
.A(n_13654),
.Y(n_14099)
);

INVx1_ASAP7_75t_L g14100 ( 
.A(n_13488),
.Y(n_14100)
);

AND2x4_ASAP7_75t_L g14101 ( 
.A(n_13585),
.B(n_10346),
.Y(n_14101)
);

AND2x2_ASAP7_75t_L g14102 ( 
.A(n_13422),
.B(n_10346),
.Y(n_14102)
);

INVx1_ASAP7_75t_L g14103 ( 
.A(n_13522),
.Y(n_14103)
);

INVx2_ASAP7_75t_L g14104 ( 
.A(n_13582),
.Y(n_14104)
);

INVx1_ASAP7_75t_L g14105 ( 
.A(n_13345),
.Y(n_14105)
);

NAND2xp5_ASAP7_75t_L g14106 ( 
.A(n_13493),
.B(n_10030),
.Y(n_14106)
);

INVx1_ASAP7_75t_L g14107 ( 
.A(n_13722),
.Y(n_14107)
);

AND2x2_ASAP7_75t_L g14108 ( 
.A(n_13420),
.B(n_10368),
.Y(n_14108)
);

INVx1_ASAP7_75t_L g14109 ( 
.A(n_13395),
.Y(n_14109)
);

NOR2xp33_ASAP7_75t_SL g14110 ( 
.A(n_13310),
.B(n_8797),
.Y(n_14110)
);

INVx3_ASAP7_75t_L g14111 ( 
.A(n_13697),
.Y(n_14111)
);

AND2x2_ASAP7_75t_L g14112 ( 
.A(n_13230),
.B(n_10368),
.Y(n_14112)
);

INVx3_ASAP7_75t_L g14113 ( 
.A(n_13697),
.Y(n_14113)
);

INVx1_ASAP7_75t_L g14114 ( 
.A(n_13410),
.Y(n_14114)
);

OR2x2_ASAP7_75t_L g14115 ( 
.A(n_13281),
.B(n_10371),
.Y(n_14115)
);

INVx1_ASAP7_75t_L g14116 ( 
.A(n_13612),
.Y(n_14116)
);

AND2x4_ASAP7_75t_L g14117 ( 
.A(n_13231),
.B(n_8200),
.Y(n_14117)
);

INVxp33_ASAP7_75t_L g14118 ( 
.A(n_13523),
.Y(n_14118)
);

INVx2_ASAP7_75t_L g14119 ( 
.A(n_13716),
.Y(n_14119)
);

INVx2_ASAP7_75t_L g14120 ( 
.A(n_13716),
.Y(n_14120)
);

NAND2xp5_ASAP7_75t_L g14121 ( 
.A(n_13496),
.B(n_10033),
.Y(n_14121)
);

INVx1_ASAP7_75t_L g14122 ( 
.A(n_13232),
.Y(n_14122)
);

INVx2_ASAP7_75t_SL g14123 ( 
.A(n_13690),
.Y(n_14123)
);

NAND2xp5_ASAP7_75t_L g14124 ( 
.A(n_13504),
.B(n_10033),
.Y(n_14124)
);

OR2x2_ASAP7_75t_L g14125 ( 
.A(n_13499),
.B(n_10371),
.Y(n_14125)
);

AND2x2_ASAP7_75t_L g14126 ( 
.A(n_13272),
.B(n_10378),
.Y(n_14126)
);

INVx1_ASAP7_75t_L g14127 ( 
.A(n_13273),
.Y(n_14127)
);

NAND3xp33_ASAP7_75t_L g14128 ( 
.A(n_13628),
.B(n_10041),
.C(n_10035),
.Y(n_14128)
);

AND2x2_ASAP7_75t_L g14129 ( 
.A(n_13660),
.B(n_10378),
.Y(n_14129)
);

INVxp67_ASAP7_75t_L g14130 ( 
.A(n_13644),
.Y(n_14130)
);

AND2x2_ASAP7_75t_L g14131 ( 
.A(n_13724),
.B(n_10100),
.Y(n_14131)
);

NAND2xp5_ASAP7_75t_L g14132 ( 
.A(n_13553),
.B(n_10035),
.Y(n_14132)
);

INVx1_ASAP7_75t_L g14133 ( 
.A(n_13705),
.Y(n_14133)
);

AND2x2_ASAP7_75t_L g14134 ( 
.A(n_13711),
.B(n_10100),
.Y(n_14134)
);

AND2x2_ASAP7_75t_L g14135 ( 
.A(n_13641),
.B(n_8291),
.Y(n_14135)
);

AND2x2_ASAP7_75t_L g14136 ( 
.A(n_13444),
.B(n_8291),
.Y(n_14136)
);

AND2x2_ASAP7_75t_L g14137 ( 
.A(n_13452),
.B(n_8291),
.Y(n_14137)
);

NAND2xp5_ASAP7_75t_L g14138 ( 
.A(n_13706),
.B(n_10041),
.Y(n_14138)
);

INVx1_ASAP7_75t_SL g14139 ( 
.A(n_13545),
.Y(n_14139)
);

INVx1_ASAP7_75t_L g14140 ( 
.A(n_13657),
.Y(n_14140)
);

AND2x4_ASAP7_75t_L g14141 ( 
.A(n_13510),
.B(n_8200),
.Y(n_14141)
);

AND2x4_ASAP7_75t_L g14142 ( 
.A(n_13714),
.B(n_8200),
.Y(n_14142)
);

NOR2xp67_ASAP7_75t_L g14143 ( 
.A(n_13454),
.B(n_10048),
.Y(n_14143)
);

AND2x2_ASAP7_75t_L g14144 ( 
.A(n_13559),
.B(n_8303),
.Y(n_14144)
);

NAND2xp5_ASAP7_75t_SL g14145 ( 
.A(n_13506),
.B(n_11172),
.Y(n_14145)
);

AND2x2_ASAP7_75t_L g14146 ( 
.A(n_13560),
.B(n_8303),
.Y(n_14146)
);

AND2x2_ASAP7_75t_L g14147 ( 
.A(n_13567),
.B(n_8303),
.Y(n_14147)
);

AND2x4_ASAP7_75t_L g14148 ( 
.A(n_13588),
.B(n_8200),
.Y(n_14148)
);

AND2x2_ASAP7_75t_L g14149 ( 
.A(n_13570),
.B(n_10381),
.Y(n_14149)
);

AND2x2_ASAP7_75t_L g14150 ( 
.A(n_13571),
.B(n_10385),
.Y(n_14150)
);

AND2x4_ASAP7_75t_L g14151 ( 
.A(n_13592),
.B(n_8200),
.Y(n_14151)
);

AND2x2_ASAP7_75t_L g14152 ( 
.A(n_13574),
.B(n_10385),
.Y(n_14152)
);

NAND2xp5_ASAP7_75t_L g14153 ( 
.A(n_13581),
.B(n_10048),
.Y(n_14153)
);

NAND2xp5_ASAP7_75t_L g14154 ( 
.A(n_13604),
.B(n_10049),
.Y(n_14154)
);

INVx2_ASAP7_75t_L g14155 ( 
.A(n_13729),
.Y(n_14155)
);

OAI22xp5_ASAP7_75t_L g14156 ( 
.A1(n_13659),
.A2(n_8893),
.B1(n_10211),
.B2(n_10064),
.Y(n_14156)
);

AND2x2_ASAP7_75t_L g14157 ( 
.A(n_13536),
.B(n_8968),
.Y(n_14157)
);

NAND2xp5_ASAP7_75t_L g14158 ( 
.A(n_13550),
.B(n_10049),
.Y(n_14158)
);

AND2x4_ASAP7_75t_L g14159 ( 
.A(n_13600),
.B(n_8203),
.Y(n_14159)
);

AND2x2_ASAP7_75t_L g14160 ( 
.A(n_13538),
.B(n_8968),
.Y(n_14160)
);

AND2x4_ASAP7_75t_SL g14161 ( 
.A(n_13546),
.B(n_5781),
.Y(n_14161)
);

HB1xp67_ASAP7_75t_L g14162 ( 
.A(n_13308),
.Y(n_14162)
);

AND4x1_ASAP7_75t_L g14163 ( 
.A(n_13432),
.B(n_10828),
.C(n_10833),
.D(n_10824),
.Y(n_14163)
);

NAND2xp5_ASAP7_75t_L g14164 ( 
.A(n_13590),
.B(n_10064),
.Y(n_14164)
);

INVx1_ASAP7_75t_L g14165 ( 
.A(n_13667),
.Y(n_14165)
);

INVx2_ASAP7_75t_L g14166 ( 
.A(n_13734),
.Y(n_14166)
);

BUFx2_ASAP7_75t_L g14167 ( 
.A(n_13539),
.Y(n_14167)
);

OR2x2_ASAP7_75t_L g14168 ( 
.A(n_13367),
.B(n_9670),
.Y(n_14168)
);

AND2x2_ASAP7_75t_L g14169 ( 
.A(n_13719),
.B(n_8984),
.Y(n_14169)
);

INVx1_ASAP7_75t_L g14170 ( 
.A(n_13451),
.Y(n_14170)
);

OR2x2_ASAP7_75t_L g14171 ( 
.A(n_13720),
.B(n_9670),
.Y(n_14171)
);

INVx2_ASAP7_75t_L g14172 ( 
.A(n_13734),
.Y(n_14172)
);

INVx2_ASAP7_75t_L g14173 ( 
.A(n_13321),
.Y(n_14173)
);

AND2x4_ASAP7_75t_L g14174 ( 
.A(n_13515),
.B(n_8203),
.Y(n_14174)
);

NAND2xp5_ASAP7_75t_L g14175 ( 
.A(n_13590),
.B(n_10065),
.Y(n_14175)
);

AND2x2_ASAP7_75t_L g14176 ( 
.A(n_13725),
.B(n_8984),
.Y(n_14176)
);

AND2x2_ASAP7_75t_L g14177 ( 
.A(n_13517),
.B(n_13521),
.Y(n_14177)
);

NAND5xp2_ASAP7_75t_SL g14178 ( 
.A(n_13741),
.B(n_11049),
.C(n_10836),
.D(n_10772),
.E(n_11138),
.Y(n_14178)
);

INVx1_ASAP7_75t_L g14179 ( 
.A(n_13449),
.Y(n_14179)
);

OR2x2_ASAP7_75t_L g14180 ( 
.A(n_13498),
.B(n_9670),
.Y(n_14180)
);

INVx1_ASAP7_75t_L g14181 ( 
.A(n_13348),
.Y(n_14181)
);

BUFx3_ASAP7_75t_L g14182 ( 
.A(n_13528),
.Y(n_14182)
);

INVx3_ASAP7_75t_L g14183 ( 
.A(n_13668),
.Y(n_14183)
);

OR2x2_ASAP7_75t_L g14184 ( 
.A(n_13670),
.B(n_9670),
.Y(n_14184)
);

BUFx2_ASAP7_75t_SL g14185 ( 
.A(n_13426),
.Y(n_14185)
);

AND2x2_ASAP7_75t_L g14186 ( 
.A(n_13431),
.B(n_8986),
.Y(n_14186)
);

AND2x2_ASAP7_75t_L g14187 ( 
.A(n_13615),
.B(n_8986),
.Y(n_14187)
);

INVx3_ASAP7_75t_L g14188 ( 
.A(n_13599),
.Y(n_14188)
);

AND2x2_ASAP7_75t_L g14189 ( 
.A(n_13579),
.B(n_8990),
.Y(n_14189)
);

NOR2xp67_ASAP7_75t_L g14190 ( 
.A(n_13360),
.B(n_10065),
.Y(n_14190)
);

NAND2xp5_ASAP7_75t_SL g14191 ( 
.A(n_13665),
.B(n_10069),
.Y(n_14191)
);

OR2x2_ASAP7_75t_L g14192 ( 
.A(n_13677),
.B(n_8216),
.Y(n_14192)
);

INVx1_ASAP7_75t_L g14193 ( 
.A(n_13564),
.Y(n_14193)
);

INVx1_ASAP7_75t_L g14194 ( 
.A(n_13742),
.Y(n_14194)
);

INVx1_ASAP7_75t_L g14195 ( 
.A(n_13985),
.Y(n_14195)
);

AND2x2_ASAP7_75t_L g14196 ( 
.A(n_13824),
.B(n_13337),
.Y(n_14196)
);

OAI211xp5_ASAP7_75t_L g14197 ( 
.A1(n_13886),
.A2(n_13563),
.B(n_13682),
.C(n_13681),
.Y(n_14197)
);

AND2x2_ASAP7_75t_L g14198 ( 
.A(n_13760),
.B(n_13343),
.Y(n_14198)
);

AND2x2_ASAP7_75t_L g14199 ( 
.A(n_13832),
.B(n_13694),
.Y(n_14199)
);

INVx2_ASAP7_75t_L g14200 ( 
.A(n_13783),
.Y(n_14200)
);

NAND2xp5_ASAP7_75t_L g14201 ( 
.A(n_13880),
.B(n_13624),
.Y(n_14201)
);

INVx1_ASAP7_75t_L g14202 ( 
.A(n_13985),
.Y(n_14202)
);

NOR2xp33_ASAP7_75t_L g14203 ( 
.A(n_14183),
.B(n_14018),
.Y(n_14203)
);

INVx2_ASAP7_75t_L g14204 ( 
.A(n_14018),
.Y(n_14204)
);

OR2x2_ASAP7_75t_L g14205 ( 
.A(n_13766),
.B(n_13699),
.Y(n_14205)
);

AND4x1_ASAP7_75t_L g14206 ( 
.A(n_13857),
.B(n_13594),
.C(n_13568),
.D(n_13589),
.Y(n_14206)
);

INVx2_ASAP7_75t_L g14207 ( 
.A(n_14026),
.Y(n_14207)
);

AND2x4_ASAP7_75t_L g14208 ( 
.A(n_13752),
.B(n_13859),
.Y(n_14208)
);

INVx1_ASAP7_75t_L g14209 ( 
.A(n_14061),
.Y(n_14209)
);

AND2x2_ASAP7_75t_L g14210 ( 
.A(n_13776),
.B(n_13687),
.Y(n_14210)
);

OR2x2_ASAP7_75t_L g14211 ( 
.A(n_13818),
.B(n_13596),
.Y(n_14211)
);

INVx1_ASAP7_75t_L g14212 ( 
.A(n_14061),
.Y(n_14212)
);

NOR2xp67_ASAP7_75t_L g14213 ( 
.A(n_13891),
.B(n_13621),
.Y(n_14213)
);

BUFx3_ASAP7_75t_L g14214 ( 
.A(n_13879),
.Y(n_14214)
);

OR2x2_ASAP7_75t_L g14215 ( 
.A(n_13959),
.B(n_13602),
.Y(n_14215)
);

INVx2_ASAP7_75t_L g14216 ( 
.A(n_14035),
.Y(n_14216)
);

INVx2_ASAP7_75t_L g14217 ( 
.A(n_13922),
.Y(n_14217)
);

AND2x2_ASAP7_75t_L g14218 ( 
.A(n_13777),
.B(n_13688),
.Y(n_14218)
);

INVx4_ASAP7_75t_L g14219 ( 
.A(n_14046),
.Y(n_14219)
);

OR2x2_ASAP7_75t_L g14220 ( 
.A(n_13788),
.B(n_13613),
.Y(n_14220)
);

INVx2_ASAP7_75t_L g14221 ( 
.A(n_13769),
.Y(n_14221)
);

INVx1_ASAP7_75t_L g14222 ( 
.A(n_14066),
.Y(n_14222)
);

NAND2xp5_ASAP7_75t_L g14223 ( 
.A(n_13790),
.B(n_13625),
.Y(n_14223)
);

INVx1_ASAP7_75t_L g14224 ( 
.A(n_14090),
.Y(n_14224)
);

INVx1_ASAP7_75t_SL g14225 ( 
.A(n_13753),
.Y(n_14225)
);

INVx1_ASAP7_75t_L g14226 ( 
.A(n_13761),
.Y(n_14226)
);

INVx1_ASAP7_75t_L g14227 ( 
.A(n_13770),
.Y(n_14227)
);

OR2x2_ASAP7_75t_L g14228 ( 
.A(n_13997),
.B(n_13616),
.Y(n_14228)
);

OR2x2_ASAP7_75t_L g14229 ( 
.A(n_14074),
.B(n_13802),
.Y(n_14229)
);

NAND2xp5_ASAP7_75t_L g14230 ( 
.A(n_14006),
.B(n_13514),
.Y(n_14230)
);

NAND2xp5_ASAP7_75t_L g14231 ( 
.A(n_14007),
.B(n_13675),
.Y(n_14231)
);

AND2x2_ASAP7_75t_L g14232 ( 
.A(n_13762),
.B(n_13529),
.Y(n_14232)
);

AND2x2_ASAP7_75t_L g14233 ( 
.A(n_13793),
.B(n_13530),
.Y(n_14233)
);

AND2x2_ASAP7_75t_L g14234 ( 
.A(n_13781),
.B(n_13534),
.Y(n_14234)
);

INVx3_ASAP7_75t_L g14235 ( 
.A(n_13800),
.Y(n_14235)
);

INVx1_ASAP7_75t_L g14236 ( 
.A(n_13808),
.Y(n_14236)
);

INVx1_ASAP7_75t_L g14237 ( 
.A(n_13808),
.Y(n_14237)
);

BUFx2_ASAP7_75t_L g14238 ( 
.A(n_14167),
.Y(n_14238)
);

AND2x2_ASAP7_75t_L g14239 ( 
.A(n_13757),
.B(n_13535),
.Y(n_14239)
);

INVx1_ASAP7_75t_L g14240 ( 
.A(n_13748),
.Y(n_14240)
);

INVx2_ASAP7_75t_L g14241 ( 
.A(n_13953),
.Y(n_14241)
);

AND2x4_ASAP7_75t_L g14242 ( 
.A(n_13797),
.B(n_13812),
.Y(n_14242)
);

AND2x2_ASAP7_75t_L g14243 ( 
.A(n_13794),
.B(n_13549),
.Y(n_14243)
);

AND2x2_ASAP7_75t_L g14244 ( 
.A(n_13771),
.B(n_13551),
.Y(n_14244)
);

INVx1_ASAP7_75t_L g14245 ( 
.A(n_13772),
.Y(n_14245)
);

OR2x2_ASAP7_75t_L g14246 ( 
.A(n_14071),
.B(n_13703),
.Y(n_14246)
);

AND2x2_ASAP7_75t_L g14247 ( 
.A(n_13773),
.B(n_13557),
.Y(n_14247)
);

AND2x4_ASAP7_75t_SL g14248 ( 
.A(n_13758),
.B(n_13558),
.Y(n_14248)
);

NAND2xp5_ASAP7_75t_L g14249 ( 
.A(n_13833),
.B(n_13666),
.Y(n_14249)
);

AND2x2_ASAP7_75t_L g14250 ( 
.A(n_13810),
.B(n_13566),
.Y(n_14250)
);

OR2x2_ASAP7_75t_L g14251 ( 
.A(n_13764),
.B(n_13713),
.Y(n_14251)
);

NAND2xp5_ASAP7_75t_L g14252 ( 
.A(n_13858),
.B(n_13642),
.Y(n_14252)
);

AND2x2_ASAP7_75t_L g14253 ( 
.A(n_13780),
.B(n_13569),
.Y(n_14253)
);

AND2x4_ASAP7_75t_L g14254 ( 
.A(n_13952),
.B(n_13573),
.Y(n_14254)
);

BUFx3_ASAP7_75t_L g14255 ( 
.A(n_13811),
.Y(n_14255)
);

INVx1_ASAP7_75t_SL g14256 ( 
.A(n_13911),
.Y(n_14256)
);

AND2x2_ASAP7_75t_L g14257 ( 
.A(n_13779),
.B(n_13575),
.Y(n_14257)
);

NAND2xp33_ASAP7_75t_R g14258 ( 
.A(n_13953),
.B(n_13727),
.Y(n_14258)
);

AND2x4_ASAP7_75t_L g14259 ( 
.A(n_13976),
.B(n_13578),
.Y(n_14259)
);

BUFx3_ASAP7_75t_L g14260 ( 
.A(n_13834),
.Y(n_14260)
);

INVx1_ASAP7_75t_L g14261 ( 
.A(n_13889),
.Y(n_14261)
);

NAND2xp5_ASAP7_75t_L g14262 ( 
.A(n_13979),
.B(n_13643),
.Y(n_14262)
);

AND2x2_ASAP7_75t_L g14263 ( 
.A(n_13822),
.B(n_13728),
.Y(n_14263)
);

INVx1_ASAP7_75t_L g14264 ( 
.A(n_14099),
.Y(n_14264)
);

AND2x2_ASAP7_75t_L g14265 ( 
.A(n_13902),
.B(n_13736),
.Y(n_14265)
);

AND2x2_ASAP7_75t_L g14266 ( 
.A(n_13978),
.B(n_13738),
.Y(n_14266)
);

HB1xp67_ASAP7_75t_L g14267 ( 
.A(n_13823),
.Y(n_14267)
);

AND2x2_ASAP7_75t_L g14268 ( 
.A(n_13951),
.B(n_13733),
.Y(n_14268)
);

INVx1_ASAP7_75t_SL g14269 ( 
.A(n_13801),
.Y(n_14269)
);

INVx1_ASAP7_75t_L g14270 ( 
.A(n_13843),
.Y(n_14270)
);

NAND2xp5_ASAP7_75t_L g14271 ( 
.A(n_13933),
.B(n_13836),
.Y(n_14271)
);

NAND2xp5_ASAP7_75t_L g14272 ( 
.A(n_13837),
.B(n_13926),
.Y(n_14272)
);

OR2x2_ASAP7_75t_L g14273 ( 
.A(n_13746),
.B(n_13617),
.Y(n_14273)
);

INVx2_ASAP7_75t_L g14274 ( 
.A(n_13863),
.Y(n_14274)
);

AND2x2_ASAP7_75t_L g14275 ( 
.A(n_13789),
.B(n_13537),
.Y(n_14275)
);

AND2x2_ASAP7_75t_L g14276 ( 
.A(n_13906),
.B(n_13731),
.Y(n_14276)
);

INVx2_ASAP7_75t_L g14277 ( 
.A(n_13895),
.Y(n_14277)
);

AND2x2_ASAP7_75t_L g14278 ( 
.A(n_13813),
.B(n_13541),
.Y(n_14278)
);

AOI21xp33_ASAP7_75t_L g14279 ( 
.A1(n_14118),
.A2(n_13629),
.B(n_13543),
.Y(n_14279)
);

INVx5_ASAP7_75t_L g14280 ( 
.A(n_14167),
.Y(n_14280)
);

AOI221xp5_ASAP7_75t_L g14281 ( 
.A1(n_14178),
.A2(n_13639),
.B1(n_13721),
.B2(n_13680),
.C(n_13737),
.Y(n_14281)
);

INVx6_ASAP7_75t_L g14282 ( 
.A(n_13823),
.Y(n_14282)
);

OAI21xp33_ASAP7_75t_L g14283 ( 
.A1(n_13820),
.A2(n_13708),
.B(n_13715),
.Y(n_14283)
);

NAND2xp5_ASAP7_75t_L g14284 ( 
.A(n_13851),
.B(n_13839),
.Y(n_14284)
);

AND2x2_ASAP7_75t_L g14285 ( 
.A(n_13805),
.B(n_13676),
.Y(n_14285)
);

INVx1_ASAP7_75t_L g14286 ( 
.A(n_13955),
.Y(n_14286)
);

NAND2xp5_ASAP7_75t_L g14287 ( 
.A(n_14084),
.B(n_13669),
.Y(n_14287)
);

NAND2xp5_ASAP7_75t_L g14288 ( 
.A(n_13803),
.B(n_13672),
.Y(n_14288)
);

INVx4_ASAP7_75t_L g14289 ( 
.A(n_14000),
.Y(n_14289)
);

INVx1_ASAP7_75t_L g14290 ( 
.A(n_13955),
.Y(n_14290)
);

AND2x2_ASAP7_75t_L g14291 ( 
.A(n_13825),
.B(n_13745),
.Y(n_14291)
);

AND2x2_ASAP7_75t_L g14292 ( 
.A(n_13831),
.B(n_13268),
.Y(n_14292)
);

HB1xp67_ASAP7_75t_L g14293 ( 
.A(n_13899),
.Y(n_14293)
);

AND2x2_ASAP7_75t_L g14294 ( 
.A(n_13910),
.B(n_9742),
.Y(n_14294)
);

INVx1_ASAP7_75t_L g14295 ( 
.A(n_13869),
.Y(n_14295)
);

INVx2_ASAP7_75t_L g14296 ( 
.A(n_13897),
.Y(n_14296)
);

INVx1_ASAP7_75t_L g14297 ( 
.A(n_13862),
.Y(n_14297)
);

NAND2xp5_ASAP7_75t_L g14298 ( 
.A(n_13841),
.B(n_10069),
.Y(n_14298)
);

INVx1_ASAP7_75t_L g14299 ( 
.A(n_13865),
.Y(n_14299)
);

AND2x2_ASAP7_75t_L g14300 ( 
.A(n_13847),
.B(n_9769),
.Y(n_14300)
);

OAI21xp5_ASAP7_75t_L g14301 ( 
.A1(n_13884),
.A2(n_13658),
.B(n_9769),
.Y(n_14301)
);

OR2x2_ASAP7_75t_L g14302 ( 
.A(n_13795),
.B(n_10075),
.Y(n_14302)
);

AND2x2_ASAP7_75t_L g14303 ( 
.A(n_14008),
.B(n_9449),
.Y(n_14303)
);

AND2x2_ASAP7_75t_L g14304 ( 
.A(n_13939),
.B(n_9449),
.Y(n_14304)
);

AND2x2_ASAP7_75t_L g14305 ( 
.A(n_13973),
.B(n_10188),
.Y(n_14305)
);

INVx2_ASAP7_75t_L g14306 ( 
.A(n_13881),
.Y(n_14306)
);

INVx1_ASAP7_75t_L g14307 ( 
.A(n_13786),
.Y(n_14307)
);

NAND2xp5_ASAP7_75t_L g14308 ( 
.A(n_13787),
.B(n_10075),
.Y(n_14308)
);

INVx4_ASAP7_75t_L g14309 ( 
.A(n_14182),
.Y(n_14309)
);

CKINVDCx5p33_ASAP7_75t_R g14310 ( 
.A(n_14139),
.Y(n_14310)
);

AND2x2_ASAP7_75t_L g14311 ( 
.A(n_14078),
.B(n_10188),
.Y(n_14311)
);

AOI22xp33_ASAP7_75t_L g14312 ( 
.A1(n_14054),
.A2(n_11152),
.B1(n_10092),
.B2(n_10081),
.Y(n_14312)
);

AND2x4_ASAP7_75t_L g14313 ( 
.A(n_14064),
.B(n_8203),
.Y(n_14313)
);

AND2x2_ASAP7_75t_L g14314 ( 
.A(n_13898),
.B(n_10193),
.Y(n_14314)
);

NAND2xp5_ASAP7_75t_L g14315 ( 
.A(n_13817),
.B(n_10076),
.Y(n_14315)
);

INVxp67_ASAP7_75t_SL g14316 ( 
.A(n_13846),
.Y(n_14316)
);

AND2x2_ASAP7_75t_L g14317 ( 
.A(n_13893),
.B(n_10193),
.Y(n_14317)
);

OAI22xp33_ASAP7_75t_L g14318 ( 
.A1(n_13919),
.A2(n_10081),
.B1(n_10076),
.B2(n_11196),
.Y(n_14318)
);

INVx2_ASAP7_75t_L g14319 ( 
.A(n_13909),
.Y(n_14319)
);

NAND2xp33_ASAP7_75t_R g14320 ( 
.A(n_13844),
.B(n_9363),
.Y(n_14320)
);

NOR2xp33_ASAP7_75t_L g14321 ( 
.A(n_13954),
.B(n_11197),
.Y(n_14321)
);

NOR2x1_ASAP7_75t_L g14322 ( 
.A(n_13888),
.B(n_13883),
.Y(n_14322)
);

INVx2_ASAP7_75t_L g14323 ( 
.A(n_14010),
.Y(n_14323)
);

BUFx12f_ASAP7_75t_L g14324 ( 
.A(n_13751),
.Y(n_14324)
);

OR2x2_ASAP7_75t_L g14325 ( 
.A(n_13917),
.B(n_8216),
.Y(n_14325)
);

INVx2_ASAP7_75t_L g14326 ( 
.A(n_14010),
.Y(n_14326)
);

AND2x2_ASAP7_75t_L g14327 ( 
.A(n_13971),
.B(n_10111),
.Y(n_14327)
);

INVx1_ASAP7_75t_L g14328 ( 
.A(n_13755),
.Y(n_14328)
);

NOR3xp33_ASAP7_75t_SL g14329 ( 
.A(n_13778),
.B(n_6829),
.C(n_8073),
.Y(n_14329)
);

NAND4xp25_ASAP7_75t_L g14330 ( 
.A(n_13785),
.B(n_8247),
.C(n_8117),
.D(n_8073),
.Y(n_14330)
);

AND2x2_ASAP7_75t_L g14331 ( 
.A(n_13977),
.B(n_10111),
.Y(n_14331)
);

INVx2_ASAP7_75t_L g14332 ( 
.A(n_13829),
.Y(n_14332)
);

AND2x2_ASAP7_75t_L g14333 ( 
.A(n_13920),
.B(n_10139),
.Y(n_14333)
);

INVx1_ASAP7_75t_L g14334 ( 
.A(n_13936),
.Y(n_14334)
);

INVx2_ASAP7_75t_L g14335 ( 
.A(n_13919),
.Y(n_14335)
);

NAND2xp5_ASAP7_75t_L g14336 ( 
.A(n_14188),
.B(n_8990),
.Y(n_14336)
);

INVx3_ASAP7_75t_SL g14337 ( 
.A(n_13948),
.Y(n_14337)
);

AND2x4_ASAP7_75t_L g14338 ( 
.A(n_13845),
.B(n_8203),
.Y(n_14338)
);

AND2x2_ASAP7_75t_L g14339 ( 
.A(n_13904),
.B(n_14135),
.Y(n_14339)
);

NOR2x1_ASAP7_75t_L g14340 ( 
.A(n_13816),
.B(n_9376),
.Y(n_14340)
);

NOR2x1_ASAP7_75t_L g14341 ( 
.A(n_13814),
.B(n_9376),
.Y(n_14341)
);

INVxp67_ASAP7_75t_SL g14342 ( 
.A(n_13807),
.Y(n_14342)
);

HB1xp67_ASAP7_75t_L g14343 ( 
.A(n_13844),
.Y(n_14343)
);

NAND4xp25_ASAP7_75t_SL g14344 ( 
.A(n_13999),
.B(n_6554),
.C(n_8223),
.D(n_8194),
.Y(n_14344)
);

NAND2xp5_ASAP7_75t_L g14345 ( 
.A(n_14086),
.B(n_8995),
.Y(n_14345)
);

INVx1_ASAP7_75t_L g14346 ( 
.A(n_13986),
.Y(n_14346)
);

OAI21xp33_ASAP7_75t_SL g14347 ( 
.A1(n_13756),
.A2(n_9932),
.B(n_10139),
.Y(n_14347)
);

AND2x4_ASAP7_75t_L g14348 ( 
.A(n_13916),
.B(n_13826),
.Y(n_14348)
);

OAI33xp33_ASAP7_75t_L g14349 ( 
.A1(n_13759),
.A2(n_9325),
.A3(n_9319),
.B1(n_9344),
.B2(n_9321),
.B3(n_9316),
.Y(n_14349)
);

NAND2xp5_ASAP7_75t_L g14350 ( 
.A(n_14037),
.B(n_8995),
.Y(n_14350)
);

AOI22xp33_ASAP7_75t_SL g14351 ( 
.A1(n_14111),
.A2(n_10067),
.B1(n_10059),
.B2(n_9431),
.Y(n_14351)
);

INVx1_ASAP7_75t_L g14352 ( 
.A(n_14162),
.Y(n_14352)
);

NAND2xp5_ASAP7_75t_L g14353 ( 
.A(n_14173),
.B(n_8996),
.Y(n_14353)
);

AND2x4_ASAP7_75t_SL g14354 ( 
.A(n_13914),
.B(n_7122),
.Y(n_14354)
);

NAND3xp33_ASAP7_75t_SL g14355 ( 
.A(n_13747),
.B(n_8893),
.C(n_9154),
.Y(n_14355)
);

INVx1_ASAP7_75t_L g14356 ( 
.A(n_13828),
.Y(n_14356)
);

INVxp67_ASAP7_75t_L g14357 ( 
.A(n_14185),
.Y(n_14357)
);

AND2x2_ASAP7_75t_L g14358 ( 
.A(n_13912),
.B(n_10145),
.Y(n_14358)
);

INVx1_ASAP7_75t_L g14359 ( 
.A(n_14036),
.Y(n_14359)
);

NAND2xp5_ASAP7_75t_L g14360 ( 
.A(n_13875),
.B(n_8996),
.Y(n_14360)
);

AND2x2_ASAP7_75t_L g14361 ( 
.A(n_13853),
.B(n_10145),
.Y(n_14361)
);

NAND2xp5_ASAP7_75t_L g14362 ( 
.A(n_14105),
.B(n_9002),
.Y(n_14362)
);

OR2x2_ASAP7_75t_L g14363 ( 
.A(n_13887),
.B(n_13890),
.Y(n_14363)
);

INVx2_ASAP7_75t_L g14364 ( 
.A(n_14041),
.Y(n_14364)
);

AND2x2_ASAP7_75t_L g14365 ( 
.A(n_13930),
.B(n_10162),
.Y(n_14365)
);

INVx1_ASAP7_75t_L g14366 ( 
.A(n_13840),
.Y(n_14366)
);

AND2x2_ASAP7_75t_L g14367 ( 
.A(n_13937),
.B(n_10162),
.Y(n_14367)
);

INVx1_ASAP7_75t_L g14368 ( 
.A(n_13994),
.Y(n_14368)
);

INVxp67_ASAP7_75t_L g14369 ( 
.A(n_13763),
.Y(n_14369)
);

AND2x2_ASAP7_75t_L g14370 ( 
.A(n_13935),
.B(n_9932),
.Y(n_14370)
);

INVx1_ASAP7_75t_L g14371 ( 
.A(n_13903),
.Y(n_14371)
);

OR2x2_ASAP7_75t_L g14372 ( 
.A(n_13799),
.B(n_8232),
.Y(n_14372)
);

NAND2xp5_ASAP7_75t_L g14373 ( 
.A(n_14155),
.B(n_9002),
.Y(n_14373)
);

AOI21xp5_ASAP7_75t_SL g14374 ( 
.A1(n_13768),
.A2(n_9431),
.B(n_9376),
.Y(n_14374)
);

AND2x2_ASAP7_75t_L g14375 ( 
.A(n_13940),
.B(n_9379),
.Y(n_14375)
);

AND2x2_ASAP7_75t_L g14376 ( 
.A(n_13894),
.B(n_9410),
.Y(n_14376)
);

AND2x2_ASAP7_75t_L g14377 ( 
.A(n_14144),
.B(n_9410),
.Y(n_14377)
);

AND2x2_ASAP7_75t_L g14378 ( 
.A(n_14146),
.B(n_9431),
.Y(n_14378)
);

AND2x4_ASAP7_75t_L g14379 ( 
.A(n_13804),
.B(n_9786),
.Y(n_14379)
);

INVx1_ASAP7_75t_L g14380 ( 
.A(n_14113),
.Y(n_14380)
);

INVx1_ASAP7_75t_L g14381 ( 
.A(n_13849),
.Y(n_14381)
);

NAND2xp5_ASAP7_75t_L g14382 ( 
.A(n_14025),
.B(n_9008),
.Y(n_14382)
);

NOR2xp33_ASAP7_75t_L g14383 ( 
.A(n_13848),
.B(n_10059),
.Y(n_14383)
);

INVx4_ASAP7_75t_L g14384 ( 
.A(n_13792),
.Y(n_14384)
);

INVx1_ASAP7_75t_SL g14385 ( 
.A(n_13798),
.Y(n_14385)
);

AND2x2_ASAP7_75t_L g14386 ( 
.A(n_14147),
.B(n_9431),
.Y(n_14386)
);

AND2x2_ASAP7_75t_L g14387 ( 
.A(n_13855),
.B(n_9788),
.Y(n_14387)
);

INVx1_ASAP7_75t_L g14388 ( 
.A(n_13850),
.Y(n_14388)
);

INVx3_ASAP7_75t_L g14389 ( 
.A(n_13901),
.Y(n_14389)
);

AND2x2_ASAP7_75t_L g14390 ( 
.A(n_13856),
.B(n_9788),
.Y(n_14390)
);

NAND2x1p5_ASAP7_75t_L g14391 ( 
.A(n_13861),
.B(n_8203),
.Y(n_14391)
);

AND2x2_ASAP7_75t_L g14392 ( 
.A(n_13872),
.B(n_9800),
.Y(n_14392)
);

AOI22xp33_ASAP7_75t_L g14393 ( 
.A1(n_13988),
.A2(n_13989),
.B1(n_13754),
.B2(n_13944),
.Y(n_14393)
);

NAND2xp5_ASAP7_75t_L g14394 ( 
.A(n_14104),
.B(n_9008),
.Y(n_14394)
);

AND2x4_ASAP7_75t_L g14395 ( 
.A(n_13854),
.B(n_9786),
.Y(n_14395)
);

INVx2_ASAP7_75t_L g14396 ( 
.A(n_14136),
.Y(n_14396)
);

INVx2_ASAP7_75t_L g14397 ( 
.A(n_14137),
.Y(n_14397)
);

INVx3_ASAP7_75t_L g14398 ( 
.A(n_14002),
.Y(n_14398)
);

OAI22xp5_ASAP7_75t_SL g14399 ( 
.A1(n_14123),
.A2(n_10067),
.B1(n_10059),
.B2(n_8893),
.Y(n_14399)
);

AND2x4_ASAP7_75t_L g14400 ( 
.A(n_13854),
.B(n_9891),
.Y(n_14400)
);

INVx2_ASAP7_75t_SL g14401 ( 
.A(n_13806),
.Y(n_14401)
);

AND2x2_ASAP7_75t_L g14402 ( 
.A(n_13782),
.B(n_9800),
.Y(n_14402)
);

INVx1_ASAP7_75t_SL g14403 ( 
.A(n_13791),
.Y(n_14403)
);

NOR3xp33_ASAP7_75t_L g14404 ( 
.A(n_13892),
.B(n_9891),
.C(n_10198),
.Y(n_14404)
);

AOI21xp5_ASAP7_75t_L g14405 ( 
.A1(n_13860),
.A2(n_10067),
.B(n_10217),
.Y(n_14405)
);

NOR3xp33_ASAP7_75t_L g14406 ( 
.A(n_14077),
.B(n_13876),
.C(n_13864),
.Y(n_14406)
);

OR2x2_ASAP7_75t_L g14407 ( 
.A(n_13821),
.B(n_8232),
.Y(n_14407)
);

OAI221xp5_ASAP7_75t_L g14408 ( 
.A1(n_14119),
.A2(n_10092),
.B1(n_8835),
.B2(n_8832),
.C(n_8827),
.Y(n_14408)
);

AND2x2_ASAP7_75t_L g14409 ( 
.A(n_13784),
.B(n_9518),
.Y(n_14409)
);

AND2x2_ASAP7_75t_L g14410 ( 
.A(n_13962),
.B(n_9518),
.Y(n_14410)
);

AND2x2_ASAP7_75t_L g14411 ( 
.A(n_13968),
.B(n_13998),
.Y(n_14411)
);

INVx1_ASAP7_75t_L g14412 ( 
.A(n_13750),
.Y(n_14412)
);

INVx1_ASAP7_75t_L g14413 ( 
.A(n_13896),
.Y(n_14413)
);

AND2x2_ASAP7_75t_L g14414 ( 
.A(n_14001),
.B(n_9528),
.Y(n_14414)
);

OR2x2_ASAP7_75t_L g14415 ( 
.A(n_14181),
.B(n_8246),
.Y(n_14415)
);

AND2x2_ASAP7_75t_L g14416 ( 
.A(n_14089),
.B(n_9528),
.Y(n_14416)
);

OAI31xp33_ASAP7_75t_L g14417 ( 
.A1(n_14156),
.A2(n_8832),
.A3(n_8835),
.B(n_9382),
.Y(n_14417)
);

NAND2xp5_ASAP7_75t_L g14418 ( 
.A(n_14194),
.B(n_9009),
.Y(n_14418)
);

INVx1_ASAP7_75t_L g14419 ( 
.A(n_13878),
.Y(n_14419)
);

INVx1_ASAP7_75t_L g14420 ( 
.A(n_14004),
.Y(n_14420)
);

INVx1_ASAP7_75t_L g14421 ( 
.A(n_13925),
.Y(n_14421)
);

INVx1_ASAP7_75t_L g14422 ( 
.A(n_13852),
.Y(n_14422)
);

INVx2_ASAP7_75t_L g14423 ( 
.A(n_13990),
.Y(n_14423)
);

AND2x2_ASAP7_75t_L g14424 ( 
.A(n_13913),
.B(n_9600),
.Y(n_14424)
);

NAND3xp33_ASAP7_75t_SL g14425 ( 
.A(n_13838),
.B(n_9158),
.C(n_9154),
.Y(n_14425)
);

INVx1_ASAP7_75t_L g14426 ( 
.A(n_14063),
.Y(n_14426)
);

INVx1_ASAP7_75t_L g14427 ( 
.A(n_14091),
.Y(n_14427)
);

OR2x2_ASAP7_75t_L g14428 ( 
.A(n_14076),
.B(n_14085),
.Y(n_14428)
);

OR2x2_ASAP7_75t_L g14429 ( 
.A(n_13809),
.B(n_8246),
.Y(n_14429)
);

INVx2_ASAP7_75t_L g14430 ( 
.A(n_13996),
.Y(n_14430)
);

INVx1_ASAP7_75t_L g14431 ( 
.A(n_14157),
.Y(n_14431)
);

AND2x2_ASAP7_75t_L g14432 ( 
.A(n_13796),
.B(n_9600),
.Y(n_14432)
);

INVx1_ASAP7_75t_L g14433 ( 
.A(n_14160),
.Y(n_14433)
);

INVx2_ASAP7_75t_L g14434 ( 
.A(n_13941),
.Y(n_14434)
);

BUFx2_ASAP7_75t_SL g14435 ( 
.A(n_14177),
.Y(n_14435)
);

HB1xp67_ASAP7_75t_L g14436 ( 
.A(n_14190),
.Y(n_14436)
);

INVx1_ASAP7_75t_L g14437 ( 
.A(n_14050),
.Y(n_14437)
);

OR2x2_ASAP7_75t_L g14438 ( 
.A(n_14053),
.B(n_8251),
.Y(n_14438)
);

OR2x6_ASAP7_75t_L g14439 ( 
.A(n_13900),
.B(n_8907),
.Y(n_14439)
);

INVx1_ASAP7_75t_L g14440 ( 
.A(n_14120),
.Y(n_14440)
);

AND2x2_ASAP7_75t_L g14441 ( 
.A(n_14140),
.B(n_9812),
.Y(n_14441)
);

NOR2xp33_ASAP7_75t_L g14442 ( 
.A(n_14056),
.B(n_9321),
.Y(n_14442)
);

AND2x2_ASAP7_75t_L g14443 ( 
.A(n_14165),
.B(n_9812),
.Y(n_14443)
);

INVx1_ASAP7_75t_SL g14444 ( 
.A(n_13827),
.Y(n_14444)
);

A2O1A1Ixp33_ASAP7_75t_L g14445 ( 
.A1(n_14168),
.A2(n_10202),
.B(n_10198),
.C(n_10217),
.Y(n_14445)
);

AND2x2_ASAP7_75t_L g14446 ( 
.A(n_13873),
.B(n_8928),
.Y(n_14446)
);

INVx2_ASAP7_75t_L g14447 ( 
.A(n_13941),
.Y(n_14447)
);

INVx1_ASAP7_75t_L g14448 ( 
.A(n_13749),
.Y(n_14448)
);

NOR3xp33_ASAP7_75t_L g14449 ( 
.A(n_13882),
.B(n_10202),
.C(n_8835),
.Y(n_14449)
);

AND2x2_ASAP7_75t_L g14450 ( 
.A(n_13992),
.B(n_8947),
.Y(n_14450)
);

AND2x2_ASAP7_75t_L g14451 ( 
.A(n_13993),
.B(n_10284),
.Y(n_14451)
);

AND2x2_ASAP7_75t_L g14452 ( 
.A(n_14087),
.B(n_10284),
.Y(n_14452)
);

OR2x2_ASAP7_75t_L g14453 ( 
.A(n_13815),
.B(n_8251),
.Y(n_14453)
);

OR2x2_ASAP7_75t_L g14454 ( 
.A(n_13819),
.B(n_8257),
.Y(n_14454)
);

AND2x4_ASAP7_75t_SL g14455 ( 
.A(n_14016),
.B(n_14003),
.Y(n_14455)
);

O2A1O1Ixp33_ASAP7_75t_L g14456 ( 
.A1(n_13835),
.A2(n_9382),
.B(n_9398),
.C(n_9395),
.Y(n_14456)
);

HB1xp67_ASAP7_75t_L g14457 ( 
.A(n_14002),
.Y(n_14457)
);

INVx1_ASAP7_75t_L g14458 ( 
.A(n_13774),
.Y(n_14458)
);

OR2x2_ASAP7_75t_L g14459 ( 
.A(n_14193),
.B(n_8257),
.Y(n_14459)
);

AND2x2_ASAP7_75t_L g14460 ( 
.A(n_14045),
.B(n_10299),
.Y(n_14460)
);

AND2x2_ASAP7_75t_L g14461 ( 
.A(n_13982),
.B(n_10299),
.Y(n_14461)
);

NAND2x1_ASAP7_75t_L g14462 ( 
.A(n_13775),
.B(n_7563),
.Y(n_14462)
);

NAND2xp5_ASAP7_75t_L g14463 ( 
.A(n_14179),
.B(n_9009),
.Y(n_14463)
);

INVx1_ASAP7_75t_L g14464 ( 
.A(n_14023),
.Y(n_14464)
);

OR2x2_ASAP7_75t_L g14465 ( 
.A(n_14116),
.B(n_8258),
.Y(n_14465)
);

INVx1_ASAP7_75t_L g14466 ( 
.A(n_13947),
.Y(n_14466)
);

INVx1_ASAP7_75t_L g14467 ( 
.A(n_13765),
.Y(n_14467)
);

AND2x2_ASAP7_75t_L g14468 ( 
.A(n_13983),
.B(n_10342),
.Y(n_14468)
);

INVx1_ASAP7_75t_L g14469 ( 
.A(n_13767),
.Y(n_14469)
);

INVx1_ASAP7_75t_L g14470 ( 
.A(n_14107),
.Y(n_14470)
);

BUFx2_ASAP7_75t_L g14471 ( 
.A(n_14067),
.Y(n_14471)
);

AND2x2_ASAP7_75t_L g14472 ( 
.A(n_14161),
.B(n_14133),
.Y(n_14472)
);

AND2x4_ASAP7_75t_L g14473 ( 
.A(n_13907),
.B(n_10342),
.Y(n_14473)
);

INVx1_ASAP7_75t_SL g14474 ( 
.A(n_13842),
.Y(n_14474)
);

OR2x2_ASAP7_75t_L g14475 ( 
.A(n_13867),
.B(n_8258),
.Y(n_14475)
);

NAND2xp5_ASAP7_75t_L g14476 ( 
.A(n_14038),
.B(n_9011),
.Y(n_14476)
);

OR2x2_ASAP7_75t_L g14477 ( 
.A(n_13874),
.B(n_8287),
.Y(n_14477)
);

AND2x2_ASAP7_75t_L g14478 ( 
.A(n_13980),
.B(n_10343),
.Y(n_14478)
);

HB1xp67_ASAP7_75t_L g14479 ( 
.A(n_13963),
.Y(n_14479)
);

AND2x2_ASAP7_75t_L g14480 ( 
.A(n_14080),
.B(n_10343),
.Y(n_14480)
);

OR2x2_ASAP7_75t_L g14481 ( 
.A(n_13981),
.B(n_8287),
.Y(n_14481)
);

OR2x2_ASAP7_75t_L g14482 ( 
.A(n_14029),
.B(n_8194),
.Y(n_14482)
);

AND2x2_ASAP7_75t_L g14483 ( 
.A(n_14014),
.B(n_10357),
.Y(n_14483)
);

HB1xp67_ASAP7_75t_L g14484 ( 
.A(n_13991),
.Y(n_14484)
);

OR2x2_ASAP7_75t_L g14485 ( 
.A(n_14103),
.B(n_8194),
.Y(n_14485)
);

INVx1_ASAP7_75t_L g14486 ( 
.A(n_14125),
.Y(n_14486)
);

O2A1O1Ixp33_ASAP7_75t_SL g14487 ( 
.A1(n_13877),
.A2(n_9344),
.B(n_9345),
.C(n_9325),
.Y(n_14487)
);

AND2x2_ASAP7_75t_L g14488 ( 
.A(n_14034),
.B(n_10357),
.Y(n_14488)
);

AND2x2_ASAP7_75t_L g14489 ( 
.A(n_13943),
.B(n_10375),
.Y(n_14489)
);

INVx1_ASAP7_75t_L g14490 ( 
.A(n_14102),
.Y(n_14490)
);

INVx1_ASAP7_75t_SL g14491 ( 
.A(n_14028),
.Y(n_14491)
);

AND2x2_ASAP7_75t_L g14492 ( 
.A(n_13870),
.B(n_10375),
.Y(n_14492)
);

INVx4_ASAP7_75t_L g14493 ( 
.A(n_14122),
.Y(n_14493)
);

NAND2xp5_ASAP7_75t_L g14494 ( 
.A(n_14075),
.B(n_9011),
.Y(n_14494)
);

AOI22xp33_ASAP7_75t_L g14495 ( 
.A1(n_13830),
.A2(n_10092),
.B1(n_9398),
.B2(n_9402),
.Y(n_14495)
);

INVx4_ASAP7_75t_L g14496 ( 
.A(n_14127),
.Y(n_14496)
);

INVx3_ASAP7_75t_L g14497 ( 
.A(n_14017),
.Y(n_14497)
);

INVx1_ASAP7_75t_SL g14498 ( 
.A(n_14115),
.Y(n_14498)
);

AND2x2_ASAP7_75t_L g14499 ( 
.A(n_14051),
.B(n_10376),
.Y(n_14499)
);

HB1xp67_ASAP7_75t_L g14500 ( 
.A(n_14143),
.Y(n_14500)
);

NAND2xp33_ASAP7_75t_SL g14501 ( 
.A(n_14032),
.B(n_6547),
.Y(n_14501)
);

INVx1_ASAP7_75t_L g14502 ( 
.A(n_14055),
.Y(n_14502)
);

NAND2xp5_ASAP7_75t_L g14503 ( 
.A(n_14052),
.B(n_9017),
.Y(n_14503)
);

NAND2x1p5_ASAP7_75t_L g14504 ( 
.A(n_14092),
.B(n_8206),
.Y(n_14504)
);

AND2x2_ASAP7_75t_SL g14505 ( 
.A(n_13885),
.B(n_7181),
.Y(n_14505)
);

NOR2x1_ASAP7_75t_L g14506 ( 
.A(n_13866),
.B(n_9345),
.Y(n_14506)
);

INVx2_ASAP7_75t_L g14507 ( 
.A(n_14013),
.Y(n_14507)
);

BUFx2_ASAP7_75t_L g14508 ( 
.A(n_13975),
.Y(n_14508)
);

NAND2x1p5_ASAP7_75t_L g14509 ( 
.A(n_14057),
.B(n_8206),
.Y(n_14509)
);

AND2x2_ASAP7_75t_L g14510 ( 
.A(n_14059),
.B(n_10376),
.Y(n_14510)
);

OAI211xp5_ASAP7_75t_SL g14511 ( 
.A1(n_14130),
.A2(n_8206),
.B(n_8279),
.C(n_8247),
.Y(n_14511)
);

AND2x2_ASAP7_75t_L g14512 ( 
.A(n_14060),
.B(n_9348),
.Y(n_14512)
);

NOR2xp33_ASAP7_75t_R g14513 ( 
.A(n_14065),
.B(n_6547),
.Y(n_14513)
);

INVx2_ASAP7_75t_L g14514 ( 
.A(n_14039),
.Y(n_14514)
);

OR2x2_ASAP7_75t_L g14515 ( 
.A(n_14081),
.B(n_8223),
.Y(n_14515)
);

AND2x2_ASAP7_75t_L g14516 ( 
.A(n_14117),
.B(n_9348),
.Y(n_14516)
);

INVx1_ASAP7_75t_L g14517 ( 
.A(n_14072),
.Y(n_14517)
);

INVx1_ASAP7_75t_L g14518 ( 
.A(n_14180),
.Y(n_14518)
);

CKINVDCx5p33_ASAP7_75t_R g14519 ( 
.A(n_14170),
.Y(n_14519)
);

INVx1_ASAP7_75t_SL g14520 ( 
.A(n_14108),
.Y(n_14520)
);

INVx4_ASAP7_75t_L g14521 ( 
.A(n_14068),
.Y(n_14521)
);

NOR3xp33_ASAP7_75t_SL g14522 ( 
.A(n_14027),
.B(n_8117),
.C(n_6554),
.Y(n_14522)
);

AND2x2_ASAP7_75t_L g14523 ( 
.A(n_14142),
.B(n_9352),
.Y(n_14523)
);

AND2x2_ASAP7_75t_L g14524 ( 
.A(n_14148),
.B(n_9352),
.Y(n_14524)
);

AND2x4_ASAP7_75t_L g14525 ( 
.A(n_13921),
.B(n_8206),
.Y(n_14525)
);

AND2x4_ASAP7_75t_L g14526 ( 
.A(n_13923),
.B(n_8206),
.Y(n_14526)
);

AND2x2_ASAP7_75t_L g14527 ( 
.A(n_14151),
.B(n_9357),
.Y(n_14527)
);

INVxp67_ASAP7_75t_L g14528 ( 
.A(n_13960),
.Y(n_14528)
);

OR2x2_ASAP7_75t_L g14529 ( 
.A(n_14094),
.B(n_8223),
.Y(n_14529)
);

AND2x2_ASAP7_75t_L g14530 ( 
.A(n_14159),
.B(n_9357),
.Y(n_14530)
);

INVx1_ASAP7_75t_L g14531 ( 
.A(n_14112),
.Y(n_14531)
);

AND2x2_ASAP7_75t_SL g14532 ( 
.A(n_14100),
.B(n_7181),
.Y(n_14532)
);

OAI21xp33_ASAP7_75t_L g14533 ( 
.A1(n_14110),
.A2(n_7956),
.B(n_7953),
.Y(n_14533)
);

NOR2xp33_ASAP7_75t_L g14534 ( 
.A(n_13946),
.B(n_9359),
.Y(n_14534)
);

INVx1_ASAP7_75t_L g14535 ( 
.A(n_14126),
.Y(n_14535)
);

AND2x2_ASAP7_75t_L g14536 ( 
.A(n_14098),
.B(n_9359),
.Y(n_14536)
);

HB1xp67_ASAP7_75t_L g14537 ( 
.A(n_14031),
.Y(n_14537)
);

AND2x2_ASAP7_75t_L g14538 ( 
.A(n_14043),
.B(n_9360),
.Y(n_14538)
);

AND2x2_ASAP7_75t_L g14539 ( 
.A(n_14129),
.B(n_9360),
.Y(n_14539)
);

INVx1_ASAP7_75t_L g14540 ( 
.A(n_14169),
.Y(n_14540)
);

INVx1_ASAP7_75t_L g14541 ( 
.A(n_14176),
.Y(n_14541)
);

INVx1_ASAP7_75t_L g14542 ( 
.A(n_13918),
.Y(n_14542)
);

NAND2xp5_ASAP7_75t_L g14543 ( 
.A(n_14040),
.B(n_9017),
.Y(n_14543)
);

NOR2xp67_ASAP7_75t_L g14544 ( 
.A(n_14128),
.B(n_9027),
.Y(n_14544)
);

INVx1_ASAP7_75t_L g14545 ( 
.A(n_13929),
.Y(n_14545)
);

NOR2xp33_ASAP7_75t_L g14546 ( 
.A(n_14033),
.B(n_9370),
.Y(n_14546)
);

INVx1_ASAP7_75t_L g14547 ( 
.A(n_13932),
.Y(n_14547)
);

INVx3_ASAP7_75t_L g14548 ( 
.A(n_14017),
.Y(n_14548)
);

INVx1_ASAP7_75t_L g14549 ( 
.A(n_13949),
.Y(n_14549)
);

OAI221xp5_ASAP7_75t_L g14550 ( 
.A1(n_14005),
.A2(n_9407),
.B1(n_9413),
.B2(n_9402),
.C(n_9395),
.Y(n_14550)
);

AND2x2_ASAP7_75t_SL g14551 ( 
.A(n_13924),
.B(n_7181),
.Y(n_14551)
);

AOI22xp33_ASAP7_75t_L g14552 ( 
.A1(n_13871),
.A2(n_9407),
.B1(n_9413),
.B2(n_9402),
.Y(n_14552)
);

AND2x4_ASAP7_75t_L g14553 ( 
.A(n_13927),
.B(n_8279),
.Y(n_14553)
);

HB1xp67_ASAP7_75t_L g14554 ( 
.A(n_14024),
.Y(n_14554)
);

INVx1_ASAP7_75t_L g14555 ( 
.A(n_13969),
.Y(n_14555)
);

INVx1_ASAP7_75t_L g14556 ( 
.A(n_13972),
.Y(n_14556)
);

AND2x2_ASAP7_75t_L g14557 ( 
.A(n_14174),
.B(n_9370),
.Y(n_14557)
);

AND2x2_ASAP7_75t_L g14558 ( 
.A(n_14047),
.B(n_9371),
.Y(n_14558)
);

HB1xp67_ASAP7_75t_L g14559 ( 
.A(n_14024),
.Y(n_14559)
);

AND2x2_ASAP7_75t_L g14560 ( 
.A(n_14048),
.B(n_9371),
.Y(n_14560)
);

NOR2xp33_ASAP7_75t_L g14561 ( 
.A(n_14062),
.B(n_9384),
.Y(n_14561)
);

OAI33xp33_ASAP7_75t_L g14562 ( 
.A1(n_13868),
.A2(n_9400),
.A3(n_9393),
.B1(n_9401),
.B2(n_9394),
.B3(n_9384),
.Y(n_14562)
);

OR2x2_ASAP7_75t_L g14563 ( 
.A(n_13938),
.B(n_8250),
.Y(n_14563)
);

NAND2xp5_ASAP7_75t_L g14564 ( 
.A(n_14141),
.B(n_9027),
.Y(n_14564)
);

INVx4_ASAP7_75t_L g14565 ( 
.A(n_13956),
.Y(n_14565)
);

AND2x2_ASAP7_75t_L g14566 ( 
.A(n_14049),
.B(n_9393),
.Y(n_14566)
);

INVx2_ASAP7_75t_L g14567 ( 
.A(n_14192),
.Y(n_14567)
);

INVx1_ASAP7_75t_SL g14568 ( 
.A(n_14009),
.Y(n_14568)
);

NOR2xp33_ASAP7_75t_L g14569 ( 
.A(n_14145),
.B(n_9394),
.Y(n_14569)
);

AND2x2_ASAP7_75t_L g14570 ( 
.A(n_14109),
.B(n_9400),
.Y(n_14570)
);

AND2x2_ASAP7_75t_L g14571 ( 
.A(n_14114),
.B(n_9401),
.Y(n_14571)
);

AND2x2_ASAP7_75t_L g14572 ( 
.A(n_13945),
.B(n_9404),
.Y(n_14572)
);

NAND2x1p5_ASAP7_75t_L g14573 ( 
.A(n_13957),
.B(n_8279),
.Y(n_14573)
);

AND2x4_ASAP7_75t_SL g14574 ( 
.A(n_13964),
.B(n_7123),
.Y(n_14574)
);

NAND2xp5_ASAP7_75t_L g14575 ( 
.A(n_14101),
.B(n_9031),
.Y(n_14575)
);

BUFx3_ASAP7_75t_L g14576 ( 
.A(n_13966),
.Y(n_14576)
);

AND2x2_ASAP7_75t_L g14577 ( 
.A(n_14079),
.B(n_9404),
.Y(n_14577)
);

INVx1_ASAP7_75t_L g14578 ( 
.A(n_14012),
.Y(n_14578)
);

INVx1_ASAP7_75t_L g14579 ( 
.A(n_14044),
.Y(n_14579)
);

INVx1_ASAP7_75t_L g14580 ( 
.A(n_14186),
.Y(n_14580)
);

AND2x2_ASAP7_75t_L g14581 ( 
.A(n_14083),
.B(n_9408),
.Y(n_14581)
);

OR2x2_ASAP7_75t_L g14582 ( 
.A(n_13958),
.B(n_8250),
.Y(n_14582)
);

OR2x2_ASAP7_75t_L g14583 ( 
.A(n_14042),
.B(n_8250),
.Y(n_14583)
);

AND2x2_ASAP7_75t_L g14584 ( 
.A(n_14095),
.B(n_9408),
.Y(n_14584)
);

NAND3xp33_ASAP7_75t_SL g14585 ( 
.A(n_14166),
.B(n_9158),
.C(n_9154),
.Y(n_14585)
);

AND2x2_ASAP7_75t_L g14586 ( 
.A(n_14097),
.B(n_9414),
.Y(n_14586)
);

AOI322xp5_ASAP7_75t_L g14587 ( 
.A1(n_14134),
.A2(n_9413),
.A3(n_9415),
.B1(n_9436),
.B2(n_9422),
.C1(n_9407),
.C2(n_9302),
.Y(n_14587)
);

AND2x2_ASAP7_75t_L g14588 ( 
.A(n_13942),
.B(n_9414),
.Y(n_14588)
);

OR2x2_ASAP7_75t_L g14589 ( 
.A(n_14020),
.B(n_8268),
.Y(n_14589)
);

NAND2xp5_ASAP7_75t_L g14590 ( 
.A(n_14101),
.B(n_9031),
.Y(n_14590)
);

OR2x2_ASAP7_75t_L g14591 ( 
.A(n_14153),
.B(n_8268),
.Y(n_14591)
);

INVx1_ASAP7_75t_L g14592 ( 
.A(n_14187),
.Y(n_14592)
);

OR2x2_ASAP7_75t_L g14593 ( 
.A(n_14154),
.B(n_8268),
.Y(n_14593)
);

AND2x4_ASAP7_75t_L g14594 ( 
.A(n_14088),
.B(n_8279),
.Y(n_14594)
);

HB1xp67_ASAP7_75t_L g14595 ( 
.A(n_14164),
.Y(n_14595)
);

INVx1_ASAP7_75t_L g14596 ( 
.A(n_14189),
.Y(n_14596)
);

INVx2_ASAP7_75t_SL g14597 ( 
.A(n_14070),
.Y(n_14597)
);

INVx2_ASAP7_75t_L g14598 ( 
.A(n_14171),
.Y(n_14598)
);

INVx1_ASAP7_75t_L g14599 ( 
.A(n_14158),
.Y(n_14599)
);

NAND2xp5_ASAP7_75t_L g14600 ( 
.A(n_13928),
.B(n_9033),
.Y(n_14600)
);

OR2x2_ASAP7_75t_L g14601 ( 
.A(n_14019),
.B(n_7953),
.Y(n_14601)
);

INVxp67_ASAP7_75t_SL g14602 ( 
.A(n_13934),
.Y(n_14602)
);

OR2x2_ASAP7_75t_L g14603 ( 
.A(n_14058),
.B(n_13908),
.Y(n_14603)
);

OR2x2_ASAP7_75t_L g14604 ( 
.A(n_13915),
.B(n_7956),
.Y(n_14604)
);

OR2x2_ASAP7_75t_L g14605 ( 
.A(n_13950),
.B(n_7992),
.Y(n_14605)
);

AND2x2_ASAP7_75t_L g14606 ( 
.A(n_14022),
.B(n_14069),
.Y(n_14606)
);

INVx2_ASAP7_75t_SL g14607 ( 
.A(n_13931),
.Y(n_14607)
);

NAND2xp5_ASAP7_75t_L g14608 ( 
.A(n_14172),
.B(n_9033),
.Y(n_14608)
);

NOR2xp33_ASAP7_75t_L g14609 ( 
.A(n_14106),
.B(n_9417),
.Y(n_14609)
);

OR2x2_ASAP7_75t_L g14610 ( 
.A(n_14225),
.B(n_14337),
.Y(n_14610)
);

INVxp67_ASAP7_75t_L g14611 ( 
.A(n_14435),
.Y(n_14611)
);

NAND2xp5_ASAP7_75t_L g14612 ( 
.A(n_14310),
.B(n_14343),
.Y(n_14612)
);

OR2x2_ASAP7_75t_L g14613 ( 
.A(n_14205),
.B(n_13995),
.Y(n_14613)
);

INVx2_ASAP7_75t_SL g14614 ( 
.A(n_14282),
.Y(n_14614)
);

INVxp67_ASAP7_75t_L g14615 ( 
.A(n_14203),
.Y(n_14615)
);

NAND2xp5_ASAP7_75t_L g14616 ( 
.A(n_14199),
.B(n_14121),
.Y(n_14616)
);

INVx1_ASAP7_75t_L g14617 ( 
.A(n_14238),
.Y(n_14617)
);

INVx3_ASAP7_75t_L g14618 ( 
.A(n_14289),
.Y(n_14618)
);

NAND2xp5_ASAP7_75t_L g14619 ( 
.A(n_14208),
.B(n_14235),
.Y(n_14619)
);

INVx1_ASAP7_75t_L g14620 ( 
.A(n_14238),
.Y(n_14620)
);

INVx2_ASAP7_75t_L g14621 ( 
.A(n_14255),
.Y(n_14621)
);

AOI22xp5_ASAP7_75t_L g14622 ( 
.A1(n_14269),
.A2(n_14131),
.B1(n_14150),
.B2(n_14149),
.Y(n_14622)
);

INVx2_ASAP7_75t_L g14623 ( 
.A(n_14260),
.Y(n_14623)
);

INVx1_ASAP7_75t_L g14624 ( 
.A(n_14363),
.Y(n_14624)
);

INVx1_ASAP7_75t_L g14625 ( 
.A(n_14239),
.Y(n_14625)
);

NOR2xp33_ASAP7_75t_L g14626 ( 
.A(n_14324),
.B(n_14124),
.Y(n_14626)
);

AND2x2_ASAP7_75t_L g14627 ( 
.A(n_14196),
.B(n_14152),
.Y(n_14627)
);

INVx1_ASAP7_75t_L g14628 ( 
.A(n_14232),
.Y(n_14628)
);

NOR2xp33_ASAP7_75t_L g14629 ( 
.A(n_14282),
.B(n_14132),
.Y(n_14629)
);

INVx1_ASAP7_75t_SL g14630 ( 
.A(n_14292),
.Y(n_14630)
);

OR2x2_ASAP7_75t_L g14631 ( 
.A(n_14385),
.B(n_14021),
.Y(n_14631)
);

NAND2xp5_ASAP7_75t_L g14632 ( 
.A(n_14278),
.B(n_14030),
.Y(n_14632)
);

AND2x4_ASAP7_75t_L g14633 ( 
.A(n_14214),
.B(n_14073),
.Y(n_14633)
);

INVx1_ASAP7_75t_L g14634 ( 
.A(n_14284),
.Y(n_14634)
);

OR3x2_ASAP7_75t_L g14635 ( 
.A(n_14229),
.B(n_14184),
.C(n_14163),
.Y(n_14635)
);

A2O1A1Ixp33_ASAP7_75t_L g14636 ( 
.A1(n_14281),
.A2(n_14138),
.B(n_14093),
.C(n_14096),
.Y(n_14636)
);

NAND2x1p5_ASAP7_75t_L g14637 ( 
.A(n_14219),
.B(n_14191),
.Y(n_14637)
);

OAI32xp33_ASAP7_75t_L g14638 ( 
.A1(n_14201),
.A2(n_13974),
.A3(n_13984),
.B1(n_13970),
.B2(n_13967),
.Y(n_14638)
);

NAND2xp5_ASAP7_75t_L g14639 ( 
.A(n_14444),
.B(n_13905),
.Y(n_14639)
);

INVx1_ASAP7_75t_L g14640 ( 
.A(n_14280),
.Y(n_14640)
);

AOI211xp5_ASAP7_75t_SL g14641 ( 
.A1(n_14197),
.A2(n_14082),
.B(n_13987),
.C(n_13965),
.Y(n_14641)
);

AND2x2_ASAP7_75t_L g14642 ( 
.A(n_14198),
.B(n_14011),
.Y(n_14642)
);

INVx1_ASAP7_75t_L g14643 ( 
.A(n_14280),
.Y(n_14643)
);

INVx1_ASAP7_75t_L g14644 ( 
.A(n_14280),
.Y(n_14644)
);

NAND2x2_ASAP7_75t_L g14645 ( 
.A(n_14401),
.B(n_14015),
.Y(n_14645)
);

INVx2_ASAP7_75t_L g14646 ( 
.A(n_14251),
.Y(n_14646)
);

INVx1_ASAP7_75t_L g14647 ( 
.A(n_14230),
.Y(n_14647)
);

CKINVDCx16_ASAP7_75t_R g14648 ( 
.A(n_14275),
.Y(n_14648)
);

OR2x2_ASAP7_75t_L g14649 ( 
.A(n_14403),
.B(n_14175),
.Y(n_14649)
);

INVx1_ASAP7_75t_L g14650 ( 
.A(n_14263),
.Y(n_14650)
);

AND2x2_ASAP7_75t_L g14651 ( 
.A(n_14233),
.B(n_14257),
.Y(n_14651)
);

INVx1_ASAP7_75t_L g14652 ( 
.A(n_14457),
.Y(n_14652)
);

NAND2xp5_ASAP7_75t_L g14653 ( 
.A(n_14285),
.B(n_13961),
.Y(n_14653)
);

AND2x4_ASAP7_75t_L g14654 ( 
.A(n_14242),
.B(n_14204),
.Y(n_14654)
);

HB1xp67_ASAP7_75t_L g14655 ( 
.A(n_14213),
.Y(n_14655)
);

NAND2xp5_ASAP7_75t_L g14656 ( 
.A(n_14286),
.B(n_14290),
.Y(n_14656)
);

INVx1_ASAP7_75t_L g14657 ( 
.A(n_14234),
.Y(n_14657)
);

NAND2xp5_ASAP7_75t_L g14658 ( 
.A(n_14520),
.B(n_14244),
.Y(n_14658)
);

INVx1_ASAP7_75t_L g14659 ( 
.A(n_14243),
.Y(n_14659)
);

AND2x4_ASAP7_75t_L g14660 ( 
.A(n_14335),
.B(n_8817),
.Y(n_14660)
);

NAND2xp5_ASAP7_75t_L g14661 ( 
.A(n_14247),
.B(n_9417),
.Y(n_14661)
);

OR2x2_ASAP7_75t_L g14662 ( 
.A(n_14474),
.B(n_7992),
.Y(n_14662)
);

NAND3xp33_ASAP7_75t_L g14663 ( 
.A(n_14206),
.B(n_7220),
.C(n_7181),
.Y(n_14663)
);

INVx1_ASAP7_75t_L g14664 ( 
.A(n_14210),
.Y(n_14664)
);

OAI33xp33_ASAP7_75t_L g14665 ( 
.A1(n_14195),
.A2(n_9427),
.A3(n_9425),
.B1(n_9433),
.B2(n_9426),
.B3(n_9424),
.Y(n_14665)
);

INVx1_ASAP7_75t_L g14666 ( 
.A(n_14218),
.Y(n_14666)
);

INVx1_ASAP7_75t_L g14667 ( 
.A(n_14253),
.Y(n_14667)
);

OAI22xp5_ASAP7_75t_L g14668 ( 
.A1(n_14413),
.A2(n_9425),
.B1(n_9426),
.B2(n_9424),
.Y(n_14668)
);

INVx1_ASAP7_75t_L g14669 ( 
.A(n_14220),
.Y(n_14669)
);

INVx1_ASAP7_75t_L g14670 ( 
.A(n_14223),
.Y(n_14670)
);

OA222x2_ASAP7_75t_L g14671 ( 
.A1(n_14202),
.A2(n_8279),
.B1(n_6271),
.B2(n_9302),
.C1(n_9324),
.C2(n_9300),
.Y(n_14671)
);

INVx1_ASAP7_75t_SL g14672 ( 
.A(n_14248),
.Y(n_14672)
);

OAI22xp33_ASAP7_75t_L g14673 ( 
.A1(n_14320),
.A2(n_9422),
.B1(n_9436),
.B2(n_9415),
.Y(n_14673)
);

INVx2_ASAP7_75t_L g14674 ( 
.A(n_14211),
.Y(n_14674)
);

AND2x4_ASAP7_75t_L g14675 ( 
.A(n_14348),
.B(n_8817),
.Y(n_14675)
);

INVx2_ASAP7_75t_L g14676 ( 
.A(n_14309),
.Y(n_14676)
);

INVx1_ASAP7_75t_L g14677 ( 
.A(n_14293),
.Y(n_14677)
);

INVx1_ASAP7_75t_L g14678 ( 
.A(n_14209),
.Y(n_14678)
);

AOI32xp33_ASAP7_75t_L g14679 ( 
.A1(n_14341),
.A2(n_8858),
.A3(n_8819),
.B1(n_7484),
.B2(n_7343),
.Y(n_14679)
);

O2A1O1Ixp5_ASAP7_75t_R g14680 ( 
.A1(n_14249),
.A2(n_7139),
.B(n_7125),
.C(n_6916),
.Y(n_14680)
);

INVx2_ASAP7_75t_L g14681 ( 
.A(n_14391),
.Y(n_14681)
);

INVx1_ASAP7_75t_L g14682 ( 
.A(n_14212),
.Y(n_14682)
);

NAND2x1_ASAP7_75t_L g14683 ( 
.A(n_14398),
.B(n_7563),
.Y(n_14683)
);

AOI22xp33_ASAP7_75t_L g14684 ( 
.A1(n_14279),
.A2(n_9422),
.B1(n_9436),
.B2(n_9415),
.Y(n_14684)
);

OAI33xp33_ASAP7_75t_L g14685 ( 
.A1(n_14236),
.A2(n_9433),
.A3(n_9435),
.B1(n_9427),
.B2(n_9057),
.B3(n_9040),
.Y(n_14685)
);

AOI22xp33_ASAP7_75t_L g14686 ( 
.A1(n_14312),
.A2(n_7220),
.B1(n_7443),
.B2(n_9300),
.Y(n_14686)
);

OR2x2_ASAP7_75t_L g14687 ( 
.A(n_14221),
.B(n_9435),
.Y(n_14687)
);

OAI22xp33_ASAP7_75t_L g14688 ( 
.A1(n_14537),
.A2(n_14568),
.B1(n_14319),
.B2(n_14428),
.Y(n_14688)
);

NAND4xp75_ASAP7_75t_L g14689 ( 
.A(n_14322),
.B(n_7498),
.C(n_8043),
.D(n_8032),
.Y(n_14689)
);

CKINVDCx5p33_ASAP7_75t_R g14690 ( 
.A(n_14519),
.Y(n_14690)
);

INVx1_ASAP7_75t_L g14691 ( 
.A(n_14500),
.Y(n_14691)
);

INVx1_ASAP7_75t_L g14692 ( 
.A(n_14271),
.Y(n_14692)
);

INVx2_ASAP7_75t_L g14693 ( 
.A(n_14508),
.Y(n_14693)
);

A2O1A1Ixp33_ASAP7_75t_L g14694 ( 
.A1(n_14383),
.A2(n_7224),
.B(n_7241),
.C(n_7167),
.Y(n_14694)
);

OR2x6_ASAP7_75t_L g14695 ( 
.A(n_14306),
.B(n_8912),
.Y(n_14695)
);

OR2x2_ASAP7_75t_L g14696 ( 
.A(n_14272),
.B(n_9037),
.Y(n_14696)
);

INVx1_ASAP7_75t_L g14697 ( 
.A(n_14266),
.Y(n_14697)
);

INVx1_ASAP7_75t_L g14698 ( 
.A(n_14231),
.Y(n_14698)
);

AND2x4_ASAP7_75t_L g14699 ( 
.A(n_14323),
.B(n_14326),
.Y(n_14699)
);

INVx2_ASAP7_75t_SL g14700 ( 
.A(n_14455),
.Y(n_14700)
);

AND2x2_ASAP7_75t_L g14701 ( 
.A(n_14332),
.B(n_9037),
.Y(n_14701)
);

AND2x2_ASAP7_75t_L g14702 ( 
.A(n_14411),
.B(n_9040),
.Y(n_14702)
);

INVx2_ASAP7_75t_L g14703 ( 
.A(n_14508),
.Y(n_14703)
);

NAND2xp5_ASAP7_75t_L g14704 ( 
.A(n_14342),
.B(n_9324),
.Y(n_14704)
);

AOI22xp5_ASAP7_75t_L g14705 ( 
.A1(n_14347),
.A2(n_7220),
.B1(n_7443),
.B2(n_7284),
.Y(n_14705)
);

INVx1_ASAP7_75t_L g14706 ( 
.A(n_14554),
.Y(n_14706)
);

INVx2_ASAP7_75t_SL g14707 ( 
.A(n_14273),
.Y(n_14707)
);

OAI31xp33_ASAP7_75t_L g14708 ( 
.A1(n_14436),
.A2(n_9158),
.A3(n_9223),
.B(n_9171),
.Y(n_14708)
);

NOR2xp33_ASAP7_75t_L g14709 ( 
.A(n_14565),
.B(n_14521),
.Y(n_14709)
);

NAND2xp5_ASAP7_75t_L g14710 ( 
.A(n_14366),
.B(n_9052),
.Y(n_14710)
);

O2A1O1Ixp33_ASAP7_75t_L g14711 ( 
.A1(n_14237),
.A2(n_7220),
.B(n_7443),
.C(n_7618),
.Y(n_14711)
);

AOI32xp33_ASAP7_75t_L g14712 ( 
.A1(n_14340),
.A2(n_8858),
.A3(n_8819),
.B1(n_7484),
.B2(n_7343),
.Y(n_14712)
);

OA222x2_ASAP7_75t_L g14713 ( 
.A1(n_14576),
.A2(n_6271),
.B1(n_9058),
.B2(n_9062),
.C1(n_9057),
.C2(n_9052),
.Y(n_14713)
);

INVx2_ASAP7_75t_L g14714 ( 
.A(n_14215),
.Y(n_14714)
);

NAND2xp5_ASAP7_75t_L g14715 ( 
.A(n_14261),
.B(n_9058),
.Y(n_14715)
);

NAND2xp5_ASAP7_75t_L g14716 ( 
.A(n_14498),
.B(n_9062),
.Y(n_14716)
);

INVx1_ASAP7_75t_L g14717 ( 
.A(n_14559),
.Y(n_14717)
);

AND2x2_ASAP7_75t_L g14718 ( 
.A(n_14339),
.B(n_9068),
.Y(n_14718)
);

AND2x2_ASAP7_75t_L g14719 ( 
.A(n_14268),
.B(n_9068),
.Y(n_14719)
);

AND2x2_ASAP7_75t_L g14720 ( 
.A(n_14291),
.B(n_9072),
.Y(n_14720)
);

OAI211xp5_ASAP7_75t_L g14721 ( 
.A1(n_14283),
.A2(n_7460),
.B(n_6197),
.C(n_9280),
.Y(n_14721)
);

INVx1_ASAP7_75t_L g14722 ( 
.A(n_14352),
.Y(n_14722)
);

INVx1_ASAP7_75t_L g14723 ( 
.A(n_14267),
.Y(n_14723)
);

OAI33xp33_ASAP7_75t_L g14724 ( 
.A1(n_14226),
.A2(n_9080),
.A3(n_9073),
.B1(n_9084),
.B2(n_9076),
.B3(n_9072),
.Y(n_14724)
);

INVx3_ASAP7_75t_L g14725 ( 
.A(n_14384),
.Y(n_14725)
);

AND2x2_ASAP7_75t_L g14726 ( 
.A(n_14250),
.B(n_9073),
.Y(n_14726)
);

NAND2x2_ASAP7_75t_L g14727 ( 
.A(n_14597),
.B(n_6706),
.Y(n_14727)
);

INVx1_ASAP7_75t_L g14728 ( 
.A(n_14316),
.Y(n_14728)
);

OAI33xp33_ASAP7_75t_L g14729 ( 
.A1(n_14227),
.A2(n_9086),
.A3(n_9080),
.B1(n_9088),
.B2(n_9084),
.B3(n_9076),
.Y(n_14729)
);

OAI31xp33_ASAP7_75t_L g14730 ( 
.A1(n_14440),
.A2(n_9171),
.A3(n_9223),
.B(n_8168),
.Y(n_14730)
);

INVx1_ASAP7_75t_L g14731 ( 
.A(n_14241),
.Y(n_14731)
);

INVx1_ASAP7_75t_SL g14732 ( 
.A(n_14228),
.Y(n_14732)
);

AOI33xp33_ASAP7_75t_L g14733 ( 
.A1(n_14393),
.A2(n_9098),
.A3(n_9088),
.B1(n_9099),
.B2(n_9094),
.B3(n_9086),
.Y(n_14733)
);

NOR3xp33_ASAP7_75t_SL g14734 ( 
.A(n_14258),
.B(n_7826),
.C(n_7801),
.Y(n_14734)
);

INVx1_ASAP7_75t_L g14735 ( 
.A(n_14246),
.Y(n_14735)
);

NOR2x1_ASAP7_75t_L g14736 ( 
.A(n_14420),
.B(n_9094),
.Y(n_14736)
);

AOI21x1_ASAP7_75t_L g14737 ( 
.A1(n_14437),
.A2(n_9099),
.B(n_9098),
.Y(n_14737)
);

AOI22xp5_ASAP7_75t_L g14738 ( 
.A1(n_14404),
.A2(n_7443),
.B1(n_7174),
.B2(n_7284),
.Y(n_14738)
);

OAI22xp33_ASAP7_75t_L g14739 ( 
.A1(n_14371),
.A2(n_9223),
.B1(n_9171),
.B2(n_7920),
.Y(n_14739)
);

INVxp67_ASAP7_75t_L g14740 ( 
.A(n_14479),
.Y(n_14740)
);

AND2x2_ASAP7_75t_L g14741 ( 
.A(n_14277),
.B(n_14200),
.Y(n_14741)
);

OR2x2_ASAP7_75t_L g14742 ( 
.A(n_14491),
.B(n_14288),
.Y(n_14742)
);

INVx1_ASAP7_75t_L g14743 ( 
.A(n_14262),
.Y(n_14743)
);

INVx3_ASAP7_75t_L g14744 ( 
.A(n_14497),
.Y(n_14744)
);

INVx2_ASAP7_75t_L g14745 ( 
.A(n_14573),
.Y(n_14745)
);

INVx2_ASAP7_75t_L g14746 ( 
.A(n_14509),
.Y(n_14746)
);

NAND2xp5_ASAP7_75t_L g14747 ( 
.A(n_14548),
.B(n_9101),
.Y(n_14747)
);

AOI22xp5_ASAP7_75t_L g14748 ( 
.A1(n_14505),
.A2(n_7443),
.B1(n_7174),
.B2(n_7284),
.Y(n_14748)
);

AOI22xp33_ASAP7_75t_SL g14749 ( 
.A1(n_14532),
.A2(n_7443),
.B1(n_7920),
.B2(n_7346),
.Y(n_14749)
);

NAND2xp5_ASAP7_75t_L g14750 ( 
.A(n_14265),
.B(n_9101),
.Y(n_14750)
);

AND2x2_ASAP7_75t_L g14751 ( 
.A(n_14217),
.B(n_9104),
.Y(n_14751)
);

INVx1_ASAP7_75t_L g14752 ( 
.A(n_14264),
.Y(n_14752)
);

OAI21xp33_ASAP7_75t_L g14753 ( 
.A1(n_14321),
.A2(n_9107),
.B(n_9104),
.Y(n_14753)
);

OA222x2_ASAP7_75t_L g14754 ( 
.A1(n_14334),
.A2(n_6271),
.B1(n_9116),
.B2(n_9118),
.C1(n_9115),
.C2(n_9107),
.Y(n_14754)
);

INVx2_ASAP7_75t_L g14755 ( 
.A(n_14504),
.Y(n_14755)
);

INVx2_ASAP7_75t_L g14756 ( 
.A(n_14302),
.Y(n_14756)
);

OAI32xp33_ASAP7_75t_L g14757 ( 
.A1(n_14256),
.A2(n_8099),
.A3(n_8174),
.B1(n_8153),
.B2(n_9115),
.Y(n_14757)
);

AOI22xp5_ASAP7_75t_L g14758 ( 
.A1(n_14449),
.A2(n_7174),
.B1(n_7284),
.B2(n_7920),
.Y(n_14758)
);

INVx1_ASAP7_75t_L g14759 ( 
.A(n_14222),
.Y(n_14759)
);

OAI332xp33_ASAP7_75t_L g14760 ( 
.A1(n_14359),
.A2(n_8174),
.A3(n_8099),
.B1(n_8153),
.B2(n_7201),
.B3(n_6537),
.C1(n_6568),
.C2(n_6575),
.Y(n_14760)
);

INVx1_ASAP7_75t_L g14761 ( 
.A(n_14224),
.Y(n_14761)
);

INVx2_ASAP7_75t_L g14762 ( 
.A(n_14507),
.Y(n_14762)
);

NAND4xp25_ASAP7_75t_L g14763 ( 
.A(n_14406),
.B(n_7768),
.C(n_7861),
.D(n_8187),
.Y(n_14763)
);

OR2x2_ASAP7_75t_L g14764 ( 
.A(n_14514),
.B(n_9116),
.Y(n_14764)
);

NAND2xp5_ASAP7_75t_L g14765 ( 
.A(n_14490),
.B(n_9118),
.Y(n_14765)
);

INVx1_ASAP7_75t_L g14766 ( 
.A(n_14346),
.Y(n_14766)
);

AND2x2_ASAP7_75t_L g14767 ( 
.A(n_14207),
.B(n_9120),
.Y(n_14767)
);

AO221x1_ASAP7_75t_L g14768 ( 
.A1(n_14357),
.A2(n_7954),
.B1(n_8033),
.B2(n_8009),
.C(n_7977),
.Y(n_14768)
);

NAND2xp5_ASAP7_75t_L g14769 ( 
.A(n_14464),
.B(n_9120),
.Y(n_14769)
);

INVx1_ASAP7_75t_L g14770 ( 
.A(n_14274),
.Y(n_14770)
);

AOI22xp5_ASAP7_75t_L g14771 ( 
.A1(n_14387),
.A2(n_14392),
.B1(n_14390),
.B2(n_14311),
.Y(n_14771)
);

AOI22xp33_ASAP7_75t_L g14772 ( 
.A1(n_14551),
.A2(n_7224),
.B1(n_7167),
.B2(n_7460),
.Y(n_14772)
);

INVx1_ASAP7_75t_L g14773 ( 
.A(n_14254),
.Y(n_14773)
);

INVx2_ASAP7_75t_L g14774 ( 
.A(n_14603),
.Y(n_14774)
);

INVx2_ASAP7_75t_SL g14775 ( 
.A(n_14259),
.Y(n_14775)
);

INVx1_ASAP7_75t_L g14776 ( 
.A(n_14502),
.Y(n_14776)
);

OR2x2_ASAP7_75t_L g14777 ( 
.A(n_14216),
.B(n_9124),
.Y(n_14777)
);

NAND2xp5_ASAP7_75t_L g14778 ( 
.A(n_14517),
.B(n_9124),
.Y(n_14778)
);

INVx2_ASAP7_75t_L g14779 ( 
.A(n_14606),
.Y(n_14779)
);

INVx2_ASAP7_75t_SL g14780 ( 
.A(n_14364),
.Y(n_14780)
);

INVx1_ASAP7_75t_L g14781 ( 
.A(n_14531),
.Y(n_14781)
);

INVx1_ASAP7_75t_L g14782 ( 
.A(n_14535),
.Y(n_14782)
);

INVxp67_ASAP7_75t_SL g14783 ( 
.A(n_14484),
.Y(n_14783)
);

NAND2xp5_ASAP7_75t_L g14784 ( 
.A(n_14567),
.B(n_9132),
.Y(n_14784)
);

INVx1_ASAP7_75t_L g14785 ( 
.A(n_14252),
.Y(n_14785)
);

AOI22xp33_ASAP7_75t_SL g14786 ( 
.A1(n_14317),
.A2(n_14300),
.B1(n_14361),
.B2(n_14365),
.Y(n_14786)
);

NOR2x1_ASAP7_75t_L g14787 ( 
.A(n_14493),
.B(n_9132),
.Y(n_14787)
);

XOR2x2_ASAP7_75t_L g14788 ( 
.A(n_14287),
.B(n_7060),
.Y(n_14788)
);

INVx1_ASAP7_75t_L g14789 ( 
.A(n_14602),
.Y(n_14789)
);

NOR2xp67_ASAP7_75t_L g14790 ( 
.A(n_14496),
.B(n_9135),
.Y(n_14790)
);

O2A1O1Ixp5_ASAP7_75t_R g14791 ( 
.A1(n_14308),
.A2(n_7139),
.B(n_7125),
.C(n_6916),
.Y(n_14791)
);

INVx2_ASAP7_75t_L g14792 ( 
.A(n_14475),
.Y(n_14792)
);

INVx2_ASAP7_75t_L g14793 ( 
.A(n_14438),
.Y(n_14793)
);

AOI22xp5_ASAP7_75t_L g14794 ( 
.A1(n_14305),
.A2(n_7284),
.B1(n_7174),
.B2(n_7920),
.Y(n_14794)
);

INVx1_ASAP7_75t_L g14795 ( 
.A(n_14295),
.Y(n_14795)
);

INVx1_ASAP7_75t_L g14796 ( 
.A(n_14270),
.Y(n_14796)
);

INVx2_ASAP7_75t_SL g14797 ( 
.A(n_14276),
.Y(n_14797)
);

AND2x2_ASAP7_75t_L g14798 ( 
.A(n_14296),
.B(n_9135),
.Y(n_14798)
);

INVx1_ASAP7_75t_L g14799 ( 
.A(n_14542),
.Y(n_14799)
);

INVx1_ASAP7_75t_L g14800 ( 
.A(n_14545),
.Y(n_14800)
);

NAND2xp5_ASAP7_75t_L g14801 ( 
.A(n_14540),
.B(n_14541),
.Y(n_14801)
);

AOI22x1_ASAP7_75t_L g14802 ( 
.A1(n_14471),
.A2(n_6687),
.B1(n_6703),
.B2(n_6547),
.Y(n_14802)
);

INVx1_ASAP7_75t_L g14803 ( 
.A(n_14547),
.Y(n_14803)
);

INVx1_ASAP7_75t_L g14804 ( 
.A(n_14549),
.Y(n_14804)
);

INVx2_ASAP7_75t_L g14805 ( 
.A(n_14477),
.Y(n_14805)
);

INVx1_ASAP7_75t_L g14806 ( 
.A(n_14555),
.Y(n_14806)
);

INVx1_ASAP7_75t_L g14807 ( 
.A(n_14556),
.Y(n_14807)
);

OAI32xp33_ASAP7_75t_L g14808 ( 
.A1(n_14240),
.A2(n_8099),
.A3(n_8174),
.B1(n_8153),
.B2(n_9137),
.Y(n_14808)
);

NAND2xp5_ASAP7_75t_L g14809 ( 
.A(n_14580),
.B(n_9137),
.Y(n_14809)
);

AND2x4_ASAP7_75t_L g14810 ( 
.A(n_14423),
.B(n_9280),
.Y(n_14810)
);

AND2x2_ASAP7_75t_L g14811 ( 
.A(n_14430),
.B(n_9141),
.Y(n_14811)
);

INVx1_ASAP7_75t_L g14812 ( 
.A(n_14578),
.Y(n_14812)
);

OA222x2_ASAP7_75t_L g14813 ( 
.A1(n_14369),
.A2(n_6271),
.B1(n_9150),
.B2(n_9157),
.C1(n_9146),
.C2(n_9141),
.Y(n_14813)
);

NAND2xp5_ASAP7_75t_L g14814 ( 
.A(n_14592),
.B(n_9146),
.Y(n_14814)
);

NAND2xp5_ASAP7_75t_L g14815 ( 
.A(n_14596),
.B(n_9150),
.Y(n_14815)
);

INVx2_ASAP7_75t_L g14816 ( 
.A(n_14396),
.Y(n_14816)
);

AND2x2_ASAP7_75t_L g14817 ( 
.A(n_14397),
.B(n_9157),
.Y(n_14817)
);

NAND2xp5_ASAP7_75t_L g14818 ( 
.A(n_14579),
.B(n_9161),
.Y(n_14818)
);

INVx2_ASAP7_75t_L g14819 ( 
.A(n_14481),
.Y(n_14819)
);

OAI32xp33_ASAP7_75t_L g14820 ( 
.A1(n_14245),
.A2(n_9182),
.A3(n_9183),
.B1(n_9179),
.B2(n_9161),
.Y(n_14820)
);

OR2x2_ASAP7_75t_L g14821 ( 
.A(n_14426),
.B(n_9179),
.Y(n_14821)
);

INVx1_ASAP7_75t_L g14822 ( 
.A(n_14421),
.Y(n_14822)
);

OR2x2_ASAP7_75t_L g14823 ( 
.A(n_14466),
.B(n_14427),
.Y(n_14823)
);

AND2x2_ASAP7_75t_L g14824 ( 
.A(n_14471),
.B(n_9182),
.Y(n_14824)
);

INVx1_ASAP7_75t_L g14825 ( 
.A(n_14595),
.Y(n_14825)
);

INVx1_ASAP7_75t_L g14826 ( 
.A(n_14563),
.Y(n_14826)
);

NAND2x1p5_ASAP7_75t_L g14827 ( 
.A(n_14486),
.B(n_8276),
.Y(n_14827)
);

NAND2xp5_ASAP7_75t_L g14828 ( 
.A(n_14458),
.B(n_9183),
.Y(n_14828)
);

OR2x2_ASAP7_75t_L g14829 ( 
.A(n_14470),
.B(n_9184),
.Y(n_14829)
);

NAND5xp2_ASAP7_75t_L g14830 ( 
.A(n_14301),
.B(n_8274),
.C(n_8269),
.D(n_8061),
.E(n_8072),
.Y(n_14830)
);

OR2x2_ASAP7_75t_L g14831 ( 
.A(n_14482),
.B(n_9184),
.Y(n_14831)
);

AND2x4_ASAP7_75t_L g14832 ( 
.A(n_14434),
.B(n_9308),
.Y(n_14832)
);

OAI211xp5_ASAP7_75t_L g14833 ( 
.A1(n_14528),
.A2(n_7460),
.B(n_6197),
.C(n_9308),
.Y(n_14833)
);

OAI32xp33_ASAP7_75t_L g14834 ( 
.A1(n_14485),
.A2(n_9193),
.A3(n_9195),
.B1(n_9190),
.B2(n_9185),
.Y(n_14834)
);

AND2x4_ASAP7_75t_L g14835 ( 
.A(n_14447),
.B(n_9051),
.Y(n_14835)
);

OR2x2_ASAP7_75t_L g14836 ( 
.A(n_14515),
.B(n_9185),
.Y(n_14836)
);

INVxp67_ASAP7_75t_L g14837 ( 
.A(n_14607),
.Y(n_14837)
);

NAND2xp5_ASAP7_75t_L g14838 ( 
.A(n_14431),
.B(n_9190),
.Y(n_14838)
);

NAND2xp5_ASAP7_75t_L g14839 ( 
.A(n_14433),
.B(n_9193),
.Y(n_14839)
);

INVx1_ASAP7_75t_SL g14840 ( 
.A(n_14513),
.Y(n_14840)
);

NAND2x1_ASAP7_75t_SL g14841 ( 
.A(n_14328),
.B(n_6547),
.Y(n_14841)
);

AND2x2_ASAP7_75t_L g14842 ( 
.A(n_14329),
.B(n_9195),
.Y(n_14842)
);

INVx2_ASAP7_75t_L g14843 ( 
.A(n_14536),
.Y(n_14843)
);

OR2x2_ASAP7_75t_L g14844 ( 
.A(n_14529),
.B(n_9197),
.Y(n_14844)
);

INVx1_ASAP7_75t_L g14845 ( 
.A(n_14429),
.Y(n_14845)
);

AOI22xp33_ASAP7_75t_L g14846 ( 
.A1(n_14370),
.A2(n_7224),
.B1(n_7460),
.B2(n_7412),
.Y(n_14846)
);

NAND2xp5_ASAP7_75t_L g14847 ( 
.A(n_14419),
.B(n_14313),
.Y(n_14847)
);

INVx1_ASAP7_75t_L g14848 ( 
.A(n_14407),
.Y(n_14848)
);

INVx1_ASAP7_75t_L g14849 ( 
.A(n_14453),
.Y(n_14849)
);

INVx1_ASAP7_75t_L g14850 ( 
.A(n_14454),
.Y(n_14850)
);

O2A1O1Ixp33_ASAP7_75t_L g14851 ( 
.A1(n_14380),
.A2(n_7618),
.B(n_7759),
.C(n_7460),
.Y(n_14851)
);

NAND2xp5_ASAP7_75t_L g14852 ( 
.A(n_14525),
.B(n_9197),
.Y(n_14852)
);

AND2x2_ASAP7_75t_L g14853 ( 
.A(n_14338),
.B(n_9202),
.Y(n_14853)
);

NAND2xp5_ASAP7_75t_L g14854 ( 
.A(n_14526),
.B(n_9202),
.Y(n_14854)
);

OR2x2_ASAP7_75t_L g14855 ( 
.A(n_14297),
.B(n_9204),
.Y(n_14855)
);

INVx1_ASAP7_75t_L g14856 ( 
.A(n_14325),
.Y(n_14856)
);

AND2x2_ASAP7_75t_L g14857 ( 
.A(n_14422),
.B(n_9204),
.Y(n_14857)
);

INVx1_ASAP7_75t_L g14858 ( 
.A(n_14459),
.Y(n_14858)
);

INVxp67_ASAP7_75t_L g14859 ( 
.A(n_14299),
.Y(n_14859)
);

INVx1_ASAP7_75t_L g14860 ( 
.A(n_14415),
.Y(n_14860)
);

INVx1_ASAP7_75t_L g14861 ( 
.A(n_14465),
.Y(n_14861)
);

INVx2_ASAP7_75t_SL g14862 ( 
.A(n_14354),
.Y(n_14862)
);

OAI33xp33_ASAP7_75t_L g14863 ( 
.A1(n_14307),
.A2(n_9234),
.A3(n_9219),
.B1(n_9239),
.B2(n_9226),
.B3(n_9206),
.Y(n_14863)
);

AOI22xp5_ASAP7_75t_L g14864 ( 
.A1(n_14304),
.A2(n_7174),
.B1(n_7920),
.B2(n_7412),
.Y(n_14864)
);

INVxp33_ASAP7_75t_L g14865 ( 
.A(n_14472),
.Y(n_14865)
);

INVx2_ASAP7_75t_L g14866 ( 
.A(n_14439),
.Y(n_14866)
);

AND2x4_ASAP7_75t_L g14867 ( 
.A(n_14356),
.B(n_9051),
.Y(n_14867)
);

INVx2_ASAP7_75t_L g14868 ( 
.A(n_14439),
.Y(n_14868)
);

INVx1_ASAP7_75t_L g14869 ( 
.A(n_14494),
.Y(n_14869)
);

INVx1_ASAP7_75t_L g14870 ( 
.A(n_14575),
.Y(n_14870)
);

OAI31xp33_ASAP7_75t_L g14871 ( 
.A1(n_14445),
.A2(n_8168),
.A3(n_8283),
.B(n_8231),
.Y(n_14871)
);

INVx1_ASAP7_75t_L g14872 ( 
.A(n_14590),
.Y(n_14872)
);

AOI32xp33_ASAP7_75t_L g14873 ( 
.A1(n_14561),
.A2(n_7484),
.A3(n_7397),
.B1(n_8418),
.B2(n_8385),
.Y(n_14873)
);

AOI22xp5_ASAP7_75t_L g14874 ( 
.A1(n_14416),
.A2(n_7920),
.B1(n_7412),
.B2(n_7460),
.Y(n_14874)
);

NAND2xp5_ASAP7_75t_L g14875 ( 
.A(n_14553),
.B(n_9206),
.Y(n_14875)
);

NAND2xp5_ASAP7_75t_L g14876 ( 
.A(n_14599),
.B(n_9219),
.Y(n_14876)
);

INVx2_ASAP7_75t_L g14877 ( 
.A(n_14376),
.Y(n_14877)
);

AOI22xp5_ASAP7_75t_L g14878 ( 
.A1(n_14598),
.A2(n_7412),
.B1(n_9234),
.B2(n_9226),
.Y(n_14878)
);

INVx2_ASAP7_75t_L g14879 ( 
.A(n_14538),
.Y(n_14879)
);

A2O1A1Ixp33_ASAP7_75t_L g14880 ( 
.A1(n_14405),
.A2(n_7248),
.B(n_7397),
.C(n_7240),
.Y(n_14880)
);

INVx1_ASAP7_75t_L g14881 ( 
.A(n_14512),
.Y(n_14881)
);

OR2x2_ASAP7_75t_L g14882 ( 
.A(n_14582),
.B(n_9239),
.Y(n_14882)
);

INVx3_ASAP7_75t_L g14883 ( 
.A(n_14594),
.Y(n_14883)
);

INVx1_ASAP7_75t_L g14884 ( 
.A(n_14601),
.Y(n_14884)
);

NAND2x1p5_ASAP7_75t_L g14885 ( 
.A(n_14368),
.B(n_8276),
.Y(n_14885)
);

AND2x2_ASAP7_75t_L g14886 ( 
.A(n_14522),
.B(n_9241),
.Y(n_14886)
);

INVx1_ASAP7_75t_L g14887 ( 
.A(n_14604),
.Y(n_14887)
);

AOI22xp5_ASAP7_75t_L g14888 ( 
.A1(n_14460),
.A2(n_7412),
.B1(n_9244),
.B2(n_9241),
.Y(n_14888)
);

AOI22xp5_ASAP7_75t_L g14889 ( 
.A1(n_14355),
.A2(n_7412),
.B1(n_9247),
.B2(n_9244),
.Y(n_14889)
);

AND2x4_ASAP7_75t_L g14890 ( 
.A(n_14389),
.B(n_9247),
.Y(n_14890)
);

INVx1_ASAP7_75t_L g14891 ( 
.A(n_14605),
.Y(n_14891)
);

OAI32xp33_ASAP7_75t_L g14892 ( 
.A1(n_14298),
.A2(n_9253),
.A3(n_9256),
.B1(n_9251),
.B2(n_9249),
.Y(n_14892)
);

NAND2xp5_ASAP7_75t_L g14893 ( 
.A(n_14539),
.B(n_9249),
.Y(n_14893)
);

INVx2_ASAP7_75t_L g14894 ( 
.A(n_14558),
.Y(n_14894)
);

NAND2xp5_ASAP7_75t_L g14895 ( 
.A(n_14570),
.B(n_9251),
.Y(n_14895)
);

NOR2x1_ASAP7_75t_L g14896 ( 
.A(n_14381),
.B(n_9253),
.Y(n_14896)
);

INVx1_ASAP7_75t_L g14897 ( 
.A(n_14572),
.Y(n_14897)
);

INVx2_ASAP7_75t_L g14898 ( 
.A(n_14560),
.Y(n_14898)
);

INVx1_ASAP7_75t_L g14899 ( 
.A(n_14571),
.Y(n_14899)
);

INVx1_ASAP7_75t_L g14900 ( 
.A(n_14506),
.Y(n_14900)
);

OAI222xp33_ASAP7_75t_L g14901 ( 
.A1(n_14583),
.A2(n_7385),
.B1(n_7200),
.B2(n_7402),
.C1(n_7281),
.C2(n_7164),
.Y(n_14901)
);

OAI22xp33_ASAP7_75t_SL g14902 ( 
.A1(n_14518),
.A2(n_7200),
.B1(n_7281),
.B2(n_7164),
.Y(n_14902)
);

INVx1_ASAP7_75t_L g14903 ( 
.A(n_14372),
.Y(n_14903)
);

NOR2x1p5_ASAP7_75t_L g14904 ( 
.A(n_14388),
.B(n_6939),
.Y(n_14904)
);

OAI33xp33_ASAP7_75t_L g14905 ( 
.A1(n_14412),
.A2(n_9260),
.A3(n_9258),
.B1(n_9263),
.B2(n_9259),
.B3(n_9256),
.Y(n_14905)
);

INVx1_ASAP7_75t_L g14906 ( 
.A(n_14476),
.Y(n_14906)
);

INVx1_ASAP7_75t_L g14907 ( 
.A(n_14543),
.Y(n_14907)
);

INVx1_ASAP7_75t_L g14908 ( 
.A(n_14373),
.Y(n_14908)
);

NAND2xp5_ASAP7_75t_L g14909 ( 
.A(n_14566),
.B(n_9258),
.Y(n_14909)
);

A2O1A1Ixp33_ASAP7_75t_L g14910 ( 
.A1(n_14480),
.A2(n_7248),
.B(n_7397),
.C(n_7240),
.Y(n_14910)
);

INVx2_ASAP7_75t_SL g14911 ( 
.A(n_14574),
.Y(n_14911)
);

NAND2xp5_ASAP7_75t_SL g14912 ( 
.A(n_14448),
.B(n_9259),
.Y(n_14912)
);

INVx1_ASAP7_75t_L g14913 ( 
.A(n_14467),
.Y(n_14913)
);

INVx1_ASAP7_75t_L g14914 ( 
.A(n_14469),
.Y(n_14914)
);

INVxp67_ASAP7_75t_L g14915 ( 
.A(n_14315),
.Y(n_14915)
);

INVx1_ASAP7_75t_L g14916 ( 
.A(n_14503),
.Y(n_14916)
);

NAND2xp5_ASAP7_75t_L g14917 ( 
.A(n_14569),
.B(n_9260),
.Y(n_14917)
);

INVx1_ASAP7_75t_L g14918 ( 
.A(n_14336),
.Y(n_14918)
);

INVx1_ASAP7_75t_L g14919 ( 
.A(n_14353),
.Y(n_14919)
);

INVx2_ASAP7_75t_L g14920 ( 
.A(n_14577),
.Y(n_14920)
);

HB1xp67_ASAP7_75t_L g14921 ( 
.A(n_14492),
.Y(n_14921)
);

OR3x2_ASAP7_75t_L g14922 ( 
.A(n_14591),
.B(n_6568),
.C(n_6537),
.Y(n_14922)
);

INVx1_ASAP7_75t_L g14923 ( 
.A(n_14487),
.Y(n_14923)
);

OR2x2_ASAP7_75t_L g14924 ( 
.A(n_14589),
.B(n_9263),
.Y(n_14924)
);

INVx1_ASAP7_75t_L g14925 ( 
.A(n_14418),
.Y(n_14925)
);

NAND2xp5_ASAP7_75t_L g14926 ( 
.A(n_14581),
.B(n_9267),
.Y(n_14926)
);

INVx1_ASAP7_75t_L g14927 ( 
.A(n_14394),
.Y(n_14927)
);

AND2x2_ASAP7_75t_L g14928 ( 
.A(n_14367),
.B(n_9267),
.Y(n_14928)
);

INVxp67_ASAP7_75t_L g14929 ( 
.A(n_14501),
.Y(n_14929)
);

AOI322xp5_ASAP7_75t_L g14930 ( 
.A1(n_14499),
.A2(n_7201),
.A3(n_7082),
.B1(n_7538),
.B2(n_7131),
.C1(n_7130),
.C2(n_8127),
.Y(n_14930)
);

INVx1_ASAP7_75t_L g14931 ( 
.A(n_14345),
.Y(n_14931)
);

XNOR2xp5_ASAP7_75t_L g14932 ( 
.A(n_14432),
.B(n_7060),
.Y(n_14932)
);

INVx1_ASAP7_75t_SL g14933 ( 
.A(n_14510),
.Y(n_14933)
);

OR2x2_ASAP7_75t_L g14934 ( 
.A(n_14593),
.B(n_9268),
.Y(n_14934)
);

INVx1_ASAP7_75t_L g14935 ( 
.A(n_14362),
.Y(n_14935)
);

AND2x2_ASAP7_75t_L g14936 ( 
.A(n_14303),
.B(n_9268),
.Y(n_14936)
);

INVx1_ASAP7_75t_L g14937 ( 
.A(n_14350),
.Y(n_14937)
);

NAND2xp5_ASAP7_75t_L g14938 ( 
.A(n_14584),
.B(n_9274),
.Y(n_14938)
);

AND2x2_ASAP7_75t_L g14939 ( 
.A(n_14402),
.B(n_9274),
.Y(n_14939)
);

AND2x4_ASAP7_75t_L g14940 ( 
.A(n_14360),
.B(n_9064),
.Y(n_14940)
);

AOI22xp5_ASAP7_75t_L g14941 ( 
.A1(n_14314),
.A2(n_9290),
.B1(n_9296),
.B2(n_9286),
.Y(n_14941)
);

AND2x2_ASAP7_75t_L g14942 ( 
.A(n_14409),
.B(n_9286),
.Y(n_14942)
);

INVxp67_ASAP7_75t_L g14943 ( 
.A(n_14463),
.Y(n_14943)
);

NOR2xp33_ASAP7_75t_L g14944 ( 
.A(n_14585),
.B(n_9290),
.Y(n_14944)
);

INVx1_ASAP7_75t_L g14945 ( 
.A(n_14600),
.Y(n_14945)
);

INVx2_ASAP7_75t_SL g14946 ( 
.A(n_14462),
.Y(n_14946)
);

INVx2_ASAP7_75t_SL g14947 ( 
.A(n_14441),
.Y(n_14947)
);

INVx1_ASAP7_75t_L g14948 ( 
.A(n_14382),
.Y(n_14948)
);

AOI22xp5_ASAP7_75t_L g14949 ( 
.A1(n_14443),
.A2(n_9310),
.B1(n_9311),
.B2(n_9296),
.Y(n_14949)
);

NOR2x1_ASAP7_75t_L g14950 ( 
.A(n_14618),
.B(n_14425),
.Y(n_14950)
);

NAND2xp5_ASAP7_75t_L g14951 ( 
.A(n_14648),
.B(n_14546),
.Y(n_14951)
);

NAND2xp33_ASAP7_75t_R g14952 ( 
.A(n_14651),
.B(n_14690),
.Y(n_14952)
);

AND2x2_ASAP7_75t_L g14953 ( 
.A(n_14700),
.B(n_14483),
.Y(n_14953)
);

INVxp33_ASAP7_75t_L g14954 ( 
.A(n_14709),
.Y(n_14954)
);

NAND2xp5_ASAP7_75t_L g14955 ( 
.A(n_14654),
.B(n_14452),
.Y(n_14955)
);

NOR2xp33_ASAP7_75t_L g14956 ( 
.A(n_14732),
.B(n_14349),
.Y(n_14956)
);

AND2x4_ASAP7_75t_L g14957 ( 
.A(n_14699),
.B(n_14608),
.Y(n_14957)
);

NAND2xp5_ASAP7_75t_L g14958 ( 
.A(n_14707),
.B(n_14488),
.Y(n_14958)
);

INVx1_ASAP7_75t_L g14959 ( 
.A(n_14655),
.Y(n_14959)
);

NAND2xp5_ASAP7_75t_L g14960 ( 
.A(n_14642),
.B(n_14609),
.Y(n_14960)
);

INVx2_ASAP7_75t_L g14961 ( 
.A(n_14742),
.Y(n_14961)
);

NAND2xp5_ASAP7_75t_SL g14962 ( 
.A(n_14688),
.B(n_14674),
.Y(n_14962)
);

INVx2_ASAP7_75t_L g14963 ( 
.A(n_14725),
.Y(n_14963)
);

INVx1_ASAP7_75t_L g14964 ( 
.A(n_14612),
.Y(n_14964)
);

OR2x2_ASAP7_75t_L g14965 ( 
.A(n_14610),
.B(n_14586),
.Y(n_14965)
);

AND2x2_ASAP7_75t_L g14966 ( 
.A(n_14627),
.B(n_14358),
.Y(n_14966)
);

AND2x2_ASAP7_75t_SL g14967 ( 
.A(n_14714),
.B(n_14442),
.Y(n_14967)
);

NAND2xp5_ASAP7_75t_L g14968 ( 
.A(n_14672),
.B(n_14516),
.Y(n_14968)
);

NOR2xp33_ASAP7_75t_L g14969 ( 
.A(n_14646),
.B(n_14562),
.Y(n_14969)
);

OR2x2_ASAP7_75t_L g14970 ( 
.A(n_14775),
.B(n_14564),
.Y(n_14970)
);

INVx1_ASAP7_75t_L g14971 ( 
.A(n_14658),
.Y(n_14971)
);

INVx5_ASAP7_75t_L g14972 ( 
.A(n_14614),
.Y(n_14972)
);

AOI21xp33_ASAP7_75t_L g14973 ( 
.A1(n_14933),
.A2(n_14417),
.B(n_14446),
.Y(n_14973)
);

AOI22xp33_ASAP7_75t_L g14974 ( 
.A1(n_14921),
.A2(n_14468),
.B1(n_14461),
.B2(n_14351),
.Y(n_14974)
);

INVx1_ASAP7_75t_L g14975 ( 
.A(n_14613),
.Y(n_14975)
);

OR2x2_ASAP7_75t_L g14976 ( 
.A(n_14797),
.B(n_14330),
.Y(n_14976)
);

HB1xp67_ASAP7_75t_L g14977 ( 
.A(n_14619),
.Y(n_14977)
);

NAND4xp25_ASAP7_75t_L g14978 ( 
.A(n_14641),
.B(n_14544),
.C(n_14534),
.D(n_14511),
.Y(n_14978)
);

AND2x4_ASAP7_75t_L g14979 ( 
.A(n_14744),
.B(n_14779),
.Y(n_14979)
);

AND2x2_ASAP7_75t_L g14980 ( 
.A(n_14741),
.B(n_14327),
.Y(n_14980)
);

NOR2xp33_ASAP7_75t_L g14981 ( 
.A(n_14630),
.B(n_14588),
.Y(n_14981)
);

INVx3_ASAP7_75t_SL g14982 ( 
.A(n_14780),
.Y(n_14982)
);

INVx1_ASAP7_75t_L g14983 ( 
.A(n_14617),
.Y(n_14983)
);

AND2x2_ASAP7_75t_L g14984 ( 
.A(n_14865),
.B(n_14331),
.Y(n_14984)
);

AOI22xp33_ASAP7_75t_L g14985 ( 
.A1(n_14635),
.A2(n_14489),
.B1(n_14451),
.B2(n_14294),
.Y(n_14985)
);

AND2x2_ASAP7_75t_L g14986 ( 
.A(n_14625),
.B(n_14333),
.Y(n_14986)
);

INVx1_ASAP7_75t_L g14987 ( 
.A(n_14620),
.Y(n_14987)
);

AND2x2_ASAP7_75t_L g14988 ( 
.A(n_14664),
.B(n_14375),
.Y(n_14988)
);

NOR2xp33_ASAP7_75t_R g14989 ( 
.A(n_14666),
.B(n_14344),
.Y(n_14989)
);

INVx1_ASAP7_75t_L g14990 ( 
.A(n_14783),
.Y(n_14990)
);

INVx2_ASAP7_75t_L g14991 ( 
.A(n_14774),
.Y(n_14991)
);

HB1xp67_ASAP7_75t_L g14992 ( 
.A(n_14624),
.Y(n_14992)
);

INVx1_ASAP7_75t_L g14993 ( 
.A(n_14616),
.Y(n_14993)
);

INVx1_ASAP7_75t_L g14994 ( 
.A(n_14823),
.Y(n_14994)
);

NAND2xp5_ASAP7_75t_L g14995 ( 
.A(n_14669),
.B(n_14523),
.Y(n_14995)
);

AND2x2_ASAP7_75t_L g14996 ( 
.A(n_14650),
.B(n_14424),
.Y(n_14996)
);

BUFx2_ASAP7_75t_L g14997 ( 
.A(n_14841),
.Y(n_14997)
);

INVx1_ASAP7_75t_L g14998 ( 
.A(n_14631),
.Y(n_14998)
);

INVx1_ASAP7_75t_L g14999 ( 
.A(n_14657),
.Y(n_14999)
);

INVx2_ASAP7_75t_L g15000 ( 
.A(n_14922),
.Y(n_15000)
);

NOR2xp33_ASAP7_75t_L g15001 ( 
.A(n_14628),
.B(n_14478),
.Y(n_15001)
);

AOI22xp5_ASAP7_75t_L g15002 ( 
.A1(n_14622),
.A2(n_14947),
.B1(n_14786),
.B2(n_14771),
.Y(n_15002)
);

INVx1_ASAP7_75t_SL g15003 ( 
.A(n_14649),
.Y(n_15003)
);

INVx1_ASAP7_75t_SL g15004 ( 
.A(n_14653),
.Y(n_15004)
);

INVx1_ASAP7_75t_L g15005 ( 
.A(n_14659),
.Y(n_15005)
);

AND2x2_ASAP7_75t_L g15006 ( 
.A(n_14816),
.B(n_14524),
.Y(n_15006)
);

AND2x2_ASAP7_75t_L g15007 ( 
.A(n_14621),
.B(n_14527),
.Y(n_15007)
);

INVx6_ASAP7_75t_L g15008 ( 
.A(n_14645),
.Y(n_15008)
);

OR2x2_ASAP7_75t_L g15009 ( 
.A(n_14706),
.B(n_14533),
.Y(n_15009)
);

NAND2xp5_ASAP7_75t_L g15010 ( 
.A(n_14667),
.B(n_14530),
.Y(n_15010)
);

AND2x2_ASAP7_75t_L g15011 ( 
.A(n_14697),
.B(n_14557),
.Y(n_15011)
);

NAND2xp5_ASAP7_75t_L g15012 ( 
.A(n_14770),
.B(n_14379),
.Y(n_15012)
);

OR2x2_ASAP7_75t_L g15013 ( 
.A(n_14717),
.B(n_14410),
.Y(n_15013)
);

AND2x2_ASAP7_75t_L g15014 ( 
.A(n_14633),
.B(n_14623),
.Y(n_15014)
);

NOR3xp33_ASAP7_75t_L g15015 ( 
.A(n_14723),
.B(n_14399),
.C(n_14408),
.Y(n_15015)
);

INVx1_ASAP7_75t_L g15016 ( 
.A(n_14632),
.Y(n_15016)
);

CKINVDCx20_ASAP7_75t_R g15017 ( 
.A(n_14615),
.Y(n_15017)
);

OR2x2_ASAP7_75t_L g15018 ( 
.A(n_14652),
.B(n_14639),
.Y(n_15018)
);

INVx1_ASAP7_75t_L g15019 ( 
.A(n_14693),
.Y(n_15019)
);

AND2x2_ASAP7_75t_L g15020 ( 
.A(n_14773),
.B(n_14414),
.Y(n_15020)
);

NOR2x1_ASAP7_75t_L g15021 ( 
.A(n_14640),
.B(n_14374),
.Y(n_15021)
);

NOR2xp33_ASAP7_75t_L g15022 ( 
.A(n_14647),
.B(n_14379),
.Y(n_15022)
);

AND2x2_ASAP7_75t_L g15023 ( 
.A(n_14735),
.B(n_14377),
.Y(n_15023)
);

NAND2xp5_ASAP7_75t_L g15024 ( 
.A(n_14819),
.B(n_14400),
.Y(n_15024)
);

AND2x2_ASAP7_75t_L g15025 ( 
.A(n_14611),
.B(n_14400),
.Y(n_15025)
);

AND2x2_ASAP7_75t_L g15026 ( 
.A(n_14676),
.B(n_14450),
.Y(n_15026)
);

INVxp67_ASAP7_75t_SL g15027 ( 
.A(n_14637),
.Y(n_15027)
);

OR2x2_ASAP7_75t_L g15028 ( 
.A(n_14762),
.B(n_14378),
.Y(n_15028)
);

OAI31xp33_ASAP7_75t_SL g15029 ( 
.A1(n_14663),
.A2(n_14473),
.A3(n_14395),
.B(n_14318),
.Y(n_15029)
);

INVx1_ASAP7_75t_L g15030 ( 
.A(n_14703),
.Y(n_15030)
);

INVx1_ASAP7_75t_L g15031 ( 
.A(n_14643),
.Y(n_15031)
);

AND2x2_ASAP7_75t_L g15032 ( 
.A(n_14837),
.B(n_14395),
.Y(n_15032)
);

NOR2xp33_ASAP7_75t_L g15033 ( 
.A(n_14728),
.B(n_14677),
.Y(n_15033)
);

HB1xp67_ASAP7_75t_L g15034 ( 
.A(n_14756),
.Y(n_15034)
);

AOI31xp33_ASAP7_75t_L g15035 ( 
.A1(n_14740),
.A2(n_14473),
.A3(n_14386),
.B(n_14495),
.Y(n_15035)
);

NAND2xp5_ASAP7_75t_L g15036 ( 
.A(n_14793),
.B(n_14456),
.Y(n_15036)
);

AND2x2_ASAP7_75t_L g15037 ( 
.A(n_14826),
.B(n_14552),
.Y(n_15037)
);

OR2x2_ASAP7_75t_L g15038 ( 
.A(n_14796),
.B(n_14550),
.Y(n_15038)
);

NOR3xp33_ASAP7_75t_L g15039 ( 
.A(n_14629),
.B(n_14587),
.C(n_7514),
.Y(n_15039)
);

AND2x2_ASAP7_75t_L g15040 ( 
.A(n_14731),
.B(n_9310),
.Y(n_15040)
);

NAND2xp5_ASAP7_75t_L g15041 ( 
.A(n_14792),
.B(n_9311),
.Y(n_15041)
);

HB1xp67_ASAP7_75t_L g15042 ( 
.A(n_14644),
.Y(n_15042)
);

INVx1_ASAP7_75t_L g15043 ( 
.A(n_14720),
.Y(n_15043)
);

INVx1_ASAP7_75t_SL g15044 ( 
.A(n_14656),
.Y(n_15044)
);

AND2x2_ASAP7_75t_L g15045 ( 
.A(n_14734),
.B(n_8276),
.Y(n_15045)
);

INVx2_ASAP7_75t_SL g15046 ( 
.A(n_14727),
.Y(n_15046)
);

INVx1_ASAP7_75t_L g15047 ( 
.A(n_14737),
.Y(n_15047)
);

CKINVDCx8_ASAP7_75t_R g15048 ( 
.A(n_14626),
.Y(n_15048)
);

NOR2xp33_ASAP7_75t_L g15049 ( 
.A(n_14638),
.B(n_5897),
.Y(n_15049)
);

AND2x2_ASAP7_75t_L g15050 ( 
.A(n_14743),
.B(n_8276),
.Y(n_15050)
);

NAND2xp5_ASAP7_75t_L g15051 ( 
.A(n_14805),
.B(n_14884),
.Y(n_15051)
);

INVx2_ASAP7_75t_SL g15052 ( 
.A(n_14904),
.Y(n_15052)
);

NAND2xp5_ASAP7_75t_L g15053 ( 
.A(n_14887),
.B(n_14891),
.Y(n_15053)
);

AND2x2_ASAP7_75t_L g15054 ( 
.A(n_14692),
.B(n_8276),
.Y(n_15054)
);

INVx1_ASAP7_75t_L g15055 ( 
.A(n_14726),
.Y(n_15055)
);

NAND2xp5_ASAP7_75t_L g15056 ( 
.A(n_14856),
.B(n_7201),
.Y(n_15056)
);

INVx2_ASAP7_75t_L g15057 ( 
.A(n_14885),
.Y(n_15057)
);

NOR2xp33_ASAP7_75t_L g15058 ( 
.A(n_14859),
.B(n_7226),
.Y(n_15058)
);

NAND3xp33_ASAP7_75t_SL g15059 ( 
.A(n_14636),
.B(n_7281),
.C(n_7164),
.Y(n_15059)
);

INVx1_ASAP7_75t_L g15060 ( 
.A(n_14824),
.Y(n_15060)
);

AND2x2_ASAP7_75t_L g15061 ( 
.A(n_14670),
.B(n_8276),
.Y(n_15061)
);

AOI22xp33_ASAP7_75t_L g15062 ( 
.A1(n_14686),
.A2(n_8224),
.B1(n_8209),
.B2(n_7358),
.Y(n_15062)
);

OR2x2_ASAP7_75t_L g15063 ( 
.A(n_14662),
.B(n_7852),
.Y(n_15063)
);

OR2x2_ASAP7_75t_L g15064 ( 
.A(n_14825),
.B(n_7852),
.Y(n_15064)
);

AND2x2_ASAP7_75t_L g15065 ( 
.A(n_14634),
.B(n_6193),
.Y(n_15065)
);

INVx1_ASAP7_75t_L g15066 ( 
.A(n_14719),
.Y(n_15066)
);

AND2x2_ASAP7_75t_L g15067 ( 
.A(n_14862),
.B(n_6193),
.Y(n_15067)
);

INVx1_ASAP7_75t_L g15068 ( 
.A(n_14845),
.Y(n_15068)
);

NAND2xp33_ASAP7_75t_SL g15069 ( 
.A(n_14911),
.B(n_6687),
.Y(n_15069)
);

HB1xp67_ASAP7_75t_L g15070 ( 
.A(n_14790),
.Y(n_15070)
);

AND2x4_ASAP7_75t_L g15071 ( 
.A(n_14879),
.B(n_9064),
.Y(n_15071)
);

AND2x2_ASAP7_75t_L g15072 ( 
.A(n_14698),
.B(n_6193),
.Y(n_15072)
);

NOR3xp33_ASAP7_75t_L g15073 ( 
.A(n_14691),
.B(n_7514),
.C(n_7503),
.Y(n_15073)
);

INVx1_ASAP7_75t_L g15074 ( 
.A(n_14858),
.Y(n_15074)
);

AND2x2_ASAP7_75t_L g15075 ( 
.A(n_14789),
.B(n_6217),
.Y(n_15075)
);

OR2x2_ASAP7_75t_L g15076 ( 
.A(n_14894),
.B(n_7852),
.Y(n_15076)
);

INVx1_ASAP7_75t_L g15077 ( 
.A(n_14860),
.Y(n_15077)
);

INVx2_ASAP7_75t_L g15078 ( 
.A(n_14827),
.Y(n_15078)
);

AND2x2_ASAP7_75t_L g15079 ( 
.A(n_14898),
.B(n_6217),
.Y(n_15079)
);

AND2x2_ASAP7_75t_L g15080 ( 
.A(n_14920),
.B(n_6217),
.Y(n_15080)
);

OAI211xp5_ASAP7_75t_SL g15081 ( 
.A1(n_14929),
.A2(n_8195),
.B(n_8199),
.C(n_8187),
.Y(n_15081)
);

NAND2xp5_ASAP7_75t_L g15082 ( 
.A(n_14861),
.B(n_7201),
.Y(n_15082)
);

NAND2xp5_ASAP7_75t_L g15083 ( 
.A(n_14903),
.B(n_7201),
.Y(n_15083)
);

OR2x2_ASAP7_75t_L g15084 ( 
.A(n_14799),
.B(n_7852),
.Y(n_15084)
);

NAND2xp5_ASAP7_75t_SL g15085 ( 
.A(n_14800),
.B(n_7173),
.Y(n_15085)
);

NAND2xp5_ASAP7_75t_L g15086 ( 
.A(n_14849),
.B(n_7201),
.Y(n_15086)
);

NAND2xp5_ASAP7_75t_L g15087 ( 
.A(n_14850),
.B(n_7201),
.Y(n_15087)
);

AND2x2_ASAP7_75t_L g15088 ( 
.A(n_14843),
.B(n_6234),
.Y(n_15088)
);

HB1xp67_ASAP7_75t_L g15089 ( 
.A(n_14900),
.Y(n_15089)
);

AND2x2_ASAP7_75t_L g15090 ( 
.A(n_14785),
.B(n_6234),
.Y(n_15090)
);

INVx1_ASAP7_75t_L g15091 ( 
.A(n_14848),
.Y(n_15091)
);

NOR2xp33_ASAP7_75t_L g15092 ( 
.A(n_14915),
.B(n_7239),
.Y(n_15092)
);

AND2x2_ASAP7_75t_L g15093 ( 
.A(n_14842),
.B(n_6234),
.Y(n_15093)
);

INVx1_ASAP7_75t_L g15094 ( 
.A(n_14718),
.Y(n_15094)
);

NAND2xp5_ASAP7_75t_L g15095 ( 
.A(n_14897),
.B(n_7201),
.Y(n_15095)
);

NAND2xp5_ASAP7_75t_L g15096 ( 
.A(n_14881),
.B(n_7852),
.Y(n_15096)
);

AND2x4_ASAP7_75t_L g15097 ( 
.A(n_14803),
.B(n_9092),
.Y(n_15097)
);

INVx2_ASAP7_75t_L g15098 ( 
.A(n_14695),
.Y(n_15098)
);

NAND4xp25_ASAP7_75t_SL g15099 ( 
.A(n_14801),
.B(n_8199),
.C(n_8249),
.D(n_8195),
.Y(n_15099)
);

INVx1_ASAP7_75t_L g15100 ( 
.A(n_14702),
.Y(n_15100)
);

CKINVDCx5p33_ASAP7_75t_R g15101 ( 
.A(n_14840),
.Y(n_15101)
);

INVx1_ASAP7_75t_L g15102 ( 
.A(n_14899),
.Y(n_15102)
);

OR2x2_ASAP7_75t_L g15103 ( 
.A(n_14804),
.B(n_7852),
.Y(n_15103)
);

AND2x2_ASAP7_75t_L g15104 ( 
.A(n_14806),
.B(n_6256),
.Y(n_15104)
);

INVx1_ASAP7_75t_L g15105 ( 
.A(n_14807),
.Y(n_15105)
);

HB1xp67_ASAP7_75t_L g15106 ( 
.A(n_14946),
.Y(n_15106)
);

NAND2xp5_ASAP7_75t_L g15107 ( 
.A(n_14943),
.B(n_7852),
.Y(n_15107)
);

AND2x2_ASAP7_75t_L g15108 ( 
.A(n_14812),
.B(n_14759),
.Y(n_15108)
);

INVxp67_ASAP7_75t_L g15109 ( 
.A(n_14678),
.Y(n_15109)
);

NAND3xp33_ASAP7_75t_SL g15110 ( 
.A(n_14682),
.B(n_7281),
.C(n_7164),
.Y(n_15110)
);

INVxp67_ASAP7_75t_L g15111 ( 
.A(n_14704),
.Y(n_15111)
);

NAND2xp5_ASAP7_75t_L g15112 ( 
.A(n_14701),
.B(n_7852),
.Y(n_15112)
);

NAND2xp5_ASAP7_75t_L g15113 ( 
.A(n_14908),
.B(n_7984),
.Y(n_15113)
);

INVxp67_ASAP7_75t_SL g15114 ( 
.A(n_14847),
.Y(n_15114)
);

NAND2xp33_ASAP7_75t_SL g15115 ( 
.A(n_14761),
.B(n_6687),
.Y(n_15115)
);

INVx2_ASAP7_75t_L g15116 ( 
.A(n_14695),
.Y(n_15116)
);

OR2x4_ASAP7_75t_L g15117 ( 
.A(n_14722),
.B(n_7173),
.Y(n_15117)
);

AND2x2_ASAP7_75t_L g15118 ( 
.A(n_14776),
.B(n_6256),
.Y(n_15118)
);

AND2x2_ASAP7_75t_L g15119 ( 
.A(n_14781),
.B(n_6256),
.Y(n_15119)
);

NAND2x1p5_ASAP7_75t_L g15120 ( 
.A(n_14752),
.B(n_14822),
.Y(n_15120)
);

AND2x2_ASAP7_75t_SL g15121 ( 
.A(n_14782),
.B(n_8023),
.Y(n_15121)
);

NAND2xp5_ASAP7_75t_L g15122 ( 
.A(n_14919),
.B(n_7984),
.Y(n_15122)
);

INVx1_ASAP7_75t_L g15123 ( 
.A(n_14787),
.Y(n_15123)
);

NAND2xp5_ASAP7_75t_L g15124 ( 
.A(n_14927),
.B(n_14857),
.Y(n_15124)
);

INVx1_ASAP7_75t_SL g15125 ( 
.A(n_14877),
.Y(n_15125)
);

INVx1_ASAP7_75t_SL g15126 ( 
.A(n_14913),
.Y(n_15126)
);

INVx2_ASAP7_75t_L g15127 ( 
.A(n_14788),
.Y(n_15127)
);

AND2x2_ASAP7_75t_L g15128 ( 
.A(n_14795),
.B(n_6257),
.Y(n_15128)
);

OR2x2_ASAP7_75t_L g15129 ( 
.A(n_14914),
.B(n_7984),
.Y(n_15129)
);

NAND2xp5_ASAP7_75t_L g15130 ( 
.A(n_14925),
.B(n_14931),
.Y(n_15130)
);

BUFx2_ASAP7_75t_L g15131 ( 
.A(n_14736),
.Y(n_15131)
);

INVx1_ASAP7_75t_L g15132 ( 
.A(n_14750),
.Y(n_15132)
);

AND2x2_ASAP7_75t_L g15133 ( 
.A(n_14883),
.B(n_6257),
.Y(n_15133)
);

INVx1_ASAP7_75t_SL g15134 ( 
.A(n_14766),
.Y(n_15134)
);

AND2x4_ASAP7_75t_SL g15135 ( 
.A(n_14681),
.B(n_7130),
.Y(n_15135)
);

OR2x2_ASAP7_75t_L g15136 ( 
.A(n_14696),
.B(n_7984),
.Y(n_15136)
);

INVx1_ASAP7_75t_L g15137 ( 
.A(n_14661),
.Y(n_15137)
);

AND2x2_ASAP7_75t_L g15138 ( 
.A(n_14886),
.B(n_6257),
.Y(n_15138)
);

NOR2xp33_ASAP7_75t_R g15139 ( 
.A(n_14945),
.B(n_6687),
.Y(n_15139)
);

NAND2xp5_ASAP7_75t_L g15140 ( 
.A(n_14935),
.B(n_7984),
.Y(n_15140)
);

INVx1_ASAP7_75t_L g15141 ( 
.A(n_14831),
.Y(n_15141)
);

INVx5_ASAP7_75t_L g15142 ( 
.A(n_14866),
.Y(n_15142)
);

INVx1_ASAP7_75t_L g15143 ( 
.A(n_14836),
.Y(n_15143)
);

NOR2xp33_ASAP7_75t_L g15144 ( 
.A(n_14724),
.B(n_14729),
.Y(n_15144)
);

NAND2xp5_ASAP7_75t_L g15145 ( 
.A(n_14937),
.B(n_14948),
.Y(n_15145)
);

NAND2xp5_ASAP7_75t_L g15146 ( 
.A(n_14798),
.B(n_7984),
.Y(n_15146)
);

NAND2xp5_ASAP7_75t_L g15147 ( 
.A(n_14811),
.B(n_7984),
.Y(n_15147)
);

INVx1_ASAP7_75t_L g15148 ( 
.A(n_14844),
.Y(n_15148)
);

AND2x2_ASAP7_75t_L g15149 ( 
.A(n_14817),
.B(n_6327),
.Y(n_15149)
);

INVx1_ASAP7_75t_L g15150 ( 
.A(n_14895),
.Y(n_15150)
);

OR2x2_ASAP7_75t_L g15151 ( 
.A(n_14716),
.B(n_7984),
.Y(n_15151)
);

OR2x2_ASAP7_75t_L g15152 ( 
.A(n_14784),
.B(n_7764),
.Y(n_15152)
);

HB1xp67_ASAP7_75t_L g15153 ( 
.A(n_14923),
.Y(n_15153)
);

INVx2_ASAP7_75t_L g15154 ( 
.A(n_14924),
.Y(n_15154)
);

INVx1_ASAP7_75t_L g15155 ( 
.A(n_14882),
.Y(n_15155)
);

AND2x2_ASAP7_75t_L g15156 ( 
.A(n_14869),
.B(n_14906),
.Y(n_15156)
);

NAND2xp33_ASAP7_75t_R g15157 ( 
.A(n_14907),
.B(n_7847),
.Y(n_15157)
);

INVx1_ASAP7_75t_L g15158 ( 
.A(n_14934),
.Y(n_15158)
);

CKINVDCx16_ASAP7_75t_R g15159 ( 
.A(n_14918),
.Y(n_15159)
);

INVx1_ASAP7_75t_L g15160 ( 
.A(n_14855),
.Y(n_15160)
);

NAND2xp5_ASAP7_75t_L g15161 ( 
.A(n_14751),
.B(n_7764),
.Y(n_15161)
);

OR2x2_ASAP7_75t_L g15162 ( 
.A(n_14777),
.B(n_7764),
.Y(n_15162)
);

NAND2xp5_ASAP7_75t_L g15163 ( 
.A(n_14767),
.B(n_14890),
.Y(n_15163)
);

AND2x2_ASAP7_75t_L g15164 ( 
.A(n_14746),
.B(n_6327),
.Y(n_15164)
);

AND2x2_ASAP7_75t_L g15165 ( 
.A(n_14755),
.B(n_6327),
.Y(n_15165)
);

NAND2xp5_ASAP7_75t_L g15166 ( 
.A(n_14745),
.B(n_7764),
.Y(n_15166)
);

INVx1_ASAP7_75t_SL g15167 ( 
.A(n_14868),
.Y(n_15167)
);

INVx2_ASAP7_75t_L g15168 ( 
.A(n_14689),
.Y(n_15168)
);

INVx1_ASAP7_75t_L g15169 ( 
.A(n_14821),
.Y(n_15169)
);

INVxp67_ASAP7_75t_L g15170 ( 
.A(n_14870),
.Y(n_15170)
);

INVx1_ASAP7_75t_L g15171 ( 
.A(n_14829),
.Y(n_15171)
);

INVx1_ASAP7_75t_L g15172 ( 
.A(n_14896),
.Y(n_15172)
);

INVx1_ASAP7_75t_L g15173 ( 
.A(n_14764),
.Y(n_15173)
);

OR2x2_ASAP7_75t_L g15174 ( 
.A(n_14687),
.B(n_7764),
.Y(n_15174)
);

OR2x6_ASAP7_75t_L g15175 ( 
.A(n_14916),
.B(n_7346),
.Y(n_15175)
);

INVx1_ASAP7_75t_L g15176 ( 
.A(n_14733),
.Y(n_15176)
);

INVx1_ASAP7_75t_L g15177 ( 
.A(n_14893),
.Y(n_15177)
);

AO21x1_ASAP7_75t_L g15178 ( 
.A1(n_14872),
.A2(n_8418),
.B(n_8385),
.Y(n_15178)
);

NAND2xp5_ASAP7_75t_L g15179 ( 
.A(n_14928),
.B(n_7764),
.Y(n_15179)
);

INVx1_ASAP7_75t_L g15180 ( 
.A(n_14909),
.Y(n_15180)
);

NAND2xp33_ASAP7_75t_SL g15181 ( 
.A(n_14683),
.B(n_6703),
.Y(n_15181)
);

INVx1_ASAP7_75t_SL g15182 ( 
.A(n_14828),
.Y(n_15182)
);

INVx1_ASAP7_75t_L g15183 ( 
.A(n_14926),
.Y(n_15183)
);

NAND2xp5_ASAP7_75t_L g15184 ( 
.A(n_14939),
.B(n_14942),
.Y(n_15184)
);

AND2x2_ASAP7_75t_L g15185 ( 
.A(n_14932),
.B(n_6348),
.Y(n_15185)
);

INVx2_ASAP7_75t_SL g15186 ( 
.A(n_14802),
.Y(n_15186)
);

INVx1_ASAP7_75t_L g15187 ( 
.A(n_14938),
.Y(n_15187)
);

AND2x2_ASAP7_75t_L g15188 ( 
.A(n_14853),
.B(n_6348),
.Y(n_15188)
);

INVx2_ASAP7_75t_L g15189 ( 
.A(n_14936),
.Y(n_15189)
);

BUFx2_ASAP7_75t_L g15190 ( 
.A(n_14747),
.Y(n_15190)
);

INVx1_ASAP7_75t_L g15191 ( 
.A(n_14917),
.Y(n_15191)
);

INVx1_ASAP7_75t_SL g15192 ( 
.A(n_14710),
.Y(n_15192)
);

HB1xp67_ASAP7_75t_L g15193 ( 
.A(n_14818),
.Y(n_15193)
);

NAND2xp5_ASAP7_75t_L g15194 ( 
.A(n_14944),
.B(n_7764),
.Y(n_15194)
);

BUFx3_ASAP7_75t_L g15195 ( 
.A(n_14876),
.Y(n_15195)
);

AND2x4_ASAP7_75t_L g15196 ( 
.A(n_14715),
.B(n_9092),
.Y(n_15196)
);

OR2x6_ASAP7_75t_L g15197 ( 
.A(n_14765),
.B(n_7346),
.Y(n_15197)
);

HB1xp67_ASAP7_75t_L g15198 ( 
.A(n_14838),
.Y(n_15198)
);

AOI21xp33_ASAP7_75t_L g15199 ( 
.A1(n_14673),
.A2(n_7263),
.B(n_7239),
.Y(n_15199)
);

NOR3xp33_ASAP7_75t_SL g15200 ( 
.A(n_14721),
.B(n_8249),
.C(n_8043),
.Y(n_15200)
);

NAND2xp5_ASAP7_75t_SL g15201 ( 
.A(n_14708),
.B(n_7173),
.Y(n_15201)
);

INVx1_ASAP7_75t_L g15202 ( 
.A(n_14839),
.Y(n_15202)
);

NOR2xp33_ASAP7_75t_R g15203 ( 
.A(n_14769),
.B(n_6703),
.Y(n_15203)
);

INVx1_ASAP7_75t_L g15204 ( 
.A(n_14778),
.Y(n_15204)
);

NOR2xp33_ASAP7_75t_L g15205 ( 
.A(n_14863),
.B(n_7239),
.Y(n_15205)
);

AND2x2_ASAP7_75t_L g15206 ( 
.A(n_14680),
.B(n_6348),
.Y(n_15206)
);

AND2x2_ASAP7_75t_L g15207 ( 
.A(n_14794),
.B(n_6350),
.Y(n_15207)
);

AND2x2_ASAP7_75t_L g15208 ( 
.A(n_14791),
.B(n_6350),
.Y(n_15208)
);

INVx2_ASAP7_75t_L g15209 ( 
.A(n_14660),
.Y(n_15209)
);

NOR3xp33_ASAP7_75t_L g15210 ( 
.A(n_14912),
.B(n_14814),
.C(n_14809),
.Y(n_15210)
);

AND2x2_ASAP7_75t_L g15211 ( 
.A(n_14768),
.B(n_6350),
.Y(n_15211)
);

INVx1_ASAP7_75t_L g15212 ( 
.A(n_14815),
.Y(n_15212)
);

INVx1_ASAP7_75t_L g15213 ( 
.A(n_14852),
.Y(n_15213)
);

NAND2xp5_ASAP7_75t_L g15214 ( 
.A(n_14753),
.B(n_14854),
.Y(n_15214)
);

OR2x2_ASAP7_75t_L g15215 ( 
.A(n_14830),
.B(n_7764),
.Y(n_15215)
);

NOR3xp33_ASAP7_75t_L g15216 ( 
.A(n_14905),
.B(n_7514),
.C(n_7503),
.Y(n_15216)
);

NOR2xp33_ASAP7_75t_R g15217 ( 
.A(n_14875),
.B(n_6703),
.Y(n_15217)
);

NAND2xp5_ASAP7_75t_L g15218 ( 
.A(n_14949),
.B(n_14760),
.Y(n_15218)
);

INVx1_ASAP7_75t_L g15219 ( 
.A(n_14820),
.Y(n_15219)
);

INVx2_ASAP7_75t_L g15220 ( 
.A(n_14660),
.Y(n_15220)
);

NAND2xp5_ASAP7_75t_L g15221 ( 
.A(n_14941),
.B(n_7816),
.Y(n_15221)
);

OAI33xp33_ASAP7_75t_L g15222 ( 
.A1(n_14668),
.A2(n_7631),
.A3(n_7647),
.B1(n_7663),
.B2(n_7651),
.B3(n_7617),
.Y(n_15222)
);

OR2x2_ASAP7_75t_L g15223 ( 
.A(n_14763),
.B(n_7816),
.Y(n_15223)
);

AND2x2_ASAP7_75t_L g15224 ( 
.A(n_14754),
.B(n_6419),
.Y(n_15224)
);

NOR2x1p5_ASAP7_75t_L g15225 ( 
.A(n_14675),
.B(n_14940),
.Y(n_15225)
);

AOI22xp33_ASAP7_75t_L g15226 ( 
.A1(n_14705),
.A2(n_8224),
.B1(n_8209),
.B2(n_7359),
.Y(n_15226)
);

OAI21x1_ASAP7_75t_L g15227 ( 
.A1(n_14711),
.A2(n_8434),
.B(n_8427),
.Y(n_15227)
);

AND2x2_ASAP7_75t_L g15228 ( 
.A(n_14758),
.B(n_6419),
.Y(n_15228)
);

AND2x2_ASAP7_75t_L g15229 ( 
.A(n_14813),
.B(n_6419),
.Y(n_15229)
);

INVx1_ASAP7_75t_L g15230 ( 
.A(n_14892),
.Y(n_15230)
);

INVx1_ASAP7_75t_SL g15231 ( 
.A(n_14889),
.Y(n_15231)
);

INVx1_ASAP7_75t_L g15232 ( 
.A(n_14834),
.Y(n_15232)
);

INVxp67_ASAP7_75t_SL g15233 ( 
.A(n_14878),
.Y(n_15233)
);

NAND2xp5_ASAP7_75t_L g15234 ( 
.A(n_14749),
.B(n_7816),
.Y(n_15234)
);

INVx1_ASAP7_75t_L g15235 ( 
.A(n_14888),
.Y(n_15235)
);

NAND2xp5_ASAP7_75t_L g15236 ( 
.A(n_14748),
.B(n_7816),
.Y(n_15236)
);

INVx1_ASAP7_75t_L g15237 ( 
.A(n_14757),
.Y(n_15237)
);

NOR2xp67_ASAP7_75t_SL g15238 ( 
.A(n_14833),
.B(n_6939),
.Y(n_15238)
);

NAND2xp5_ASAP7_75t_L g15239 ( 
.A(n_14738),
.B(n_7816),
.Y(n_15239)
);

INVx2_ASAP7_75t_L g15240 ( 
.A(n_14675),
.Y(n_15240)
);

INVx1_ASAP7_75t_L g15241 ( 
.A(n_14808),
.Y(n_15241)
);

INVx1_ASAP7_75t_SL g15242 ( 
.A(n_14864),
.Y(n_15242)
);

OR2x2_ASAP7_75t_L g15243 ( 
.A(n_14874),
.B(n_7816),
.Y(n_15243)
);

AND2x2_ASAP7_75t_L g15244 ( 
.A(n_14671),
.B(n_6423),
.Y(n_15244)
);

AND2x2_ASAP7_75t_L g15245 ( 
.A(n_14713),
.B(n_6423),
.Y(n_15245)
);

BUFx2_ASAP7_75t_L g15246 ( 
.A(n_14810),
.Y(n_15246)
);

INVxp67_ASAP7_75t_SL g15247 ( 
.A(n_14851),
.Y(n_15247)
);

OAI21xp33_ASAP7_75t_SL g15248 ( 
.A1(n_14679),
.A2(n_8434),
.B(n_8427),
.Y(n_15248)
);

NOR2xp33_ASAP7_75t_L g15249 ( 
.A(n_14685),
.B(n_14665),
.Y(n_15249)
);

BUFx2_ASAP7_75t_L g15250 ( 
.A(n_14940),
.Y(n_15250)
);

OAI21xp5_ASAP7_75t_L g15251 ( 
.A1(n_14880),
.A2(n_8618),
.B(n_8540),
.Y(n_15251)
);

NOR2xp33_ASAP7_75t_L g15252 ( 
.A(n_14739),
.B(n_7239),
.Y(n_15252)
);

AND2x2_ASAP7_75t_L g15253 ( 
.A(n_14930),
.B(n_6423),
.Y(n_15253)
);

NAND2xp5_ASAP7_75t_L g15254 ( 
.A(n_14871),
.B(n_7816),
.Y(n_15254)
);

NAND2xp5_ASAP7_75t_SL g15255 ( 
.A(n_14902),
.B(n_7173),
.Y(n_15255)
);

AND2x2_ASAP7_75t_L g15256 ( 
.A(n_14867),
.B(n_6480),
.Y(n_15256)
);

INVx1_ASAP7_75t_L g15257 ( 
.A(n_14694),
.Y(n_15257)
);

AND2x2_ASAP7_75t_L g15258 ( 
.A(n_14867),
.B(n_6480),
.Y(n_15258)
);

INVx2_ASAP7_75t_L g15259 ( 
.A(n_14835),
.Y(n_15259)
);

INVx2_ASAP7_75t_L g15260 ( 
.A(n_14835),
.Y(n_15260)
);

INVx1_ASAP7_75t_L g15261 ( 
.A(n_14684),
.Y(n_15261)
);

AND2x2_ASAP7_75t_L g15262 ( 
.A(n_14832),
.B(n_6480),
.Y(n_15262)
);

BUFx2_ASAP7_75t_L g15263 ( 
.A(n_14832),
.Y(n_15263)
);

INVx1_ASAP7_75t_L g15264 ( 
.A(n_14772),
.Y(n_15264)
);

BUFx2_ASAP7_75t_L g15265 ( 
.A(n_14910),
.Y(n_15265)
);

AND4x1_ASAP7_75t_L g15266 ( 
.A(n_14730),
.B(n_8032),
.C(n_8072),
.D(n_8061),
.Y(n_15266)
);

NAND2xp5_ASAP7_75t_L g15267 ( 
.A(n_14712),
.B(n_7816),
.Y(n_15267)
);

NOR2xp33_ASAP7_75t_L g15268 ( 
.A(n_14901),
.B(n_7263),
.Y(n_15268)
);

INVx1_ASAP7_75t_L g15269 ( 
.A(n_14846),
.Y(n_15269)
);

AND2x2_ASAP7_75t_L g15270 ( 
.A(n_14873),
.B(n_6504),
.Y(n_15270)
);

INVx4_ASAP7_75t_L g15271 ( 
.A(n_14972),
.Y(n_15271)
);

AND2x2_ASAP7_75t_L g15272 ( 
.A(n_14982),
.B(n_7171),
.Y(n_15272)
);

INVx1_ASAP7_75t_SL g15273 ( 
.A(n_15003),
.Y(n_15273)
);

AND2x2_ASAP7_75t_L g15274 ( 
.A(n_14972),
.B(n_14979),
.Y(n_15274)
);

NAND2xp5_ASAP7_75t_L g15275 ( 
.A(n_14972),
.B(n_7418),
.Y(n_15275)
);

INVx1_ASAP7_75t_L g15276 ( 
.A(n_15034),
.Y(n_15276)
);

NAND2xp5_ASAP7_75t_L g15277 ( 
.A(n_14957),
.B(n_7418),
.Y(n_15277)
);

INVx3_ASAP7_75t_L g15278 ( 
.A(n_14957),
.Y(n_15278)
);

NAND2xp5_ASAP7_75t_L g15279 ( 
.A(n_14979),
.B(n_15044),
.Y(n_15279)
);

INVx1_ASAP7_75t_SL g15280 ( 
.A(n_15017),
.Y(n_15280)
);

AOI22xp33_ASAP7_75t_L g15281 ( 
.A1(n_15039),
.A2(n_7359),
.B1(n_7358),
.B2(n_7263),
.Y(n_15281)
);

NAND3x1_ASAP7_75t_L g15282 ( 
.A(n_14950),
.B(n_14951),
.C(n_15014),
.Y(n_15282)
);

AOI22xp5_ASAP7_75t_L g15283 ( 
.A1(n_15244),
.A2(n_7358),
.B1(n_7359),
.B2(n_5044),
.Y(n_15283)
);

AND2x2_ASAP7_75t_L g15284 ( 
.A(n_14961),
.B(n_7171),
.Y(n_15284)
);

NAND2xp5_ASAP7_75t_L g15285 ( 
.A(n_14977),
.B(n_7418),
.Y(n_15285)
);

CKINVDCx16_ASAP7_75t_R g15286 ( 
.A(n_14952),
.Y(n_15286)
);

AND2x2_ASAP7_75t_L g15287 ( 
.A(n_14980),
.B(n_7171),
.Y(n_15287)
);

INVx1_ASAP7_75t_L g15288 ( 
.A(n_14992),
.Y(n_15288)
);

OR2x2_ASAP7_75t_L g15289 ( 
.A(n_14991),
.B(n_7131),
.Y(n_15289)
);

NAND3x1_ASAP7_75t_L g15290 ( 
.A(n_14958),
.B(n_7082),
.C(n_6540),
.Y(n_15290)
);

AND2x2_ASAP7_75t_L g15291 ( 
.A(n_14966),
.B(n_7171),
.Y(n_15291)
);

INVx1_ASAP7_75t_L g15292 ( 
.A(n_15004),
.Y(n_15292)
);

INVx1_ASAP7_75t_L g15293 ( 
.A(n_14994),
.Y(n_15293)
);

INVxp67_ASAP7_75t_L g15294 ( 
.A(n_15106),
.Y(n_15294)
);

OAI21x1_ASAP7_75t_L g15295 ( 
.A1(n_14962),
.A2(n_8618),
.B(n_8540),
.Y(n_15295)
);

INVx1_ASAP7_75t_L g15296 ( 
.A(n_15263),
.Y(n_15296)
);

INVx1_ASAP7_75t_L g15297 ( 
.A(n_15051),
.Y(n_15297)
);

INVx1_ASAP7_75t_L g15298 ( 
.A(n_15131),
.Y(n_15298)
);

INVx1_ASAP7_75t_L g15299 ( 
.A(n_14975),
.Y(n_15299)
);

NAND3x1_ASAP7_75t_L g15300 ( 
.A(n_14960),
.B(n_6540),
.C(n_6504),
.Y(n_15300)
);

AND2x4_ASAP7_75t_L g15301 ( 
.A(n_15027),
.B(n_9166),
.Y(n_15301)
);

INVx1_ASAP7_75t_L g15302 ( 
.A(n_15120),
.Y(n_15302)
);

NAND2xp5_ASAP7_75t_L g15303 ( 
.A(n_15159),
.B(n_7263),
.Y(n_15303)
);

AND2x2_ASAP7_75t_L g15304 ( 
.A(n_14953),
.B(n_7171),
.Y(n_15304)
);

AOI22xp33_ASAP7_75t_L g15305 ( 
.A1(n_15224),
.A2(n_7359),
.B1(n_7358),
.B2(n_7267),
.Y(n_15305)
);

NAND2xp5_ASAP7_75t_L g15306 ( 
.A(n_14998),
.B(n_7267),
.Y(n_15306)
);

AOI22xp33_ASAP7_75t_SL g15307 ( 
.A1(n_14984),
.A2(n_15000),
.B1(n_15245),
.B2(n_15020),
.Y(n_15307)
);

INVx2_ASAP7_75t_L g15308 ( 
.A(n_14967),
.Y(n_15308)
);

OR2x2_ASAP7_75t_L g15309 ( 
.A(n_15018),
.B(n_8127),
.Y(n_15309)
);

NAND2xp5_ASAP7_75t_L g15310 ( 
.A(n_15114),
.B(n_7267),
.Y(n_15310)
);

NAND2xp5_ASAP7_75t_SL g15311 ( 
.A(n_15002),
.B(n_7173),
.Y(n_15311)
);

AND2x2_ASAP7_75t_L g15312 ( 
.A(n_15023),
.B(n_15006),
.Y(n_15312)
);

NOR2x1_ASAP7_75t_L g15313 ( 
.A(n_14965),
.B(n_7768),
.Y(n_15313)
);

OR2x2_ASAP7_75t_L g15314 ( 
.A(n_15028),
.B(n_8127),
.Y(n_15314)
);

OR2x2_ASAP7_75t_L g15315 ( 
.A(n_15125),
.B(n_8127),
.Y(n_15315)
);

OR2x2_ASAP7_75t_L g15316 ( 
.A(n_14955),
.B(n_8127),
.Y(n_15316)
);

INVx1_ASAP7_75t_L g15317 ( 
.A(n_15042),
.Y(n_15317)
);

CKINVDCx16_ASAP7_75t_R g15318 ( 
.A(n_14989),
.Y(n_15318)
);

INVx1_ASAP7_75t_L g15319 ( 
.A(n_15053),
.Y(n_15319)
);

INVx1_ASAP7_75t_L g15320 ( 
.A(n_15108),
.Y(n_15320)
);

AND2x2_ASAP7_75t_L g15321 ( 
.A(n_15133),
.B(n_7178),
.Y(n_15321)
);

INVx2_ASAP7_75t_L g15322 ( 
.A(n_15229),
.Y(n_15322)
);

AND2x2_ASAP7_75t_L g15323 ( 
.A(n_14986),
.B(n_7178),
.Y(n_15323)
);

INVx3_ASAP7_75t_L g15324 ( 
.A(n_15048),
.Y(n_15324)
);

INVx2_ASAP7_75t_SL g15325 ( 
.A(n_15008),
.Y(n_15325)
);

NAND2xp5_ASAP7_75t_L g15326 ( 
.A(n_14993),
.B(n_7267),
.Y(n_15326)
);

INVx1_ASAP7_75t_L g15327 ( 
.A(n_15250),
.Y(n_15327)
);

INVx1_ASAP7_75t_L g15328 ( 
.A(n_15153),
.Y(n_15328)
);

AND2x2_ASAP7_75t_L g15329 ( 
.A(n_14996),
.B(n_7178),
.Y(n_15329)
);

AND2x2_ASAP7_75t_L g15330 ( 
.A(n_15118),
.B(n_7178),
.Y(n_15330)
);

INVx1_ASAP7_75t_L g15331 ( 
.A(n_14990),
.Y(n_15331)
);

OR2x2_ASAP7_75t_L g15332 ( 
.A(n_15134),
.B(n_8127),
.Y(n_15332)
);

INVx1_ASAP7_75t_L g15333 ( 
.A(n_15070),
.Y(n_15333)
);

INVx1_ASAP7_75t_L g15334 ( 
.A(n_15047),
.Y(n_15334)
);

INVx1_ASAP7_75t_SL g15335 ( 
.A(n_15013),
.Y(n_15335)
);

BUFx6f_ASAP7_75t_L g15336 ( 
.A(n_14963),
.Y(n_15336)
);

INVx2_ASAP7_75t_L g15337 ( 
.A(n_15195),
.Y(n_15337)
);

NAND2xp5_ASAP7_75t_L g15338 ( 
.A(n_15016),
.B(n_7318),
.Y(n_15338)
);

OR2x2_ASAP7_75t_L g15339 ( 
.A(n_15126),
.B(n_8127),
.Y(n_15339)
);

INVx1_ASAP7_75t_L g15340 ( 
.A(n_15089),
.Y(n_15340)
);

INVx1_ASAP7_75t_SL g15341 ( 
.A(n_15032),
.Y(n_15341)
);

INVx1_ASAP7_75t_SL g15342 ( 
.A(n_14988),
.Y(n_15342)
);

INVxp67_ASAP7_75t_SL g15343 ( 
.A(n_14981),
.Y(n_15343)
);

OR2x2_ASAP7_75t_L g15344 ( 
.A(n_15024),
.B(n_8127),
.Y(n_15344)
);

AND2x2_ASAP7_75t_L g15345 ( 
.A(n_15119),
.B(n_15104),
.Y(n_15345)
);

NAND2xp5_ASAP7_75t_L g15346 ( 
.A(n_15182),
.B(n_7318),
.Y(n_15346)
);

INVx2_ASAP7_75t_L g15347 ( 
.A(n_15156),
.Y(n_15347)
);

BUFx2_ASAP7_75t_L g15348 ( 
.A(n_14997),
.Y(n_15348)
);

INVx3_ASAP7_75t_L g15349 ( 
.A(n_15197),
.Y(n_15349)
);

NAND2xp5_ASAP7_75t_L g15350 ( 
.A(n_15192),
.B(n_15193),
.Y(n_15350)
);

NAND2xp5_ASAP7_75t_L g15351 ( 
.A(n_15198),
.B(n_15154),
.Y(n_15351)
);

CKINVDCx14_ASAP7_75t_R g15352 ( 
.A(n_15101),
.Y(n_15352)
);

INVx1_ASAP7_75t_L g15353 ( 
.A(n_15019),
.Y(n_15353)
);

INVx1_ASAP7_75t_SL g15354 ( 
.A(n_14970),
.Y(n_15354)
);

AND2x4_ASAP7_75t_L g15355 ( 
.A(n_15030),
.B(n_9166),
.Y(n_15355)
);

OR2x2_ASAP7_75t_L g15356 ( 
.A(n_15012),
.B(n_7002),
.Y(n_15356)
);

AND2x2_ASAP7_75t_L g15357 ( 
.A(n_15121),
.B(n_7178),
.Y(n_15357)
);

INVx2_ASAP7_75t_L g15358 ( 
.A(n_15008),
.Y(n_15358)
);

AND2x2_ASAP7_75t_L g15359 ( 
.A(n_15128),
.B(n_7207),
.Y(n_15359)
);

NAND2xp5_ASAP7_75t_L g15360 ( 
.A(n_15060),
.B(n_7318),
.Y(n_15360)
);

INVx1_ASAP7_75t_L g15361 ( 
.A(n_15184),
.Y(n_15361)
);

NOR2xp33_ASAP7_75t_L g15362 ( 
.A(n_14978),
.B(n_7318),
.Y(n_15362)
);

INVx2_ASAP7_75t_SL g15363 ( 
.A(n_15026),
.Y(n_15363)
);

INVx1_ASAP7_75t_L g15364 ( 
.A(n_15124),
.Y(n_15364)
);

INVx1_ASAP7_75t_L g15365 ( 
.A(n_15065),
.Y(n_15365)
);

INVx2_ASAP7_75t_L g15366 ( 
.A(n_15225),
.Y(n_15366)
);

INVx1_ASAP7_75t_L g15367 ( 
.A(n_15246),
.Y(n_15367)
);

INVx1_ASAP7_75t_L g15368 ( 
.A(n_15072),
.Y(n_15368)
);

OR2x2_ASAP7_75t_L g15369 ( 
.A(n_14968),
.B(n_15091),
.Y(n_15369)
);

INVx1_ASAP7_75t_L g15370 ( 
.A(n_15142),
.Y(n_15370)
);

INVx1_ASAP7_75t_L g15371 ( 
.A(n_15142),
.Y(n_15371)
);

INVx2_ASAP7_75t_L g15372 ( 
.A(n_15190),
.Y(n_15372)
);

INVx1_ASAP7_75t_L g15373 ( 
.A(n_15142),
.Y(n_15373)
);

AND2x4_ASAP7_75t_L g15374 ( 
.A(n_15007),
.B(n_9168),
.Y(n_15374)
);

INVx1_ASAP7_75t_L g15375 ( 
.A(n_15090),
.Y(n_15375)
);

AND2x2_ASAP7_75t_L g15376 ( 
.A(n_15079),
.B(n_7207),
.Y(n_15376)
);

AOI22xp33_ASAP7_75t_L g15377 ( 
.A1(n_15264),
.A2(n_7359),
.B1(n_7358),
.B2(n_7326),
.Y(n_15377)
);

AOI21xp5_ASAP7_75t_SL g15378 ( 
.A1(n_15022),
.A2(n_7975),
.B(n_7963),
.Y(n_15378)
);

AND2x2_ASAP7_75t_L g15379 ( 
.A(n_15080),
.B(n_15088),
.Y(n_15379)
);

BUFx2_ASAP7_75t_L g15380 ( 
.A(n_15117),
.Y(n_15380)
);

INVx1_ASAP7_75t_L g15381 ( 
.A(n_14971),
.Y(n_15381)
);

INVx1_ASAP7_75t_L g15382 ( 
.A(n_15075),
.Y(n_15382)
);

INVx1_ASAP7_75t_L g15383 ( 
.A(n_14959),
.Y(n_15383)
);

NAND2xp5_ASAP7_75t_L g15384 ( 
.A(n_15160),
.B(n_7326),
.Y(n_15384)
);

INVx2_ASAP7_75t_L g15385 ( 
.A(n_15197),
.Y(n_15385)
);

HB1xp67_ASAP7_75t_L g15386 ( 
.A(n_15021),
.Y(n_15386)
);

CKINVDCx16_ASAP7_75t_R g15387 ( 
.A(n_14976),
.Y(n_15387)
);

INVx1_ASAP7_75t_L g15388 ( 
.A(n_15068),
.Y(n_15388)
);

AND2x2_ASAP7_75t_L g15389 ( 
.A(n_15067),
.B(n_7207),
.Y(n_15389)
);

NAND2xp5_ASAP7_75t_L g15390 ( 
.A(n_15171),
.B(n_7326),
.Y(n_15390)
);

INVx2_ASAP7_75t_L g15391 ( 
.A(n_15175),
.Y(n_15391)
);

OAI22xp5_ASAP7_75t_L g15392 ( 
.A1(n_14974),
.A2(n_8139),
.B1(n_8006),
.B2(n_7187),
.Y(n_15392)
);

AND2x4_ASAP7_75t_L g15393 ( 
.A(n_15011),
.B(n_9168),
.Y(n_15393)
);

INVx1_ASAP7_75t_L g15394 ( 
.A(n_15074),
.Y(n_15394)
);

INVx2_ASAP7_75t_L g15395 ( 
.A(n_15175),
.Y(n_15395)
);

AND2x2_ASAP7_75t_L g15396 ( 
.A(n_15149),
.B(n_7207),
.Y(n_15396)
);

NOR2xp33_ASAP7_75t_L g15397 ( 
.A(n_15109),
.B(n_7326),
.Y(n_15397)
);

HB1xp67_ASAP7_75t_L g15398 ( 
.A(n_15077),
.Y(n_15398)
);

NAND2xp5_ASAP7_75t_L g15399 ( 
.A(n_15169),
.B(n_7329),
.Y(n_15399)
);

INVx1_ASAP7_75t_L g15400 ( 
.A(n_15035),
.Y(n_15400)
);

INVx1_ASAP7_75t_SL g15401 ( 
.A(n_15025),
.Y(n_15401)
);

INVx2_ASAP7_75t_L g15402 ( 
.A(n_15189),
.Y(n_15402)
);

INVx3_ASAP7_75t_L g15403 ( 
.A(n_15135),
.Y(n_15403)
);

AND2x2_ASAP7_75t_L g15404 ( 
.A(n_15093),
.B(n_7207),
.Y(n_15404)
);

INVx2_ASAP7_75t_L g15405 ( 
.A(n_15155),
.Y(n_15405)
);

OR2x2_ASAP7_75t_L g15406 ( 
.A(n_15241),
.B(n_7002),
.Y(n_15406)
);

INVx1_ASAP7_75t_L g15407 ( 
.A(n_14983),
.Y(n_15407)
);

INVx1_ASAP7_75t_SL g15408 ( 
.A(n_15009),
.Y(n_15408)
);

NOR2xp33_ASAP7_75t_L g15409 ( 
.A(n_15158),
.B(n_15141),
.Y(n_15409)
);

INVx1_ASAP7_75t_L g15410 ( 
.A(n_14987),
.Y(n_15410)
);

NOR2xp33_ASAP7_75t_SL g15411 ( 
.A(n_15033),
.B(n_14964),
.Y(n_15411)
);

NAND2x1_ASAP7_75t_L g15412 ( 
.A(n_15172),
.B(n_7977),
.Y(n_15412)
);

INVx2_ASAP7_75t_L g15413 ( 
.A(n_15173),
.Y(n_15413)
);

INVx1_ASAP7_75t_L g15414 ( 
.A(n_14995),
.Y(n_15414)
);

CKINVDCx16_ASAP7_75t_R g15415 ( 
.A(n_15167),
.Y(n_15415)
);

AND2x2_ASAP7_75t_L g15416 ( 
.A(n_15211),
.B(n_7233),
.Y(n_15416)
);

NOR2xp33_ASAP7_75t_L g15417 ( 
.A(n_15143),
.B(n_7329),
.Y(n_15417)
);

AND2x2_ASAP7_75t_L g15418 ( 
.A(n_15164),
.B(n_7233),
.Y(n_15418)
);

NOR2xp33_ASAP7_75t_L g15419 ( 
.A(n_15148),
.B(n_15043),
.Y(n_15419)
);

INVx2_ASAP7_75t_SL g15420 ( 
.A(n_15094),
.Y(n_15420)
);

INVx1_ASAP7_75t_L g15421 ( 
.A(n_15130),
.Y(n_15421)
);

HB1xp67_ASAP7_75t_L g15422 ( 
.A(n_15237),
.Y(n_15422)
);

INVxp67_ASAP7_75t_SL g15423 ( 
.A(n_15163),
.Y(n_15423)
);

INVxp67_ASAP7_75t_L g15424 ( 
.A(n_15001),
.Y(n_15424)
);

AOI22xp33_ASAP7_75t_L g15425 ( 
.A1(n_15269),
.A2(n_7359),
.B1(n_7358),
.B2(n_7329),
.Y(n_15425)
);

AO22x1_ASAP7_75t_L g15426 ( 
.A1(n_14954),
.A2(n_7132),
.B1(n_6992),
.B2(n_6080),
.Y(n_15426)
);

INVx1_ASAP7_75t_L g15427 ( 
.A(n_15145),
.Y(n_15427)
);

AND2x2_ASAP7_75t_L g15428 ( 
.A(n_15165),
.B(n_7233),
.Y(n_15428)
);

AND2x2_ASAP7_75t_L g15429 ( 
.A(n_15138),
.B(n_7233),
.Y(n_15429)
);

INVx2_ASAP7_75t_L g15430 ( 
.A(n_15066),
.Y(n_15430)
);

INVx1_ASAP7_75t_L g15431 ( 
.A(n_15105),
.Y(n_15431)
);

INVxp67_ASAP7_75t_L g15432 ( 
.A(n_14956),
.Y(n_15432)
);

NAND4xp75_ASAP7_75t_L g15433 ( 
.A(n_14999),
.B(n_7498),
.C(n_7861),
.D(n_7133),
.Y(n_15433)
);

INVx1_ASAP7_75t_L g15434 ( 
.A(n_15259),
.Y(n_15434)
);

NOR2x1_ASAP7_75t_L g15435 ( 
.A(n_15005),
.B(n_7963),
.Y(n_15435)
);

INVx1_ASAP7_75t_L g15436 ( 
.A(n_15260),
.Y(n_15436)
);

AOI22xp33_ASAP7_75t_L g15437 ( 
.A1(n_15231),
.A2(n_7329),
.B1(n_7372),
.B2(n_7340),
.Y(n_15437)
);

OR2x2_ASAP7_75t_L g15438 ( 
.A(n_15100),
.B(n_7036),
.Y(n_15438)
);

AOI222xp33_ASAP7_75t_SL g15439 ( 
.A1(n_15102),
.A2(n_8067),
.B1(n_7977),
.B2(n_8114),
.C1(n_8033),
.C2(n_8009),
.Y(n_15439)
);

NAND2xp5_ASAP7_75t_L g15440 ( 
.A(n_15055),
.B(n_7340),
.Y(n_15440)
);

INVx1_ASAP7_75t_L g15441 ( 
.A(n_15123),
.Y(n_15441)
);

AND2x2_ASAP7_75t_L g15442 ( 
.A(n_15206),
.B(n_7233),
.Y(n_15442)
);

INVx1_ASAP7_75t_L g15443 ( 
.A(n_15037),
.Y(n_15443)
);

OR2x2_ASAP7_75t_L g15444 ( 
.A(n_15010),
.B(n_7036),
.Y(n_15444)
);

INVx1_ASAP7_75t_L g15445 ( 
.A(n_15036),
.Y(n_15445)
);

BUFx3_ASAP7_75t_L g15446 ( 
.A(n_15150),
.Y(n_15446)
);

INVx1_ASAP7_75t_L g15447 ( 
.A(n_15209),
.Y(n_15447)
);

INVx1_ASAP7_75t_SL g15448 ( 
.A(n_15069),
.Y(n_15448)
);

NAND2xp5_ASAP7_75t_L g15449 ( 
.A(n_15029),
.B(n_7340),
.Y(n_15449)
);

INVx1_ASAP7_75t_L g15450 ( 
.A(n_15220),
.Y(n_15450)
);

AND2x2_ASAP7_75t_L g15451 ( 
.A(n_15208),
.B(n_15262),
.Y(n_15451)
);

OAI22xp5_ASAP7_75t_L g15452 ( 
.A1(n_14985),
.A2(n_8139),
.B1(n_8006),
.B2(n_7187),
.Y(n_15452)
);

OR2x2_ASAP7_75t_L g15453 ( 
.A(n_15218),
.B(n_7047),
.Y(n_15453)
);

NAND2xp5_ASAP7_75t_L g15454 ( 
.A(n_15040),
.B(n_15210),
.Y(n_15454)
);

AND2x2_ASAP7_75t_L g15455 ( 
.A(n_15200),
.B(n_7313),
.Y(n_15455)
);

CKINVDCx16_ASAP7_75t_R g15456 ( 
.A(n_15127),
.Y(n_15456)
);

INVx1_ASAP7_75t_L g15457 ( 
.A(n_15240),
.Y(n_15457)
);

INVx1_ASAP7_75t_L g15458 ( 
.A(n_15038),
.Y(n_15458)
);

AND2x2_ASAP7_75t_L g15459 ( 
.A(n_15188),
.B(n_7313),
.Y(n_15459)
);

INVx2_ASAP7_75t_L g15460 ( 
.A(n_15054),
.Y(n_15460)
);

AOI22xp33_ASAP7_75t_L g15461 ( 
.A1(n_15235),
.A2(n_7340),
.B1(n_7373),
.B2(n_7372),
.Y(n_15461)
);

CKINVDCx16_ASAP7_75t_R g15462 ( 
.A(n_15052),
.Y(n_15462)
);

INVx1_ASAP7_75t_L g15463 ( 
.A(n_15041),
.Y(n_15463)
);

NAND2xp5_ASAP7_75t_L g15464 ( 
.A(n_15045),
.B(n_7372),
.Y(n_15464)
);

INVx1_ASAP7_75t_SL g15465 ( 
.A(n_15115),
.Y(n_15465)
);

INVx1_ASAP7_75t_L g15466 ( 
.A(n_15132),
.Y(n_15466)
);

INVx1_ASAP7_75t_L g15467 ( 
.A(n_15031),
.Y(n_15467)
);

NAND2xp5_ASAP7_75t_L g15468 ( 
.A(n_15202),
.B(n_7372),
.Y(n_15468)
);

AND2x2_ASAP7_75t_L g15469 ( 
.A(n_15256),
.B(n_7313),
.Y(n_15469)
);

AND2x4_ASAP7_75t_SL g15470 ( 
.A(n_15046),
.B(n_6422),
.Y(n_15470)
);

INVx1_ASAP7_75t_L g15471 ( 
.A(n_15204),
.Y(n_15471)
);

HB1xp67_ASAP7_75t_L g15472 ( 
.A(n_15170),
.Y(n_15472)
);

OR2x2_ASAP7_75t_L g15473 ( 
.A(n_15232),
.B(n_7047),
.Y(n_15473)
);

INVx1_ASAP7_75t_L g15474 ( 
.A(n_15212),
.Y(n_15474)
);

INVx1_ASAP7_75t_L g15475 ( 
.A(n_15056),
.Y(n_15475)
);

OA21x2_ASAP7_75t_L g15476 ( 
.A1(n_15219),
.A2(n_8925),
.B(n_8870),
.Y(n_15476)
);

AND2x2_ASAP7_75t_L g15477 ( 
.A(n_15258),
.B(n_7313),
.Y(n_15477)
);

INVx1_ASAP7_75t_L g15478 ( 
.A(n_15086),
.Y(n_15478)
);

OAI22xp5_ASAP7_75t_SL g15479 ( 
.A1(n_14969),
.A2(n_7132),
.B1(n_6992),
.B2(n_8006),
.Y(n_15479)
);

AND2x2_ASAP7_75t_L g15480 ( 
.A(n_15185),
.B(n_7313),
.Y(n_15480)
);

INVx1_ASAP7_75t_SL g15481 ( 
.A(n_15139),
.Y(n_15481)
);

AOI22xp5_ASAP7_75t_L g15482 ( 
.A1(n_15233),
.A2(n_7975),
.B1(n_8064),
.B2(n_7963),
.Y(n_15482)
);

NAND2xp5_ASAP7_75t_L g15483 ( 
.A(n_15137),
.B(n_7373),
.Y(n_15483)
);

NAND2xp5_ASAP7_75t_L g15484 ( 
.A(n_15177),
.B(n_7373),
.Y(n_15484)
);

INVx4_ASAP7_75t_L g15485 ( 
.A(n_15186),
.Y(n_15485)
);

NOR2x1_ASAP7_75t_L g15486 ( 
.A(n_15180),
.B(n_7963),
.Y(n_15486)
);

BUFx12f_ASAP7_75t_L g15487 ( 
.A(n_15111),
.Y(n_15487)
);

OAI22xp5_ASAP7_75t_L g15488 ( 
.A1(n_15230),
.A2(n_8139),
.B1(n_8006),
.B2(n_7187),
.Y(n_15488)
);

NOR2xp33_ASAP7_75t_L g15489 ( 
.A(n_15242),
.B(n_7373),
.Y(n_15489)
);

AND2x2_ASAP7_75t_L g15490 ( 
.A(n_15049),
.B(n_7445),
.Y(n_15490)
);

INVx1_ASAP7_75t_L g15491 ( 
.A(n_15087),
.Y(n_15491)
);

INVx3_ASAP7_75t_SL g15492 ( 
.A(n_15098),
.Y(n_15492)
);

AND2x2_ASAP7_75t_L g15493 ( 
.A(n_15253),
.B(n_7445),
.Y(n_15493)
);

OR2x2_ASAP7_75t_L g15494 ( 
.A(n_15214),
.B(n_7067),
.Y(n_15494)
);

AND2x2_ASAP7_75t_L g15495 ( 
.A(n_15270),
.B(n_7445),
.Y(n_15495)
);

INVx1_ASAP7_75t_L g15496 ( 
.A(n_15183),
.Y(n_15496)
);

AND2x2_ASAP7_75t_L g15497 ( 
.A(n_15061),
.B(n_7445),
.Y(n_15497)
);

INVx2_ASAP7_75t_L g15498 ( 
.A(n_15050),
.Y(n_15498)
);

AND2x2_ASAP7_75t_SL g15499 ( 
.A(n_15015),
.B(n_8023),
.Y(n_15499)
);

NOR2x1_ASAP7_75t_L g15500 ( 
.A(n_15187),
.B(n_7963),
.Y(n_15500)
);

INVx1_ASAP7_75t_L g15501 ( 
.A(n_15082),
.Y(n_15501)
);

OR2x2_ASAP7_75t_L g15502 ( 
.A(n_15085),
.B(n_7067),
.Y(n_15502)
);

NAND4xp75_ASAP7_75t_L g15503 ( 
.A(n_15191),
.B(n_7133),
.C(n_6627),
.D(n_6638),
.Y(n_15503)
);

INVx2_ASAP7_75t_L g15504 ( 
.A(n_15215),
.Y(n_15504)
);

INVx1_ASAP7_75t_SL g15505 ( 
.A(n_15203),
.Y(n_15505)
);

NOR2xp33_ASAP7_75t_L g15506 ( 
.A(n_15116),
.B(n_7386),
.Y(n_15506)
);

AND2x2_ASAP7_75t_L g15507 ( 
.A(n_15168),
.B(n_7445),
.Y(n_15507)
);

OR2x2_ASAP7_75t_L g15508 ( 
.A(n_15099),
.B(n_7930),
.Y(n_15508)
);

INVx2_ASAP7_75t_L g15509 ( 
.A(n_15084),
.Y(n_15509)
);

INVx1_ASAP7_75t_SL g15510 ( 
.A(n_15217),
.Y(n_15510)
);

HB1xp67_ASAP7_75t_L g15511 ( 
.A(n_15265),
.Y(n_15511)
);

INVx2_ASAP7_75t_L g15512 ( 
.A(n_15103),
.Y(n_15512)
);

INVx2_ASAP7_75t_L g15513 ( 
.A(n_15129),
.Y(n_15513)
);

INVx1_ASAP7_75t_L g15514 ( 
.A(n_15083),
.Y(n_15514)
);

OAI22xp5_ASAP7_75t_L g15515 ( 
.A1(n_15176),
.A2(n_8139),
.B1(n_8006),
.B2(n_7187),
.Y(n_15515)
);

INVx1_ASAP7_75t_L g15516 ( 
.A(n_15095),
.Y(n_15516)
);

NAND2xp5_ASAP7_75t_SL g15517 ( 
.A(n_14973),
.B(n_7173),
.Y(n_15517)
);

NAND3xp33_ASAP7_75t_L g15518 ( 
.A(n_15257),
.B(n_7390),
.C(n_7386),
.Y(n_15518)
);

NAND2xp5_ASAP7_75t_L g15519 ( 
.A(n_15092),
.B(n_7386),
.Y(n_15519)
);

INVx2_ASAP7_75t_L g15520 ( 
.A(n_15063),
.Y(n_15520)
);

INVx1_ASAP7_75t_L g15521 ( 
.A(n_15247),
.Y(n_15521)
);

INVx1_ASAP7_75t_L g15522 ( 
.A(n_15057),
.Y(n_15522)
);

INVx1_ASAP7_75t_SL g15523 ( 
.A(n_15181),
.Y(n_15523)
);

INVx3_ASAP7_75t_L g15524 ( 
.A(n_15078),
.Y(n_15524)
);

CKINVDCx16_ASAP7_75t_R g15525 ( 
.A(n_15213),
.Y(n_15525)
);

AND2x2_ASAP7_75t_L g15526 ( 
.A(n_15207),
.B(n_15228),
.Y(n_15526)
);

AND2x2_ASAP7_75t_L g15527 ( 
.A(n_15144),
.B(n_7454),
.Y(n_15527)
);

AND2x2_ASAP7_75t_L g15528 ( 
.A(n_15249),
.B(n_7454),
.Y(n_15528)
);

AOI22xp33_ASAP7_75t_L g15529 ( 
.A1(n_15261),
.A2(n_7386),
.B1(n_7396),
.B2(n_7390),
.Y(n_15529)
);

AND2x2_ASAP7_75t_L g15530 ( 
.A(n_15058),
.B(n_7454),
.Y(n_15530)
);

OR2x2_ASAP7_75t_L g15531 ( 
.A(n_15112),
.B(n_7930),
.Y(n_15531)
);

AND2x2_ASAP7_75t_L g15532 ( 
.A(n_15238),
.B(n_7454),
.Y(n_15532)
);

NOR2xp33_ASAP7_75t_L g15533 ( 
.A(n_15266),
.B(n_7390),
.Y(n_15533)
);

INVx1_ASAP7_75t_L g15534 ( 
.A(n_15113),
.Y(n_15534)
);

INVx1_ASAP7_75t_SL g15535 ( 
.A(n_15122),
.Y(n_15535)
);

A2O1A1Ixp33_ASAP7_75t_L g15536 ( 
.A1(n_15521),
.A2(n_15205),
.B(n_15248),
.C(n_15140),
.Y(n_15536)
);

AOI21xp33_ASAP7_75t_L g15537 ( 
.A1(n_15511),
.A2(n_15157),
.B(n_15107),
.Y(n_15537)
);

INVx1_ASAP7_75t_L g15538 ( 
.A(n_15415),
.Y(n_15538)
);

INVx1_ASAP7_75t_L g15539 ( 
.A(n_15274),
.Y(n_15539)
);

NAND2xp5_ASAP7_75t_L g15540 ( 
.A(n_15280),
.B(n_15096),
.Y(n_15540)
);

OAI222xp33_ASAP7_75t_L g15541 ( 
.A1(n_15273),
.A2(n_15201),
.B1(n_15166),
.B2(n_15064),
.C1(n_15151),
.C2(n_15243),
.Y(n_15541)
);

OAI32xp33_ASAP7_75t_SL g15542 ( 
.A1(n_15352),
.A2(n_15152),
.A3(n_15222),
.B1(n_15136),
.B2(n_15194),
.Y(n_15542)
);

INVx1_ASAP7_75t_SL g15543 ( 
.A(n_15312),
.Y(n_15543)
);

A2O1A1Ixp33_ASAP7_75t_L g15544 ( 
.A1(n_15432),
.A2(n_15162),
.B(n_15174),
.C(n_15267),
.Y(n_15544)
);

A2O1A1Ixp33_ASAP7_75t_SL g15545 ( 
.A1(n_15324),
.A2(n_15252),
.B(n_15268),
.C(n_15216),
.Y(n_15545)
);

OAI222xp33_ASAP7_75t_L g15546 ( 
.A1(n_15335),
.A2(n_15255),
.B1(n_15223),
.B2(n_15254),
.C1(n_15076),
.C2(n_15161),
.Y(n_15546)
);

NAND2x1p5_ASAP7_75t_L g15547 ( 
.A(n_15278),
.B(n_15097),
.Y(n_15547)
);

OAI221xp5_ASAP7_75t_L g15548 ( 
.A1(n_15307),
.A2(n_15147),
.B1(n_15146),
.B2(n_15179),
.C(n_15221),
.Y(n_15548)
);

AOI21xp5_ASAP7_75t_L g15549 ( 
.A1(n_15279),
.A2(n_15234),
.B(n_15059),
.Y(n_15549)
);

NAND2xp5_ASAP7_75t_L g15550 ( 
.A(n_15456),
.B(n_15073),
.Y(n_15550)
);

INVx1_ASAP7_75t_L g15551 ( 
.A(n_15422),
.Y(n_15551)
);

INVx1_ASAP7_75t_L g15552 ( 
.A(n_15348),
.Y(n_15552)
);

INVx1_ASAP7_75t_L g15553 ( 
.A(n_15271),
.Y(n_15553)
);

OR2x2_ASAP7_75t_L g15554 ( 
.A(n_15286),
.B(n_15236),
.Y(n_15554)
);

AND2x2_ASAP7_75t_L g15555 ( 
.A(n_15318),
.B(n_15071),
.Y(n_15555)
);

AOI21xp33_ASAP7_75t_L g15556 ( 
.A1(n_15322),
.A2(n_15239),
.B(n_15226),
.Y(n_15556)
);

NAND2xp33_ASAP7_75t_SL g15557 ( 
.A(n_15336),
.B(n_15071),
.Y(n_15557)
);

AO22x1_ASAP7_75t_L g15558 ( 
.A1(n_15343),
.A2(n_15196),
.B1(n_15251),
.B2(n_15081),
.Y(n_15558)
);

NAND4xp25_ASAP7_75t_L g15559 ( 
.A(n_15411),
.B(n_15110),
.C(n_15062),
.D(n_15196),
.Y(n_15559)
);

OAI22xp33_ASAP7_75t_L g15560 ( 
.A1(n_15283),
.A2(n_15199),
.B1(n_15178),
.B2(n_15227),
.Y(n_15560)
);

OR2x2_ASAP7_75t_L g15561 ( 
.A(n_15342),
.B(n_6295),
.Y(n_15561)
);

AOI221xp5_ASAP7_75t_L g15562 ( 
.A1(n_15479),
.A2(n_7759),
.B1(n_7618),
.B2(n_7396),
.C(n_7432),
.Y(n_15562)
);

AOI332xp33_ASAP7_75t_L g15563 ( 
.A1(n_15276),
.A2(n_7651),
.A3(n_7631),
.B1(n_7664),
.B2(n_7663),
.B3(n_7812),
.C1(n_7647),
.C2(n_7617),
.Y(n_15563)
);

INVxp67_ASAP7_75t_L g15564 ( 
.A(n_15398),
.Y(n_15564)
);

OAI221xp5_ASAP7_75t_L g15565 ( 
.A1(n_15305),
.A2(n_7411),
.B1(n_7510),
.B2(n_7402),
.C(n_7385),
.Y(n_15565)
);

INVx1_ASAP7_75t_L g15566 ( 
.A(n_15370),
.Y(n_15566)
);

A2O1A1Ixp33_ASAP7_75t_L g15567 ( 
.A1(n_15371),
.A2(n_7248),
.B(n_7186),
.C(n_7198),
.Y(n_15567)
);

INVx1_ASAP7_75t_L g15568 ( 
.A(n_15373),
.Y(n_15568)
);

OR2x2_ASAP7_75t_L g15569 ( 
.A(n_15408),
.B(n_6344),
.Y(n_15569)
);

INVx1_ASAP7_75t_L g15570 ( 
.A(n_15292),
.Y(n_15570)
);

INVx2_ASAP7_75t_L g15571 ( 
.A(n_15336),
.Y(n_15571)
);

INVx1_ASAP7_75t_L g15572 ( 
.A(n_15347),
.Y(n_15572)
);

INVx1_ASAP7_75t_L g15573 ( 
.A(n_15369),
.Y(n_15573)
);

OAI32xp33_ASAP7_75t_L g15574 ( 
.A1(n_15462),
.A2(n_8274),
.A3(n_8269),
.B1(n_7411),
.B2(n_7510),
.Y(n_15574)
);

AOI211x1_ASAP7_75t_SL g15575 ( 
.A1(n_15488),
.A2(n_7005),
.B(n_7013),
.C(n_6638),
.Y(n_15575)
);

AOI22xp5_ASAP7_75t_L g15576 ( 
.A1(n_15527),
.A2(n_15528),
.B1(n_15451),
.B2(n_15498),
.Y(n_15576)
);

NAND2xp5_ASAP7_75t_L g15577 ( 
.A(n_15354),
.B(n_7390),
.Y(n_15577)
);

AOI22xp5_ASAP7_75t_L g15578 ( 
.A1(n_15460),
.A2(n_8064),
.B1(n_8126),
.B2(n_7975),
.Y(n_15578)
);

OAI22xp33_ASAP7_75t_L g15579 ( 
.A1(n_15288),
.A2(n_7187),
.B1(n_7206),
.B2(n_7173),
.Y(n_15579)
);

OR2x2_ASAP7_75t_L g15580 ( 
.A(n_15363),
.B(n_6344),
.Y(n_15580)
);

INVx1_ASAP7_75t_L g15581 ( 
.A(n_15472),
.Y(n_15581)
);

NAND2x1p5_ASAP7_75t_L g15582 ( 
.A(n_15302),
.B(n_9187),
.Y(n_15582)
);

NAND2xp5_ASAP7_75t_L g15583 ( 
.A(n_15525),
.B(n_7396),
.Y(n_15583)
);

NAND2xp33_ASAP7_75t_SL g15584 ( 
.A(n_15386),
.B(n_6992),
.Y(n_15584)
);

AOI21xp5_ASAP7_75t_L g15585 ( 
.A1(n_15350),
.A2(n_7188),
.B(n_7186),
.Y(n_15585)
);

OAI22xp33_ASAP7_75t_L g15586 ( 
.A1(n_15296),
.A2(n_7187),
.B1(n_7206),
.B2(n_7173),
.Y(n_15586)
);

INVx1_ASAP7_75t_L g15587 ( 
.A(n_15317),
.Y(n_15587)
);

AOI221x1_ASAP7_75t_L g15588 ( 
.A1(n_15400),
.A2(n_15334),
.B1(n_15327),
.B2(n_15328),
.C(n_15298),
.Y(n_15588)
);

NAND2xp5_ASAP7_75t_L g15589 ( 
.A(n_15341),
.B(n_15401),
.Y(n_15589)
);

INVx1_ASAP7_75t_L g15590 ( 
.A(n_15351),
.Y(n_15590)
);

NAND2xp5_ASAP7_75t_L g15591 ( 
.A(n_15294),
.B(n_7396),
.Y(n_15591)
);

OR2x2_ASAP7_75t_L g15592 ( 
.A(n_15320),
.B(n_6408),
.Y(n_15592)
);

INVx1_ASAP7_75t_L g15593 ( 
.A(n_15443),
.Y(n_15593)
);

NOR2x1_ASAP7_75t_L g15594 ( 
.A(n_15340),
.B(n_7975),
.Y(n_15594)
);

INVx1_ASAP7_75t_L g15595 ( 
.A(n_15345),
.Y(n_15595)
);

OAI22xp5_ASAP7_75t_L g15596 ( 
.A1(n_15297),
.A2(n_8139),
.B1(n_8006),
.B2(n_7206),
.Y(n_15596)
);

NAND2xp5_ASAP7_75t_L g15597 ( 
.A(n_15387),
.B(n_7426),
.Y(n_15597)
);

INVx1_ASAP7_75t_SL g15598 ( 
.A(n_15282),
.Y(n_15598)
);

INVx1_ASAP7_75t_L g15599 ( 
.A(n_15379),
.Y(n_15599)
);

INVx1_ASAP7_75t_L g15600 ( 
.A(n_15372),
.Y(n_15600)
);

OAI32xp33_ASAP7_75t_L g15601 ( 
.A1(n_15353),
.A2(n_8274),
.A3(n_8269),
.B1(n_7411),
.B2(n_7510),
.Y(n_15601)
);

OAI211xp5_ASAP7_75t_L g15602 ( 
.A1(n_15424),
.A2(n_6197),
.B(n_9187),
.C(n_6426),
.Y(n_15602)
);

NAND2xp5_ASAP7_75t_L g15603 ( 
.A(n_15458),
.B(n_7426),
.Y(n_15603)
);

INVx1_ASAP7_75t_L g15604 ( 
.A(n_15299),
.Y(n_15604)
);

NAND2xp5_ASAP7_75t_L g15605 ( 
.A(n_15445),
.B(n_7426),
.Y(n_15605)
);

INVx1_ASAP7_75t_L g15606 ( 
.A(n_15405),
.Y(n_15606)
);

AND2x4_ASAP7_75t_L g15607 ( 
.A(n_15402),
.B(n_8870),
.Y(n_15607)
);

INVx1_ASAP7_75t_L g15608 ( 
.A(n_15423),
.Y(n_15608)
);

AOI221xp5_ASAP7_75t_L g15609 ( 
.A1(n_15380),
.A2(n_7759),
.B1(n_7447),
.B2(n_7475),
.C(n_7432),
.Y(n_15609)
);

INVxp67_ASAP7_75t_L g15610 ( 
.A(n_15409),
.Y(n_15610)
);

OR2x2_ASAP7_75t_L g15611 ( 
.A(n_15308),
.B(n_6408),
.Y(n_15611)
);

OAI21xp5_ASAP7_75t_L g15612 ( 
.A1(n_15419),
.A2(n_7503),
.B(n_7959),
.Y(n_15612)
);

OAI211xp5_ASAP7_75t_SL g15613 ( 
.A1(n_15367),
.A2(n_7005),
.B(n_7013),
.C(n_7631),
.Y(n_15613)
);

INVx1_ASAP7_75t_L g15614 ( 
.A(n_15319),
.Y(n_15614)
);

NAND2xp5_ASAP7_75t_L g15615 ( 
.A(n_15421),
.B(n_7426),
.Y(n_15615)
);

AOI21xp33_ASAP7_75t_SL g15616 ( 
.A1(n_15325),
.A2(n_7959),
.B(n_7402),
.Y(n_15616)
);

INVx1_ASAP7_75t_L g15617 ( 
.A(n_15413),
.Y(n_15617)
);

AOI22xp5_ASAP7_75t_L g15618 ( 
.A1(n_15487),
.A2(n_8064),
.B1(n_8126),
.B2(n_7975),
.Y(n_15618)
);

INVx2_ASAP7_75t_SL g15619 ( 
.A(n_15435),
.Y(n_15619)
);

INVx1_ASAP7_75t_L g15620 ( 
.A(n_15293),
.Y(n_15620)
);

OAI221xp5_ASAP7_75t_SL g15621 ( 
.A1(n_15523),
.A2(n_6931),
.B1(n_6998),
.B2(n_6989),
.C(n_6967),
.Y(n_15621)
);

INVxp67_ASAP7_75t_SL g15622 ( 
.A(n_15454),
.Y(n_15622)
);

OAI221xp5_ASAP7_75t_L g15623 ( 
.A1(n_15281),
.A2(n_7411),
.B1(n_7510),
.B2(n_7402),
.C(n_7385),
.Y(n_15623)
);

INVx1_ASAP7_75t_SL g15624 ( 
.A(n_15446),
.Y(n_15624)
);

AOI21xp5_ASAP7_75t_L g15625 ( 
.A1(n_15517),
.A2(n_15311),
.B(n_15420),
.Y(n_15625)
);

OAI21xp5_ASAP7_75t_SL g15626 ( 
.A1(n_15465),
.A2(n_8274),
.B(n_8269),
.Y(n_15626)
);

INVx1_ASAP7_75t_L g15627 ( 
.A(n_15337),
.Y(n_15627)
);

OAI22xp33_ASAP7_75t_L g15628 ( 
.A1(n_15303),
.A2(n_7206),
.B1(n_7365),
.B2(n_7187),
.Y(n_15628)
);

OAI31xp33_ASAP7_75t_L g15629 ( 
.A1(n_15535),
.A2(n_7385),
.A3(n_7513),
.B(n_7512),
.Y(n_15629)
);

NAND2xp5_ASAP7_75t_L g15630 ( 
.A(n_15427),
.B(n_7432),
.Y(n_15630)
);

INVx1_ASAP7_75t_L g15631 ( 
.A(n_15467),
.Y(n_15631)
);

INVx1_ASAP7_75t_SL g15632 ( 
.A(n_15448),
.Y(n_15632)
);

OAI22xp5_ASAP7_75t_SL g15633 ( 
.A1(n_15383),
.A2(n_7132),
.B1(n_6992),
.B2(n_6964),
.Y(n_15633)
);

OAI21xp5_ASAP7_75t_L g15634 ( 
.A1(n_15449),
.A2(n_7240),
.B(n_8925),
.Y(n_15634)
);

O2A1O1Ixp33_ASAP7_75t_L g15635 ( 
.A1(n_15366),
.A2(n_8033),
.B(n_8067),
.C(n_8009),
.Y(n_15635)
);

INVx1_ASAP7_75t_L g15636 ( 
.A(n_15407),
.Y(n_15636)
);

OAI322xp33_ASAP7_75t_L g15637 ( 
.A1(n_15406),
.A2(n_7664),
.A3(n_7651),
.B1(n_7812),
.B2(n_7819),
.C1(n_7663),
.C2(n_7647),
.Y(n_15637)
);

NAND2xp5_ASAP7_75t_L g15638 ( 
.A(n_15323),
.B(n_7432),
.Y(n_15638)
);

NAND3xp33_ASAP7_75t_L g15639 ( 
.A(n_15457),
.B(n_7475),
.C(n_7447),
.Y(n_15639)
);

NOR2xp33_ASAP7_75t_L g15640 ( 
.A(n_15524),
.B(n_7447),
.Y(n_15640)
);

NAND2xp5_ASAP7_75t_L g15641 ( 
.A(n_15329),
.B(n_7447),
.Y(n_15641)
);

INVx1_ASAP7_75t_L g15642 ( 
.A(n_15410),
.Y(n_15642)
);

AOI22xp33_ASAP7_75t_SL g15643 ( 
.A1(n_15333),
.A2(n_8139),
.B1(n_7187),
.B2(n_7365),
.Y(n_15643)
);

AOI22xp33_ASAP7_75t_L g15644 ( 
.A1(n_15504),
.A2(n_7488),
.B1(n_7496),
.B2(n_7475),
.Y(n_15644)
);

OAI32xp33_ASAP7_75t_L g15645 ( 
.A1(n_15485),
.A2(n_7635),
.A3(n_7513),
.B1(n_7512),
.B2(n_6426),
.Y(n_15645)
);

HB1xp67_ASAP7_75t_L g15646 ( 
.A(n_15430),
.Y(n_15646)
);

AND2x2_ASAP7_75t_L g15647 ( 
.A(n_15291),
.B(n_7454),
.Y(n_15647)
);

NAND2xp5_ASAP7_75t_SL g15648 ( 
.A(n_15499),
.B(n_7206),
.Y(n_15648)
);

AOI22xp5_ASAP7_75t_L g15649 ( 
.A1(n_15522),
.A2(n_8126),
.B1(n_8151),
.B2(n_8064),
.Y(n_15649)
);

INVx1_ASAP7_75t_L g15650 ( 
.A(n_15388),
.Y(n_15650)
);

A2O1A1Ixp33_ASAP7_75t_L g15651 ( 
.A1(n_15397),
.A2(n_7188),
.B(n_7198),
.C(n_7186),
.Y(n_15651)
);

NOR2xp67_ASAP7_75t_L g15652 ( 
.A(n_15403),
.B(n_6939),
.Y(n_15652)
);

INVx1_ASAP7_75t_L g15653 ( 
.A(n_15394),
.Y(n_15653)
);

OAI21xp5_ASAP7_75t_SL g15654 ( 
.A1(n_15481),
.A2(n_15505),
.B(n_15331),
.Y(n_15654)
);

AOI322xp5_ASAP7_75t_L g15655 ( 
.A1(n_15434),
.A2(n_7538),
.A3(n_7557),
.B1(n_7620),
.B2(n_7685),
.C1(n_7542),
.C2(n_7507),
.Y(n_15655)
);

AND2x2_ASAP7_75t_L g15656 ( 
.A(n_15287),
.B(n_7519),
.Y(n_15656)
);

INVx1_ASAP7_75t_L g15657 ( 
.A(n_15284),
.Y(n_15657)
);

NAND2x1_ASAP7_75t_SL g15658 ( 
.A(n_15381),
.B(n_7132),
.Y(n_15658)
);

OR2x2_ASAP7_75t_L g15659 ( 
.A(n_15431),
.B(n_15414),
.Y(n_15659)
);

INVx1_ASAP7_75t_L g15660 ( 
.A(n_15364),
.Y(n_15660)
);

AND2x2_ASAP7_75t_L g15661 ( 
.A(n_15272),
.B(n_7519),
.Y(n_15661)
);

INVx1_ASAP7_75t_L g15662 ( 
.A(n_15436),
.Y(n_15662)
);

OR2x2_ASAP7_75t_L g15663 ( 
.A(n_15289),
.B(n_6429),
.Y(n_15663)
);

INVx1_ASAP7_75t_L g15664 ( 
.A(n_15447),
.Y(n_15664)
);

AND2x2_ASAP7_75t_L g15665 ( 
.A(n_15304),
.B(n_7519),
.Y(n_15665)
);

OAI22xp5_ASAP7_75t_SL g15666 ( 
.A1(n_15382),
.A2(n_6964),
.B1(n_7023),
.B2(n_6939),
.Y(n_15666)
);

AOI221x1_ASAP7_75t_L g15667 ( 
.A1(n_15441),
.A2(n_7954),
.B1(n_8114),
.B2(n_8067),
.C(n_7819),
.Y(n_15667)
);

O2A1O1Ixp33_ASAP7_75t_SL g15668 ( 
.A1(n_15361),
.A2(n_6476),
.B(n_6534),
.C(n_6429),
.Y(n_15668)
);

INVx2_ASAP7_75t_L g15669 ( 
.A(n_15455),
.Y(n_15669)
);

INVxp67_ASAP7_75t_L g15670 ( 
.A(n_15450),
.Y(n_15670)
);

AOI22xp5_ASAP7_75t_L g15671 ( 
.A1(n_15533),
.A2(n_8126),
.B1(n_8151),
.B2(n_8064),
.Y(n_15671)
);

AOI321xp33_ASAP7_75t_L g15672 ( 
.A1(n_15362),
.A2(n_7709),
.A3(n_7705),
.B1(n_7700),
.B2(n_8296),
.C(n_8151),
.Y(n_15672)
);

NAND2xp5_ASAP7_75t_L g15673 ( 
.A(n_15365),
.B(n_7475),
.Y(n_15673)
);

NAND2xp5_ASAP7_75t_L g15674 ( 
.A(n_15368),
.B(n_7488),
.Y(n_15674)
);

OAI21xp5_ASAP7_75t_L g15675 ( 
.A1(n_15358),
.A2(n_15375),
.B(n_15466),
.Y(n_15675)
);

INVxp67_ASAP7_75t_SL g15676 ( 
.A(n_15349),
.Y(n_15676)
);

INVx1_ASAP7_75t_L g15677 ( 
.A(n_15310),
.Y(n_15677)
);

INVx1_ASAP7_75t_L g15678 ( 
.A(n_15346),
.Y(n_15678)
);

NAND2xp5_ASAP7_75t_L g15679 ( 
.A(n_15496),
.B(n_7488),
.Y(n_15679)
);

INVx1_ASAP7_75t_L g15680 ( 
.A(n_15486),
.Y(n_15680)
);

OAI21xp5_ASAP7_75t_SL g15681 ( 
.A1(n_15510),
.A2(n_15500),
.B(n_15526),
.Y(n_15681)
);

INVx1_ASAP7_75t_L g15682 ( 
.A(n_15471),
.Y(n_15682)
);

NAND2x1p5_ASAP7_75t_L g15683 ( 
.A(n_15474),
.B(n_15463),
.Y(n_15683)
);

NAND3xp33_ASAP7_75t_L g15684 ( 
.A(n_15385),
.B(n_7496),
.C(n_7488),
.Y(n_15684)
);

OAI22xp5_ASAP7_75t_L g15685 ( 
.A1(n_15508),
.A2(n_7365),
.B1(n_7369),
.B2(n_7206),
.Y(n_15685)
);

AOI222xp33_ASAP7_75t_L g15686 ( 
.A1(n_15492),
.A2(n_7162),
.B1(n_7506),
.B2(n_7534),
.C1(n_7507),
.C2(n_7501),
.Y(n_15686)
);

INVx2_ASAP7_75t_SL g15687 ( 
.A(n_15313),
.Y(n_15687)
);

NAND2xp5_ASAP7_75t_SL g15688 ( 
.A(n_15391),
.B(n_7206),
.Y(n_15688)
);

AOI211xp5_ASAP7_75t_L g15689 ( 
.A1(n_15473),
.A2(n_9012),
.B(n_9041),
.C(n_7162),
.Y(n_15689)
);

OAI21xp5_ASAP7_75t_SL g15690 ( 
.A1(n_15507),
.A2(n_7513),
.B(n_7512),
.Y(n_15690)
);

INVx1_ASAP7_75t_L g15691 ( 
.A(n_15306),
.Y(n_15691)
);

AOI22xp5_ASAP7_75t_L g15692 ( 
.A1(n_15497),
.A2(n_8151),
.B1(n_8164),
.B2(n_8126),
.Y(n_15692)
);

AND2x4_ASAP7_75t_L g15693 ( 
.A(n_15395),
.B(n_9012),
.Y(n_15693)
);

OAI22xp33_ASAP7_75t_L g15694 ( 
.A1(n_15285),
.A2(n_15344),
.B1(n_15453),
.B2(n_15316),
.Y(n_15694)
);

OAI31xp33_ASAP7_75t_L g15695 ( 
.A1(n_15516),
.A2(n_7512),
.A3(n_7635),
.B(n_7513),
.Y(n_15695)
);

INVx2_ASAP7_75t_L g15696 ( 
.A(n_15295),
.Y(n_15696)
);

NAND2xp33_ASAP7_75t_SL g15697 ( 
.A(n_15356),
.B(n_7206),
.Y(n_15697)
);

OAI31xp33_ASAP7_75t_L g15698 ( 
.A1(n_15534),
.A2(n_7635),
.A3(n_7740),
.B(n_7106),
.Y(n_15698)
);

INVx2_ASAP7_75t_SL g15699 ( 
.A(n_15412),
.Y(n_15699)
);

NOR2xp33_ASAP7_75t_L g15700 ( 
.A(n_15489),
.B(n_7496),
.Y(n_15700)
);

OAI22xp5_ASAP7_75t_L g15701 ( 
.A1(n_15290),
.A2(n_15300),
.B1(n_15425),
.B2(n_15377),
.Y(n_15701)
);

INVx1_ASAP7_75t_L g15702 ( 
.A(n_15326),
.Y(n_15702)
);

NAND2xp5_ASAP7_75t_L g15703 ( 
.A(n_15416),
.B(n_7496),
.Y(n_15703)
);

OAI221xp5_ASAP7_75t_L g15704 ( 
.A1(n_15464),
.A2(n_7635),
.B1(n_7369),
.B2(n_7493),
.C(n_7478),
.Y(n_15704)
);

NOR3xp33_ASAP7_75t_L g15705 ( 
.A(n_15475),
.B(n_7740),
.C(n_7495),
.Y(n_15705)
);

BUFx2_ASAP7_75t_L g15706 ( 
.A(n_15476),
.Y(n_15706)
);

AOI21xp33_ASAP7_75t_L g15707 ( 
.A1(n_15478),
.A2(n_7506),
.B(n_7501),
.Y(n_15707)
);

AOI221xp5_ASAP7_75t_SL g15708 ( 
.A1(n_15515),
.A2(n_15275),
.B1(n_15392),
.B2(n_15490),
.C(n_15452),
.Y(n_15708)
);

INVx1_ASAP7_75t_L g15709 ( 
.A(n_15338),
.Y(n_15709)
);

AOI211xp5_ASAP7_75t_L g15710 ( 
.A1(n_15491),
.A2(n_9041),
.B(n_7162),
.C(n_8631),
.Y(n_15710)
);

OAI22xp33_ASAP7_75t_L g15711 ( 
.A1(n_15309),
.A2(n_7369),
.B1(n_7478),
.B2(n_7365),
.Y(n_15711)
);

INVx1_ASAP7_75t_L g15712 ( 
.A(n_15384),
.Y(n_15712)
);

INVxp67_ASAP7_75t_L g15713 ( 
.A(n_15501),
.Y(n_15713)
);

NAND2xp5_ASAP7_75t_L g15714 ( 
.A(n_15442),
.B(n_15417),
.Y(n_15714)
);

OAI21xp33_ASAP7_75t_SL g15715 ( 
.A1(n_15378),
.A2(n_8631),
.B(n_8629),
.Y(n_15715)
);

OAI22xp5_ASAP7_75t_L g15716 ( 
.A1(n_15495),
.A2(n_15438),
.B1(n_15277),
.B2(n_15494),
.Y(n_15716)
);

AOI21xp33_ASAP7_75t_SL g15717 ( 
.A1(n_15514),
.A2(n_7847),
.B(n_8629),
.Y(n_15717)
);

AND2x2_ASAP7_75t_L g15718 ( 
.A(n_15357),
.B(n_7519),
.Y(n_15718)
);

OAI22xp33_ASAP7_75t_L g15719 ( 
.A1(n_15314),
.A2(n_7369),
.B1(n_7478),
.B2(n_7365),
.Y(n_15719)
);

OAI21xp5_ASAP7_75t_L g15720 ( 
.A1(n_15483),
.A2(n_7354),
.B(n_8635),
.Y(n_15720)
);

NAND4xp25_ASAP7_75t_SL g15721 ( 
.A(n_15444),
.B(n_7812),
.C(n_7819),
.D(n_7664),
.Y(n_15721)
);

OAI22xp5_ASAP7_75t_L g15722 ( 
.A1(n_15476),
.A2(n_7369),
.B1(n_7478),
.B2(n_7365),
.Y(n_15722)
);

XOR2x2_ASAP7_75t_L g15723 ( 
.A(n_15506),
.B(n_6654),
.Y(n_15723)
);

NAND3xp33_ASAP7_75t_L g15724 ( 
.A(n_15509),
.B(n_7506),
.C(n_7501),
.Y(n_15724)
);

INVx1_ASAP7_75t_L g15725 ( 
.A(n_15390),
.Y(n_15725)
);

INVx1_ASAP7_75t_L g15726 ( 
.A(n_15399),
.Y(n_15726)
);

OAI22xp5_ASAP7_75t_L g15727 ( 
.A1(n_15374),
.A2(n_7369),
.B1(n_7478),
.B2(n_7365),
.Y(n_15727)
);

OR2x2_ASAP7_75t_L g15728 ( 
.A(n_15440),
.B(n_6476),
.Y(n_15728)
);

NAND4xp25_ASAP7_75t_SL g15729 ( 
.A(n_15502),
.B(n_15493),
.C(n_15532),
.D(n_15360),
.Y(n_15729)
);

O2A1O1Ixp33_ASAP7_75t_L g15730 ( 
.A1(n_15512),
.A2(n_8114),
.B(n_7954),
.C(n_7506),
.Y(n_15730)
);

O2A1O1Ixp33_ASAP7_75t_L g15731 ( 
.A1(n_15513),
.A2(n_7507),
.B(n_7534),
.C(n_7501),
.Y(n_15731)
);

NAND2xp5_ASAP7_75t_L g15732 ( 
.A(n_15480),
.B(n_7507),
.Y(n_15732)
);

NAND2xp5_ASAP7_75t_L g15733 ( 
.A(n_15530),
.B(n_7534),
.Y(n_15733)
);

INVx2_ASAP7_75t_L g15734 ( 
.A(n_15301),
.Y(n_15734)
);

A2O1A1Ixp33_ASAP7_75t_L g15735 ( 
.A1(n_15315),
.A2(n_7198),
.B(n_7188),
.C(n_7272),
.Y(n_15735)
);

INVx1_ASAP7_75t_L g15736 ( 
.A(n_15484),
.Y(n_15736)
);

AOI21xp5_ASAP7_75t_L g15737 ( 
.A1(n_15468),
.A2(n_7321),
.B(n_7831),
.Y(n_15737)
);

INVx2_ASAP7_75t_L g15738 ( 
.A(n_15301),
.Y(n_15738)
);

INVx1_ASAP7_75t_L g15739 ( 
.A(n_15332),
.Y(n_15739)
);

OAI21xp33_ASAP7_75t_SL g15740 ( 
.A1(n_15389),
.A2(n_8635),
.B(n_7894),
.Y(n_15740)
);

NAND2xp5_ASAP7_75t_L g15741 ( 
.A(n_15330),
.B(n_7534),
.Y(n_15741)
);

AND2x2_ASAP7_75t_L g15742 ( 
.A(n_15359),
.B(n_7519),
.Y(n_15742)
);

O2A1O1Ixp33_ASAP7_75t_SL g15743 ( 
.A1(n_15339),
.A2(n_6594),
.B(n_6639),
.C(n_6534),
.Y(n_15743)
);

INVx1_ASAP7_75t_L g15744 ( 
.A(n_15520),
.Y(n_15744)
);

NAND2xp33_ASAP7_75t_SL g15745 ( 
.A(n_15321),
.B(n_7365),
.Y(n_15745)
);

OAI21xp5_ASAP7_75t_SL g15746 ( 
.A1(n_15470),
.A2(n_15531),
.B(n_15428),
.Y(n_15746)
);

OAI21xp5_ASAP7_75t_L g15747 ( 
.A1(n_15518),
.A2(n_7354),
.B(n_7294),
.Y(n_15747)
);

NAND3xp33_ASAP7_75t_SL g15748 ( 
.A(n_15519),
.B(n_7550),
.C(n_7542),
.Y(n_15748)
);

AOI21xp5_ASAP7_75t_L g15749 ( 
.A1(n_15426),
.A2(n_7321),
.B(n_7831),
.Y(n_15749)
);

INVx1_ASAP7_75t_L g15750 ( 
.A(n_15376),
.Y(n_15750)
);

NAND2xp5_ASAP7_75t_L g15751 ( 
.A(n_15418),
.B(n_7542),
.Y(n_15751)
);

INVx1_ASAP7_75t_L g15752 ( 
.A(n_15404),
.Y(n_15752)
);

OAI22xp5_ASAP7_75t_L g15753 ( 
.A1(n_15393),
.A2(n_7478),
.B1(n_7493),
.B2(n_7369),
.Y(n_15753)
);

NAND2xp5_ASAP7_75t_L g15754 ( 
.A(n_15429),
.B(n_7542),
.Y(n_15754)
);

INVx1_ASAP7_75t_L g15755 ( 
.A(n_15396),
.Y(n_15755)
);

AND2x4_ASAP7_75t_SL g15756 ( 
.A(n_15469),
.B(n_6570),
.Y(n_15756)
);

INVx2_ASAP7_75t_L g15757 ( 
.A(n_15355),
.Y(n_15757)
);

AOI322xp5_ASAP7_75t_L g15758 ( 
.A1(n_15437),
.A2(n_8138),
.A3(n_7744),
.B1(n_8220),
.B2(n_8275),
.C1(n_7773),
.C2(n_7690),
.Y(n_15758)
);

NOR2xp33_ASAP7_75t_L g15759 ( 
.A(n_15477),
.B(n_7550),
.Y(n_15759)
);

OAI221xp5_ASAP7_75t_L g15760 ( 
.A1(n_15538),
.A2(n_15482),
.B1(n_15529),
.B2(n_15461),
.C(n_15459),
.Y(n_15760)
);

NAND4xp25_ASAP7_75t_SL g15761 ( 
.A(n_15543),
.B(n_15439),
.C(n_15503),
.D(n_15433),
.Y(n_15761)
);

AND2x2_ASAP7_75t_L g15762 ( 
.A(n_15646),
.B(n_7646),
.Y(n_15762)
);

INVx1_ASAP7_75t_SL g15763 ( 
.A(n_15624),
.Y(n_15763)
);

AOI22xp33_ASAP7_75t_L g15764 ( 
.A1(n_15706),
.A2(n_8298),
.B1(n_8275),
.B2(n_7553),
.Y(n_15764)
);

NOR2xp33_ASAP7_75t_L g15765 ( 
.A(n_15551),
.B(n_15564),
.Y(n_15765)
);

AOI21xp33_ASAP7_75t_L g15766 ( 
.A1(n_15545),
.A2(n_15550),
.B(n_15554),
.Y(n_15766)
);

OAI21xp5_ASAP7_75t_L g15767 ( 
.A1(n_15670),
.A2(n_7388),
.B(n_7384),
.Y(n_15767)
);

OAI211xp5_ASAP7_75t_SL g15768 ( 
.A1(n_15598),
.A2(n_7831),
.B(n_7980),
.C(n_7973),
.Y(n_15768)
);

OAI22xp33_ASAP7_75t_SL g15769 ( 
.A1(n_15552),
.A2(n_7550),
.B1(n_7557),
.B2(n_7553),
.Y(n_15769)
);

AOI31xp33_ASAP7_75t_L g15770 ( 
.A1(n_15589),
.A2(n_6816),
.A3(n_6847),
.B(n_6658),
.Y(n_15770)
);

INVx1_ASAP7_75t_L g15771 ( 
.A(n_15573),
.Y(n_15771)
);

NAND2xp5_ASAP7_75t_L g15772 ( 
.A(n_15622),
.B(n_7550),
.Y(n_15772)
);

INVx1_ASAP7_75t_L g15773 ( 
.A(n_15676),
.Y(n_15773)
);

INVx1_ASAP7_75t_L g15774 ( 
.A(n_15599),
.Y(n_15774)
);

NAND2xp5_ASAP7_75t_L g15775 ( 
.A(n_15555),
.B(n_7553),
.Y(n_15775)
);

NAND2xp5_ASAP7_75t_L g15776 ( 
.A(n_15619),
.B(n_7553),
.Y(n_15776)
);

AOI211xp5_ASAP7_75t_L g15777 ( 
.A1(n_15681),
.A2(n_15694),
.B(n_15556),
.C(n_15581),
.Y(n_15777)
);

OAI332xp33_ASAP7_75t_L g15778 ( 
.A1(n_15632),
.A2(n_7106),
.A3(n_7108),
.B1(n_7138),
.B2(n_6568),
.B3(n_6537),
.C1(n_6648),
.C2(n_6575),
.Y(n_15778)
);

OAI211xp5_ASAP7_75t_SL g15779 ( 
.A1(n_15537),
.A2(n_7973),
.B(n_8004),
.C(n_7980),
.Y(n_15779)
);

OAI22xp5_ASAP7_75t_L g15780 ( 
.A1(n_15608),
.A2(n_7478),
.B1(n_7493),
.B2(n_7369),
.Y(n_15780)
);

NOR3xp33_ASAP7_75t_SL g15781 ( 
.A(n_15557),
.B(n_6904),
.C(n_7973),
.Y(n_15781)
);

NAND2xp5_ASAP7_75t_L g15782 ( 
.A(n_15595),
.B(n_7557),
.Y(n_15782)
);

OR2x2_ASAP7_75t_L g15783 ( 
.A(n_15547),
.B(n_6594),
.Y(n_15783)
);

INVx1_ASAP7_75t_SL g15784 ( 
.A(n_15659),
.Y(n_15784)
);

HB1xp67_ASAP7_75t_L g15785 ( 
.A(n_15593),
.Y(n_15785)
);

OAI221xp5_ASAP7_75t_SL g15786 ( 
.A1(n_15654),
.A2(n_6967),
.B1(n_6998),
.B2(n_6989),
.C(n_6931),
.Y(n_15786)
);

NAND2xp5_ASAP7_75t_L g15787 ( 
.A(n_15539),
.B(n_7557),
.Y(n_15787)
);

AND2x2_ASAP7_75t_L g15788 ( 
.A(n_15571),
.B(n_7533),
.Y(n_15788)
);

AOI21xp33_ASAP7_75t_L g15789 ( 
.A1(n_15744),
.A2(n_8298),
.B(n_7587),
.Y(n_15789)
);

INVx1_ASAP7_75t_L g15790 ( 
.A(n_15683),
.Y(n_15790)
);

OAI21xp33_ASAP7_75t_L g15791 ( 
.A1(n_15600),
.A2(n_7548),
.B(n_7533),
.Y(n_15791)
);

INVx2_ASAP7_75t_L g15792 ( 
.A(n_15658),
.Y(n_15792)
);

AOI22xp5_ASAP7_75t_L g15793 ( 
.A1(n_15576),
.A2(n_8164),
.B1(n_8197),
.B2(n_8151),
.Y(n_15793)
);

OA21x2_ASAP7_75t_L g15794 ( 
.A1(n_15588),
.A2(n_7321),
.B(n_7847),
.Y(n_15794)
);

AOI221xp5_ASAP7_75t_L g15795 ( 
.A1(n_15542),
.A2(n_7607),
.B1(n_7659),
.B2(n_7587),
.C(n_7566),
.Y(n_15795)
);

INVx2_ASAP7_75t_L g15796 ( 
.A(n_15590),
.Y(n_15796)
);

INVx1_ASAP7_75t_L g15797 ( 
.A(n_15662),
.Y(n_15797)
);

INVx2_ASAP7_75t_SL g15798 ( 
.A(n_15594),
.Y(n_15798)
);

O2A1O1Ixp33_ASAP7_75t_L g15799 ( 
.A1(n_15610),
.A2(n_7587),
.B(n_7607),
.C(n_7566),
.Y(n_15799)
);

NAND2xp5_ASAP7_75t_L g15800 ( 
.A(n_15558),
.B(n_7566),
.Y(n_15800)
);

NAND2x1_ASAP7_75t_L g15801 ( 
.A(n_15680),
.B(n_7271),
.Y(n_15801)
);

OR2x2_ASAP7_75t_L g15802 ( 
.A(n_15597),
.B(n_6639),
.Y(n_15802)
);

INVx1_ASAP7_75t_SL g15803 ( 
.A(n_15664),
.Y(n_15803)
);

INVx1_ASAP7_75t_L g15804 ( 
.A(n_15606),
.Y(n_15804)
);

INVx1_ASAP7_75t_L g15805 ( 
.A(n_15617),
.Y(n_15805)
);

NAND2xp5_ASAP7_75t_L g15806 ( 
.A(n_15699),
.B(n_15640),
.Y(n_15806)
);

NAND2xp5_ASAP7_75t_L g15807 ( 
.A(n_15750),
.B(n_7566),
.Y(n_15807)
);

INVx1_ASAP7_75t_L g15808 ( 
.A(n_15572),
.Y(n_15808)
);

INVx1_ASAP7_75t_L g15809 ( 
.A(n_15627),
.Y(n_15809)
);

OR2x2_ASAP7_75t_L g15810 ( 
.A(n_15559),
.B(n_15569),
.Y(n_15810)
);

OAI21xp33_ASAP7_75t_L g15811 ( 
.A1(n_15675),
.A2(n_7548),
.B(n_7533),
.Y(n_15811)
);

INVx1_ASAP7_75t_L g15812 ( 
.A(n_15604),
.Y(n_15812)
);

AND2x2_ASAP7_75t_L g15813 ( 
.A(n_15661),
.B(n_7564),
.Y(n_15813)
);

INVx1_ASAP7_75t_L g15814 ( 
.A(n_15620),
.Y(n_15814)
);

OAI221xp5_ASAP7_75t_L g15815 ( 
.A1(n_15536),
.A2(n_7493),
.B1(n_7543),
.B2(n_7541),
.C(n_7478),
.Y(n_15815)
);

INVx1_ASAP7_75t_L g15816 ( 
.A(n_15682),
.Y(n_15816)
);

INVx1_ASAP7_75t_L g15817 ( 
.A(n_15660),
.Y(n_15817)
);

INVxp67_ASAP7_75t_L g15818 ( 
.A(n_15752),
.Y(n_15818)
);

OR2x2_ASAP7_75t_L g15819 ( 
.A(n_15583),
.B(n_6658),
.Y(n_15819)
);

NAND2xp5_ASAP7_75t_L g15820 ( 
.A(n_15614),
.B(n_7587),
.Y(n_15820)
);

INVxp67_ASAP7_75t_L g15821 ( 
.A(n_15755),
.Y(n_15821)
);

NOR2xp33_ASAP7_75t_L g15822 ( 
.A(n_15669),
.B(n_7607),
.Y(n_15822)
);

OAI22xp33_ASAP7_75t_L g15823 ( 
.A1(n_15714),
.A2(n_15587),
.B1(n_15540),
.B2(n_15631),
.Y(n_15823)
);

NAND2xp33_ASAP7_75t_SL g15824 ( 
.A(n_15570),
.B(n_7493),
.Y(n_15824)
);

AND2x4_ASAP7_75t_L g15825 ( 
.A(n_15652),
.B(n_7533),
.Y(n_15825)
);

INVx2_ASAP7_75t_L g15826 ( 
.A(n_15723),
.Y(n_15826)
);

OAI31xp33_ASAP7_75t_L g15827 ( 
.A1(n_15560),
.A2(n_7548),
.A3(n_7564),
.B(n_7533),
.Y(n_15827)
);

OAI21xp5_ASAP7_75t_L g15828 ( 
.A1(n_15549),
.A2(n_15713),
.B(n_15625),
.Y(n_15828)
);

NAND2xp5_ASAP7_75t_L g15829 ( 
.A(n_15718),
.B(n_7620),
.Y(n_15829)
);

INVx1_ASAP7_75t_SL g15830 ( 
.A(n_15636),
.Y(n_15830)
);

INVx2_ASAP7_75t_L g15831 ( 
.A(n_15582),
.Y(n_15831)
);

OAI21xp5_ASAP7_75t_L g15832 ( 
.A1(n_15577),
.A2(n_7388),
.B(n_7384),
.Y(n_15832)
);

INVx1_ASAP7_75t_L g15833 ( 
.A(n_15642),
.Y(n_15833)
);

OR2x2_ASAP7_75t_L g15834 ( 
.A(n_15553),
.B(n_6676),
.Y(n_15834)
);

AOI22xp5_ASAP7_75t_L g15835 ( 
.A1(n_15696),
.A2(n_8197),
.B1(n_8198),
.B2(n_8164),
.Y(n_15835)
);

AOI22xp33_ASAP7_75t_L g15836 ( 
.A1(n_15739),
.A2(n_8298),
.B1(n_7620),
.B2(n_7656),
.Y(n_15836)
);

NAND2xp5_ASAP7_75t_L g15837 ( 
.A(n_15657),
.B(n_7620),
.Y(n_15837)
);

NAND2xp5_ASAP7_75t_L g15838 ( 
.A(n_15650),
.B(n_7656),
.Y(n_15838)
);

OAI32xp33_ASAP7_75t_L g15839 ( 
.A1(n_15653),
.A2(n_6704),
.A3(n_6731),
.B1(n_6726),
.B2(n_6676),
.Y(n_15839)
);

OAI322xp33_ASAP7_75t_L g15840 ( 
.A1(n_15734),
.A2(n_8128),
.A3(n_8004),
.B1(n_8129),
.B2(n_8133),
.C1(n_8085),
.C2(n_7980),
.Y(n_15840)
);

OAI22xp33_ASAP7_75t_L g15841 ( 
.A1(n_15757),
.A2(n_7541),
.B1(n_7543),
.B2(n_7493),
.Y(n_15841)
);

AOI22xp5_ASAP7_75t_L g15842 ( 
.A1(n_15701),
.A2(n_8197),
.B1(n_8198),
.B2(n_8164),
.Y(n_15842)
);

INVx2_ASAP7_75t_L g15843 ( 
.A(n_15738),
.Y(n_15843)
);

AOI332xp33_ASAP7_75t_L g15844 ( 
.A1(n_15566),
.A2(n_8085),
.A3(n_8133),
.B1(n_8129),
.B2(n_8128),
.B3(n_8234),
.C1(n_8225),
.C2(n_8004),
.Y(n_15844)
);

AOI221xp5_ASAP7_75t_L g15845 ( 
.A1(n_15546),
.A2(n_7659),
.B1(n_7670),
.B2(n_7668),
.C(n_7607),
.Y(n_15845)
);

OAI322xp33_ASAP7_75t_L g15846 ( 
.A1(n_15611),
.A2(n_15548),
.A3(n_15568),
.B1(n_15687),
.B2(n_15561),
.C1(n_15688),
.C2(n_15716),
.Y(n_15846)
);

AOI22xp5_ASAP7_75t_L g15847 ( 
.A1(n_15729),
.A2(n_8197),
.B1(n_8198),
.B2(n_8164),
.Y(n_15847)
);

AOI32xp33_ASAP7_75t_L g15848 ( 
.A1(n_15584),
.A2(n_7849),
.A3(n_7853),
.B1(n_7294),
.B2(n_7946),
.Y(n_15848)
);

CKINVDCx6p67_ASAP7_75t_R g15849 ( 
.A(n_15677),
.Y(n_15849)
);

INVx1_ASAP7_75t_L g15850 ( 
.A(n_15605),
.Y(n_15850)
);

A2O1A1Ixp33_ASAP7_75t_SL g15851 ( 
.A1(n_15702),
.A2(n_8128),
.B(n_8129),
.C(n_8085),
.Y(n_15851)
);

AOI22xp33_ASAP7_75t_SL g15852 ( 
.A1(n_15678),
.A2(n_7541),
.B1(n_7543),
.B2(n_7493),
.Y(n_15852)
);

OAI222xp33_ASAP7_75t_L g15853 ( 
.A1(n_15648),
.A2(n_7548),
.B1(n_7592),
.B2(n_7646),
.C1(n_7568),
.C2(n_7564),
.Y(n_15853)
);

NOR2x1_ASAP7_75t_L g15854 ( 
.A(n_15709),
.B(n_7155),
.Y(n_15854)
);

AOI22xp5_ASAP7_75t_L g15855 ( 
.A1(n_15746),
.A2(n_8198),
.B1(n_8244),
.B2(n_8197),
.Y(n_15855)
);

INVx1_ASAP7_75t_L g15856 ( 
.A(n_15603),
.Y(n_15856)
);

NAND2xp5_ASAP7_75t_L g15857 ( 
.A(n_15691),
.B(n_7656),
.Y(n_15857)
);

INVx1_ASAP7_75t_L g15858 ( 
.A(n_15580),
.Y(n_15858)
);

INVx1_ASAP7_75t_L g15859 ( 
.A(n_15679),
.Y(n_15859)
);

OAI22xp5_ASAP7_75t_L g15860 ( 
.A1(n_15591),
.A2(n_7541),
.B1(n_7543),
.B2(n_7493),
.Y(n_15860)
);

INVx1_ASAP7_75t_L g15861 ( 
.A(n_15615),
.Y(n_15861)
);

OR2x2_ASAP7_75t_L g15862 ( 
.A(n_15592),
.B(n_6704),
.Y(n_15862)
);

INVx1_ASAP7_75t_L g15863 ( 
.A(n_15630),
.Y(n_15863)
);

OAI21xp33_ASAP7_75t_L g15864 ( 
.A1(n_15673),
.A2(n_7564),
.B(n_7548),
.Y(n_15864)
);

XOR2xp5_ASAP7_75t_L g15865 ( 
.A(n_15666),
.B(n_7700),
.Y(n_15865)
);

OR2x2_ASAP7_75t_L g15866 ( 
.A(n_15663),
.B(n_6726),
.Y(n_15866)
);

OAI211xp5_ASAP7_75t_L g15867 ( 
.A1(n_15736),
.A2(n_6741),
.B(n_6787),
.C(n_6731),
.Y(n_15867)
);

INVx2_ASAP7_75t_L g15868 ( 
.A(n_15756),
.Y(n_15868)
);

OAI21xp5_ASAP7_75t_SL g15869 ( 
.A1(n_15541),
.A2(n_8244),
.B(n_8198),
.Y(n_15869)
);

NOR2x1_ASAP7_75t_L g15870 ( 
.A(n_15712),
.B(n_15725),
.Y(n_15870)
);

AOI211xp5_ASAP7_75t_L g15871 ( 
.A1(n_15544),
.A2(n_7272),
.B(n_7249),
.C(n_7255),
.Y(n_15871)
);

AOI22xp5_ASAP7_75t_L g15872 ( 
.A1(n_15703),
.A2(n_15726),
.B1(n_15745),
.B2(n_15697),
.Y(n_15872)
);

INVx1_ASAP7_75t_L g15873 ( 
.A(n_15674),
.Y(n_15873)
);

INVxp33_ASAP7_75t_L g15874 ( 
.A(n_15633),
.Y(n_15874)
);

AND2x2_ASAP7_75t_L g15875 ( 
.A(n_15665),
.B(n_7568),
.Y(n_15875)
);

INVx1_ASAP7_75t_L g15876 ( 
.A(n_15728),
.Y(n_15876)
);

AND2x4_ASAP7_75t_L g15877 ( 
.A(n_15647),
.B(n_8244),
.Y(n_15877)
);

OAI21xp5_ASAP7_75t_L g15878 ( 
.A1(n_15708),
.A2(n_7388),
.B(n_7384),
.Y(n_15878)
);

INVx1_ASAP7_75t_L g15879 ( 
.A(n_15668),
.Y(n_15879)
);

INVx1_ASAP7_75t_L g15880 ( 
.A(n_15743),
.Y(n_15880)
);

OAI22xp33_ASAP7_75t_L g15881 ( 
.A1(n_15638),
.A2(n_7543),
.B1(n_7555),
.B2(n_7541),
.Y(n_15881)
);

OAI22xp5_ASAP7_75t_L g15882 ( 
.A1(n_15643),
.A2(n_7543),
.B1(n_7555),
.B2(n_7541),
.Y(n_15882)
);

AND2x2_ASAP7_75t_L g15883 ( 
.A(n_15656),
.B(n_7564),
.Y(n_15883)
);

INVx2_ASAP7_75t_L g15884 ( 
.A(n_15641),
.Y(n_15884)
);

INVx1_ASAP7_75t_L g15885 ( 
.A(n_15751),
.Y(n_15885)
);

AOI22xp33_ASAP7_75t_SL g15886 ( 
.A1(n_15700),
.A2(n_7543),
.B1(n_7555),
.B2(n_7541),
.Y(n_15886)
);

NAND2x1_ASAP7_75t_L g15887 ( 
.A(n_15742),
.B(n_7271),
.Y(n_15887)
);

OAI21xp33_ASAP7_75t_SL g15888 ( 
.A1(n_15618),
.A2(n_15721),
.B(n_15649),
.Y(n_15888)
);

NOR4xp25_ASAP7_75t_L g15889 ( 
.A(n_15731),
.B(n_7656),
.C(n_7668),
.D(n_7659),
.Y(n_15889)
);

AND2x2_ASAP7_75t_L g15890 ( 
.A(n_15759),
.B(n_7568),
.Y(n_15890)
);

NAND2xp5_ASAP7_75t_SL g15891 ( 
.A(n_15586),
.B(n_7541),
.Y(n_15891)
);

OAI21xp5_ASAP7_75t_L g15892 ( 
.A1(n_15715),
.A2(n_7294),
.B(n_7354),
.Y(n_15892)
);

AOI22xp33_ASAP7_75t_L g15893 ( 
.A1(n_15705),
.A2(n_8298),
.B1(n_7668),
.B2(n_7670),
.Y(n_15893)
);

OAI22xp5_ASAP7_75t_SL g15894 ( 
.A1(n_15732),
.A2(n_15741),
.B1(n_15754),
.B2(n_15733),
.Y(n_15894)
);

INVx1_ASAP7_75t_L g15895 ( 
.A(n_15575),
.Y(n_15895)
);

NOR3xp33_ASAP7_75t_L g15896 ( 
.A(n_15602),
.B(n_7495),
.C(n_6678),
.Y(n_15896)
);

AOI211x1_ASAP7_75t_SL g15897 ( 
.A1(n_15685),
.A2(n_15749),
.B(n_15737),
.C(n_15634),
.Y(n_15897)
);

AND2x2_ASAP7_75t_L g15898 ( 
.A(n_15578),
.B(n_7568),
.Y(n_15898)
);

INVx1_ASAP7_75t_L g15899 ( 
.A(n_15639),
.Y(n_15899)
);

NAND4xp25_ASAP7_75t_SL g15900 ( 
.A(n_15563),
.B(n_8225),
.C(n_8234),
.D(n_8133),
.Y(n_15900)
);

AOI22xp5_ASAP7_75t_L g15901 ( 
.A1(n_15719),
.A2(n_8290),
.B1(n_8296),
.B2(n_8244),
.Y(n_15901)
);

OAI31xp33_ASAP7_75t_SL g15902 ( 
.A1(n_15711),
.A2(n_7849),
.A3(n_7853),
.B(n_7520),
.Y(n_15902)
);

INVx1_ASAP7_75t_L g15903 ( 
.A(n_15724),
.Y(n_15903)
);

NOR2xp33_ASAP7_75t_L g15904 ( 
.A(n_15707),
.B(n_7659),
.Y(n_15904)
);

OA21x2_ASAP7_75t_L g15905 ( 
.A1(n_15735),
.A2(n_7177),
.B(n_7175),
.Y(n_15905)
);

AOI22xp5_ASAP7_75t_L g15906 ( 
.A1(n_15740),
.A2(n_8290),
.B1(n_8296),
.B2(n_8244),
.Y(n_15906)
);

INVx1_ASAP7_75t_L g15907 ( 
.A(n_15684),
.Y(n_15907)
);

OAI21xp33_ASAP7_75t_L g15908 ( 
.A1(n_15596),
.A2(n_7592),
.B(n_7568),
.Y(n_15908)
);

OAI21xp5_ASAP7_75t_L g15909 ( 
.A1(n_15585),
.A2(n_7391),
.B(n_7272),
.Y(n_15909)
);

INVx1_ASAP7_75t_L g15910 ( 
.A(n_15637),
.Y(n_15910)
);

A2O1A1Ixp33_ASAP7_75t_L g15911 ( 
.A1(n_15717),
.A2(n_7254),
.B(n_7255),
.C(n_7249),
.Y(n_15911)
);

NAND2xp5_ASAP7_75t_L g15912 ( 
.A(n_15607),
.B(n_7668),
.Y(n_15912)
);

AOI32xp33_ASAP7_75t_L g15913 ( 
.A1(n_15613),
.A2(n_7853),
.A3(n_7849),
.B1(n_7957),
.B2(n_7946),
.Y(n_15913)
);

AOI21xp5_ASAP7_75t_L g15914 ( 
.A1(n_15579),
.A2(n_8234),
.B(n_8225),
.Y(n_15914)
);

INVx2_ASAP7_75t_L g15915 ( 
.A(n_15607),
.Y(n_15915)
);

XNOR2x2_ASAP7_75t_L g15916 ( 
.A(n_15612),
.B(n_7205),
.Y(n_15916)
);

INVx1_ASAP7_75t_SL g15917 ( 
.A(n_15671),
.Y(n_15917)
);

INVx1_ASAP7_75t_L g15918 ( 
.A(n_15748),
.Y(n_15918)
);

NAND2xp5_ASAP7_75t_L g15919 ( 
.A(n_15698),
.B(n_7670),
.Y(n_15919)
);

OR2x2_ASAP7_75t_L g15920 ( 
.A(n_15621),
.B(n_6741),
.Y(n_15920)
);

AOI322xp5_ASAP7_75t_L g15921 ( 
.A1(n_15644),
.A2(n_7678),
.A3(n_7685),
.B1(n_7690),
.B2(n_7710),
.C1(n_7697),
.C2(n_7670),
.Y(n_15921)
);

AOI322xp5_ASAP7_75t_L g15922 ( 
.A1(n_15609),
.A2(n_15628),
.A3(n_15562),
.B1(n_15693),
.B2(n_15651),
.C1(n_15567),
.C2(n_15692),
.Y(n_15922)
);

INVx1_ASAP7_75t_L g15923 ( 
.A(n_15672),
.Y(n_15923)
);

INVxp67_ASAP7_75t_L g15924 ( 
.A(n_15623),
.Y(n_15924)
);

AOI22xp5_ASAP7_75t_L g15925 ( 
.A1(n_15565),
.A2(n_8290),
.B1(n_8296),
.B2(n_7785),
.Y(n_15925)
);

INVx1_ASAP7_75t_L g15926 ( 
.A(n_15730),
.Y(n_15926)
);

AOI21xp33_ASAP7_75t_R g15927 ( 
.A1(n_15710),
.A2(n_8241),
.B(n_8239),
.Y(n_15927)
);

NAND4xp25_ASAP7_75t_L g15928 ( 
.A(n_15629),
.B(n_8296),
.C(n_8290),
.D(n_6709),
.Y(n_15928)
);

INVx1_ASAP7_75t_L g15929 ( 
.A(n_15747),
.Y(n_15929)
);

INVx2_ASAP7_75t_L g15930 ( 
.A(n_15693),
.Y(n_15930)
);

OAI21xp5_ASAP7_75t_L g15931 ( 
.A1(n_15655),
.A2(n_7391),
.B(n_7254),
.Y(n_15931)
);

OAI22xp5_ASAP7_75t_L g15932 ( 
.A1(n_15689),
.A2(n_7555),
.B1(n_7589),
.B2(n_7543),
.Y(n_15932)
);

INVx2_ASAP7_75t_L g15933 ( 
.A(n_15722),
.Y(n_15933)
);

INVx1_ASAP7_75t_L g15934 ( 
.A(n_15686),
.Y(n_15934)
);

OR2x2_ASAP7_75t_L g15935 ( 
.A(n_15690),
.B(n_6787),
.Y(n_15935)
);

NAND2xp5_ASAP7_75t_L g15936 ( 
.A(n_15758),
.B(n_7685),
.Y(n_15936)
);

AOI21xp5_ASAP7_75t_L g15937 ( 
.A1(n_15626),
.A2(n_8241),
.B(n_8239),
.Y(n_15937)
);

OAI322xp33_ASAP7_75t_L g15938 ( 
.A1(n_15616),
.A2(n_8241),
.A3(n_8242),
.B1(n_8239),
.B2(n_6967),
.C1(n_6931),
.C2(n_6989),
.Y(n_15938)
);

INVx1_ASAP7_75t_L g15939 ( 
.A(n_15720),
.Y(n_15939)
);

NOR2xp33_ASAP7_75t_L g15940 ( 
.A(n_15704),
.B(n_7678),
.Y(n_15940)
);

AOI32xp33_ASAP7_75t_L g15941 ( 
.A1(n_15727),
.A2(n_7957),
.A3(n_7946),
.B1(n_8290),
.B2(n_7311),
.Y(n_15941)
);

NAND2xp5_ASAP7_75t_L g15942 ( 
.A(n_15695),
.B(n_15753),
.Y(n_15942)
);

INVx2_ASAP7_75t_L g15943 ( 
.A(n_15667),
.Y(n_15943)
);

AND2x2_ASAP7_75t_L g15944 ( 
.A(n_15635),
.B(n_7592),
.Y(n_15944)
);

INVx2_ASAP7_75t_L g15945 ( 
.A(n_15645),
.Y(n_15945)
);

INVx2_ASAP7_75t_L g15946 ( 
.A(n_15601),
.Y(n_15946)
);

OAI221xp5_ASAP7_75t_SL g15947 ( 
.A1(n_15574),
.A2(n_7066),
.B1(n_6998),
.B2(n_6904),
.C(n_7191),
.Y(n_15947)
);

OAI21xp5_ASAP7_75t_L g15948 ( 
.A1(n_15564),
.A2(n_7391),
.B(n_7254),
.Y(n_15948)
);

HB1xp67_ASAP7_75t_L g15949 ( 
.A(n_15646),
.Y(n_15949)
);

INVxp67_ASAP7_75t_SL g15950 ( 
.A(n_15646),
.Y(n_15950)
);

NAND2xp5_ASAP7_75t_L g15951 ( 
.A(n_15543),
.B(n_7678),
.Y(n_15951)
);

NAND4xp25_ASAP7_75t_L g15952 ( 
.A(n_15588),
.B(n_6709),
.C(n_6735),
.D(n_6706),
.Y(n_15952)
);

NOR2xp33_ASAP7_75t_L g15953 ( 
.A(n_15538),
.B(n_7678),
.Y(n_15953)
);

INVx1_ASAP7_75t_L g15954 ( 
.A(n_15706),
.Y(n_15954)
);

INVx1_ASAP7_75t_L g15955 ( 
.A(n_15706),
.Y(n_15955)
);

AOI22xp5_ASAP7_75t_L g15956 ( 
.A1(n_15581),
.A2(n_7785),
.B1(n_7805),
.B2(n_7777),
.Y(n_15956)
);

AOI321xp33_ASAP7_75t_L g15957 ( 
.A1(n_15676),
.A2(n_7700),
.A3(n_7709),
.B1(n_7705),
.B2(n_7785),
.C(n_7777),
.Y(n_15957)
);

OR2x2_ASAP7_75t_L g15958 ( 
.A(n_15543),
.B(n_6788),
.Y(n_15958)
);

OR2x6_ASAP7_75t_L g15959 ( 
.A(n_15538),
.B(n_5952),
.Y(n_15959)
);

OR2x2_ASAP7_75t_L g15960 ( 
.A(n_15949),
.B(n_6788),
.Y(n_15960)
);

NAND2xp5_ASAP7_75t_L g15961 ( 
.A(n_15950),
.B(n_7685),
.Y(n_15961)
);

NAND2xp5_ASAP7_75t_L g15962 ( 
.A(n_15784),
.B(n_7690),
.Y(n_15962)
);

AND2x2_ASAP7_75t_L g15963 ( 
.A(n_15762),
.B(n_7592),
.Y(n_15963)
);

NAND2xp5_ASAP7_75t_L g15964 ( 
.A(n_15773),
.B(n_7690),
.Y(n_15964)
);

NOR2xp33_ASAP7_75t_L g15965 ( 
.A(n_15785),
.B(n_7697),
.Y(n_15965)
);

AND2x2_ASAP7_75t_L g15966 ( 
.A(n_15763),
.B(n_7592),
.Y(n_15966)
);

INVx2_ASAP7_75t_L g15967 ( 
.A(n_15796),
.Y(n_15967)
);

INVxp67_ASAP7_75t_L g15968 ( 
.A(n_15790),
.Y(n_15968)
);

AND2x2_ASAP7_75t_L g15969 ( 
.A(n_15803),
.B(n_7646),
.Y(n_15969)
);

OR2x2_ASAP7_75t_L g15970 ( 
.A(n_15830),
.B(n_6816),
.Y(n_15970)
);

NAND2xp5_ASAP7_75t_L g15971 ( 
.A(n_15798),
.B(n_7697),
.Y(n_15971)
);

NAND2xp5_ASAP7_75t_SL g15972 ( 
.A(n_15823),
.B(n_7555),
.Y(n_15972)
);

NAND2xp5_ASAP7_75t_L g15973 ( 
.A(n_15849),
.B(n_7697),
.Y(n_15973)
);

NAND2xp5_ASAP7_75t_L g15974 ( 
.A(n_15777),
.B(n_7710),
.Y(n_15974)
);

INVx2_ASAP7_75t_L g15975 ( 
.A(n_15771),
.Y(n_15975)
);

INVx1_ASAP7_75t_L g15976 ( 
.A(n_15809),
.Y(n_15976)
);

AND2x2_ASAP7_75t_L g15977 ( 
.A(n_15875),
.B(n_7646),
.Y(n_15977)
);

AND2x4_ASAP7_75t_L g15978 ( 
.A(n_15870),
.B(n_7646),
.Y(n_15978)
);

NOR2x1_ASAP7_75t_L g15979 ( 
.A(n_15954),
.B(n_7155),
.Y(n_15979)
);

INVx1_ASAP7_75t_SL g15980 ( 
.A(n_15808),
.Y(n_15980)
);

INVx1_ASAP7_75t_L g15981 ( 
.A(n_15955),
.Y(n_15981)
);

INVx1_ASAP7_75t_SL g15982 ( 
.A(n_15774),
.Y(n_15982)
);

AOI22xp5_ASAP7_75t_L g15983 ( 
.A1(n_15765),
.A2(n_7785),
.B1(n_7805),
.B2(n_7777),
.Y(n_15983)
);

NOR3xp33_ASAP7_75t_L g15984 ( 
.A(n_15766),
.B(n_6678),
.C(n_7495),
.Y(n_15984)
);

OR2x2_ASAP7_75t_L g15985 ( 
.A(n_15783),
.B(n_6846),
.Y(n_15985)
);

NAND2xp5_ASAP7_75t_L g15986 ( 
.A(n_15843),
.B(n_7710),
.Y(n_15986)
);

AND2x2_ASAP7_75t_L g15987 ( 
.A(n_15883),
.B(n_7671),
.Y(n_15987)
);

NAND2xp5_ASAP7_75t_L g15988 ( 
.A(n_15792),
.B(n_7710),
.Y(n_15988)
);

NAND2xp5_ASAP7_75t_L g15989 ( 
.A(n_15930),
.B(n_7711),
.Y(n_15989)
);

AND2x2_ASAP7_75t_L g15990 ( 
.A(n_15813),
.B(n_7671),
.Y(n_15990)
);

INVx1_ASAP7_75t_L g15991 ( 
.A(n_15804),
.Y(n_15991)
);

INVxp67_ASAP7_75t_L g15992 ( 
.A(n_15805),
.Y(n_15992)
);

AO21x1_ASAP7_75t_L g15993 ( 
.A1(n_15828),
.A2(n_8242),
.B(n_8051),
.Y(n_15993)
);

NAND2xp5_ASAP7_75t_L g15994 ( 
.A(n_15880),
.B(n_7711),
.Y(n_15994)
);

INVx1_ASAP7_75t_L g15995 ( 
.A(n_15797),
.Y(n_15995)
);

INVx1_ASAP7_75t_SL g15996 ( 
.A(n_15817),
.Y(n_15996)
);

AND2x2_ASAP7_75t_L g15997 ( 
.A(n_15788),
.B(n_7671),
.Y(n_15997)
);

INVx2_ASAP7_75t_SL g15998 ( 
.A(n_15854),
.Y(n_15998)
);

INVx1_ASAP7_75t_L g15999 ( 
.A(n_15812),
.Y(n_15999)
);

AND2x2_ASAP7_75t_L g16000 ( 
.A(n_15825),
.B(n_7671),
.Y(n_16000)
);

NAND2xp5_ASAP7_75t_L g16001 ( 
.A(n_15923),
.B(n_7711),
.Y(n_16001)
);

INVx1_ASAP7_75t_SL g16002 ( 
.A(n_15814),
.Y(n_16002)
);

INVx1_ASAP7_75t_L g16003 ( 
.A(n_15816),
.Y(n_16003)
);

INVx1_ASAP7_75t_L g16004 ( 
.A(n_15833),
.Y(n_16004)
);

INVxp67_ASAP7_75t_L g16005 ( 
.A(n_15879),
.Y(n_16005)
);

HB1xp67_ASAP7_75t_L g16006 ( 
.A(n_15818),
.Y(n_16006)
);

INVx1_ASAP7_75t_L g16007 ( 
.A(n_15821),
.Y(n_16007)
);

NAND2xp5_ASAP7_75t_L g16008 ( 
.A(n_15884),
.B(n_7711),
.Y(n_16008)
);

NAND2xp5_ASAP7_75t_L g16009 ( 
.A(n_15825),
.B(n_15943),
.Y(n_16009)
);

NAND2xp5_ASAP7_75t_L g16010 ( 
.A(n_15831),
.B(n_7719),
.Y(n_16010)
);

AND2x2_ASAP7_75t_L g16011 ( 
.A(n_15877),
.B(n_7671),
.Y(n_16011)
);

INVx1_ASAP7_75t_L g16012 ( 
.A(n_15772),
.Y(n_16012)
);

NOR2x1_ASAP7_75t_L g16013 ( 
.A(n_15846),
.B(n_7155),
.Y(n_16013)
);

OR2x2_ASAP7_75t_L g16014 ( 
.A(n_15952),
.B(n_6846),
.Y(n_16014)
);

INVx1_ASAP7_75t_L g16015 ( 
.A(n_15958),
.Y(n_16015)
);

INVx1_ASAP7_75t_L g16016 ( 
.A(n_15951),
.Y(n_16016)
);

INVx1_ASAP7_75t_L g16017 ( 
.A(n_15915),
.Y(n_16017)
);

AND2x2_ASAP7_75t_SL g16018 ( 
.A(n_15810),
.B(n_8023),
.Y(n_16018)
);

HB1xp67_ASAP7_75t_L g16019 ( 
.A(n_15858),
.Y(n_16019)
);

INVxp67_ASAP7_75t_L g16020 ( 
.A(n_15806),
.Y(n_16020)
);

NAND2xp5_ASAP7_75t_L g16021 ( 
.A(n_15872),
.B(n_15907),
.Y(n_16021)
);

INVx1_ASAP7_75t_L g16022 ( 
.A(n_15820),
.Y(n_16022)
);

AND2x2_ASAP7_75t_L g16023 ( 
.A(n_15890),
.B(n_6504),
.Y(n_16023)
);

NOR2xp33_ASAP7_75t_L g16024 ( 
.A(n_15934),
.B(n_7719),
.Y(n_16024)
);

AOI22xp5_ASAP7_75t_L g16025 ( 
.A1(n_15929),
.A2(n_7785),
.B1(n_7805),
.B2(n_7777),
.Y(n_16025)
);

NAND2xp5_ASAP7_75t_L g16026 ( 
.A(n_15903),
.B(n_7719),
.Y(n_16026)
);

AND2x2_ASAP7_75t_L g16027 ( 
.A(n_15944),
.B(n_6540),
.Y(n_16027)
);

AND2x2_ASAP7_75t_L g16028 ( 
.A(n_15959),
.B(n_6546),
.Y(n_16028)
);

INVx1_ASAP7_75t_L g16029 ( 
.A(n_15894),
.Y(n_16029)
);

NOR2x1_ASAP7_75t_L g16030 ( 
.A(n_15876),
.B(n_6142),
.Y(n_16030)
);

INVx1_ASAP7_75t_L g16031 ( 
.A(n_15800),
.Y(n_16031)
);

INVxp67_ASAP7_75t_L g16032 ( 
.A(n_15859),
.Y(n_16032)
);

INVx2_ASAP7_75t_L g16033 ( 
.A(n_15916),
.Y(n_16033)
);

INVx1_ASAP7_75t_L g16034 ( 
.A(n_15838),
.Y(n_16034)
);

INVx1_ASAP7_75t_SL g16035 ( 
.A(n_15917),
.Y(n_16035)
);

NAND2xp5_ASAP7_75t_SL g16036 ( 
.A(n_15946),
.B(n_7555),
.Y(n_16036)
);

OR2x2_ASAP7_75t_L g16037 ( 
.A(n_15775),
.B(n_6847),
.Y(n_16037)
);

INVx1_ASAP7_75t_L g16038 ( 
.A(n_15787),
.Y(n_16038)
);

NAND2xp5_ASAP7_75t_L g16039 ( 
.A(n_15781),
.B(n_7719),
.Y(n_16039)
);

INVx1_ASAP7_75t_L g16040 ( 
.A(n_15782),
.Y(n_16040)
);

OR2x2_ASAP7_75t_L g16041 ( 
.A(n_15776),
.B(n_7930),
.Y(n_16041)
);

NOR3xp33_ASAP7_75t_L g16042 ( 
.A(n_15856),
.B(n_15873),
.C(n_15861),
.Y(n_16042)
);

NAND2xp5_ASAP7_75t_L g16043 ( 
.A(n_15850),
.B(n_7723),
.Y(n_16043)
);

AND2x2_ASAP7_75t_L g16044 ( 
.A(n_15959),
.B(n_6546),
.Y(n_16044)
);

INVx2_ASAP7_75t_L g16045 ( 
.A(n_15794),
.Y(n_16045)
);

NAND2xp5_ASAP7_75t_L g16046 ( 
.A(n_15863),
.B(n_7723),
.Y(n_16046)
);

NOR2xp67_ASAP7_75t_L g16047 ( 
.A(n_15761),
.B(n_6964),
.Y(n_16047)
);

NOR2xp33_ASAP7_75t_L g16048 ( 
.A(n_15760),
.B(n_7723),
.Y(n_16048)
);

NAND2xp5_ASAP7_75t_L g16049 ( 
.A(n_15899),
.B(n_7723),
.Y(n_16049)
);

INVx1_ASAP7_75t_L g16050 ( 
.A(n_15807),
.Y(n_16050)
);

NAND2xp5_ASAP7_75t_L g16051 ( 
.A(n_15918),
.B(n_7725),
.Y(n_16051)
);

NAND2xp5_ASAP7_75t_L g16052 ( 
.A(n_15895),
.B(n_7725),
.Y(n_16052)
);

INVx1_ASAP7_75t_SL g16053 ( 
.A(n_15885),
.Y(n_16053)
);

INVx1_ASAP7_75t_L g16054 ( 
.A(n_15837),
.Y(n_16054)
);

NOR2xp33_ASAP7_75t_L g16055 ( 
.A(n_15910),
.B(n_7725),
.Y(n_16055)
);

AND2x2_ASAP7_75t_L g16056 ( 
.A(n_15898),
.B(n_6546),
.Y(n_16056)
);

AND2x2_ASAP7_75t_L g16057 ( 
.A(n_15811),
.B(n_6564),
.Y(n_16057)
);

AOI22xp5_ASAP7_75t_L g16058 ( 
.A1(n_15939),
.A2(n_7805),
.B1(n_7896),
.B2(n_7777),
.Y(n_16058)
);

INVx2_ASAP7_75t_L g16059 ( 
.A(n_15794),
.Y(n_16059)
);

AOI222xp33_ASAP7_75t_L g16060 ( 
.A1(n_15824),
.A2(n_7725),
.B1(n_7738),
.B2(n_7746),
.C1(n_7744),
.C2(n_7734),
.Y(n_16060)
);

INVx1_ASAP7_75t_L g16061 ( 
.A(n_15857),
.Y(n_16061)
);

NAND2xp5_ASAP7_75t_SL g16062 ( 
.A(n_15945),
.B(n_7555),
.Y(n_16062)
);

OR2x2_ASAP7_75t_L g16063 ( 
.A(n_15829),
.B(n_7930),
.Y(n_16063)
);

OAI222xp33_ASAP7_75t_L g16064 ( 
.A1(n_15924),
.A2(n_7746),
.B1(n_7738),
.B2(n_7773),
.C1(n_7744),
.C2(n_7734),
.Y(n_16064)
);

INVx2_ASAP7_75t_L g16065 ( 
.A(n_15862),
.Y(n_16065)
);

INVx2_ASAP7_75t_L g16066 ( 
.A(n_15866),
.Y(n_16066)
);

NAND2xp5_ASAP7_75t_L g16067 ( 
.A(n_15822),
.B(n_7734),
.Y(n_16067)
);

INVx2_ASAP7_75t_L g16068 ( 
.A(n_15834),
.Y(n_16068)
);

INVxp67_ASAP7_75t_L g16069 ( 
.A(n_15953),
.Y(n_16069)
);

NOR2xp33_ASAP7_75t_SL g16070 ( 
.A(n_15826),
.B(n_6002),
.Y(n_16070)
);

OR2x2_ASAP7_75t_L g16071 ( 
.A(n_15920),
.B(n_7930),
.Y(n_16071)
);

INVx1_ASAP7_75t_L g16072 ( 
.A(n_15933),
.Y(n_16072)
);

NAND2x1_ASAP7_75t_SL g16073 ( 
.A(n_15926),
.B(n_8242),
.Y(n_16073)
);

INVx1_ASAP7_75t_L g16074 ( 
.A(n_15819),
.Y(n_16074)
);

INVx2_ASAP7_75t_L g16075 ( 
.A(n_15802),
.Y(n_16075)
);

INVx1_ASAP7_75t_L g16076 ( 
.A(n_15897),
.Y(n_16076)
);

AOI22xp33_ASAP7_75t_L g16077 ( 
.A1(n_15893),
.A2(n_7738),
.B1(n_7744),
.B2(n_7734),
.Y(n_16077)
);

NAND2x1_ASAP7_75t_L g16078 ( 
.A(n_15868),
.B(n_15770),
.Y(n_16078)
);

NOR2xp33_ASAP7_75t_L g16079 ( 
.A(n_15779),
.B(n_8275),
.Y(n_16079)
);

INVx1_ASAP7_75t_L g16080 ( 
.A(n_15900),
.Y(n_16080)
);

OR2x2_ASAP7_75t_L g16081 ( 
.A(n_15935),
.B(n_7930),
.Y(n_16081)
);

NAND2xp5_ASAP7_75t_L g16082 ( 
.A(n_15827),
.B(n_7738),
.Y(n_16082)
);

HB1xp67_ASAP7_75t_L g16083 ( 
.A(n_15888),
.Y(n_16083)
);

AOI22xp33_ASAP7_75t_L g16084 ( 
.A1(n_15896),
.A2(n_7773),
.B1(n_7775),
.B2(n_7746),
.Y(n_16084)
);

AND2x2_ASAP7_75t_L g16085 ( 
.A(n_15791),
.B(n_6564),
.Y(n_16085)
);

INVx1_ASAP7_75t_L g16086 ( 
.A(n_15768),
.Y(n_16086)
);

AND2x2_ASAP7_75t_L g16087 ( 
.A(n_15874),
.B(n_6564),
.Y(n_16087)
);

NAND2x1_ASAP7_75t_SL g16088 ( 
.A(n_15842),
.B(n_7805),
.Y(n_16088)
);

INVx1_ASAP7_75t_L g16089 ( 
.A(n_15912),
.Y(n_16089)
);

NAND2xp5_ASAP7_75t_L g16090 ( 
.A(n_15927),
.B(n_7746),
.Y(n_16090)
);

NAND2xp5_ASAP7_75t_L g16091 ( 
.A(n_15922),
.B(n_7773),
.Y(n_16091)
);

INVx1_ASAP7_75t_L g16092 ( 
.A(n_15919),
.Y(n_16092)
);

INVx1_ASAP7_75t_L g16093 ( 
.A(n_15942),
.Y(n_16093)
);

BUFx2_ASAP7_75t_SL g16094 ( 
.A(n_15847),
.Y(n_16094)
);

INVx1_ASAP7_75t_L g16095 ( 
.A(n_15865),
.Y(n_16095)
);

NOR2x1_ASAP7_75t_L g16096 ( 
.A(n_15869),
.B(n_15928),
.Y(n_16096)
);

NAND2xp5_ASAP7_75t_L g16097 ( 
.A(n_15851),
.B(n_7775),
.Y(n_16097)
);

NOR2xp33_ASAP7_75t_L g16098 ( 
.A(n_15801),
.B(n_7775),
.Y(n_16098)
);

NOR2xp33_ASAP7_75t_L g16099 ( 
.A(n_15789),
.B(n_7775),
.Y(n_16099)
);

NAND2xp5_ASAP7_75t_L g16100 ( 
.A(n_15889),
.B(n_7794),
.Y(n_16100)
);

OR2x2_ASAP7_75t_L g16101 ( 
.A(n_15878),
.B(n_7930),
.Y(n_16101)
);

NAND2xp5_ASAP7_75t_L g16102 ( 
.A(n_15904),
.B(n_7794),
.Y(n_16102)
);

INVx1_ASAP7_75t_L g16103 ( 
.A(n_15936),
.Y(n_16103)
);

NAND2xp5_ASAP7_75t_L g16104 ( 
.A(n_15871),
.B(n_7794),
.Y(n_16104)
);

NAND2xp5_ASAP7_75t_L g16105 ( 
.A(n_15940),
.B(n_7794),
.Y(n_16105)
);

AND2x2_ASAP7_75t_L g16106 ( 
.A(n_15793),
.B(n_6610),
.Y(n_16106)
);

INVxp33_ASAP7_75t_L g16107 ( 
.A(n_15887),
.Y(n_16107)
);

INVxp67_ASAP7_75t_SL g16108 ( 
.A(n_15769),
.Y(n_16108)
);

NAND2xp5_ASAP7_75t_L g16109 ( 
.A(n_15909),
.B(n_7803),
.Y(n_16109)
);

NAND2xp5_ASAP7_75t_L g16110 ( 
.A(n_15764),
.B(n_7803),
.Y(n_16110)
);

NAND2xp5_ASAP7_75t_L g16111 ( 
.A(n_15795),
.B(n_7803),
.Y(n_16111)
);

INVx1_ASAP7_75t_L g16112 ( 
.A(n_15867),
.Y(n_16112)
);

NAND2xp5_ASAP7_75t_L g16113 ( 
.A(n_15767),
.B(n_7803),
.Y(n_16113)
);

NOR2xp33_ASAP7_75t_L g16114 ( 
.A(n_15947),
.B(n_15938),
.Y(n_16114)
);

INVx1_ASAP7_75t_L g16115 ( 
.A(n_15839),
.Y(n_16115)
);

NOR2xp33_ASAP7_75t_L g16116 ( 
.A(n_15778),
.B(n_7840),
.Y(n_16116)
);

AND2x2_ASAP7_75t_L g16117 ( 
.A(n_15855),
.B(n_6610),
.Y(n_16117)
);

INVx1_ASAP7_75t_L g16118 ( 
.A(n_15799),
.Y(n_16118)
);

OAI22xp5_ASAP7_75t_L g16119 ( 
.A1(n_15815),
.A2(n_7555),
.B1(n_7837),
.B2(n_7589),
.Y(n_16119)
);

INVx2_ASAP7_75t_L g16120 ( 
.A(n_15891),
.Y(n_16120)
);

INVx2_ASAP7_75t_SL g16121 ( 
.A(n_15780),
.Y(n_16121)
);

AND2x2_ASAP7_75t_L g16122 ( 
.A(n_15956),
.B(n_6610),
.Y(n_16122)
);

INVx1_ASAP7_75t_SL g16123 ( 
.A(n_15852),
.Y(n_16123)
);

INVx1_ASAP7_75t_SL g16124 ( 
.A(n_15937),
.Y(n_16124)
);

OAI22xp5_ASAP7_75t_L g16125 ( 
.A1(n_15835),
.A2(n_7589),
.B1(n_7862),
.B2(n_7837),
.Y(n_16125)
);

OR2x2_ASAP7_75t_L g16126 ( 
.A(n_15786),
.B(n_15864),
.Y(n_16126)
);

INVx1_ASAP7_75t_L g16127 ( 
.A(n_15840),
.Y(n_16127)
);

AND2x2_ASAP7_75t_L g16128 ( 
.A(n_15906),
.B(n_6624),
.Y(n_16128)
);

INVx1_ASAP7_75t_L g16129 ( 
.A(n_15832),
.Y(n_16129)
);

NOR2xp67_ASAP7_75t_L g16130 ( 
.A(n_15914),
.B(n_6964),
.Y(n_16130)
);

INVx1_ASAP7_75t_SL g16131 ( 
.A(n_15948),
.Y(n_16131)
);

INVx1_ASAP7_75t_L g16132 ( 
.A(n_15836),
.Y(n_16132)
);

NAND2xp5_ASAP7_75t_L g16133 ( 
.A(n_15845),
.B(n_7840),
.Y(n_16133)
);

BUFx2_ASAP7_75t_L g16134 ( 
.A(n_15892),
.Y(n_16134)
);

OR2x2_ASAP7_75t_L g16135 ( 
.A(n_15911),
.B(n_7930),
.Y(n_16135)
);

INVx1_ASAP7_75t_L g16136 ( 
.A(n_15931),
.Y(n_16136)
);

INVx1_ASAP7_75t_L g16137 ( 
.A(n_15905),
.Y(n_16137)
);

NAND2x1_ASAP7_75t_L g16138 ( 
.A(n_15905),
.B(n_7271),
.Y(n_16138)
);

INVx1_ASAP7_75t_L g16139 ( 
.A(n_15841),
.Y(n_16139)
);

BUFx4f_ASAP7_75t_SL g16140 ( 
.A(n_15957),
.Y(n_16140)
);

NAND2xp5_ASAP7_75t_L g16141 ( 
.A(n_15902),
.B(n_7840),
.Y(n_16141)
);

AND2x2_ASAP7_75t_L g16142 ( 
.A(n_15908),
.B(n_6624),
.Y(n_16142)
);

AND2x2_ASAP7_75t_L g16143 ( 
.A(n_15925),
.B(n_6624),
.Y(n_16143)
);

NAND2xp5_ASAP7_75t_L g16144 ( 
.A(n_15913),
.B(n_7840),
.Y(n_16144)
);

NAND2xp5_ASAP7_75t_L g16145 ( 
.A(n_15921),
.B(n_7846),
.Y(n_16145)
);

INVx1_ASAP7_75t_SL g16146 ( 
.A(n_15886),
.Y(n_16146)
);

OR2x2_ASAP7_75t_L g16147 ( 
.A(n_15932),
.B(n_15860),
.Y(n_16147)
);

NAND2xp5_ASAP7_75t_L g16148 ( 
.A(n_15848),
.B(n_15941),
.Y(n_16148)
);

NAND2xp5_ASAP7_75t_L g16149 ( 
.A(n_15881),
.B(n_7846),
.Y(n_16149)
);

INVx1_ASAP7_75t_L g16150 ( 
.A(n_15882),
.Y(n_16150)
);

AOI22xp33_ASAP7_75t_L g16151 ( 
.A1(n_15901),
.A2(n_7850),
.B1(n_7875),
.B2(n_7846),
.Y(n_16151)
);

NAND2xp5_ASAP7_75t_L g16152 ( 
.A(n_15844),
.B(n_7846),
.Y(n_16152)
);

AND2x4_ASAP7_75t_L g16153 ( 
.A(n_15853),
.B(n_7589),
.Y(n_16153)
);

OR2x2_ASAP7_75t_L g16154 ( 
.A(n_15949),
.B(n_8046),
.Y(n_16154)
);

INVx1_ASAP7_75t_L g16155 ( 
.A(n_15949),
.Y(n_16155)
);

INVx1_ASAP7_75t_SL g16156 ( 
.A(n_15784),
.Y(n_16156)
);

INVx1_ASAP7_75t_L g16157 ( 
.A(n_15949),
.Y(n_16157)
);

NAND2xp5_ASAP7_75t_L g16158 ( 
.A(n_15950),
.B(n_7850),
.Y(n_16158)
);

AOI22xp5_ASAP7_75t_L g16159 ( 
.A1(n_15950),
.A2(n_7900),
.B1(n_7908),
.B2(n_7896),
.Y(n_16159)
);

AND2x2_ASAP7_75t_L g16160 ( 
.A(n_15950),
.B(n_6673),
.Y(n_16160)
);

NOR2xp33_ASAP7_75t_L g16161 ( 
.A(n_15949),
.B(n_8275),
.Y(n_16161)
);

NAND2xp5_ASAP7_75t_L g16162 ( 
.A(n_15950),
.B(n_7850),
.Y(n_16162)
);

NAND2xp5_ASAP7_75t_L g16163 ( 
.A(n_15950),
.B(n_7850),
.Y(n_16163)
);

INVx1_ASAP7_75t_L g16164 ( 
.A(n_15949),
.Y(n_16164)
);

AND2x2_ASAP7_75t_L g16165 ( 
.A(n_15950),
.B(n_6673),
.Y(n_16165)
);

OR2x2_ASAP7_75t_L g16166 ( 
.A(n_16156),
.B(n_8046),
.Y(n_16166)
);

NOR2x1_ASAP7_75t_L g16167 ( 
.A(n_16155),
.B(n_7896),
.Y(n_16167)
);

NAND2xp5_ASAP7_75t_L g16168 ( 
.A(n_16083),
.B(n_7902),
.Y(n_16168)
);

INVx1_ASAP7_75t_SL g16169 ( 
.A(n_15982),
.Y(n_16169)
);

INVx1_ASAP7_75t_L g16170 ( 
.A(n_16019),
.Y(n_16170)
);

OAI21xp5_ASAP7_75t_L g16171 ( 
.A1(n_16157),
.A2(n_7473),
.B(n_7255),
.Y(n_16171)
);

OAI22xp5_ASAP7_75t_L g16172 ( 
.A1(n_16005),
.A2(n_16164),
.B1(n_15981),
.B2(n_16140),
.Y(n_16172)
);

NAND2xp5_ASAP7_75t_L g16173 ( 
.A(n_15978),
.B(n_7936),
.Y(n_16173)
);

INVx1_ASAP7_75t_L g16174 ( 
.A(n_16006),
.Y(n_16174)
);

INVx1_ASAP7_75t_L g16175 ( 
.A(n_16160),
.Y(n_16175)
);

INVx2_ASAP7_75t_L g16176 ( 
.A(n_15978),
.Y(n_16176)
);

NOR3xp33_ASAP7_75t_SL g16177 ( 
.A(n_16076),
.B(n_6080),
.C(n_6002),
.Y(n_16177)
);

INVx1_ASAP7_75t_L g16178 ( 
.A(n_16165),
.Y(n_16178)
);

NAND2xp5_ASAP7_75t_SL g16179 ( 
.A(n_15967),
.B(n_7589),
.Y(n_16179)
);

INVx1_ASAP7_75t_L g16180 ( 
.A(n_16035),
.Y(n_16180)
);

AND2x2_ASAP7_75t_L g16181 ( 
.A(n_15966),
.B(n_6673),
.Y(n_16181)
);

BUFx2_ASAP7_75t_L g16182 ( 
.A(n_16013),
.Y(n_16182)
);

OR2x2_ASAP7_75t_L g16183 ( 
.A(n_15996),
.B(n_16002),
.Y(n_16183)
);

OAI211xp5_ASAP7_75t_L g16184 ( 
.A1(n_15968),
.A2(n_7589),
.B(n_7862),
.C(n_7837),
.Y(n_16184)
);

AND2x2_ASAP7_75t_L g16185 ( 
.A(n_15969),
.B(n_6675),
.Y(n_16185)
);

AOI22xp33_ASAP7_75t_L g16186 ( 
.A1(n_15975),
.A2(n_7888),
.B1(n_7902),
.B2(n_7875),
.Y(n_16186)
);

NAND2xp5_ASAP7_75t_L g16187 ( 
.A(n_15980),
.B(n_16053),
.Y(n_16187)
);

NAND2xp5_ASAP7_75t_SL g16188 ( 
.A(n_15976),
.B(n_7589),
.Y(n_16188)
);

INVxp67_ASAP7_75t_L g16189 ( 
.A(n_16009),
.Y(n_16189)
);

INVx1_ASAP7_75t_L g16190 ( 
.A(n_16072),
.Y(n_16190)
);

XOR2xp5_ASAP7_75t_L g16191 ( 
.A(n_16093),
.B(n_7700),
.Y(n_16191)
);

INVx1_ASAP7_75t_L g16192 ( 
.A(n_16045),
.Y(n_16192)
);

INVx1_ASAP7_75t_L g16193 ( 
.A(n_16059),
.Y(n_16193)
);

INVx1_ASAP7_75t_L g16194 ( 
.A(n_16137),
.Y(n_16194)
);

XNOR2xp5_ASAP7_75t_L g16195 ( 
.A(n_16047),
.B(n_7700),
.Y(n_16195)
);

INVx1_ASAP7_75t_L g16196 ( 
.A(n_16073),
.Y(n_16196)
);

INVx1_ASAP7_75t_L g16197 ( 
.A(n_15991),
.Y(n_16197)
);

NAND2xp5_ASAP7_75t_SL g16198 ( 
.A(n_15995),
.B(n_7589),
.Y(n_16198)
);

NAND2x1_ASAP7_75t_L g16199 ( 
.A(n_15979),
.B(n_7271),
.Y(n_16199)
);

OAI322xp33_ASAP7_75t_L g16200 ( 
.A1(n_16070),
.A2(n_7066),
.A3(n_6648),
.B1(n_6575),
.B2(n_7906),
.C1(n_7862),
.C2(n_7837),
.Y(n_16200)
);

INVx1_ASAP7_75t_L g16201 ( 
.A(n_15999),
.Y(n_16201)
);

NOR3xp33_ASAP7_75t_SL g16202 ( 
.A(n_16021),
.B(n_6080),
.C(n_6002),
.Y(n_16202)
);

AND2x2_ASAP7_75t_L g16203 ( 
.A(n_15963),
.B(n_6675),
.Y(n_16203)
);

INVx1_ASAP7_75t_L g16204 ( 
.A(n_16003),
.Y(n_16204)
);

AOI21xp5_ASAP7_75t_L g16205 ( 
.A1(n_16036),
.A2(n_7261),
.B(n_7249),
.Y(n_16205)
);

INVx1_ASAP7_75t_L g16206 ( 
.A(n_16004),
.Y(n_16206)
);

NOR3xp33_ASAP7_75t_L g16207 ( 
.A(n_16020),
.B(n_6678),
.C(n_7465),
.Y(n_16207)
);

INVx1_ASAP7_75t_L g16208 ( 
.A(n_15960),
.Y(n_16208)
);

XNOR2xp5_ASAP7_75t_L g16209 ( 
.A(n_16018),
.B(n_7705),
.Y(n_16209)
);

NAND2xp5_ASAP7_75t_SL g16210 ( 
.A(n_15992),
.B(n_7837),
.Y(n_16210)
);

AOI311xp33_ASAP7_75t_L g16211 ( 
.A1(n_16115),
.A2(n_6498),
.A3(n_6510),
.B(n_6482),
.C(n_6477),
.Y(n_16211)
);

INVx1_ASAP7_75t_L g16212 ( 
.A(n_16007),
.Y(n_16212)
);

AOI22xp33_ASAP7_75t_L g16213 ( 
.A1(n_16033),
.A2(n_7888),
.B1(n_7902),
.B2(n_7875),
.Y(n_16213)
);

NAND2xp5_ASAP7_75t_SL g16214 ( 
.A(n_16029),
.B(n_7837),
.Y(n_16214)
);

NAND2xp5_ASAP7_75t_L g16215 ( 
.A(n_16108),
.B(n_7962),
.Y(n_16215)
);

NAND2xp5_ASAP7_75t_L g16216 ( 
.A(n_15998),
.B(n_7962),
.Y(n_16216)
);

INVx1_ASAP7_75t_L g16217 ( 
.A(n_16087),
.Y(n_16217)
);

CKINVDCx5p33_ASAP7_75t_R g16218 ( 
.A(n_16017),
.Y(n_16218)
);

AOI322xp5_ASAP7_75t_L g16219 ( 
.A1(n_16042),
.A2(n_7875),
.A3(n_7909),
.B1(n_7902),
.B2(n_7936),
.C1(n_7916),
.C2(n_7888),
.Y(n_16219)
);

AOI21xp5_ASAP7_75t_L g16220 ( 
.A1(n_16078),
.A2(n_7261),
.B(n_7211),
.Y(n_16220)
);

AND2x2_ASAP7_75t_L g16221 ( 
.A(n_15977),
.B(n_6675),
.Y(n_16221)
);

XOR2x2_ASAP7_75t_L g16222 ( 
.A(n_16096),
.B(n_6141),
.Y(n_16222)
);

NAND2xp5_ASAP7_75t_L g16223 ( 
.A(n_16134),
.B(n_7940),
.Y(n_16223)
);

OR2x2_ASAP7_75t_L g16224 ( 
.A(n_15973),
.B(n_8046),
.Y(n_16224)
);

NOR4xp25_ASAP7_75t_SL g16225 ( 
.A(n_16015),
.B(n_6891),
.C(n_6932),
.D(n_6862),
.Y(n_16225)
);

INVx1_ASAP7_75t_L g16226 ( 
.A(n_15970),
.Y(n_16226)
);

INVx2_ASAP7_75t_L g16227 ( 
.A(n_16068),
.Y(n_16227)
);

INVx2_ASAP7_75t_L g16228 ( 
.A(n_16065),
.Y(n_16228)
);

NAND2xp5_ASAP7_75t_L g16229 ( 
.A(n_15965),
.B(n_7940),
.Y(n_16229)
);

NAND2xp5_ASAP7_75t_SL g16230 ( 
.A(n_16032),
.B(n_7837),
.Y(n_16230)
);

INVx2_ASAP7_75t_L g16231 ( 
.A(n_16066),
.Y(n_16231)
);

NAND2xp5_ASAP7_75t_L g16232 ( 
.A(n_16161),
.B(n_7940),
.Y(n_16232)
);

INVx1_ASAP7_75t_L g16233 ( 
.A(n_15986),
.Y(n_16233)
);

INVx1_ASAP7_75t_SL g16234 ( 
.A(n_16094),
.Y(n_16234)
);

NAND2xp5_ASAP7_75t_L g16235 ( 
.A(n_16131),
.B(n_7940),
.Y(n_16235)
);

NOR4xp25_ASAP7_75t_SL g16236 ( 
.A(n_16074),
.B(n_6891),
.C(n_6932),
.D(n_6862),
.Y(n_16236)
);

INVx1_ASAP7_75t_L g16237 ( 
.A(n_15962),
.Y(n_16237)
);

INVxp67_ASAP7_75t_L g16238 ( 
.A(n_15974),
.Y(n_16238)
);

NOR3xp33_ASAP7_75t_L g16239 ( 
.A(n_16012),
.B(n_7465),
.C(n_7485),
.Y(n_16239)
);

INVx2_ASAP7_75t_L g16240 ( 
.A(n_16088),
.Y(n_16240)
);

NAND2xp5_ASAP7_75t_L g16241 ( 
.A(n_16123),
.B(n_7909),
.Y(n_16241)
);

HB1xp67_ASAP7_75t_L g16242 ( 
.A(n_16030),
.Y(n_16242)
);

AOI221xp5_ASAP7_75t_L g16243 ( 
.A1(n_16136),
.A2(n_7888),
.B1(n_7936),
.B2(n_7916),
.C(n_7909),
.Y(n_16243)
);

INVx1_ASAP7_75t_SL g16244 ( 
.A(n_16146),
.Y(n_16244)
);

NAND2xp5_ASAP7_75t_L g16245 ( 
.A(n_16086),
.B(n_8010),
.Y(n_16245)
);

INVx2_ASAP7_75t_L g16246 ( 
.A(n_16075),
.Y(n_16246)
);

NOR2xp33_ASAP7_75t_L g16247 ( 
.A(n_16107),
.B(n_16069),
.Y(n_16247)
);

OAI21xp5_ASAP7_75t_L g16248 ( 
.A1(n_16055),
.A2(n_7473),
.B(n_7261),
.Y(n_16248)
);

NOR2xp33_ASAP7_75t_L g16249 ( 
.A(n_16092),
.B(n_7909),
.Y(n_16249)
);

INVx2_ASAP7_75t_L g16250 ( 
.A(n_16154),
.Y(n_16250)
);

NAND2xp5_ASAP7_75t_L g16251 ( 
.A(n_16130),
.B(n_7962),
.Y(n_16251)
);

OA22x2_ASAP7_75t_SL g16252 ( 
.A1(n_16112),
.A2(n_7039),
.B1(n_7081),
.B2(n_7023),
.Y(n_16252)
);

NAND2xp5_ASAP7_75t_SL g16253 ( 
.A(n_16120),
.B(n_7837),
.Y(n_16253)
);

INVx1_ASAP7_75t_L g16254 ( 
.A(n_15961),
.Y(n_16254)
);

AND2x2_ASAP7_75t_L g16255 ( 
.A(n_15987),
.B(n_7896),
.Y(n_16255)
);

NOR2xp33_ASAP7_75t_L g16256 ( 
.A(n_16127),
.B(n_7916),
.Y(n_16256)
);

AND2x2_ASAP7_75t_L g16257 ( 
.A(n_15990),
.B(n_7896),
.Y(n_16257)
);

INVx1_ASAP7_75t_SL g16258 ( 
.A(n_15972),
.Y(n_16258)
);

INVx2_ASAP7_75t_SL g16259 ( 
.A(n_16158),
.Y(n_16259)
);

INVxp67_ASAP7_75t_L g16260 ( 
.A(n_16031),
.Y(n_16260)
);

AND2x2_ASAP7_75t_L g16261 ( 
.A(n_16000),
.B(n_7900),
.Y(n_16261)
);

AND2x2_ASAP7_75t_L g16262 ( 
.A(n_15997),
.B(n_7900),
.Y(n_16262)
);

INVx1_ASAP7_75t_L g16263 ( 
.A(n_16162),
.Y(n_16263)
);

INVxp67_ASAP7_75t_L g16264 ( 
.A(n_16024),
.Y(n_16264)
);

AOI21xp33_ASAP7_75t_SL g16265 ( 
.A1(n_16103),
.A2(n_7465),
.B(n_7218),
.Y(n_16265)
);

OAI21xp5_ASAP7_75t_SL g16266 ( 
.A1(n_16091),
.A2(n_7908),
.B(n_7900),
.Y(n_16266)
);

NAND2xp5_ASAP7_75t_L g16267 ( 
.A(n_16016),
.B(n_7936),
.Y(n_16267)
);

INVx2_ASAP7_75t_L g16268 ( 
.A(n_16153),
.Y(n_16268)
);

INVx1_ASAP7_75t_L g16269 ( 
.A(n_16163),
.Y(n_16269)
);

AOI21xp5_ASAP7_75t_L g16270 ( 
.A1(n_16062),
.A2(n_7211),
.B(n_7205),
.Y(n_16270)
);

NOR3xp33_ASAP7_75t_SL g16271 ( 
.A(n_16095),
.B(n_6080),
.C(n_6002),
.Y(n_16271)
);

INVx2_ASAP7_75t_SL g16272 ( 
.A(n_15971),
.Y(n_16272)
);

BUFx8_ASAP7_75t_SL g16273 ( 
.A(n_16022),
.Y(n_16273)
);

CKINVDCx16_ASAP7_75t_R g16274 ( 
.A(n_16038),
.Y(n_16274)
);

INVx1_ASAP7_75t_L g16275 ( 
.A(n_16008),
.Y(n_16275)
);

INVx1_ASAP7_75t_L g16276 ( 
.A(n_16043),
.Y(n_16276)
);

NAND2xp5_ASAP7_75t_L g16277 ( 
.A(n_16034),
.B(n_8057),
.Y(n_16277)
);

INVxp67_ASAP7_75t_L g16278 ( 
.A(n_16061),
.Y(n_16278)
);

AOI221x1_ASAP7_75t_L g16279 ( 
.A1(n_16080),
.A2(n_7862),
.B1(n_8002),
.B2(n_7955),
.C(n_7906),
.Y(n_16279)
);

OAI22xp5_ASAP7_75t_L g16280 ( 
.A1(n_16126),
.A2(n_7862),
.B1(n_7955),
.B2(n_7906),
.Y(n_16280)
);

AND2x2_ASAP7_75t_L g16281 ( 
.A(n_16023),
.B(n_7900),
.Y(n_16281)
);

NOR2xp33_ASAP7_75t_L g16282 ( 
.A(n_15994),
.B(n_7916),
.Y(n_16282)
);

NAND2xp5_ASAP7_75t_L g16283 ( 
.A(n_16027),
.B(n_8010),
.Y(n_16283)
);

NAND2xp5_ASAP7_75t_L g16284 ( 
.A(n_16129),
.B(n_8010),
.Y(n_16284)
);

INVx2_ASAP7_75t_L g16285 ( 
.A(n_16153),
.Y(n_16285)
);

NAND2xp5_ASAP7_75t_L g16286 ( 
.A(n_16040),
.B(n_8010),
.Y(n_16286)
);

AND2x2_ASAP7_75t_L g16287 ( 
.A(n_16056),
.B(n_7908),
.Y(n_16287)
);

INVx1_ASAP7_75t_L g16288 ( 
.A(n_16046),
.Y(n_16288)
);

OR2x2_ASAP7_75t_L g16289 ( 
.A(n_16141),
.B(n_8046),
.Y(n_16289)
);

NAND2xp5_ASAP7_75t_L g16290 ( 
.A(n_16050),
.B(n_8102),
.Y(n_16290)
);

NOR2xp33_ASAP7_75t_R g16291 ( 
.A(n_16121),
.B(n_7023),
.Y(n_16291)
);

AOI211xp5_ASAP7_75t_L g16292 ( 
.A1(n_16124),
.A2(n_7957),
.B(n_7218),
.C(n_7211),
.Y(n_16292)
);

AND2x2_ASAP7_75t_L g16293 ( 
.A(n_16011),
.B(n_7908),
.Y(n_16293)
);

INVx1_ASAP7_75t_SL g16294 ( 
.A(n_16054),
.Y(n_16294)
);

NOR2xp33_ASAP7_75t_L g16295 ( 
.A(n_16132),
.B(n_7962),
.Y(n_16295)
);

INVx1_ASAP7_75t_SL g16296 ( 
.A(n_15964),
.Y(n_16296)
);

INVx1_ASAP7_75t_L g16297 ( 
.A(n_15985),
.Y(n_16297)
);

INVx2_ASAP7_75t_L g16298 ( 
.A(n_16138),
.Y(n_16298)
);

NOR2xp67_ASAP7_75t_L g16299 ( 
.A(n_16139),
.B(n_7023),
.Y(n_16299)
);

OAI21xp5_ASAP7_75t_L g16300 ( 
.A1(n_16001),
.A2(n_7473),
.B(n_7218),
.Y(n_16300)
);

AOI22xp5_ASAP7_75t_L g16301 ( 
.A1(n_16114),
.A2(n_7911),
.B1(n_7908),
.B2(n_7862),
.Y(n_16301)
);

INVx2_ASAP7_75t_L g16302 ( 
.A(n_16097),
.Y(n_16302)
);

INVx1_ASAP7_75t_L g16303 ( 
.A(n_16152),
.Y(n_16303)
);

INVx1_ASAP7_75t_L g16304 ( 
.A(n_16026),
.Y(n_16304)
);

INVx1_ASAP7_75t_L g16305 ( 
.A(n_16049),
.Y(n_16305)
);

NAND2xp5_ASAP7_75t_L g16306 ( 
.A(n_16089),
.B(n_8038),
.Y(n_16306)
);

INVx1_ASAP7_75t_L g16307 ( 
.A(n_15989),
.Y(n_16307)
);

INVx1_ASAP7_75t_L g16308 ( 
.A(n_16014),
.Y(n_16308)
);

INVxp67_ASAP7_75t_L g16309 ( 
.A(n_16118),
.Y(n_16309)
);

INVx1_ASAP7_75t_L g16310 ( 
.A(n_15988),
.Y(n_16310)
);

INVx1_ASAP7_75t_SL g16311 ( 
.A(n_16052),
.Y(n_16311)
);

INVxp67_ASAP7_75t_L g16312 ( 
.A(n_16150),
.Y(n_16312)
);

AND2x2_ASAP7_75t_L g16313 ( 
.A(n_16028),
.B(n_7911),
.Y(n_16313)
);

INVxp67_ASAP7_75t_L g16314 ( 
.A(n_16048),
.Y(n_16314)
);

NOR2xp33_ASAP7_75t_L g16315 ( 
.A(n_16064),
.B(n_7998),
.Y(n_16315)
);

NOR4xp25_ASAP7_75t_SL g16316 ( 
.A(n_15993),
.B(n_6932),
.C(n_6951),
.D(n_6891),
.Y(n_16316)
);

INVx1_ASAP7_75t_L g16317 ( 
.A(n_16051),
.Y(n_16317)
);

INVx1_ASAP7_75t_L g16318 ( 
.A(n_16010),
.Y(n_16318)
);

CKINVDCx5p33_ASAP7_75t_R g16319 ( 
.A(n_16148),
.Y(n_16319)
);

AND2x2_ASAP7_75t_L g16320 ( 
.A(n_16044),
.B(n_7911),
.Y(n_16320)
);

INVx2_ASAP7_75t_L g16321 ( 
.A(n_16100),
.Y(n_16321)
);

NAND2xp5_ASAP7_75t_L g16322 ( 
.A(n_16116),
.B(n_16039),
.Y(n_16322)
);

AND2x2_ASAP7_75t_L g16323 ( 
.A(n_16085),
.B(n_16128),
.Y(n_16323)
);

NAND2xp5_ASAP7_75t_L g16324 ( 
.A(n_16098),
.B(n_7998),
.Y(n_16324)
);

AOI31xp33_ASAP7_75t_L g16325 ( 
.A1(n_16147),
.A2(n_7138),
.A3(n_7108),
.B(n_7066),
.Y(n_16325)
);

NOR2xp33_ASAP7_75t_R g16326 ( 
.A(n_16071),
.B(n_7039),
.Y(n_16326)
);

NAND2xp5_ASAP7_75t_L g16327 ( 
.A(n_16090),
.B(n_7998),
.Y(n_16327)
);

INVx2_ASAP7_75t_SL g16328 ( 
.A(n_16037),
.Y(n_16328)
);

NOR2xp33_ASAP7_75t_L g16329 ( 
.A(n_16144),
.B(n_7998),
.Y(n_16329)
);

OR2x2_ASAP7_75t_L g16330 ( 
.A(n_16101),
.B(n_8046),
.Y(n_16330)
);

NAND2xp5_ASAP7_75t_L g16331 ( 
.A(n_16099),
.B(n_8167),
.Y(n_16331)
);

NAND2xp5_ASAP7_75t_L g16332 ( 
.A(n_16079),
.B(n_8167),
.Y(n_16332)
);

AOI21xp33_ASAP7_75t_L g16333 ( 
.A1(n_16081),
.A2(n_8057),
.B(n_8038),
.Y(n_16333)
);

NOR2xp33_ASAP7_75t_SL g16334 ( 
.A(n_15984),
.B(n_6002),
.Y(n_16334)
);

INVx1_ASAP7_75t_L g16335 ( 
.A(n_16067),
.Y(n_16335)
);

INVxp67_ASAP7_75t_L g16336 ( 
.A(n_16102),
.Y(n_16336)
);

INVx2_ASAP7_75t_L g16337 ( 
.A(n_16063),
.Y(n_16337)
);

INVxp33_ASAP7_75t_L g16338 ( 
.A(n_16105),
.Y(n_16338)
);

NOR3xp33_ASAP7_75t_L g16339 ( 
.A(n_16274),
.B(n_16104),
.C(n_16082),
.Y(n_16339)
);

NAND2xp5_ASAP7_75t_SL g16340 ( 
.A(n_16234),
.B(n_16084),
.Y(n_16340)
);

O2A1O1Ixp5_ASAP7_75t_L g16341 ( 
.A1(n_16187),
.A2(n_16109),
.B(n_16113),
.C(n_16111),
.Y(n_16341)
);

NOR2x1_ASAP7_75t_L g16342 ( 
.A(n_16183),
.B(n_16041),
.Y(n_16342)
);

AOI211xp5_ASAP7_75t_L g16343 ( 
.A1(n_16172),
.A2(n_16145),
.B(n_16135),
.C(n_16133),
.Y(n_16343)
);

AOI21xp5_ASAP7_75t_L g16344 ( 
.A1(n_16169),
.A2(n_16149),
.B(n_16110),
.Y(n_16344)
);

NOR3xp33_ASAP7_75t_L g16345 ( 
.A(n_16170),
.B(n_16143),
.C(n_16122),
.Y(n_16345)
);

AOI22xp5_ASAP7_75t_L g16346 ( 
.A1(n_16174),
.A2(n_16057),
.B1(n_16142),
.B2(n_16117),
.Y(n_16346)
);

INVx1_ASAP7_75t_L g16347 ( 
.A(n_16218),
.Y(n_16347)
);

INVx2_ASAP7_75t_SL g16348 ( 
.A(n_16246),
.Y(n_16348)
);

NAND3xp33_ASAP7_75t_L g16349 ( 
.A(n_16180),
.B(n_16151),
.C(n_16106),
.Y(n_16349)
);

HB1xp67_ASAP7_75t_L g16350 ( 
.A(n_16273),
.Y(n_16350)
);

AOI21xp5_ASAP7_75t_L g16351 ( 
.A1(n_16192),
.A2(n_16060),
.B(n_16125),
.Y(n_16351)
);

NAND3xp33_ASAP7_75t_L g16352 ( 
.A(n_16189),
.B(n_16159),
.C(n_15983),
.Y(n_16352)
);

NOR2xp33_ASAP7_75t_L g16353 ( 
.A(n_16244),
.B(n_16025),
.Y(n_16353)
);

OAI211xp5_ASAP7_75t_SL g16354 ( 
.A1(n_16312),
.A2(n_16058),
.B(n_16077),
.C(n_16119),
.Y(n_16354)
);

NOR2xp33_ASAP7_75t_L g16355 ( 
.A(n_16309),
.B(n_16176),
.Y(n_16355)
);

NAND2xp5_ASAP7_75t_L g16356 ( 
.A(n_16299),
.B(n_8038),
.Y(n_16356)
);

NOR2xp67_ASAP7_75t_L g16357 ( 
.A(n_16240),
.B(n_7039),
.Y(n_16357)
);

NAND2xp5_ASAP7_75t_L g16358 ( 
.A(n_16228),
.B(n_8038),
.Y(n_16358)
);

AOI211xp5_ASAP7_75t_L g16359 ( 
.A1(n_16193),
.A2(n_8170),
.B(n_8002),
.C(n_7906),
.Y(n_16359)
);

AOI22xp5_ASAP7_75t_L g16360 ( 
.A1(n_16319),
.A2(n_7862),
.B1(n_7955),
.B2(n_7906),
.Y(n_16360)
);

INVx1_ASAP7_75t_SL g16361 ( 
.A(n_16231),
.Y(n_16361)
);

INVx2_ASAP7_75t_L g16362 ( 
.A(n_16252),
.Y(n_16362)
);

OAI22xp33_ASAP7_75t_L g16363 ( 
.A1(n_16268),
.A2(n_7906),
.B1(n_7955),
.B2(n_7862),
.Y(n_16363)
);

INVx1_ASAP7_75t_L g16364 ( 
.A(n_16167),
.Y(n_16364)
);

NOR2xp67_ASAP7_75t_L g16365 ( 
.A(n_16242),
.B(n_7039),
.Y(n_16365)
);

AOI22xp33_ASAP7_75t_SL g16366 ( 
.A1(n_16182),
.A2(n_6080),
.B1(n_7081),
.B2(n_7906),
.Y(n_16366)
);

INVx1_ASAP7_75t_L g16367 ( 
.A(n_16167),
.Y(n_16367)
);

AOI21xp5_ASAP7_75t_L g16368 ( 
.A1(n_16194),
.A2(n_16196),
.B(n_16285),
.Y(n_16368)
);

OR2x2_ASAP7_75t_L g16369 ( 
.A(n_16227),
.B(n_16190),
.Y(n_16369)
);

NAND2xp5_ASAP7_75t_SL g16370 ( 
.A(n_16294),
.B(n_16197),
.Y(n_16370)
);

OAI211xp5_ASAP7_75t_SL g16371 ( 
.A1(n_16260),
.A2(n_8057),
.B(n_8138),
.C(n_8102),
.Y(n_16371)
);

INVx1_ASAP7_75t_L g16372 ( 
.A(n_16168),
.Y(n_16372)
);

AND2x2_ASAP7_75t_L g16373 ( 
.A(n_16221),
.B(n_7911),
.Y(n_16373)
);

NAND2xp5_ASAP7_75t_L g16374 ( 
.A(n_16296),
.B(n_8057),
.Y(n_16374)
);

INVx1_ASAP7_75t_L g16375 ( 
.A(n_16201),
.Y(n_16375)
);

NOR3xp33_ASAP7_75t_L g16376 ( 
.A(n_16212),
.B(n_16278),
.C(n_16206),
.Y(n_16376)
);

AOI211x1_ASAP7_75t_L g16377 ( 
.A1(n_16179),
.A2(n_6482),
.B(n_6498),
.C(n_6477),
.Y(n_16377)
);

AND2x2_ASAP7_75t_L g16378 ( 
.A(n_16203),
.B(n_7911),
.Y(n_16378)
);

AND2x2_ASAP7_75t_L g16379 ( 
.A(n_16185),
.B(n_16181),
.Y(n_16379)
);

NAND2xp5_ASAP7_75t_L g16380 ( 
.A(n_16259),
.B(n_8102),
.Y(n_16380)
);

AOI21xp5_ASAP7_75t_L g16381 ( 
.A1(n_16214),
.A2(n_8138),
.B(n_8102),
.Y(n_16381)
);

NOR3x1_ASAP7_75t_L g16382 ( 
.A(n_16328),
.B(n_7608),
.C(n_7606),
.Y(n_16382)
);

AND2x2_ASAP7_75t_L g16383 ( 
.A(n_16262),
.B(n_6131),
.Y(n_16383)
);

AOI221xp5_ASAP7_75t_L g16384 ( 
.A1(n_16303),
.A2(n_8165),
.B1(n_8167),
.B2(n_8145),
.C(n_8138),
.Y(n_16384)
);

AOI211xp5_ASAP7_75t_L g16385 ( 
.A1(n_16247),
.A2(n_8170),
.B(n_7955),
.C(n_8002),
.Y(n_16385)
);

AOI21xp5_ASAP7_75t_L g16386 ( 
.A1(n_16322),
.A2(n_8165),
.B(n_8145),
.Y(n_16386)
);

OA22x2_ASAP7_75t_L g16387 ( 
.A1(n_16191),
.A2(n_8051),
.B1(n_8183),
.B2(n_8023),
.Y(n_16387)
);

AND2x2_ASAP7_75t_L g16388 ( 
.A(n_16255),
.B(n_6131),
.Y(n_16388)
);

AOI211x1_ASAP7_75t_L g16389 ( 
.A1(n_16230),
.A2(n_6498),
.B(n_6510),
.C(n_6482),
.Y(n_16389)
);

AOI21xp5_ASAP7_75t_L g16390 ( 
.A1(n_16175),
.A2(n_8165),
.B(n_8145),
.Y(n_16390)
);

BUFx2_ASAP7_75t_L g16391 ( 
.A(n_16291),
.Y(n_16391)
);

NOR2x1p5_ASAP7_75t_SL g16392 ( 
.A(n_16178),
.B(n_6285),
.Y(n_16392)
);

NAND2xp5_ASAP7_75t_SL g16393 ( 
.A(n_16204),
.B(n_7906),
.Y(n_16393)
);

OAI211xp5_ASAP7_75t_SL g16394 ( 
.A1(n_16238),
.A2(n_8145),
.B(n_8167),
.C(n_8165),
.Y(n_16394)
);

AOI21xp5_ASAP7_75t_L g16395 ( 
.A1(n_16208),
.A2(n_8188),
.B(n_8172),
.Y(n_16395)
);

O2A1O1Ixp33_ASAP7_75t_L g16396 ( 
.A1(n_16302),
.A2(n_16297),
.B(n_16226),
.C(n_16308),
.Y(n_16396)
);

AOI211x1_ASAP7_75t_L g16397 ( 
.A1(n_16210),
.A2(n_6511),
.B(n_6512),
.C(n_6510),
.Y(n_16397)
);

OAI21xp33_ASAP7_75t_L g16398 ( 
.A1(n_16217),
.A2(n_16338),
.B(n_16311),
.Y(n_16398)
);

CKINVDCx16_ASAP7_75t_R g16399 ( 
.A(n_16272),
.Y(n_16399)
);

OAI21xp33_ASAP7_75t_L g16400 ( 
.A1(n_16222),
.A2(n_8183),
.B(n_8051),
.Y(n_16400)
);

OAI21xp5_ASAP7_75t_L g16401 ( 
.A1(n_16256),
.A2(n_7487),
.B(n_7485),
.Y(n_16401)
);

NAND2xp5_ASAP7_75t_SL g16402 ( 
.A(n_16258),
.B(n_7955),
.Y(n_16402)
);

AOI21xp5_ASAP7_75t_L g16403 ( 
.A1(n_16188),
.A2(n_8188),
.B(n_8172),
.Y(n_16403)
);

NOR3xp33_ASAP7_75t_L g16404 ( 
.A(n_16264),
.B(n_7487),
.C(n_7485),
.Y(n_16404)
);

INVx1_ASAP7_75t_L g16405 ( 
.A(n_16323),
.Y(n_16405)
);

INVx2_ASAP7_75t_L g16406 ( 
.A(n_16321),
.Y(n_16406)
);

OAI222xp33_ASAP7_75t_L g16407 ( 
.A1(n_16215),
.A2(n_8172),
.B1(n_8193),
.B2(n_8208),
.C1(n_8205),
.C2(n_8188),
.Y(n_16407)
);

OAI21xp33_ASAP7_75t_L g16408 ( 
.A1(n_16271),
.A2(n_8183),
.B(n_8051),
.Y(n_16408)
);

OAI22xp33_ASAP7_75t_L g16409 ( 
.A1(n_16334),
.A2(n_8002),
.B1(n_8125),
.B2(n_7955),
.Y(n_16409)
);

AOI21xp5_ASAP7_75t_L g16410 ( 
.A1(n_16198),
.A2(n_8188),
.B(n_8172),
.Y(n_16410)
);

NOR2xp33_ASAP7_75t_L g16411 ( 
.A(n_16336),
.B(n_8193),
.Y(n_16411)
);

AOI21xp5_ASAP7_75t_L g16412 ( 
.A1(n_16310),
.A2(n_8205),
.B(n_8193),
.Y(n_16412)
);

NOR2xp33_ASAP7_75t_L g16413 ( 
.A(n_16298),
.B(n_16241),
.Y(n_16413)
);

NAND2xp5_ASAP7_75t_L g16414 ( 
.A(n_16213),
.B(n_8193),
.Y(n_16414)
);

NOR2xp33_ASAP7_75t_L g16415 ( 
.A(n_16237),
.B(n_8205),
.Y(n_16415)
);

AOI31xp33_ASAP7_75t_L g16416 ( 
.A1(n_16314),
.A2(n_7138),
.A3(n_7927),
.B(n_7925),
.Y(n_16416)
);

OA22x2_ASAP7_75t_L g16417 ( 
.A1(n_16195),
.A2(n_8183),
.B1(n_7520),
.B2(n_7894),
.Y(n_16417)
);

INVx1_ASAP7_75t_L g16418 ( 
.A(n_16223),
.Y(n_16418)
);

AOI22xp5_ASAP7_75t_L g16419 ( 
.A1(n_16250),
.A2(n_7955),
.B1(n_8125),
.B2(n_8002),
.Y(n_16419)
);

HB1xp67_ASAP7_75t_L g16420 ( 
.A(n_16254),
.Y(n_16420)
);

NAND2xp5_ASAP7_75t_L g16421 ( 
.A(n_16249),
.B(n_8205),
.Y(n_16421)
);

AO22x2_ASAP7_75t_L g16422 ( 
.A1(n_16263),
.A2(n_8212),
.B1(n_8220),
.B2(n_8208),
.Y(n_16422)
);

INVx1_ASAP7_75t_L g16423 ( 
.A(n_16216),
.Y(n_16423)
);

INVx1_ASAP7_75t_L g16424 ( 
.A(n_16235),
.Y(n_16424)
);

OAI211xp5_ASAP7_75t_L g16425 ( 
.A1(n_16269),
.A2(n_6066),
.B(n_8125),
.C(n_8002),
.Y(n_16425)
);

INVx2_ASAP7_75t_L g16426 ( 
.A(n_16199),
.Y(n_16426)
);

NOR2x1_ASAP7_75t_L g16427 ( 
.A(n_16276),
.B(n_7925),
.Y(n_16427)
);

OA22x2_ASAP7_75t_L g16428 ( 
.A1(n_16301),
.A2(n_7520),
.B1(n_7894),
.B2(n_7608),
.Y(n_16428)
);

AOI21xp5_ASAP7_75t_L g16429 ( 
.A1(n_16288),
.A2(n_8212),
.B(n_8208),
.Y(n_16429)
);

OA22x2_ASAP7_75t_L g16430 ( 
.A1(n_16304),
.A2(n_7608),
.B1(n_7606),
.B2(n_7572),
.Y(n_16430)
);

INVx1_ASAP7_75t_L g16431 ( 
.A(n_16305),
.Y(n_16431)
);

NOR2xp67_ASAP7_75t_L g16432 ( 
.A(n_16233),
.B(n_7081),
.Y(n_16432)
);

AOI211xp5_ASAP7_75t_L g16433 ( 
.A1(n_16318),
.A2(n_8125),
.B(n_8170),
.C(n_8002),
.Y(n_16433)
);

NAND2xp5_ASAP7_75t_SL g16434 ( 
.A(n_16317),
.B(n_8002),
.Y(n_16434)
);

AOI211xp5_ASAP7_75t_L g16435 ( 
.A1(n_16275),
.A2(n_8170),
.B(n_8125),
.C(n_7213),
.Y(n_16435)
);

OA22x2_ASAP7_75t_L g16436 ( 
.A1(n_16307),
.A2(n_7606),
.B1(n_7572),
.B2(n_7571),
.Y(n_16436)
);

OAI21xp33_ASAP7_75t_SL g16437 ( 
.A1(n_16253),
.A2(n_7623),
.B(n_7622),
.Y(n_16437)
);

OA22x2_ASAP7_75t_L g16438 ( 
.A1(n_16335),
.A2(n_7572),
.B1(n_7571),
.B2(n_7925),
.Y(n_16438)
);

AOI21xp5_ASAP7_75t_L g16439 ( 
.A1(n_16337),
.A2(n_8212),
.B(n_8208),
.Y(n_16439)
);

HB1xp67_ASAP7_75t_L g16440 ( 
.A(n_16284),
.Y(n_16440)
);

OAI21xp33_ASAP7_75t_SL g16441 ( 
.A1(n_16261),
.A2(n_7623),
.B(n_7622),
.Y(n_16441)
);

AOI211xp5_ASAP7_75t_L g16442 ( 
.A1(n_16326),
.A2(n_8170),
.B(n_8125),
.C(n_7213),
.Y(n_16442)
);

NOR2xp33_ASAP7_75t_L g16443 ( 
.A(n_16295),
.B(n_8212),
.Y(n_16443)
);

CKINVDCx5p33_ASAP7_75t_R g16444 ( 
.A(n_16177),
.Y(n_16444)
);

AOI22xp5_ASAP7_75t_L g16445 ( 
.A1(n_16329),
.A2(n_16173),
.B1(n_16282),
.B2(n_16209),
.Y(n_16445)
);

INVx1_ASAP7_75t_L g16446 ( 
.A(n_16277),
.Y(n_16446)
);

INVx1_ASAP7_75t_L g16447 ( 
.A(n_16286),
.Y(n_16447)
);

INVx1_ASAP7_75t_L g16448 ( 
.A(n_16290),
.Y(n_16448)
);

NAND4xp25_ASAP7_75t_L g16449 ( 
.A(n_16245),
.B(n_16267),
.C(n_16306),
.D(n_16211),
.Y(n_16449)
);

INVx1_ASAP7_75t_L g16450 ( 
.A(n_16251),
.Y(n_16450)
);

OA22x2_ASAP7_75t_L g16451 ( 
.A1(n_16327),
.A2(n_7571),
.B1(n_7927),
.B2(n_7925),
.Y(n_16451)
);

NOR3xp33_ASAP7_75t_L g16452 ( 
.A(n_16330),
.B(n_7487),
.C(n_7474),
.Y(n_16452)
);

AOI31xp33_ASAP7_75t_L g16453 ( 
.A1(n_16293),
.A2(n_16257),
.A3(n_16166),
.B(n_16283),
.Y(n_16453)
);

NAND2xp5_ASAP7_75t_L g16454 ( 
.A(n_16315),
.B(n_8220),
.Y(n_16454)
);

AOI22x1_ASAP7_75t_L g16455 ( 
.A1(n_16313),
.A2(n_6980),
.B1(n_6142),
.B2(n_6496),
.Y(n_16455)
);

OA22x2_ASAP7_75t_L g16456 ( 
.A1(n_16266),
.A2(n_7927),
.B1(n_7925),
.B2(n_7177),
.Y(n_16456)
);

AOI22xp5_ASAP7_75t_L g16457 ( 
.A1(n_16289),
.A2(n_8125),
.B1(n_8170),
.B2(n_8220),
.Y(n_16457)
);

NAND2xp5_ASAP7_75t_L g16458 ( 
.A(n_16316),
.B(n_8248),
.Y(n_16458)
);

NOR2xp33_ASAP7_75t_L g16459 ( 
.A(n_16332),
.B(n_8248),
.Y(n_16459)
);

AOI211x1_ASAP7_75t_L g16460 ( 
.A1(n_16331),
.A2(n_6512),
.B(n_6521),
.C(n_6511),
.Y(n_16460)
);

OAI22xp5_ASAP7_75t_L g16461 ( 
.A1(n_16202),
.A2(n_16224),
.B1(n_16220),
.B2(n_16287),
.Y(n_16461)
);

AND2x2_ASAP7_75t_L g16462 ( 
.A(n_16281),
.B(n_6131),
.Y(n_16462)
);

INVx1_ASAP7_75t_SL g16463 ( 
.A(n_16229),
.Y(n_16463)
);

AOI21xp5_ASAP7_75t_L g16464 ( 
.A1(n_16324),
.A2(n_8248),
.B(n_7213),
.Y(n_16464)
);

INVx2_ASAP7_75t_SL g16465 ( 
.A(n_16320),
.Y(n_16465)
);

AOI211xp5_ASAP7_75t_L g16466 ( 
.A1(n_16200),
.A2(n_8125),
.B(n_8170),
.C(n_7205),
.Y(n_16466)
);

AOI221xp5_ASAP7_75t_L g16467 ( 
.A1(n_16232),
.A2(n_16333),
.B1(n_16325),
.B2(n_16171),
.C(n_16207),
.Y(n_16467)
);

NAND3xp33_ASAP7_75t_L g16468 ( 
.A(n_16279),
.B(n_8248),
.C(n_8170),
.Y(n_16468)
);

INVx2_ASAP7_75t_L g16469 ( 
.A(n_16280),
.Y(n_16469)
);

AOI21xp5_ASAP7_75t_L g16470 ( 
.A1(n_16225),
.A2(n_7177),
.B(n_7175),
.Y(n_16470)
);

NOR2x1_ASAP7_75t_L g16471 ( 
.A(n_16184),
.B(n_7927),
.Y(n_16471)
);

AOI221x1_ASAP7_75t_SL g16472 ( 
.A1(n_16236),
.A2(n_7705),
.B1(n_7709),
.B2(n_7927),
.C(n_6522),
.Y(n_16472)
);

NAND2xp5_ASAP7_75t_L g16473 ( 
.A(n_16186),
.B(n_7474),
.Y(n_16473)
);

OAI211xp5_ASAP7_75t_SL g16474 ( 
.A1(n_16219),
.A2(n_16248),
.B(n_16300),
.C(n_16239),
.Y(n_16474)
);

NAND2xp5_ASAP7_75t_L g16475 ( 
.A(n_16205),
.B(n_7474),
.Y(n_16475)
);

AND2x2_ASAP7_75t_L g16476 ( 
.A(n_16265),
.B(n_6155),
.Y(n_16476)
);

OAI211xp5_ASAP7_75t_SL g16477 ( 
.A1(n_16243),
.A2(n_6648),
.B(n_6669),
.C(n_6663),
.Y(n_16477)
);

INVx1_ASAP7_75t_L g16478 ( 
.A(n_16270),
.Y(n_16478)
);

NAND2xp5_ASAP7_75t_L g16479 ( 
.A(n_16292),
.B(n_8046),
.Y(n_16479)
);

AND2x2_ASAP7_75t_L g16480 ( 
.A(n_16170),
.B(n_6155),
.Y(n_16480)
);

AOI211xp5_ASAP7_75t_L g16481 ( 
.A1(n_16172),
.A2(n_7175),
.B(n_7296),
.C(n_7968),
.Y(n_16481)
);

AO22x1_ASAP7_75t_L g16482 ( 
.A1(n_16180),
.A2(n_7271),
.B1(n_6522),
.B2(n_6438),
.Y(n_16482)
);

NOR3xp33_ASAP7_75t_L g16483 ( 
.A(n_16274),
.B(n_7296),
.C(n_7305),
.Y(n_16483)
);

NAND2xp5_ASAP7_75t_L g16484 ( 
.A(n_16274),
.B(n_8046),
.Y(n_16484)
);

NAND2xp5_ASAP7_75t_L g16485 ( 
.A(n_16350),
.B(n_8299),
.Y(n_16485)
);

A2O1A1Ixp33_ASAP7_75t_SL g16486 ( 
.A1(n_16376),
.A2(n_6536),
.B(n_6544),
.C(n_6532),
.Y(n_16486)
);

XOR2x2_ASAP7_75t_L g16487 ( 
.A(n_16370),
.B(n_6141),
.Y(n_16487)
);

OAI21xp33_ASAP7_75t_L g16488 ( 
.A1(n_16361),
.A2(n_16348),
.B(n_16398),
.Y(n_16488)
);

AOI221xp5_ASAP7_75t_L g16489 ( 
.A1(n_16405),
.A2(n_6521),
.B1(n_6524),
.B2(n_6512),
.C(n_6511),
.Y(n_16489)
);

OAI32xp33_ASAP7_75t_L g16490 ( 
.A1(n_16369),
.A2(n_6668),
.A3(n_6744),
.B1(n_6826),
.B2(n_6764),
.Y(n_16490)
);

AND2x4_ASAP7_75t_L g16491 ( 
.A(n_16365),
.B(n_8008),
.Y(n_16491)
);

AOI31xp33_ASAP7_75t_L g16492 ( 
.A1(n_16347),
.A2(n_6668),
.A3(n_6764),
.B(n_6744),
.Y(n_16492)
);

NAND2xp5_ASAP7_75t_L g16493 ( 
.A(n_16399),
.B(n_8299),
.Y(n_16493)
);

XNOR2x1_ASAP7_75t_L g16494 ( 
.A(n_16342),
.B(n_16444),
.Y(n_16494)
);

NAND4xp25_ASAP7_75t_L g16495 ( 
.A(n_16396),
.B(n_7709),
.C(n_7705),
.D(n_6709),
.Y(n_16495)
);

NAND2xp5_ASAP7_75t_SL g16496 ( 
.A(n_16375),
.B(n_7754),
.Y(n_16496)
);

A2O1A1Ixp33_ASAP7_75t_L g16497 ( 
.A1(n_16368),
.A2(n_7296),
.B(n_7311),
.C(n_7305),
.Y(n_16497)
);

INVx1_ASAP7_75t_L g16498 ( 
.A(n_16420),
.Y(n_16498)
);

AOI21xp5_ASAP7_75t_L g16499 ( 
.A1(n_16340),
.A2(n_6669),
.B(n_6663),
.Y(n_16499)
);

OAI22xp33_ASAP7_75t_SL g16500 ( 
.A1(n_16364),
.A2(n_6600),
.B1(n_6762),
.B2(n_6248),
.Y(n_16500)
);

OAI211xp5_ASAP7_75t_L g16501 ( 
.A1(n_16343),
.A2(n_6066),
.B(n_6983),
.C(n_6935),
.Y(n_16501)
);

CKINVDCx5p33_ASAP7_75t_R g16502 ( 
.A(n_16355),
.Y(n_16502)
);

AO21x1_ASAP7_75t_L g16503 ( 
.A1(n_16367),
.A2(n_6990),
.B(n_6927),
.Y(n_16503)
);

AOI221xp5_ASAP7_75t_L g16504 ( 
.A1(n_16453),
.A2(n_6529),
.B1(n_6548),
.B2(n_6524),
.C(n_6521),
.Y(n_16504)
);

OAI211xp5_ASAP7_75t_L g16505 ( 
.A1(n_16344),
.A2(n_6066),
.B(n_6983),
.C(n_6935),
.Y(n_16505)
);

AOI221xp5_ASAP7_75t_L g16506 ( 
.A1(n_16339),
.A2(n_6548),
.B1(n_6551),
.B2(n_6529),
.C(n_6524),
.Y(n_16506)
);

A2O1A1Ixp33_ASAP7_75t_L g16507 ( 
.A1(n_16353),
.A2(n_7305),
.B(n_7311),
.C(n_7968),
.Y(n_16507)
);

CKINVDCx5p33_ASAP7_75t_R g16508 ( 
.A(n_16391),
.Y(n_16508)
);

AOI22xp33_ASAP7_75t_SL g16509 ( 
.A1(n_16465),
.A2(n_7081),
.B1(n_5077),
.B2(n_7709),
.Y(n_16509)
);

NAND3xp33_ASAP7_75t_SL g16510 ( 
.A(n_16463),
.B(n_6141),
.C(n_6255),
.Y(n_16510)
);

AOI21xp5_ASAP7_75t_L g16511 ( 
.A1(n_16351),
.A2(n_7419),
.B(n_6066),
.Y(n_16511)
);

OAI221xp5_ASAP7_75t_L g16512 ( 
.A1(n_16357),
.A2(n_6548),
.B1(n_6553),
.B2(n_6551),
.C(n_6529),
.Y(n_16512)
);

INVx1_ASAP7_75t_L g16513 ( 
.A(n_16379),
.Y(n_16513)
);

NAND4xp75_ASAP7_75t_L g16514 ( 
.A(n_16413),
.B(n_5979),
.C(n_6022),
.D(n_5977),
.Y(n_16514)
);

AOI21xp33_ASAP7_75t_L g16515 ( 
.A1(n_16406),
.A2(n_8299),
.B(n_8202),
.Y(n_16515)
);

AOI21xp33_ASAP7_75t_L g16516 ( 
.A1(n_16431),
.A2(n_8299),
.B(n_8202),
.Y(n_16516)
);

A2O1A1Ixp33_ASAP7_75t_SL g16517 ( 
.A1(n_16362),
.A2(n_6544),
.B(n_6562),
.C(n_6536),
.Y(n_16517)
);

NAND2xp5_ASAP7_75t_L g16518 ( 
.A(n_16432),
.B(n_8299),
.Y(n_16518)
);

AOI221xp5_ASAP7_75t_L g16519 ( 
.A1(n_16461),
.A2(n_6571),
.B1(n_6573),
.B2(n_6553),
.C(n_6551),
.Y(n_16519)
);

NAND2xp5_ASAP7_75t_L g16520 ( 
.A(n_16440),
.B(n_8154),
.Y(n_16520)
);

AOI31xp33_ASAP7_75t_L g16521 ( 
.A1(n_16372),
.A2(n_6668),
.A3(n_6764),
.B(n_6744),
.Y(n_16521)
);

NOR4xp25_ASAP7_75t_L g16522 ( 
.A(n_16424),
.B(n_6571),
.C(n_6573),
.D(n_6553),
.Y(n_16522)
);

INVx3_ASAP7_75t_L g16523 ( 
.A(n_16426),
.Y(n_16523)
);

INVx2_ASAP7_75t_SL g16524 ( 
.A(n_16427),
.Y(n_16524)
);

INVxp67_ASAP7_75t_L g16525 ( 
.A(n_16450),
.Y(n_16525)
);

INVx1_ASAP7_75t_L g16526 ( 
.A(n_16374),
.Y(n_16526)
);

AOI21xp5_ASAP7_75t_L g16527 ( 
.A1(n_16349),
.A2(n_7419),
.B(n_6066),
.Y(n_16527)
);

INVx1_ASAP7_75t_L g16528 ( 
.A(n_16480),
.Y(n_16528)
);

AOI21xp33_ASAP7_75t_L g16529 ( 
.A1(n_16418),
.A2(n_8215),
.B(n_8202),
.Y(n_16529)
);

O2A1O1Ixp33_ASAP7_75t_SL g16530 ( 
.A1(n_16393),
.A2(n_6848),
.B(n_6857),
.C(n_6826),
.Y(n_16530)
);

OAI322xp33_ASAP7_75t_SL g16531 ( 
.A1(n_16484),
.A2(n_6573),
.A3(n_6588),
.B1(n_6587),
.B2(n_6603),
.C1(n_6593),
.C2(n_6571),
.Y(n_16531)
);

AOI22xp5_ASAP7_75t_L g16532 ( 
.A1(n_16345),
.A2(n_7271),
.B1(n_8182),
.B2(n_7754),
.Y(n_16532)
);

AOI221x1_ASAP7_75t_L g16533 ( 
.A1(n_16478),
.A2(n_6438),
.B1(n_6522),
.B2(n_6588),
.C(n_6587),
.Y(n_16533)
);

AOI21xp5_ASAP7_75t_L g16534 ( 
.A1(n_16449),
.A2(n_7419),
.B(n_6066),
.Y(n_16534)
);

CKINVDCx20_ASAP7_75t_R g16535 ( 
.A(n_16346),
.Y(n_16535)
);

OAI21xp5_ASAP7_75t_L g16536 ( 
.A1(n_16341),
.A2(n_7467),
.B(n_7423),
.Y(n_16536)
);

OAI22xp5_ASAP7_75t_L g16537 ( 
.A1(n_16352),
.A2(n_6826),
.B1(n_6857),
.B2(n_6848),
.Y(n_16537)
);

INVx1_ASAP7_75t_L g16538 ( 
.A(n_16380),
.Y(n_16538)
);

INVx2_ASAP7_75t_L g16539 ( 
.A(n_16446),
.Y(n_16539)
);

OAI21xp5_ASAP7_75t_L g16540 ( 
.A1(n_16445),
.A2(n_7467),
.B(n_7423),
.Y(n_16540)
);

AOI221xp5_ASAP7_75t_L g16541 ( 
.A1(n_16474),
.A2(n_6593),
.B1(n_6603),
.B2(n_6588),
.C(n_6587),
.Y(n_16541)
);

OAI22xp5_ASAP7_75t_L g16542 ( 
.A1(n_16402),
.A2(n_6848),
.B1(n_6880),
.B2(n_6857),
.Y(n_16542)
);

OAI211xp5_ASAP7_75t_SL g16543 ( 
.A1(n_16423),
.A2(n_6603),
.B(n_6604),
.C(n_6593),
.Y(n_16543)
);

NAND2xp33_ASAP7_75t_R g16544 ( 
.A(n_16447),
.B(n_6438),
.Y(n_16544)
);

AOI21xp5_ASAP7_75t_L g16545 ( 
.A1(n_16354),
.A2(n_7467),
.B(n_7968),
.Y(n_16545)
);

AOI21xp33_ASAP7_75t_L g16546 ( 
.A1(n_16448),
.A2(n_8215),
.B(n_8202),
.Y(n_16546)
);

INVx1_ASAP7_75t_SL g16547 ( 
.A(n_16358),
.Y(n_16547)
);

HB1xp67_ASAP7_75t_L g16548 ( 
.A(n_16415),
.Y(n_16548)
);

AOI211xp5_ASAP7_75t_L g16549 ( 
.A1(n_16469),
.A2(n_7976),
.B(n_7424),
.C(n_7428),
.Y(n_16549)
);

AOI221xp5_ASAP7_75t_L g16550 ( 
.A1(n_16467),
.A2(n_6612),
.B1(n_6618),
.B2(n_6609),
.C(n_6604),
.Y(n_16550)
);

AOI22xp5_ASAP7_75t_L g16551 ( 
.A1(n_16476),
.A2(n_7271),
.B1(n_8182),
.B2(n_7754),
.Y(n_16551)
);

HB1xp67_ASAP7_75t_L g16552 ( 
.A(n_16434),
.Y(n_16552)
);

NAND2xp33_ASAP7_75t_SL g16553 ( 
.A(n_16458),
.B(n_6927),
.Y(n_16553)
);

AOI221xp5_ASAP7_75t_L g16554 ( 
.A1(n_16411),
.A2(n_6612),
.B1(n_6618),
.B2(n_6609),
.C(n_6604),
.Y(n_16554)
);

INVx2_ASAP7_75t_L g16555 ( 
.A(n_16356),
.Y(n_16555)
);

NAND5xp2_ASAP7_75t_L g16556 ( 
.A(n_16366),
.B(n_16359),
.C(n_16385),
.D(n_16466),
.E(n_16439),
.Y(n_16556)
);

NOR2xp33_ASAP7_75t_L g16557 ( 
.A(n_16454),
.B(n_16479),
.Y(n_16557)
);

AOI22xp5_ASAP7_75t_SL g16558 ( 
.A1(n_16387),
.A2(n_7271),
.B1(n_6319),
.B2(n_6496),
.Y(n_16558)
);

AOI322xp5_ASAP7_75t_L g16559 ( 
.A1(n_16409),
.A2(n_6210),
.A3(n_6171),
.B1(n_6155),
.B2(n_6730),
.C1(n_6729),
.C2(n_6707),
.Y(n_16559)
);

NAND2xp5_ASAP7_75t_L g16560 ( 
.A(n_16392),
.B(n_8202),
.Y(n_16560)
);

AOI221x1_ASAP7_75t_L g16561 ( 
.A1(n_16400),
.A2(n_6438),
.B1(n_6522),
.B2(n_6612),
.C(n_6609),
.Y(n_16561)
);

A2O1A1Ixp33_ASAP7_75t_L g16562 ( 
.A1(n_16459),
.A2(n_7976),
.B(n_7789),
.C(n_7788),
.Y(n_16562)
);

BUFx12f_ASAP7_75t_L g16563 ( 
.A(n_16383),
.Y(n_16563)
);

O2A1O1Ixp33_ASAP7_75t_L g16564 ( 
.A1(n_16421),
.A2(n_6062),
.B(n_6026),
.C(n_6706),
.Y(n_16564)
);

OAI21xp5_ASAP7_75t_L g16565 ( 
.A1(n_16443),
.A2(n_7423),
.B(n_7976),
.Y(n_16565)
);

OAI21xp33_ASAP7_75t_L g16566 ( 
.A1(n_16360),
.A2(n_6522),
.B(n_6438),
.Y(n_16566)
);

CKINVDCx20_ASAP7_75t_R g16567 ( 
.A(n_16388),
.Y(n_16567)
);

OAI211xp5_ASAP7_75t_SL g16568 ( 
.A1(n_16475),
.A2(n_6621),
.B(n_6622),
.C(n_6618),
.Y(n_16568)
);

INVxp67_ASAP7_75t_SL g16569 ( 
.A(n_16471),
.Y(n_16569)
);

AOI222xp33_ASAP7_75t_L g16570 ( 
.A1(n_16441),
.A2(n_8182),
.B1(n_7754),
.B2(n_6628),
.C1(n_6622),
.C2(n_6632),
.Y(n_16570)
);

AOI21xp5_ASAP7_75t_L g16571 ( 
.A1(n_16414),
.A2(n_6622),
.B(n_6621),
.Y(n_16571)
);

OAI21xp5_ASAP7_75t_L g16572 ( 
.A1(n_16395),
.A2(n_8091),
.B(n_8076),
.Y(n_16572)
);

AOI221xp5_ASAP7_75t_L g16573 ( 
.A1(n_16452),
.A2(n_6628),
.B1(n_6632),
.B2(n_6626),
.C(n_6621),
.Y(n_16573)
);

NAND2xp5_ASAP7_75t_L g16574 ( 
.A(n_16462),
.B(n_8215),
.Y(n_16574)
);

NAND4xp25_ASAP7_75t_L g16575 ( 
.A(n_16472),
.B(n_6735),
.C(n_6757),
.D(n_6709),
.Y(n_16575)
);

INVx1_ASAP7_75t_L g16576 ( 
.A(n_16389),
.Y(n_16576)
);

INVx2_ASAP7_75t_L g16577 ( 
.A(n_16422),
.Y(n_16577)
);

INVx1_ASAP7_75t_L g16578 ( 
.A(n_16397),
.Y(n_16578)
);

INVx1_ASAP7_75t_L g16579 ( 
.A(n_16377),
.Y(n_16579)
);

HB1xp67_ASAP7_75t_L g16580 ( 
.A(n_16373),
.Y(n_16580)
);

AOI21xp5_ASAP7_75t_L g16581 ( 
.A1(n_16473),
.A2(n_6628),
.B(n_6626),
.Y(n_16581)
);

AOI21xp5_ASAP7_75t_L g16582 ( 
.A1(n_16390),
.A2(n_6632),
.B(n_6626),
.Y(n_16582)
);

INVx2_ASAP7_75t_L g16583 ( 
.A(n_16422),
.Y(n_16583)
);

NAND5xp2_ASAP7_75t_L g16584 ( 
.A(n_16433),
.B(n_6141),
.C(n_6347),
.D(n_6352),
.E(n_6255),
.Y(n_16584)
);

INVx2_ASAP7_75t_L g16585 ( 
.A(n_16417),
.Y(n_16585)
);

OAI22xp5_ASAP7_75t_L g16586 ( 
.A1(n_16419),
.A2(n_6880),
.B1(n_6921),
.B2(n_7113),
.Y(n_16586)
);

AOI21xp5_ASAP7_75t_L g16587 ( 
.A1(n_16386),
.A2(n_6644),
.B(n_6642),
.Y(n_16587)
);

OAI221xp5_ASAP7_75t_L g16588 ( 
.A1(n_16408),
.A2(n_6642),
.B1(n_6659),
.B2(n_6653),
.C(n_6644),
.Y(n_16588)
);

BUFx2_ASAP7_75t_L g16589 ( 
.A(n_16378),
.Y(n_16589)
);

NAND2xp5_ASAP7_75t_L g16590 ( 
.A(n_16429),
.B(n_8215),
.Y(n_16590)
);

INVx1_ASAP7_75t_L g16591 ( 
.A(n_16460),
.Y(n_16591)
);

NOR5xp2_ASAP7_75t_L g16592 ( 
.A(n_16425),
.B(n_6653),
.C(n_6659),
.D(n_6644),
.E(n_6642),
.Y(n_16592)
);

NAND2xp5_ASAP7_75t_L g16593 ( 
.A(n_16412),
.B(n_8264),
.Y(n_16593)
);

AOI22xp33_ASAP7_75t_L g16594 ( 
.A1(n_16371),
.A2(n_6463),
.B1(n_6630),
.B2(n_8215),
.Y(n_16594)
);

OAI211xp5_ASAP7_75t_SL g16595 ( 
.A1(n_16442),
.A2(n_6659),
.B(n_6661),
.C(n_6653),
.Y(n_16595)
);

INVx1_ASAP7_75t_SL g16596 ( 
.A(n_16456),
.Y(n_16596)
);

AOI222xp33_ASAP7_75t_L g16597 ( 
.A1(n_16437),
.A2(n_8182),
.B1(n_7754),
.B2(n_6684),
.C1(n_6672),
.C2(n_6688),
.Y(n_16597)
);

OAI21xp33_ASAP7_75t_SL g16598 ( 
.A1(n_16457),
.A2(n_7623),
.B(n_7622),
.Y(n_16598)
);

NOR3xp33_ASAP7_75t_L g16599 ( 
.A(n_16394),
.B(n_6041),
.C(n_6029),
.Y(n_16599)
);

HB1xp67_ASAP7_75t_L g16600 ( 
.A(n_16455),
.Y(n_16600)
);

NAND5xp2_ASAP7_75t_L g16601 ( 
.A(n_16470),
.B(n_6141),
.C(n_6347),
.D(n_6352),
.E(n_6255),
.Y(n_16601)
);

AOI22xp5_ASAP7_75t_L g16602 ( 
.A1(n_16477),
.A2(n_7754),
.B1(n_8182),
.B2(n_5077),
.Y(n_16602)
);

AOI221xp5_ASAP7_75t_L g16603 ( 
.A1(n_16464),
.A2(n_6680),
.B1(n_6684),
.B2(n_6672),
.C(n_6661),
.Y(n_16603)
);

AOI221xp5_ASAP7_75t_L g16604 ( 
.A1(n_16363),
.A2(n_6680),
.B1(n_6684),
.B2(n_6672),
.C(n_6661),
.Y(n_16604)
);

INVx1_ASAP7_75t_L g16605 ( 
.A(n_16468),
.Y(n_16605)
);

NAND2xp5_ASAP7_75t_L g16606 ( 
.A(n_16381),
.B(n_8240),
.Y(n_16606)
);

AOI22xp5_ASAP7_75t_L g16607 ( 
.A1(n_16451),
.A2(n_8182),
.B1(n_7754),
.B2(n_6213),
.Y(n_16607)
);

OAI211xp5_ASAP7_75t_SL g16608 ( 
.A1(n_16488),
.A2(n_16401),
.B(n_16435),
.C(n_16410),
.Y(n_16608)
);

NOR2x1_ASAP7_75t_L g16609 ( 
.A(n_16498),
.B(n_16407),
.Y(n_16609)
);

AOI22xp5_ASAP7_75t_L g16610 ( 
.A1(n_16508),
.A2(n_16428),
.B1(n_16482),
.B2(n_16403),
.Y(n_16610)
);

NAND2xp5_ASAP7_75t_SL g16611 ( 
.A(n_16502),
.B(n_16384),
.Y(n_16611)
);

AOI221xp5_ASAP7_75t_L g16612 ( 
.A1(n_16569),
.A2(n_16416),
.B1(n_16483),
.B2(n_16404),
.C(n_16481),
.Y(n_16612)
);

NOR2xp67_ASAP7_75t_SL g16613 ( 
.A(n_16513),
.B(n_16382),
.Y(n_16613)
);

AND4x1_ASAP7_75t_L g16614 ( 
.A(n_16526),
.B(n_16528),
.C(n_16538),
.D(n_16557),
.Y(n_16614)
);

NAND2xp5_ASAP7_75t_L g16615 ( 
.A(n_16494),
.B(n_16438),
.Y(n_16615)
);

AOI311xp33_ASAP7_75t_L g16616 ( 
.A1(n_16605),
.A2(n_16579),
.A3(n_16578),
.B(n_16576),
.C(n_16591),
.Y(n_16616)
);

NOR3xp33_ASAP7_75t_L g16617 ( 
.A(n_16525),
.B(n_16436),
.C(n_16430),
.Y(n_16617)
);

AOI221xp5_ASAP7_75t_L g16618 ( 
.A1(n_16524),
.A2(n_6690),
.B1(n_6692),
.B2(n_6688),
.C(n_6680),
.Y(n_16618)
);

AND4x1_ASAP7_75t_L g16619 ( 
.A(n_16535),
.B(n_6912),
.C(n_6902),
.D(n_6910),
.Y(n_16619)
);

OAI221xp5_ASAP7_75t_L g16620 ( 
.A1(n_16589),
.A2(n_6762),
.B1(n_6783),
.B2(n_6600),
.C(n_6248),
.Y(n_16620)
);

A2O1A1Ixp33_ASAP7_75t_L g16621 ( 
.A1(n_16596),
.A2(n_7532),
.B(n_7539),
.C(n_7788),
.Y(n_16621)
);

NOR2xp33_ASAP7_75t_L g16622 ( 
.A(n_16523),
.B(n_8182),
.Y(n_16622)
);

O2A1O1Ixp33_ASAP7_75t_L g16623 ( 
.A1(n_16580),
.A2(n_6757),
.B(n_6822),
.C(n_6735),
.Y(n_16623)
);

AND4x2_ASAP7_75t_L g16624 ( 
.A(n_16511),
.B(n_6319),
.C(n_6496),
.D(n_6142),
.Y(n_16624)
);

NAND4xp25_ASAP7_75t_L g16625 ( 
.A(n_16523),
.B(n_6757),
.C(n_6822),
.D(n_6735),
.Y(n_16625)
);

INVx1_ASAP7_75t_L g16626 ( 
.A(n_16563),
.Y(n_16626)
);

NAND4xp75_ASAP7_75t_L g16627 ( 
.A(n_16539),
.B(n_6463),
.C(n_6630),
.D(n_6913),
.Y(n_16627)
);

AOI22xp33_ASAP7_75t_L g16628 ( 
.A1(n_16585),
.A2(n_6463),
.B1(n_6630),
.B2(n_8240),
.Y(n_16628)
);

NAND4xp25_ASAP7_75t_L g16629 ( 
.A(n_16547),
.B(n_6822),
.C(n_6853),
.D(n_6757),
.Y(n_16629)
);

INVx1_ASAP7_75t_L g16630 ( 
.A(n_16567),
.Y(n_16630)
);

AOI221xp5_ASAP7_75t_SL g16631 ( 
.A1(n_16485),
.A2(n_6980),
.B1(n_6987),
.B2(n_6515),
.C(n_6319),
.Y(n_16631)
);

AOI221x1_ASAP7_75t_L g16632 ( 
.A1(n_16555),
.A2(n_6522),
.B1(n_6438),
.B2(n_6690),
.C(n_6688),
.Y(n_16632)
);

OAI221xp5_ASAP7_75t_L g16633 ( 
.A1(n_16553),
.A2(n_6248),
.B1(n_6783),
.B2(n_6762),
.C(n_6600),
.Y(n_16633)
);

XNOR2xp5_ASAP7_75t_L g16634 ( 
.A(n_16487),
.B(n_7191),
.Y(n_16634)
);

NOR2xp33_ASAP7_75t_R g16635 ( 
.A(n_16544),
.B(n_6935),
.Y(n_16635)
);

OAI221xp5_ASAP7_75t_L g16636 ( 
.A1(n_16600),
.A2(n_6248),
.B1(n_6783),
.B2(n_6762),
.C(n_6600),
.Y(n_16636)
);

INVx1_ASAP7_75t_L g16637 ( 
.A(n_16548),
.Y(n_16637)
);

INVx1_ASAP7_75t_L g16638 ( 
.A(n_16577),
.Y(n_16638)
);

NOR2xp33_ASAP7_75t_L g16639 ( 
.A(n_16493),
.B(n_6463),
.Y(n_16639)
);

AOI21xp5_ASAP7_75t_L g16640 ( 
.A1(n_16583),
.A2(n_6983),
.B(n_6935),
.Y(n_16640)
);

AOI211xp5_ASAP7_75t_SL g16641 ( 
.A1(n_16552),
.A2(n_6544),
.B(n_6562),
.C(n_6536),
.Y(n_16641)
);

AOI22xp5_ASAP7_75t_L g16642 ( 
.A1(n_16496),
.A2(n_6215),
.B1(n_6267),
.B2(n_6213),
.Y(n_16642)
);

AOI221xp5_ASAP7_75t_L g16643 ( 
.A1(n_16556),
.A2(n_6710),
.B1(n_6712),
.B2(n_6692),
.C(n_6690),
.Y(n_16643)
);

NAND4xp25_ASAP7_75t_L g16644 ( 
.A(n_16520),
.B(n_6853),
.C(n_6822),
.D(n_6927),
.Y(n_16644)
);

AOI221x1_ASAP7_75t_L g16645 ( 
.A1(n_16568),
.A2(n_6710),
.B1(n_6716),
.B2(n_6712),
.C(n_6692),
.Y(n_16645)
);

AOI221xp5_ASAP7_75t_L g16646 ( 
.A1(n_16518),
.A2(n_6716),
.B1(n_6717),
.B2(n_6712),
.C(n_6710),
.Y(n_16646)
);

NAND2xp5_ASAP7_75t_L g16647 ( 
.A(n_16581),
.B(n_8046),
.Y(n_16647)
);

NOR3xp33_ASAP7_75t_L g16648 ( 
.A(n_16501),
.B(n_6990),
.C(n_6927),
.Y(n_16648)
);

OAI211xp5_ASAP7_75t_SL g16649 ( 
.A1(n_16570),
.A2(n_16597),
.B(n_16541),
.C(n_16519),
.Y(n_16649)
);

AOI222xp33_ASAP7_75t_L g16650 ( 
.A1(n_16560),
.A2(n_6732),
.B1(n_6717),
.B2(n_6734),
.C1(n_6728),
.C2(n_6716),
.Y(n_16650)
);

OAI21xp33_ASAP7_75t_SL g16651 ( 
.A1(n_16575),
.A2(n_7789),
.B(n_7788),
.Y(n_16651)
);

NAND4xp25_ASAP7_75t_L g16652 ( 
.A(n_16534),
.B(n_6853),
.C(n_6990),
.D(n_6927),
.Y(n_16652)
);

AOI211xp5_ASAP7_75t_L g16653 ( 
.A1(n_16505),
.A2(n_7462),
.B(n_7425),
.C(n_7428),
.Y(n_16653)
);

AOI221xp5_ASAP7_75t_L g16654 ( 
.A1(n_16531),
.A2(n_16516),
.B1(n_16546),
.B2(n_16529),
.C(n_16515),
.Y(n_16654)
);

NAND2xp5_ASAP7_75t_SL g16655 ( 
.A(n_16503),
.B(n_16491),
.Y(n_16655)
);

AOI221x1_ASAP7_75t_L g16656 ( 
.A1(n_16527),
.A2(n_6728),
.B1(n_6734),
.B2(n_6732),
.C(n_6717),
.Y(n_16656)
);

AND2x2_ASAP7_75t_L g16657 ( 
.A(n_16558),
.B(n_6171),
.Y(n_16657)
);

A2O1A1Ixp33_ASAP7_75t_L g16658 ( 
.A1(n_16573),
.A2(n_7532),
.B(n_7539),
.C(n_7789),
.Y(n_16658)
);

AOI221xp5_ASAP7_75t_L g16659 ( 
.A1(n_16590),
.A2(n_6734),
.B1(n_6742),
.B2(n_6732),
.C(n_6728),
.Y(n_16659)
);

AOI211xp5_ASAP7_75t_L g16660 ( 
.A1(n_16595),
.A2(n_7462),
.B(n_7425),
.C(n_7428),
.Y(n_16660)
);

OAI22xp5_ASAP7_75t_L g16661 ( 
.A1(n_16551),
.A2(n_6880),
.B1(n_6921),
.B2(n_7113),
.Y(n_16661)
);

AOI211xp5_ASAP7_75t_L g16662 ( 
.A1(n_16588),
.A2(n_7462),
.B(n_7425),
.C(n_7448),
.Y(n_16662)
);

HB1xp67_ASAP7_75t_L g16663 ( 
.A(n_16593),
.Y(n_16663)
);

AND2x4_ASAP7_75t_L g16664 ( 
.A(n_16561),
.B(n_8008),
.Y(n_16664)
);

AOI22xp33_ASAP7_75t_L g16665 ( 
.A1(n_16491),
.A2(n_6463),
.B1(n_6630),
.B2(n_8240),
.Y(n_16665)
);

NAND2xp5_ASAP7_75t_L g16666 ( 
.A(n_16504),
.B(n_8053),
.Y(n_16666)
);

AOI21xp33_ASAP7_75t_SL g16667 ( 
.A1(n_16574),
.A2(n_6983),
.B(n_6935),
.Y(n_16667)
);

OAI321xp33_ASAP7_75t_L g16668 ( 
.A1(n_16540),
.A2(n_6921),
.A3(n_7140),
.B1(n_7124),
.B2(n_7113),
.C(n_6777),
.Y(n_16668)
);

OAI221xp5_ASAP7_75t_SL g16669 ( 
.A1(n_16606),
.A2(n_16598),
.B1(n_16545),
.B2(n_16564),
.C(n_16607),
.Y(n_16669)
);

A2O1A1Ixp33_ASAP7_75t_L g16670 ( 
.A1(n_16592),
.A2(n_7532),
.B(n_7539),
.C(n_7303),
.Y(n_16670)
);

NAND4xp75_ASAP7_75t_L g16671 ( 
.A(n_16533),
.B(n_6463),
.C(n_6913),
.D(n_6747),
.Y(n_16671)
);

AOI221xp5_ASAP7_75t_L g16672 ( 
.A1(n_16603),
.A2(n_16522),
.B1(n_16517),
.B2(n_16512),
.C(n_16495),
.Y(n_16672)
);

OAI211xp5_ASAP7_75t_L g16673 ( 
.A1(n_16536),
.A2(n_16509),
.B(n_16486),
.C(n_16499),
.Y(n_16673)
);

AOI211xp5_ASAP7_75t_SL g16674 ( 
.A1(n_16500),
.A2(n_6562),
.B(n_6566),
.C(n_6544),
.Y(n_16674)
);

AOI211xp5_ASAP7_75t_SL g16675 ( 
.A1(n_16530),
.A2(n_6562),
.B(n_6566),
.C(n_6544),
.Y(n_16675)
);

OAI22xp5_ASAP7_75t_L g16676 ( 
.A1(n_16514),
.A2(n_7124),
.B1(n_7140),
.B2(n_6718),
.Y(n_16676)
);

OAI22xp5_ASAP7_75t_L g16677 ( 
.A1(n_16532),
.A2(n_7124),
.B1(n_7140),
.B2(n_6718),
.Y(n_16677)
);

AOI322xp5_ASAP7_75t_L g16678 ( 
.A1(n_16510),
.A2(n_6210),
.A3(n_6635),
.B1(n_6171),
.B2(n_6252),
.C1(n_6219),
.C2(n_6304),
.Y(n_16678)
);

NOR2xp33_ASAP7_75t_R g16679 ( 
.A(n_16601),
.B(n_6935),
.Y(n_16679)
);

AOI221xp5_ASAP7_75t_L g16680 ( 
.A1(n_16550),
.A2(n_6750),
.B1(n_6777),
.B2(n_6747),
.C(n_6742),
.Y(n_16680)
);

NAND2xp5_ASAP7_75t_L g16681 ( 
.A(n_16571),
.B(n_16506),
.Y(n_16681)
);

O2A1O1Ixp33_ASAP7_75t_L g16682 ( 
.A1(n_16537),
.A2(n_6853),
.B(n_6747),
.C(n_6750),
.Y(n_16682)
);

AOI221x1_ASAP7_75t_L g16683 ( 
.A1(n_16543),
.A2(n_6750),
.B1(n_6781),
.B2(n_6777),
.C(n_6742),
.Y(n_16683)
);

NOR3x1_ASAP7_75t_L g16684 ( 
.A(n_16572),
.B(n_7827),
.C(n_7822),
.Y(n_16684)
);

NAND2xp33_ASAP7_75t_SL g16685 ( 
.A(n_16542),
.B(n_6927),
.Y(n_16685)
);

INVx1_ASAP7_75t_L g16686 ( 
.A(n_16587),
.Y(n_16686)
);

NAND4xp25_ASAP7_75t_SL g16687 ( 
.A(n_16599),
.B(n_6718),
.C(n_6912),
.D(n_6910),
.Y(n_16687)
);

A2O1A1Ixp33_ASAP7_75t_L g16688 ( 
.A1(n_16582),
.A2(n_7303),
.B(n_7448),
.C(n_7424),
.Y(n_16688)
);

OAI21xp5_ASAP7_75t_L g16689 ( 
.A1(n_16594),
.A2(n_8091),
.B(n_8076),
.Y(n_16689)
);

OAI21xp5_ASAP7_75t_SL g16690 ( 
.A1(n_16602),
.A2(n_6134),
.B(n_6210),
.Y(n_16690)
);

OAI22xp33_ASAP7_75t_L g16691 ( 
.A1(n_16492),
.A2(n_6999),
.B1(n_7030),
.B2(n_6990),
.Y(n_16691)
);

NAND2xp33_ASAP7_75t_R g16692 ( 
.A(n_16565),
.B(n_7865),
.Y(n_16692)
);

AOI21xp5_ASAP7_75t_SL g16693 ( 
.A1(n_16604),
.A2(n_7102),
.B(n_7098),
.Y(n_16693)
);

AOI221xp5_ASAP7_75t_L g16694 ( 
.A1(n_16490),
.A2(n_6793),
.B1(n_6808),
.B2(n_6784),
.C(n_6781),
.Y(n_16694)
);

OAI21xp33_ASAP7_75t_SL g16695 ( 
.A1(n_16559),
.A2(n_7627),
.B(n_7624),
.Y(n_16695)
);

NOR3xp33_ASAP7_75t_L g16696 ( 
.A(n_16584),
.B(n_6999),
.C(n_6990),
.Y(n_16696)
);

AOI221xp5_ASAP7_75t_L g16697 ( 
.A1(n_16489),
.A2(n_6793),
.B1(n_6808),
.B2(n_6784),
.C(n_6781),
.Y(n_16697)
);

AOI221xp5_ASAP7_75t_L g16698 ( 
.A1(n_16521),
.A2(n_6808),
.B1(n_6811),
.B2(n_6793),
.C(n_6784),
.Y(n_16698)
);

NAND3xp33_ASAP7_75t_SL g16699 ( 
.A(n_16549),
.B(n_6347),
.C(n_6255),
.Y(n_16699)
);

OAI21xp5_ASAP7_75t_L g16700 ( 
.A1(n_16554),
.A2(n_8091),
.B(n_8076),
.Y(n_16700)
);

NOR2xp33_ASAP7_75t_R g16701 ( 
.A(n_16566),
.B(n_6935),
.Y(n_16701)
);

OR2x2_ASAP7_75t_L g16702 ( 
.A(n_16586),
.B(n_8053),
.Y(n_16702)
);

NOR5xp2_ASAP7_75t_L g16703 ( 
.A(n_16562),
.B(n_6830),
.C(n_6832),
.D(n_6812),
.E(n_6811),
.Y(n_16703)
);

AOI31xp33_ASAP7_75t_L g16704 ( 
.A1(n_16497),
.A2(n_6255),
.A3(n_6352),
.B(n_6347),
.Y(n_16704)
);

AOI211xp5_ASAP7_75t_L g16705 ( 
.A1(n_16507),
.A2(n_7448),
.B(n_7456),
.C(n_7424),
.Y(n_16705)
);

NAND4xp25_ASAP7_75t_L g16706 ( 
.A(n_16488),
.B(n_6999),
.C(n_7030),
.D(n_6990),
.Y(n_16706)
);

OAI211xp5_ASAP7_75t_SL g16707 ( 
.A1(n_16488),
.A2(n_6812),
.B(n_6830),
.C(n_6811),
.Y(n_16707)
);

AND2x2_ASAP7_75t_L g16708 ( 
.A(n_16498),
.B(n_6210),
.Y(n_16708)
);

OAI22xp5_ASAP7_75t_L g16709 ( 
.A1(n_16569),
.A2(n_6179),
.B1(n_6192),
.B2(n_6177),
.Y(n_16709)
);

NOR4xp25_ASAP7_75t_L g16710 ( 
.A(n_16488),
.B(n_6830),
.C(n_6832),
.D(n_6812),
.Y(n_16710)
);

AOI21xp5_ASAP7_75t_L g16711 ( 
.A1(n_16494),
.A2(n_7026),
.B(n_6983),
.Y(n_16711)
);

OAI22xp5_ASAP7_75t_L g16712 ( 
.A1(n_16569),
.A2(n_6179),
.B1(n_6192),
.B2(n_6177),
.Y(n_16712)
);

NAND2xp5_ASAP7_75t_L g16713 ( 
.A(n_16494),
.B(n_8053),
.Y(n_16713)
);

AOI211x1_ASAP7_75t_SL g16714 ( 
.A1(n_16585),
.A2(n_7129),
.B(n_7128),
.C(n_7136),
.Y(n_16714)
);

A2O1A1Ixp33_ASAP7_75t_L g16715 ( 
.A1(n_16569),
.A2(n_7303),
.B(n_7456),
.C(n_7624),
.Y(n_16715)
);

AOI211xp5_ASAP7_75t_L g16716 ( 
.A1(n_16498),
.A2(n_7456),
.B(n_8095),
.C(n_8094),
.Y(n_16716)
);

OAI22xp5_ASAP7_75t_L g16717 ( 
.A1(n_16569),
.A2(n_6179),
.B1(n_6192),
.B2(n_6177),
.Y(n_16717)
);

OAI21xp5_ASAP7_75t_L g16718 ( 
.A1(n_16494),
.A2(n_8095),
.B(n_8094),
.Y(n_16718)
);

AOI221xp5_ASAP7_75t_L g16719 ( 
.A1(n_16498),
.A2(n_6836),
.B1(n_6843),
.B2(n_6833),
.C(n_6832),
.Y(n_16719)
);

OAI211xp5_ASAP7_75t_L g16720 ( 
.A1(n_16488),
.A2(n_7026),
.B(n_7137),
.C(n_6983),
.Y(n_16720)
);

NOR3xp33_ASAP7_75t_L g16721 ( 
.A(n_16498),
.B(n_7030),
.C(n_6999),
.Y(n_16721)
);

OA21x2_ASAP7_75t_L g16722 ( 
.A1(n_16630),
.A2(n_7865),
.B(n_7827),
.Y(n_16722)
);

INVx1_ASAP7_75t_L g16723 ( 
.A(n_16626),
.Y(n_16723)
);

HB1xp67_ASAP7_75t_L g16724 ( 
.A(n_16637),
.Y(n_16724)
);

NOR3xp33_ASAP7_75t_SL g16725 ( 
.A(n_16615),
.B(n_6836),
.C(n_6833),
.Y(n_16725)
);

NAND3xp33_ASAP7_75t_L g16726 ( 
.A(n_16613),
.B(n_5188),
.C(n_5127),
.Y(n_16726)
);

NAND3xp33_ASAP7_75t_SL g16727 ( 
.A(n_16614),
.B(n_6352),
.C(n_6347),
.Y(n_16727)
);

NAND3xp33_ASAP7_75t_L g16728 ( 
.A(n_16616),
.B(n_5188),
.C(n_5127),
.Y(n_16728)
);

NOR3xp33_ASAP7_75t_L g16729 ( 
.A(n_16638),
.B(n_16663),
.C(n_16611),
.Y(n_16729)
);

NAND3xp33_ASAP7_75t_SL g16730 ( 
.A(n_16617),
.B(n_16612),
.C(n_16610),
.Y(n_16730)
);

NAND2xp5_ASAP7_75t_L g16731 ( 
.A(n_16609),
.B(n_8053),
.Y(n_16731)
);

NAND4xp75_ASAP7_75t_L g16732 ( 
.A(n_16655),
.B(n_6913),
.C(n_6836),
.D(n_6843),
.Y(n_16732)
);

NOR2xp33_ASAP7_75t_L g16733 ( 
.A(n_16713),
.B(n_7191),
.Y(n_16733)
);

NAND2xp5_ASAP7_75t_L g16734 ( 
.A(n_16622),
.B(n_8053),
.Y(n_16734)
);

NOR2x1_ASAP7_75t_L g16735 ( 
.A(n_16686),
.B(n_7191),
.Y(n_16735)
);

NAND2xp5_ASAP7_75t_L g16736 ( 
.A(n_16708),
.B(n_8053),
.Y(n_16736)
);

AND4x2_ASAP7_75t_L g16737 ( 
.A(n_16654),
.B(n_8053),
.C(n_7991),
.D(n_7989),
.Y(n_16737)
);

NAND2x1_ASAP7_75t_SL g16738 ( 
.A(n_16657),
.B(n_6999),
.Y(n_16738)
);

INVx1_ASAP7_75t_L g16739 ( 
.A(n_16681),
.Y(n_16739)
);

NOR2x1_ASAP7_75t_L g16740 ( 
.A(n_16608),
.B(n_7191),
.Y(n_16740)
);

NAND2xp5_ASAP7_75t_L g16741 ( 
.A(n_16714),
.B(n_8053),
.Y(n_16741)
);

INVx1_ASAP7_75t_L g16742 ( 
.A(n_16673),
.Y(n_16742)
);

BUFx3_ASAP7_75t_L g16743 ( 
.A(n_16634),
.Y(n_16743)
);

INVx1_ASAP7_75t_L g16744 ( 
.A(n_16649),
.Y(n_16744)
);

NOR2x1_ASAP7_75t_L g16745 ( 
.A(n_16711),
.B(n_7191),
.Y(n_16745)
);

INVxp67_ASAP7_75t_L g16746 ( 
.A(n_16639),
.Y(n_16746)
);

NOR2x1_ASAP7_75t_L g16747 ( 
.A(n_16652),
.B(n_7191),
.Y(n_16747)
);

HB1xp67_ASAP7_75t_L g16748 ( 
.A(n_16635),
.Y(n_16748)
);

NAND4xp75_ASAP7_75t_L g16749 ( 
.A(n_16672),
.B(n_6913),
.C(n_6843),
.D(n_6851),
.Y(n_16749)
);

AND2x2_ASAP7_75t_L g16750 ( 
.A(n_16679),
.B(n_6819),
.Y(n_16750)
);

INVx2_ASAP7_75t_SL g16751 ( 
.A(n_16701),
.Y(n_16751)
);

INVx1_ASAP7_75t_L g16752 ( 
.A(n_16669),
.Y(n_16752)
);

INVx1_ASAP7_75t_L g16753 ( 
.A(n_16702),
.Y(n_16753)
);

NOR2xp67_ASAP7_75t_L g16754 ( 
.A(n_16640),
.B(n_6999),
.Y(n_16754)
);

INVx1_ASAP7_75t_L g16755 ( 
.A(n_16647),
.Y(n_16755)
);

NOR3xp33_ASAP7_75t_L g16756 ( 
.A(n_16667),
.B(n_7048),
.C(n_7030),
.Y(n_16756)
);

NAND2xp5_ASAP7_75t_L g16757 ( 
.A(n_16646),
.B(n_7989),
.Y(n_16757)
);

INVx1_ASAP7_75t_L g16758 ( 
.A(n_16666),
.Y(n_16758)
);

NOR4xp75_ASAP7_75t_L g16759 ( 
.A(n_16671),
.B(n_6566),
.C(n_6596),
.D(n_6562),
.Y(n_16759)
);

NOR2x1_ASAP7_75t_L g16760 ( 
.A(n_16644),
.B(n_7221),
.Y(n_16760)
);

NOR2xp67_ASAP7_75t_L g16761 ( 
.A(n_16625),
.B(n_16629),
.Y(n_16761)
);

INVx1_ASAP7_75t_L g16762 ( 
.A(n_16656),
.Y(n_16762)
);

NAND4xp75_ASAP7_75t_L g16763 ( 
.A(n_16695),
.B(n_16631),
.C(n_16684),
.D(n_16651),
.Y(n_16763)
);

NAND2xp5_ASAP7_75t_SL g16764 ( 
.A(n_16623),
.B(n_6213),
.Y(n_16764)
);

OR2x2_ASAP7_75t_L g16765 ( 
.A(n_16699),
.B(n_7989),
.Y(n_16765)
);

INVx2_ASAP7_75t_SL g16766 ( 
.A(n_16664),
.Y(n_16766)
);

NAND2x1_ASAP7_75t_L g16767 ( 
.A(n_16693),
.B(n_7151),
.Y(n_16767)
);

INVx1_ASAP7_75t_L g16768 ( 
.A(n_16624),
.Y(n_16768)
);

AND2x4_ASAP7_75t_L g16769 ( 
.A(n_16696),
.B(n_8008),
.Y(n_16769)
);

NOR2x1_ASAP7_75t_L g16770 ( 
.A(n_16690),
.B(n_7221),
.Y(n_16770)
);

INVx1_ASAP7_75t_SL g16771 ( 
.A(n_16685),
.Y(n_16771)
);

NOR2xp33_ASAP7_75t_L g16772 ( 
.A(n_16682),
.B(n_7221),
.Y(n_16772)
);

INVx1_ASAP7_75t_L g16773 ( 
.A(n_16659),
.Y(n_16773)
);

NOR2xp33_ASAP7_75t_L g16774 ( 
.A(n_16720),
.B(n_7221),
.Y(n_16774)
);

INVx2_ASAP7_75t_L g16775 ( 
.A(n_16664),
.Y(n_16775)
);

INVx1_ASAP7_75t_L g16776 ( 
.A(n_16650),
.Y(n_16776)
);

INVx1_ASAP7_75t_L g16777 ( 
.A(n_16645),
.Y(n_16777)
);

NAND2xp5_ASAP7_75t_L g16778 ( 
.A(n_16674),
.B(n_7989),
.Y(n_16778)
);

NAND4xp25_ASAP7_75t_L g16779 ( 
.A(n_16675),
.B(n_7048),
.C(n_7051),
.D(n_7030),
.Y(n_16779)
);

NOR3x2_ASAP7_75t_L g16780 ( 
.A(n_16627),
.B(n_16703),
.C(n_16692),
.Y(n_16780)
);

NAND2xp5_ASAP7_75t_SL g16781 ( 
.A(n_16718),
.B(n_6213),
.Y(n_16781)
);

INVx1_ASAP7_75t_L g16782 ( 
.A(n_16689),
.Y(n_16782)
);

INVx1_ASAP7_75t_L g16783 ( 
.A(n_16683),
.Y(n_16783)
);

INVx1_ASAP7_75t_L g16784 ( 
.A(n_16707),
.Y(n_16784)
);

AND2x2_ASAP7_75t_L g16785 ( 
.A(n_16619),
.B(n_6819),
.Y(n_16785)
);

AOI22xp5_ASAP7_75t_L g16786 ( 
.A1(n_16687),
.A2(n_6215),
.B1(n_6267),
.B2(n_6213),
.Y(n_16786)
);

NOR2x1_ASAP7_75t_L g16787 ( 
.A(n_16620),
.B(n_7221),
.Y(n_16787)
);

AND2x4_ASAP7_75t_L g16788 ( 
.A(n_16721),
.B(n_8063),
.Y(n_16788)
);

NAND4xp25_ASAP7_75t_L g16789 ( 
.A(n_16678),
.B(n_7048),
.C(n_7051),
.D(n_7030),
.Y(n_16789)
);

INVx2_ASAP7_75t_L g16790 ( 
.A(n_16633),
.Y(n_16790)
);

NOR3xp33_ASAP7_75t_L g16791 ( 
.A(n_16668),
.B(n_7051),
.C(n_7048),
.Y(n_16791)
);

NOR2x1_ASAP7_75t_L g16792 ( 
.A(n_16700),
.B(n_16691),
.Y(n_16792)
);

OR2x2_ASAP7_75t_L g16793 ( 
.A(n_16710),
.B(n_7989),
.Y(n_16793)
);

AND2x2_ASAP7_75t_L g16794 ( 
.A(n_16648),
.B(n_6819),
.Y(n_16794)
);

INVx1_ASAP7_75t_L g16795 ( 
.A(n_16632),
.Y(n_16795)
);

NOR2xp67_ASAP7_75t_SL g16796 ( 
.A(n_16636),
.B(n_16706),
.Y(n_16796)
);

NAND4xp75_ASAP7_75t_L g16797 ( 
.A(n_16643),
.B(n_6913),
.C(n_6851),
.D(n_6861),
.Y(n_16797)
);

AND2x4_ASAP7_75t_L g16798 ( 
.A(n_16642),
.B(n_8063),
.Y(n_16798)
);

NOR3xp33_ASAP7_75t_L g16799 ( 
.A(n_16698),
.B(n_7051),
.C(n_7048),
.Y(n_16799)
);

NOR2x1p5_ASAP7_75t_L g16800 ( 
.A(n_16653),
.B(n_7098),
.Y(n_16800)
);

NAND2xp5_ASAP7_75t_L g16801 ( 
.A(n_16694),
.B(n_7989),
.Y(n_16801)
);

NOR4xp75_ASAP7_75t_L g16802 ( 
.A(n_16709),
.B(n_6596),
.C(n_6713),
.D(n_6566),
.Y(n_16802)
);

NAND2xp5_ASAP7_75t_L g16803 ( 
.A(n_16641),
.B(n_7989),
.Y(n_16803)
);

INVx1_ASAP7_75t_L g16804 ( 
.A(n_16677),
.Y(n_16804)
);

NAND2xp5_ASAP7_75t_L g16805 ( 
.A(n_16680),
.B(n_7989),
.Y(n_16805)
);

AND2x4_ASAP7_75t_L g16806 ( 
.A(n_16628),
.B(n_8092),
.Y(n_16806)
);

INVx1_ASAP7_75t_L g16807 ( 
.A(n_16661),
.Y(n_16807)
);

NAND4xp25_ASAP7_75t_L g16808 ( 
.A(n_16660),
.B(n_7051),
.C(n_7071),
.D(n_7048),
.Y(n_16808)
);

OR2x2_ASAP7_75t_L g16809 ( 
.A(n_16712),
.B(n_7991),
.Y(n_16809)
);

INVx1_ASAP7_75t_L g16810 ( 
.A(n_16717),
.Y(n_16810)
);

NOR2x1_ASAP7_75t_L g16811 ( 
.A(n_16704),
.B(n_7221),
.Y(n_16811)
);

AND2x4_ASAP7_75t_L g16812 ( 
.A(n_16688),
.B(n_8063),
.Y(n_16812)
);

NAND3xp33_ASAP7_75t_L g16813 ( 
.A(n_16662),
.B(n_5188),
.C(n_5127),
.Y(n_16813)
);

HB1xp67_ASAP7_75t_L g16814 ( 
.A(n_16705),
.Y(n_16814)
);

NOR3xp33_ASAP7_75t_L g16815 ( 
.A(n_16697),
.B(n_7071),
.C(n_7051),
.Y(n_16815)
);

NOR3xp33_ASAP7_75t_L g16816 ( 
.A(n_16724),
.B(n_16723),
.C(n_16730),
.Y(n_16816)
);

AOI221xp5_ASAP7_75t_L g16817 ( 
.A1(n_16729),
.A2(n_16719),
.B1(n_16618),
.B2(n_16665),
.C(n_16676),
.Y(n_16817)
);

NAND3xp33_ASAP7_75t_SL g16818 ( 
.A(n_16744),
.B(n_16716),
.C(n_16621),
.Y(n_16818)
);

NAND4xp75_ASAP7_75t_L g16819 ( 
.A(n_16742),
.B(n_16658),
.C(n_16670),
.D(n_16715),
.Y(n_16819)
);

NAND3xp33_ASAP7_75t_SL g16820 ( 
.A(n_16752),
.B(n_16775),
.C(n_16739),
.Y(n_16820)
);

OAI221xp5_ASAP7_75t_SL g16821 ( 
.A1(n_16768),
.A2(n_7109),
.B1(n_7110),
.B2(n_7102),
.C(n_7098),
.Y(n_16821)
);

NOR2x1_ASAP7_75t_L g16822 ( 
.A(n_16743),
.B(n_6860),
.Y(n_16822)
);

NAND2xp5_ASAP7_75t_L g16823 ( 
.A(n_16766),
.B(n_7991),
.Y(n_16823)
);

NAND4xp25_ASAP7_75t_L g16824 ( 
.A(n_16761),
.B(n_7071),
.C(n_7102),
.D(n_7098),
.Y(n_16824)
);

NAND3xp33_ASAP7_75t_SL g16825 ( 
.A(n_16758),
.B(n_6352),
.C(n_6041),
.Y(n_16825)
);

AND2x2_ASAP7_75t_L g16826 ( 
.A(n_16740),
.B(n_8092),
.Y(n_16826)
);

OAI22xp33_ASAP7_75t_L g16827 ( 
.A1(n_16731),
.A2(n_16795),
.B1(n_16771),
.B2(n_16748),
.Y(n_16827)
);

NAND2xp5_ASAP7_75t_L g16828 ( 
.A(n_16753),
.B(n_7991),
.Y(n_16828)
);

NAND3xp33_ASAP7_75t_SL g16829 ( 
.A(n_16755),
.B(n_16746),
.C(n_16790),
.Y(n_16829)
);

A2O1A1Ixp33_ASAP7_75t_SL g16830 ( 
.A1(n_16776),
.A2(n_6566),
.B(n_6713),
.C(n_6596),
.Y(n_16830)
);

NAND2xp5_ASAP7_75t_L g16831 ( 
.A(n_16751),
.B(n_7991),
.Y(n_16831)
);

NAND2xp5_ASAP7_75t_L g16832 ( 
.A(n_16782),
.B(n_7991),
.Y(n_16832)
);

AND2x2_ASAP7_75t_L g16833 ( 
.A(n_16750),
.B(n_16785),
.Y(n_16833)
);

HB1xp67_ASAP7_75t_L g16834 ( 
.A(n_16814),
.Y(n_16834)
);

AND2x2_ASAP7_75t_L g16835 ( 
.A(n_16760),
.B(n_8092),
.Y(n_16835)
);

OR2x2_ASAP7_75t_L g16836 ( 
.A(n_16767),
.B(n_7991),
.Y(n_16836)
);

AOI322xp5_ASAP7_75t_L g16837 ( 
.A1(n_16783),
.A2(n_6696),
.A3(n_6635),
.B1(n_6216),
.B2(n_6219),
.C1(n_6304),
.C2(n_6313),
.Y(n_16837)
);

NOR3xp33_ASAP7_75t_L g16838 ( 
.A(n_16810),
.B(n_7071),
.C(n_6041),
.Y(n_16838)
);

AOI21xp5_ASAP7_75t_L g16839 ( 
.A1(n_16762),
.A2(n_7026),
.B(n_6983),
.Y(n_16839)
);

OAI211xp5_ASAP7_75t_L g16840 ( 
.A1(n_16773),
.A2(n_7137),
.B(n_7026),
.C(n_7071),
.Y(n_16840)
);

NAND5xp2_ASAP7_75t_L g16841 ( 
.A(n_16804),
.B(n_6987),
.C(n_6980),
.D(n_6515),
.E(n_4758),
.Y(n_16841)
);

AND4x1_ASAP7_75t_L g16842 ( 
.A(n_16796),
.B(n_6833),
.C(n_6861),
.D(n_6851),
.Y(n_16842)
);

A2O1A1Ixp33_ASAP7_75t_L g16843 ( 
.A1(n_16777),
.A2(n_7627),
.B(n_7624),
.C(n_8146),
.Y(n_16843)
);

NAND2xp5_ASAP7_75t_L g16844 ( 
.A(n_16763),
.B(n_7991),
.Y(n_16844)
);

NAND3xp33_ASAP7_75t_SL g16845 ( 
.A(n_16807),
.B(n_6041),
.C(n_6029),
.Y(n_16845)
);

NAND5xp2_ASAP7_75t_L g16846 ( 
.A(n_16784),
.B(n_6987),
.C(n_6515),
.D(n_4758),
.E(n_4594),
.Y(n_16846)
);

OAI211xp5_ASAP7_75t_SL g16847 ( 
.A1(n_16792),
.A2(n_6863),
.B(n_6864),
.C(n_6861),
.Y(n_16847)
);

NAND4xp25_ASAP7_75t_L g16848 ( 
.A(n_16728),
.B(n_7071),
.C(n_7109),
.D(n_7102),
.Y(n_16848)
);

NAND3xp33_ASAP7_75t_SL g16849 ( 
.A(n_16725),
.B(n_6029),
.C(n_5762),
.Y(n_16849)
);

NAND2x1_ASAP7_75t_L g16850 ( 
.A(n_16754),
.B(n_7151),
.Y(n_16850)
);

NOR2x1_ASAP7_75t_SL g16851 ( 
.A(n_16764),
.B(n_16726),
.Y(n_16851)
);

OAI21xp33_ASAP7_75t_L g16852 ( 
.A1(n_16738),
.A2(n_7627),
.B(n_5182),
.Y(n_16852)
);

OAI221xp5_ASAP7_75t_L g16853 ( 
.A1(n_16733),
.A2(n_6600),
.B1(n_6783),
.B2(n_6762),
.C(n_6248),
.Y(n_16853)
);

INVx1_ASAP7_75t_L g16854 ( 
.A(n_16780),
.Y(n_16854)
);

AOI21x1_ASAP7_75t_L g16855 ( 
.A1(n_16741),
.A2(n_16781),
.B(n_16778),
.Y(n_16855)
);

OR2x2_ASAP7_75t_L g16856 ( 
.A(n_16736),
.B(n_7221),
.Y(n_16856)
);

O2A1O1Ixp33_ASAP7_75t_L g16857 ( 
.A1(n_16734),
.A2(n_7110),
.B(n_7120),
.C(n_7109),
.Y(n_16857)
);

OAI211xp5_ASAP7_75t_SL g16858 ( 
.A1(n_16809),
.A2(n_6864),
.B(n_6878),
.C(n_6863),
.Y(n_16858)
);

OAI211xp5_ASAP7_75t_SL g16859 ( 
.A1(n_16765),
.A2(n_6864),
.B(n_6878),
.C(n_6863),
.Y(n_16859)
);

NAND3xp33_ASAP7_75t_SL g16860 ( 
.A(n_16759),
.B(n_5762),
.C(n_5732),
.Y(n_16860)
);

NAND2xp5_ASAP7_75t_SL g16861 ( 
.A(n_16769),
.B(n_6213),
.Y(n_16861)
);

OAI211xp5_ASAP7_75t_L g16862 ( 
.A1(n_16747),
.A2(n_7137),
.B(n_7026),
.C(n_7110),
.Y(n_16862)
);

NOR3xp33_ASAP7_75t_L g16863 ( 
.A(n_16774),
.B(n_5762),
.C(n_5732),
.Y(n_16863)
);

AOI211xp5_ASAP7_75t_L g16864 ( 
.A1(n_16772),
.A2(n_7154),
.B(n_7136),
.C(n_6215),
.Y(n_16864)
);

NOR3xp33_ASAP7_75t_L g16865 ( 
.A(n_16745),
.B(n_16787),
.C(n_16813),
.Y(n_16865)
);

NAND2xp5_ASAP7_75t_L g16866 ( 
.A(n_16800),
.B(n_6878),
.Y(n_16866)
);

AND4x1_ASAP7_75t_L g16867 ( 
.A(n_16811),
.B(n_6885),
.C(n_6889),
.D(n_6887),
.Y(n_16867)
);

NAND4xp25_ASAP7_75t_L g16868 ( 
.A(n_16770),
.B(n_7110),
.C(n_7120),
.D(n_7109),
.Y(n_16868)
);

OAI221xp5_ASAP7_75t_SL g16869 ( 
.A1(n_16791),
.A2(n_7120),
.B1(n_6962),
.B2(n_6978),
.C(n_6961),
.Y(n_16869)
);

NOR5xp2_ASAP7_75t_L g16870 ( 
.A(n_16808),
.B(n_6889),
.C(n_6890),
.D(n_6887),
.E(n_6885),
.Y(n_16870)
);

OAI211xp5_ASAP7_75t_SL g16871 ( 
.A1(n_16757),
.A2(n_6887),
.B(n_6889),
.C(n_6885),
.Y(n_16871)
);

AOI211xp5_ASAP7_75t_L g16872 ( 
.A1(n_16801),
.A2(n_7154),
.B(n_7136),
.C(n_6215),
.Y(n_16872)
);

AOI322xp5_ASAP7_75t_L g16873 ( 
.A1(n_16769),
.A2(n_6696),
.A3(n_6635),
.B1(n_6216),
.B2(n_6219),
.C1(n_6304),
.C2(n_6313),
.Y(n_16873)
);

AOI211xp5_ASAP7_75t_L g16874 ( 
.A1(n_16793),
.A2(n_7154),
.B(n_7136),
.C(n_6215),
.Y(n_16874)
);

OAI311xp33_ASAP7_75t_L g16875 ( 
.A1(n_16789),
.A2(n_6713),
.A3(n_6765),
.B1(n_6736),
.C1(n_6596),
.Y(n_16875)
);

OAI211xp5_ASAP7_75t_SL g16876 ( 
.A1(n_16805),
.A2(n_6901),
.B(n_6908),
.C(n_6890),
.Y(n_16876)
);

NAND2xp5_ASAP7_75t_L g16877 ( 
.A(n_16794),
.B(n_6890),
.Y(n_16877)
);

NAND4xp25_ASAP7_75t_L g16878 ( 
.A(n_16735),
.B(n_7120),
.C(n_6961),
.D(n_6962),
.Y(n_16878)
);

INVx1_ASAP7_75t_L g16879 ( 
.A(n_16803),
.Y(n_16879)
);

AOI221xp5_ASAP7_75t_L g16880 ( 
.A1(n_16812),
.A2(n_6267),
.B1(n_6297),
.B2(n_6215),
.C(n_6213),
.Y(n_16880)
);

OR2x2_ASAP7_75t_L g16881 ( 
.A(n_16749),
.B(n_16806),
.Y(n_16881)
);

NOR2x1p5_ASAP7_75t_L g16882 ( 
.A(n_16797),
.B(n_6596),
.Y(n_16882)
);

NAND2x1p5_ASAP7_75t_SL g16883 ( 
.A(n_16737),
.B(n_5336),
.Y(n_16883)
);

NOR2x1_ASAP7_75t_L g16884 ( 
.A(n_16727),
.B(n_6860),
.Y(n_16884)
);

INVx1_ASAP7_75t_L g16885 ( 
.A(n_16802),
.Y(n_16885)
);

NAND2xp5_ASAP7_75t_L g16886 ( 
.A(n_16806),
.B(n_6901),
.Y(n_16886)
);

NAND5xp2_ASAP7_75t_L g16887 ( 
.A(n_16756),
.B(n_4594),
.C(n_5549),
.D(n_5611),
.E(n_5533),
.Y(n_16887)
);

NOR4xp25_ASAP7_75t_L g16888 ( 
.A(n_16779),
.B(n_16732),
.C(n_16812),
.D(n_16799),
.Y(n_16888)
);

NAND4xp25_ASAP7_75t_L g16889 ( 
.A(n_16815),
.B(n_6961),
.C(n_6962),
.D(n_6951),
.Y(n_16889)
);

OAI221xp5_ASAP7_75t_L g16890 ( 
.A1(n_16786),
.A2(n_6600),
.B1(n_6783),
.B2(n_6762),
.C(n_6248),
.Y(n_16890)
);

AND3x1_ASAP7_75t_L g16891 ( 
.A(n_16788),
.B(n_6736),
.C(n_6713),
.Y(n_16891)
);

NOR2x1_ASAP7_75t_L g16892 ( 
.A(n_16788),
.B(n_6860),
.Y(n_16892)
);

NAND3xp33_ASAP7_75t_SL g16893 ( 
.A(n_16798),
.B(n_5762),
.C(n_5732),
.Y(n_16893)
);

AOI211x1_ASAP7_75t_SL g16894 ( 
.A1(n_16798),
.A2(n_6444),
.B(n_6449),
.C(n_6441),
.Y(n_16894)
);

AOI21xp5_ASAP7_75t_L g16895 ( 
.A1(n_16722),
.A2(n_7137),
.B(n_7026),
.Y(n_16895)
);

NOR3xp33_ASAP7_75t_L g16896 ( 
.A(n_16722),
.B(n_5762),
.C(n_5732),
.Y(n_16896)
);

INVx2_ASAP7_75t_L g16897 ( 
.A(n_16834),
.Y(n_16897)
);

NOR2xp67_ASAP7_75t_L g16898 ( 
.A(n_16820),
.B(n_4809),
.Y(n_16898)
);

NOR3xp33_ASAP7_75t_L g16899 ( 
.A(n_16816),
.B(n_5795),
.C(n_5732),
.Y(n_16899)
);

NAND2xp5_ASAP7_75t_SL g16900 ( 
.A(n_16854),
.B(n_6213),
.Y(n_16900)
);

AND2x4_ASAP7_75t_L g16901 ( 
.A(n_16833),
.B(n_16865),
.Y(n_16901)
);

OAI22xp5_ASAP7_75t_L g16902 ( 
.A1(n_16844),
.A2(n_6248),
.B1(n_6762),
.B2(n_6600),
.Y(n_16902)
);

INVx2_ASAP7_75t_L g16903 ( 
.A(n_16885),
.Y(n_16903)
);

NAND4xp25_ASAP7_75t_L g16904 ( 
.A(n_16829),
.B(n_16818),
.C(n_16879),
.D(n_16817),
.Y(n_16904)
);

BUFx12f_ASAP7_75t_L g16905 ( 
.A(n_16881),
.Y(n_16905)
);

NOR2xp33_ASAP7_75t_SL g16906 ( 
.A(n_16827),
.B(n_16819),
.Y(n_16906)
);

AND2x2_ASAP7_75t_L g16907 ( 
.A(n_16826),
.B(n_7552),
.Y(n_16907)
);

NOR2x1_ASAP7_75t_L g16908 ( 
.A(n_16822),
.B(n_7552),
.Y(n_16908)
);

INVx1_ASAP7_75t_L g16909 ( 
.A(n_16855),
.Y(n_16909)
);

NAND2xp5_ASAP7_75t_L g16910 ( 
.A(n_16874),
.B(n_8121),
.Y(n_16910)
);

XNOR2x1_ASAP7_75t_L g16911 ( 
.A(n_16856),
.B(n_7552),
.Y(n_16911)
);

NAND3x1_ASAP7_75t_L g16912 ( 
.A(n_16892),
.B(n_6908),
.C(n_6901),
.Y(n_16912)
);

INVx2_ASAP7_75t_SL g16913 ( 
.A(n_16850),
.Y(n_16913)
);

NOR2x1p5_ASAP7_75t_L g16914 ( 
.A(n_16866),
.B(n_16828),
.Y(n_16914)
);

XNOR2xp5_ASAP7_75t_L g16915 ( 
.A(n_16872),
.B(n_7552),
.Y(n_16915)
);

AND2x4_ASAP7_75t_L g16916 ( 
.A(n_16851),
.B(n_6696),
.Y(n_16916)
);

NAND4xp75_ASAP7_75t_L g16917 ( 
.A(n_16884),
.B(n_6912),
.C(n_6930),
.D(n_6910),
.Y(n_16917)
);

INVx1_ASAP7_75t_L g16918 ( 
.A(n_16876),
.Y(n_16918)
);

XNOR2xp5_ASAP7_75t_L g16919 ( 
.A(n_16888),
.B(n_7552),
.Y(n_16919)
);

NOR3xp33_ASAP7_75t_L g16920 ( 
.A(n_16871),
.B(n_5811),
.C(n_5795),
.Y(n_16920)
);

NAND2xp5_ASAP7_75t_L g16921 ( 
.A(n_16835),
.B(n_7949),
.Y(n_16921)
);

INVx1_ASAP7_75t_L g16922 ( 
.A(n_16858),
.Y(n_16922)
);

AOI22xp33_ASAP7_75t_L g16923 ( 
.A1(n_16859),
.A2(n_7154),
.B1(n_7136),
.B2(n_7129),
.Y(n_16923)
);

NAND2xp5_ASAP7_75t_L g16924 ( 
.A(n_16864),
.B(n_7949),
.Y(n_16924)
);

INVx1_ASAP7_75t_L g16925 ( 
.A(n_16883),
.Y(n_16925)
);

INVxp67_ASAP7_75t_L g16926 ( 
.A(n_16832),
.Y(n_16926)
);

AO22x1_ASAP7_75t_L g16927 ( 
.A1(n_16863),
.A2(n_5188),
.B1(n_5127),
.B2(n_6696),
.Y(n_16927)
);

OAI22xp5_ASAP7_75t_SL g16928 ( 
.A1(n_16891),
.A2(n_16877),
.B1(n_16831),
.B2(n_16823),
.Y(n_16928)
);

AND2x4_ASAP7_75t_L g16929 ( 
.A(n_16839),
.B(n_6696),
.Y(n_16929)
);

NOR2x1_ASAP7_75t_SL g16930 ( 
.A(n_16862),
.B(n_16849),
.Y(n_16930)
);

INVx3_ASAP7_75t_L g16931 ( 
.A(n_16867),
.Y(n_16931)
);

NOR2x1p5_ASAP7_75t_L g16932 ( 
.A(n_16878),
.B(n_5107),
.Y(n_16932)
);

INVx1_ASAP7_75t_L g16933 ( 
.A(n_16886),
.Y(n_16933)
);

NAND3xp33_ASAP7_75t_L g16934 ( 
.A(n_16861),
.B(n_7154),
.C(n_7136),
.Y(n_16934)
);

INVx1_ASAP7_75t_SL g16935 ( 
.A(n_16836),
.Y(n_16935)
);

OR2x2_ASAP7_75t_L g16936 ( 
.A(n_16868),
.B(n_16830),
.Y(n_16936)
);

AND2x4_ASAP7_75t_L g16937 ( 
.A(n_16882),
.B(n_16895),
.Y(n_16937)
);

AND2x2_ASAP7_75t_L g16938 ( 
.A(n_16857),
.B(n_7552),
.Y(n_16938)
);

NAND2x1p5_ASAP7_75t_L g16939 ( 
.A(n_16842),
.B(n_4809),
.Y(n_16939)
);

INVx1_ASAP7_75t_L g16940 ( 
.A(n_16894),
.Y(n_16940)
);

CKINVDCx5p33_ASAP7_75t_R g16941 ( 
.A(n_16860),
.Y(n_16941)
);

NOR2x1p5_ASAP7_75t_L g16942 ( 
.A(n_16848),
.B(n_5107),
.Y(n_16942)
);

AND2x2_ASAP7_75t_L g16943 ( 
.A(n_16838),
.B(n_7552),
.Y(n_16943)
);

NOR2x1_ASAP7_75t_L g16944 ( 
.A(n_16889),
.B(n_7636),
.Y(n_16944)
);

OR2x2_ASAP7_75t_L g16945 ( 
.A(n_16869),
.B(n_16893),
.Y(n_16945)
);

INVx3_ASAP7_75t_L g16946 ( 
.A(n_16875),
.Y(n_16946)
);

NOR2xp33_ASAP7_75t_L g16947 ( 
.A(n_16852),
.B(n_6177),
.Y(n_16947)
);

INVx1_ASAP7_75t_L g16948 ( 
.A(n_16847),
.Y(n_16948)
);

INVx2_ASAP7_75t_L g16949 ( 
.A(n_16853),
.Y(n_16949)
);

INVxp67_ASAP7_75t_SL g16950 ( 
.A(n_16870),
.Y(n_16950)
);

OA22x2_ASAP7_75t_L g16951 ( 
.A1(n_16840),
.A2(n_8146),
.B1(n_7945),
.B2(n_7865),
.Y(n_16951)
);

INVx2_ASAP7_75t_SL g16952 ( 
.A(n_16845),
.Y(n_16952)
);

AND2x2_ASAP7_75t_L g16953 ( 
.A(n_16896),
.B(n_7636),
.Y(n_16953)
);

AND2x2_ASAP7_75t_L g16954 ( 
.A(n_16837),
.B(n_7636),
.Y(n_16954)
);

INVxp67_ASAP7_75t_SL g16955 ( 
.A(n_16821),
.Y(n_16955)
);

AND2x4_ASAP7_75t_L g16956 ( 
.A(n_16825),
.B(n_6696),
.Y(n_16956)
);

OR2x2_ASAP7_75t_L g16957 ( 
.A(n_16887),
.B(n_7636),
.Y(n_16957)
);

NAND4xp75_ASAP7_75t_L g16958 ( 
.A(n_16880),
.B(n_6940),
.C(n_6956),
.D(n_6930),
.Y(n_16958)
);

NOR3xp33_ASAP7_75t_SL g16959 ( 
.A(n_16841),
.B(n_6909),
.C(n_6908),
.Y(n_16959)
);

AOI22xp5_ASAP7_75t_L g16960 ( 
.A1(n_16824),
.A2(n_6783),
.B1(n_7111),
.B2(n_6267),
.Y(n_16960)
);

O2A1O1Ixp33_ASAP7_75t_L g16961 ( 
.A1(n_16897),
.A2(n_16890),
.B(n_16846),
.C(n_16843),
.Y(n_16961)
);

INVx3_ASAP7_75t_L g16962 ( 
.A(n_16901),
.Y(n_16962)
);

NOR3xp33_ASAP7_75t_L g16963 ( 
.A(n_16909),
.B(n_16873),
.C(n_5811),
.Y(n_16963)
);

NOR2x2_ASAP7_75t_L g16964 ( 
.A(n_16903),
.B(n_7636),
.Y(n_16964)
);

NAND4xp25_ASAP7_75t_L g16965 ( 
.A(n_16906),
.B(n_4303),
.C(n_4308),
.D(n_4278),
.Y(n_16965)
);

AND2x4_ASAP7_75t_L g16966 ( 
.A(n_16913),
.B(n_6635),
.Y(n_16966)
);

NAND2xp5_ASAP7_75t_SL g16967 ( 
.A(n_16925),
.B(n_6215),
.Y(n_16967)
);

NAND2xp5_ASAP7_75t_SL g16968 ( 
.A(n_16905),
.B(n_6215),
.Y(n_16968)
);

NAND2xp5_ASAP7_75t_L g16969 ( 
.A(n_16935),
.B(n_7089),
.Y(n_16969)
);

NOR4xp75_ASAP7_75t_L g16970 ( 
.A(n_16900),
.B(n_16931),
.C(n_16946),
.D(n_16904),
.Y(n_16970)
);

NAND2xp5_ASAP7_75t_L g16971 ( 
.A(n_16914),
.B(n_7089),
.Y(n_16971)
);

AND2x2_ASAP7_75t_L g16972 ( 
.A(n_16907),
.B(n_7636),
.Y(n_16972)
);

OAI211xp5_ASAP7_75t_SL g16973 ( 
.A1(n_16926),
.A2(n_6917),
.B(n_6925),
.C(n_6909),
.Y(n_16973)
);

INVx2_ASAP7_75t_L g16974 ( 
.A(n_16940),
.Y(n_16974)
);

INVx2_ASAP7_75t_L g16975 ( 
.A(n_16936),
.Y(n_16975)
);

NAND5xp2_ASAP7_75t_L g16976 ( 
.A(n_16955),
.B(n_5611),
.C(n_5649),
.D(n_5637),
.E(n_5549),
.Y(n_16976)
);

NAND3xp33_ASAP7_75t_SL g16977 ( 
.A(n_16933),
.B(n_5811),
.C(n_5795),
.Y(n_16977)
);

NOR2xp67_ASAP7_75t_L g16978 ( 
.A(n_16937),
.B(n_4809),
.Y(n_16978)
);

AND2x4_ASAP7_75t_L g16979 ( 
.A(n_16916),
.B(n_8146),
.Y(n_16979)
);

NAND2xp5_ASAP7_75t_L g16980 ( 
.A(n_16928),
.B(n_7089),
.Y(n_16980)
);

NOR3xp33_ASAP7_75t_L g16981 ( 
.A(n_16949),
.B(n_5811),
.C(n_5795),
.Y(n_16981)
);

AND2x4_ASAP7_75t_L g16982 ( 
.A(n_16938),
.B(n_6635),
.Y(n_16982)
);

AOI22xp33_ASAP7_75t_L g16983 ( 
.A1(n_16919),
.A2(n_7129),
.B1(n_7128),
.B2(n_7136),
.Y(n_16983)
);

NAND4xp75_ASAP7_75t_L g16984 ( 
.A(n_16918),
.B(n_5020),
.C(n_5045),
.D(n_4947),
.Y(n_16984)
);

NOR3xp33_ASAP7_75t_SL g16985 ( 
.A(n_16941),
.B(n_6917),
.C(n_6909),
.Y(n_16985)
);

NOR4xp25_ASAP7_75t_L g16986 ( 
.A(n_16922),
.B(n_6925),
.C(n_6928),
.D(n_6917),
.Y(n_16986)
);

INVx1_ASAP7_75t_L g16987 ( 
.A(n_16948),
.Y(n_16987)
);

OAI211xp5_ASAP7_75t_SL g16988 ( 
.A1(n_16950),
.A2(n_6928),
.B(n_6929),
.C(n_6925),
.Y(n_16988)
);

AND2x2_ASAP7_75t_L g16989 ( 
.A(n_16921),
.B(n_7636),
.Y(n_16989)
);

NAND5xp2_ASAP7_75t_L g16990 ( 
.A(n_16959),
.B(n_5649),
.C(n_5677),
.D(n_5653),
.E(n_5637),
.Y(n_16990)
);

NAND4xp25_ASAP7_75t_SL g16991 ( 
.A(n_16945),
.B(n_16899),
.C(n_16944),
.D(n_16910),
.Y(n_16991)
);

NOR2x1_ASAP7_75t_L g16992 ( 
.A(n_16898),
.B(n_7776),
.Y(n_16992)
);

OR2x2_ASAP7_75t_L g16993 ( 
.A(n_16911),
.B(n_7776),
.Y(n_16993)
);

AOI211xp5_ASAP7_75t_L g16994 ( 
.A1(n_16952),
.A2(n_7129),
.B(n_7128),
.C(n_7136),
.Y(n_16994)
);

NAND4xp75_ASAP7_75t_L g16995 ( 
.A(n_16908),
.B(n_5020),
.C(n_5045),
.D(n_4947),
.Y(n_16995)
);

NAND4xp25_ASAP7_75t_L g16996 ( 
.A(n_16954),
.B(n_4303),
.C(n_4308),
.D(n_4278),
.Y(n_16996)
);

NAND3xp33_ASAP7_75t_SL g16997 ( 
.A(n_16939),
.B(n_5811),
.C(n_5795),
.Y(n_16997)
);

CKINVDCx5p33_ASAP7_75t_R g16998 ( 
.A(n_16942),
.Y(n_16998)
);

NAND3xp33_ASAP7_75t_SL g16999 ( 
.A(n_16947),
.B(n_5818),
.C(n_5813),
.Y(n_16999)
);

INVx2_ASAP7_75t_L g17000 ( 
.A(n_16930),
.Y(n_17000)
);

NOR4xp25_ASAP7_75t_L g17001 ( 
.A(n_16912),
.B(n_6929),
.C(n_6955),
.D(n_6928),
.Y(n_17001)
);

INVx1_ASAP7_75t_L g17002 ( 
.A(n_16932),
.Y(n_17002)
);

NOR3x1_ASAP7_75t_L g17003 ( 
.A(n_16924),
.B(n_7945),
.C(n_7827),
.Y(n_17003)
);

AND3x1_ASAP7_75t_L g17004 ( 
.A(n_16953),
.B(n_6736),
.C(n_6713),
.Y(n_17004)
);

NAND4xp25_ASAP7_75t_L g17005 ( 
.A(n_16957),
.B(n_4303),
.C(n_4308),
.D(n_4278),
.Y(n_17005)
);

O2A1O1Ixp33_ASAP7_75t_L g17006 ( 
.A1(n_16943),
.A2(n_7949),
.B(n_8097),
.C(n_7776),
.Y(n_17006)
);

INVx3_ASAP7_75t_L g17007 ( 
.A(n_16929),
.Y(n_17007)
);

NAND3xp33_ASAP7_75t_L g17008 ( 
.A(n_16915),
.B(n_5188),
.C(n_7154),
.Y(n_17008)
);

AND2x4_ASAP7_75t_L g17009 ( 
.A(n_16956),
.B(n_6635),
.Y(n_17009)
);

NOR2x1_ASAP7_75t_L g17010 ( 
.A(n_16902),
.B(n_7776),
.Y(n_17010)
);

OR4x1_ASAP7_75t_L g17011 ( 
.A(n_16917),
.B(n_6955),
.C(n_6958),
.D(n_6929),
.Y(n_17011)
);

AND2x2_ASAP7_75t_SL g17012 ( 
.A(n_16960),
.B(n_4961),
.Y(n_17012)
);

OAI22xp5_ASAP7_75t_L g17013 ( 
.A1(n_16958),
.A2(n_6783),
.B1(n_7151),
.B2(n_7154),
.Y(n_17013)
);

AOI211xp5_ASAP7_75t_L g17014 ( 
.A1(n_16927),
.A2(n_7129),
.B(n_7128),
.C(n_7154),
.Y(n_17014)
);

OAI211xp5_ASAP7_75t_SL g17015 ( 
.A1(n_16934),
.A2(n_16923),
.B(n_16920),
.C(n_16951),
.Y(n_17015)
);

NOR4xp25_ASAP7_75t_L g17016 ( 
.A(n_16897),
.B(n_6958),
.C(n_6963),
.D(n_6955),
.Y(n_17016)
);

NOR3xp33_ASAP7_75t_L g17017 ( 
.A(n_16897),
.B(n_5818),
.C(n_5813),
.Y(n_17017)
);

NAND3xp33_ASAP7_75t_L g17018 ( 
.A(n_16897),
.B(n_7129),
.C(n_7128),
.Y(n_17018)
);

OR2x2_ASAP7_75t_L g17019 ( 
.A(n_16974),
.B(n_7949),
.Y(n_17019)
);

INVxp67_ASAP7_75t_SL g17020 ( 
.A(n_16962),
.Y(n_17020)
);

OAI211xp5_ASAP7_75t_SL g17021 ( 
.A1(n_17000),
.A2(n_6963),
.B(n_6968),
.C(n_6958),
.Y(n_17021)
);

AOI21xp5_ASAP7_75t_L g17022 ( 
.A1(n_16975),
.A2(n_7137),
.B(n_7026),
.Y(n_17022)
);

INVx1_ASAP7_75t_L g17023 ( 
.A(n_16970),
.Y(n_17023)
);

OAI31xp33_ASAP7_75t_L g17024 ( 
.A1(n_16987),
.A2(n_6134),
.A3(n_5854),
.B(n_5880),
.Y(n_17024)
);

INVx1_ASAP7_75t_L g17025 ( 
.A(n_17007),
.Y(n_17025)
);

NAND2xp5_ASAP7_75t_L g17026 ( 
.A(n_16998),
.B(n_7089),
.Y(n_17026)
);

NAND5xp2_ASAP7_75t_L g17027 ( 
.A(n_17002),
.B(n_5734),
.C(n_5737),
.D(n_5677),
.E(n_5653),
.Y(n_17027)
);

NOR2x1p5_ASAP7_75t_L g17028 ( 
.A(n_16980),
.B(n_16971),
.Y(n_17028)
);

AOI211xp5_ASAP7_75t_L g17029 ( 
.A1(n_16991),
.A2(n_7129),
.B(n_7128),
.C(n_7945),
.Y(n_17029)
);

AND3x4_ASAP7_75t_L g17030 ( 
.A(n_16963),
.B(n_4320),
.C(n_4303),
.Y(n_17030)
);

NOR2xp33_ASAP7_75t_L g17031 ( 
.A(n_16968),
.B(n_7128),
.Y(n_17031)
);

AOI211xp5_ASAP7_75t_L g17032 ( 
.A1(n_16961),
.A2(n_17015),
.B(n_16969),
.C(n_16967),
.Y(n_17032)
);

OA22x2_ASAP7_75t_L g17033 ( 
.A1(n_16966),
.A2(n_7822),
.B1(n_7526),
.B2(n_7530),
.Y(n_17033)
);

OAI22xp5_ASAP7_75t_SL g17034 ( 
.A1(n_17012),
.A2(n_7151),
.B1(n_6097),
.B2(n_4915),
.Y(n_17034)
);

NOR2x1p5_ASAP7_75t_L g17035 ( 
.A(n_16996),
.B(n_4278),
.Y(n_17035)
);

AOI21xp5_ASAP7_75t_L g17036 ( 
.A1(n_16993),
.A2(n_16989),
.B(n_17004),
.Y(n_17036)
);

OAI22xp5_ASAP7_75t_L g17037 ( 
.A1(n_16983),
.A2(n_7151),
.B1(n_7129),
.B2(n_7128),
.Y(n_17037)
);

INVx1_ASAP7_75t_L g17038 ( 
.A(n_16982),
.Y(n_17038)
);

NAND2xp5_ASAP7_75t_L g17039 ( 
.A(n_16972),
.B(n_7089),
.Y(n_17039)
);

NOR4xp25_ASAP7_75t_L g17040 ( 
.A(n_17005),
.B(n_6968),
.C(n_6969),
.D(n_6963),
.Y(n_17040)
);

INVx1_ASAP7_75t_L g17041 ( 
.A(n_17009),
.Y(n_17041)
);

INVx1_ASAP7_75t_L g17042 ( 
.A(n_17009),
.Y(n_17042)
);

AND2x4_ASAP7_75t_L g17043 ( 
.A(n_17008),
.B(n_16981),
.Y(n_17043)
);

AOI22xp33_ASAP7_75t_SL g17044 ( 
.A1(n_17018),
.A2(n_7137),
.B1(n_7151),
.B2(n_7129),
.Y(n_17044)
);

NAND5xp2_ASAP7_75t_L g17045 ( 
.A(n_17017),
.B(n_5806),
.C(n_5842),
.D(n_5737),
.E(n_5734),
.Y(n_17045)
);

NOR4xp25_ASAP7_75t_L g17046 ( 
.A(n_16997),
.B(n_6969),
.C(n_6973),
.D(n_6968),
.Y(n_17046)
);

INVx1_ASAP7_75t_L g17047 ( 
.A(n_16985),
.Y(n_17047)
);

NOR4xp25_ASAP7_75t_L g17048 ( 
.A(n_16965),
.B(n_6973),
.C(n_6974),
.D(n_6969),
.Y(n_17048)
);

AND2x4_ASAP7_75t_L g17049 ( 
.A(n_16992),
.B(n_6695),
.Y(n_17049)
);

NOR3xp33_ASAP7_75t_L g17050 ( 
.A(n_16990),
.B(n_5818),
.C(n_5813),
.Y(n_17050)
);

AOI21xp5_ASAP7_75t_L g17051 ( 
.A1(n_16978),
.A2(n_7137),
.B(n_4965),
.Y(n_17051)
);

NOR3xp33_ASAP7_75t_L g17052 ( 
.A(n_16999),
.B(n_5818),
.C(n_5813),
.Y(n_17052)
);

AOI221xp5_ASAP7_75t_L g17053 ( 
.A1(n_17001),
.A2(n_7128),
.B1(n_6192),
.B2(n_6250),
.C(n_6179),
.Y(n_17053)
);

NAND4xp25_ASAP7_75t_L g17054 ( 
.A(n_16976),
.B(n_4320),
.C(n_4324),
.D(n_4308),
.Y(n_17054)
);

OAI221xp5_ASAP7_75t_R g17055 ( 
.A1(n_17011),
.A2(n_6640),
.B1(n_6516),
.B2(n_6135),
.C(n_7822),
.Y(n_17055)
);

INVx2_ASAP7_75t_L g17056 ( 
.A(n_16964),
.Y(n_17056)
);

NAND2xp5_ASAP7_75t_L g17057 ( 
.A(n_16995),
.B(n_7089),
.Y(n_17057)
);

AOI22xp5_ASAP7_75t_L g17058 ( 
.A1(n_17010),
.A2(n_17014),
.B1(n_16977),
.B2(n_16994),
.Y(n_17058)
);

NOR3xp33_ASAP7_75t_SL g17059 ( 
.A(n_16988),
.B(n_6974),
.C(n_6973),
.Y(n_17059)
);

OAI222xp33_ASAP7_75t_L g17060 ( 
.A1(n_16979),
.A2(n_8121),
.B1(n_7949),
.B2(n_8169),
.C1(n_8097),
.C2(n_7776),
.Y(n_17060)
);

OAI21xp5_ASAP7_75t_L g17061 ( 
.A1(n_16984),
.A2(n_8036),
.B(n_8031),
.Y(n_17061)
);

OAI21xp33_ASAP7_75t_L g17062 ( 
.A1(n_16986),
.A2(n_5200),
.B(n_5196),
.Y(n_17062)
);

AOI22xp5_ASAP7_75t_L g17063 ( 
.A1(n_16979),
.A2(n_7111),
.B1(n_7151),
.B2(n_6177),
.Y(n_17063)
);

CKINVDCx20_ASAP7_75t_R g17064 ( 
.A(n_17023),
.Y(n_17064)
);

INVx1_ASAP7_75t_L g17065 ( 
.A(n_17020),
.Y(n_17065)
);

OAI22xp33_ASAP7_75t_R g17066 ( 
.A1(n_17025),
.A2(n_17003),
.B1(n_17006),
.B2(n_16973),
.Y(n_17066)
);

INVx2_ASAP7_75t_L g17067 ( 
.A(n_17056),
.Y(n_17067)
);

NOR2x1_ASAP7_75t_L g17068 ( 
.A(n_17041),
.B(n_17013),
.Y(n_17068)
);

INVx3_ASAP7_75t_L g17069 ( 
.A(n_17042),
.Y(n_17069)
);

OAI21xp33_ASAP7_75t_L g17070 ( 
.A1(n_17038),
.A2(n_17016),
.B(n_7949),
.Y(n_17070)
);

INVx1_ASAP7_75t_L g17071 ( 
.A(n_17047),
.Y(n_17071)
);

INVx2_ASAP7_75t_L g17072 ( 
.A(n_17028),
.Y(n_17072)
);

OR2x6_ASAP7_75t_L g17073 ( 
.A(n_17036),
.B(n_4320),
.Y(n_17073)
);

INVx1_ASAP7_75t_L g17074 ( 
.A(n_17032),
.Y(n_17074)
);

OAI22x1_ASAP7_75t_L g17075 ( 
.A1(n_17058),
.A2(n_4894),
.B1(n_4955),
.B2(n_4809),
.Y(n_17075)
);

NOR2xp67_ASAP7_75t_L g17076 ( 
.A(n_17043),
.B(n_4894),
.Y(n_17076)
);

BUFx2_ASAP7_75t_L g17077 ( 
.A(n_17049),
.Y(n_17077)
);

INVx1_ASAP7_75t_L g17078 ( 
.A(n_17026),
.Y(n_17078)
);

OAI22x1_ASAP7_75t_L g17079 ( 
.A1(n_17030),
.A2(n_4955),
.B1(n_4894),
.B2(n_6974),
.Y(n_17079)
);

A2O1A1Ixp33_ASAP7_75t_L g17080 ( 
.A1(n_17022),
.A2(n_7621),
.B(n_7851),
.C(n_7828),
.Y(n_17080)
);

OAI211xp5_ASAP7_75t_SL g17081 ( 
.A1(n_17039),
.A2(n_6736),
.B(n_6770),
.C(n_6765),
.Y(n_17081)
);

NOR4xp75_ASAP7_75t_L g17082 ( 
.A(n_17057),
.B(n_6736),
.C(n_6770),
.D(n_6765),
.Y(n_17082)
);

CKINVDCx20_ASAP7_75t_R g17083 ( 
.A(n_17059),
.Y(n_17083)
);

AOI22x1_ASAP7_75t_L g17084 ( 
.A1(n_17035),
.A2(n_5818),
.B1(n_5885),
.B2(n_5813),
.Y(n_17084)
);

INVx1_ASAP7_75t_L g17085 ( 
.A(n_17031),
.Y(n_17085)
);

NOR4xp25_ASAP7_75t_L g17086 ( 
.A(n_17054),
.B(n_6991),
.C(n_6994),
.D(n_6977),
.Y(n_17086)
);

NOR2x1_ASAP7_75t_L g17087 ( 
.A(n_17045),
.B(n_7776),
.Y(n_17087)
);

O2A1O1Ixp33_ASAP7_75t_L g17088 ( 
.A1(n_17050),
.A2(n_7949),
.B(n_8097),
.C(n_7776),
.Y(n_17088)
);

AND2x2_ASAP7_75t_L g17089 ( 
.A(n_17040),
.B(n_8097),
.Y(n_17089)
);

AOI21xp5_ASAP7_75t_L g17090 ( 
.A1(n_17051),
.A2(n_4961),
.B(n_4965),
.Y(n_17090)
);

NAND2xp5_ASAP7_75t_L g17091 ( 
.A(n_17048),
.B(n_8097),
.Y(n_17091)
);

INVx1_ASAP7_75t_L g17092 ( 
.A(n_17052),
.Y(n_17092)
);

INVx1_ASAP7_75t_L g17093 ( 
.A(n_17037),
.Y(n_17093)
);

NAND2xp5_ASAP7_75t_L g17094 ( 
.A(n_17046),
.B(n_8097),
.Y(n_17094)
);

INVx2_ASAP7_75t_L g17095 ( 
.A(n_17019),
.Y(n_17095)
);

NAND2xp5_ASAP7_75t_L g17096 ( 
.A(n_17062),
.B(n_8097),
.Y(n_17096)
);

HB1xp67_ASAP7_75t_L g17097 ( 
.A(n_17034),
.Y(n_17097)
);

XNOR2x1_ASAP7_75t_L g17098 ( 
.A(n_17055),
.B(n_8121),
.Y(n_17098)
);

AOI22xp5_ASAP7_75t_L g17099 ( 
.A1(n_17044),
.A2(n_17021),
.B1(n_17063),
.B2(n_17053),
.Y(n_17099)
);

NAND5xp2_ASAP7_75t_L g17100 ( 
.A(n_17024),
.B(n_5889),
.C(n_5920),
.D(n_5842),
.E(n_5806),
.Y(n_17100)
);

NOR2x1p5_ASAP7_75t_L g17101 ( 
.A(n_17027),
.B(n_4320),
.Y(n_17101)
);

INVx1_ASAP7_75t_L g17102 ( 
.A(n_17061),
.Y(n_17102)
);

INVx1_ASAP7_75t_SL g17103 ( 
.A(n_17033),
.Y(n_17103)
);

AOI22xp5_ASAP7_75t_L g17104 ( 
.A1(n_17064),
.A2(n_17029),
.B1(n_17060),
.B2(n_7111),
.Y(n_17104)
);

INVx2_ASAP7_75t_L g17105 ( 
.A(n_17065),
.Y(n_17105)
);

XOR2xp5_ASAP7_75t_L g17106 ( 
.A(n_17074),
.B(n_4942),
.Y(n_17106)
);

INVx2_ASAP7_75t_L g17107 ( 
.A(n_17072),
.Y(n_17107)
);

INVx1_ASAP7_75t_L g17108 ( 
.A(n_17069),
.Y(n_17108)
);

INVx1_ASAP7_75t_L g17109 ( 
.A(n_17077),
.Y(n_17109)
);

INVx1_ASAP7_75t_L g17110 ( 
.A(n_17067),
.Y(n_17110)
);

INVx2_ASAP7_75t_L g17111 ( 
.A(n_17083),
.Y(n_17111)
);

INVx1_ASAP7_75t_L g17112 ( 
.A(n_17071),
.Y(n_17112)
);

AOI22xp33_ASAP7_75t_L g17113 ( 
.A1(n_17095),
.A2(n_6179),
.B1(n_6192),
.B2(n_6177),
.Y(n_17113)
);

INVx1_ASAP7_75t_L g17114 ( 
.A(n_17068),
.Y(n_17114)
);

INVx2_ASAP7_75t_L g17115 ( 
.A(n_17103),
.Y(n_17115)
);

OR3x1_ASAP7_75t_L g17116 ( 
.A(n_17085),
.B(n_6991),
.C(n_6977),
.Y(n_17116)
);

INVx1_ASAP7_75t_L g17117 ( 
.A(n_17097),
.Y(n_17117)
);

XNOR2xp5_ASAP7_75t_SL g17118 ( 
.A(n_17078),
.B(n_4942),
.Y(n_17118)
);

XOR2xp5_ASAP7_75t_L g17119 ( 
.A(n_17102),
.B(n_4942),
.Y(n_17119)
);

XNOR2x1_ASAP7_75t_L g17120 ( 
.A(n_17093),
.B(n_17092),
.Y(n_17120)
);

INVx1_ASAP7_75t_L g17121 ( 
.A(n_17066),
.Y(n_17121)
);

INVx1_ASAP7_75t_L g17122 ( 
.A(n_17099),
.Y(n_17122)
);

INVx1_ASAP7_75t_L g17123 ( 
.A(n_17098),
.Y(n_17123)
);

INVx1_ASAP7_75t_L g17124 ( 
.A(n_17073),
.Y(n_17124)
);

INVx1_ASAP7_75t_L g17125 ( 
.A(n_17073),
.Y(n_17125)
);

INVx1_ASAP7_75t_L g17126 ( 
.A(n_17101),
.Y(n_17126)
);

INVx2_ASAP7_75t_L g17127 ( 
.A(n_17114),
.Y(n_17127)
);

INVxp67_ASAP7_75t_L g17128 ( 
.A(n_17108),
.Y(n_17128)
);

OAI22xp33_ASAP7_75t_L g17129 ( 
.A1(n_17109),
.A2(n_17091),
.B1(n_17094),
.B2(n_17096),
.Y(n_17129)
);

AND2x2_ASAP7_75t_L g17130 ( 
.A(n_17110),
.B(n_17089),
.Y(n_17130)
);

AND2x2_ASAP7_75t_L g17131 ( 
.A(n_17105),
.B(n_17087),
.Y(n_17131)
);

INVx1_ASAP7_75t_L g17132 ( 
.A(n_17112),
.Y(n_17132)
);

INVx1_ASAP7_75t_L g17133 ( 
.A(n_17117),
.Y(n_17133)
);

CKINVDCx20_ASAP7_75t_R g17134 ( 
.A(n_17122),
.Y(n_17134)
);

AO21x2_ASAP7_75t_L g17135 ( 
.A1(n_17107),
.A2(n_17090),
.B(n_17070),
.Y(n_17135)
);

NAND3xp33_ASAP7_75t_L g17136 ( 
.A(n_17120),
.B(n_17115),
.C(n_17121),
.Y(n_17136)
);

NOR2xp33_ASAP7_75t_L g17137 ( 
.A(n_17111),
.B(n_17100),
.Y(n_17137)
);

XOR2xp5_ASAP7_75t_L g17138 ( 
.A(n_17123),
.B(n_17079),
.Y(n_17138)
);

INVx2_ASAP7_75t_L g17139 ( 
.A(n_17126),
.Y(n_17139)
);

INVx4_ASAP7_75t_L g17140 ( 
.A(n_17124),
.Y(n_17140)
);

AND2x2_ASAP7_75t_SL g17141 ( 
.A(n_17125),
.B(n_17086),
.Y(n_17141)
);

OR2x2_ASAP7_75t_L g17142 ( 
.A(n_17133),
.B(n_17106),
.Y(n_17142)
);

NOR3xp33_ASAP7_75t_SL g17143 ( 
.A(n_17136),
.B(n_17118),
.C(n_17104),
.Y(n_17143)
);

OR2x2_ASAP7_75t_L g17144 ( 
.A(n_17127),
.B(n_17119),
.Y(n_17144)
);

INVx2_ASAP7_75t_L g17145 ( 
.A(n_17134),
.Y(n_17145)
);

OAI221xp5_ASAP7_75t_L g17146 ( 
.A1(n_17128),
.A2(n_17076),
.B1(n_17088),
.B2(n_17084),
.C(n_17081),
.Y(n_17146)
);

OR2x2_ASAP7_75t_L g17147 ( 
.A(n_17132),
.B(n_17113),
.Y(n_17147)
);

INVx1_ASAP7_75t_L g17148 ( 
.A(n_17140),
.Y(n_17148)
);

AOI22xp5_ASAP7_75t_L g17149 ( 
.A1(n_17131),
.A2(n_17116),
.B1(n_17082),
.B2(n_17075),
.Y(n_17149)
);

INVx3_ASAP7_75t_L g17150 ( 
.A(n_17139),
.Y(n_17150)
);

OR3x1_ASAP7_75t_L g17151 ( 
.A(n_17137),
.B(n_17080),
.C(n_6994),
.Y(n_17151)
);

AOI22xp5_ASAP7_75t_L g17152 ( 
.A1(n_17130),
.A2(n_8169),
.B1(n_8185),
.B2(n_8121),
.Y(n_17152)
);

NAND3x1_ASAP7_75t_L g17153 ( 
.A(n_17141),
.B(n_17138),
.C(n_17129),
.Y(n_17153)
);

NOR4xp25_ASAP7_75t_SL g17154 ( 
.A(n_17135),
.B(n_5920),
.C(n_5960),
.D(n_5889),
.Y(n_17154)
);

OAI22xp5_ASAP7_75t_SL g17155 ( 
.A1(n_17145),
.A2(n_4988),
.B1(n_4915),
.B2(n_6097),
.Y(n_17155)
);

INVx1_ASAP7_75t_L g17156 ( 
.A(n_17150),
.Y(n_17156)
);

INVx2_ASAP7_75t_SL g17157 ( 
.A(n_17148),
.Y(n_17157)
);

OAI22xp5_ASAP7_75t_L g17158 ( 
.A1(n_17153),
.A2(n_8169),
.B1(n_8185),
.B2(n_8121),
.Y(n_17158)
);

BUFx2_ASAP7_75t_L g17159 ( 
.A(n_17143),
.Y(n_17159)
);

INVx1_ASAP7_75t_SL g17160 ( 
.A(n_17144),
.Y(n_17160)
);

INVx2_ASAP7_75t_L g17161 ( 
.A(n_17142),
.Y(n_17161)
);

AO22x2_ASAP7_75t_L g17162 ( 
.A1(n_17147),
.A2(n_6991),
.B1(n_6994),
.B2(n_6977),
.Y(n_17162)
);

INVx1_ASAP7_75t_L g17163 ( 
.A(n_17156),
.Y(n_17163)
);

NOR2x1p5_ASAP7_75t_L g17164 ( 
.A(n_17161),
.B(n_17149),
.Y(n_17164)
);

BUFx2_ASAP7_75t_L g17165 ( 
.A(n_17157),
.Y(n_17165)
);

XNOR2xp5_ASAP7_75t_L g17166 ( 
.A(n_17160),
.B(n_17146),
.Y(n_17166)
);

NAND2xp5_ASAP7_75t_SL g17167 ( 
.A(n_17159),
.B(n_17151),
.Y(n_17167)
);

AOI22xp33_ASAP7_75t_L g17168 ( 
.A1(n_17155),
.A2(n_17154),
.B1(n_17152),
.B2(n_8169),
.Y(n_17168)
);

OAI22xp5_ASAP7_75t_SL g17169 ( 
.A1(n_17165),
.A2(n_17158),
.B1(n_17162),
.B2(n_4988),
.Y(n_17169)
);

INVx3_ASAP7_75t_SL g17170 ( 
.A(n_17167),
.Y(n_17170)
);

AOI21xp5_ASAP7_75t_L g17171 ( 
.A1(n_17163),
.A2(n_17162),
.B(n_4965),
.Y(n_17171)
);

AOI21xp5_ASAP7_75t_L g17172 ( 
.A1(n_17166),
.A2(n_4965),
.B(n_4961),
.Y(n_17172)
);

AOI21xp5_ASAP7_75t_L g17173 ( 
.A1(n_17170),
.A2(n_17164),
.B(n_17168),
.Y(n_17173)
);

OAI21x1_ASAP7_75t_SL g17174 ( 
.A1(n_17171),
.A2(n_5055),
.B(n_5045),
.Y(n_17174)
);

NOR2xp33_ASAP7_75t_L g17175 ( 
.A(n_17173),
.B(n_17169),
.Y(n_17175)
);

AOI21xp33_ASAP7_75t_SL g17176 ( 
.A1(n_17175),
.A2(n_17174),
.B(n_17172),
.Y(n_17176)
);

INVxp67_ASAP7_75t_L g17177 ( 
.A(n_17176),
.Y(n_17177)
);

AOI21xp5_ASAP7_75t_SL g17178 ( 
.A1(n_17177),
.A2(n_4590),
.B(n_4563),
.Y(n_17178)
);

OAI221xp5_ASAP7_75t_R g17179 ( 
.A1(n_17178),
.A2(n_6135),
.B1(n_6640),
.B2(n_6516),
.C(n_7575),
.Y(n_17179)
);

AOI21xp33_ASAP7_75t_L g17180 ( 
.A1(n_17179),
.A2(n_6179),
.B(n_6177),
.Y(n_17180)
);

AOI22xp5_ASAP7_75t_L g17181 ( 
.A1(n_17180),
.A2(n_4274),
.B1(n_7111),
.B2(n_4590),
.Y(n_17181)
);


endmodule