module fake_jpeg_21204_n_301 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_14),
.B(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_7),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_1),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_15),
.C(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_14),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_32),
.A2(n_29),
.B1(n_31),
.B2(n_27),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_51),
.B1(n_54),
.B2(n_35),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_36),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_28),
.B1(n_23),
.B2(n_26),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_32),
.A2(n_28),
.B1(n_16),
.B2(n_27),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_59),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_65),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_71),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_37),
.C(n_39),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_77),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_74),
.B1(n_75),
.B2(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_73),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_35),
.B1(n_36),
.B2(n_34),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_39),
.B(n_33),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_37),
.Y(n_77)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_52),
.A2(n_34),
.B1(n_53),
.B2(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_37),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_84),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_44),
.B1(n_17),
.B2(n_26),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_88),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_70),
.B1(n_81),
.B2(n_75),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_102),
.B1(n_107),
.B2(n_76),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_91),
.B(n_97),
.Y(n_128)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_53),
.B1(n_50),
.B2(n_52),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_105),
.B1(n_83),
.B2(n_66),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_60),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_SL g100 ( 
.A1(n_71),
.A2(n_16),
.B(n_22),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_22),
.B(n_20),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_52),
.B1(n_39),
.B2(n_17),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_40),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_52),
.B1(n_28),
.B2(n_25),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_68),
.A2(n_42),
.B1(n_33),
.B2(n_40),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_76),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_126),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_114),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_115),
.A2(n_129),
.B1(n_88),
.B2(n_106),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_77),
.C(n_46),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_125),
.C(n_136),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_77),
.B1(n_61),
.B2(n_73),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_118),
.B1(n_133),
.B2(n_140),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_17),
.B1(n_26),
.B2(n_25),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_41),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_121),
.B(n_123),
.Y(n_167)
);

NOR3xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_19),
.C(n_23),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_19),
.Y(n_123)
);

NOR2xp67_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_104),
.Y(n_124)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_124),
.A2(n_135),
.B(n_109),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_42),
.C(n_40),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_72),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_15),
.Y(n_127)
);

FAx1_ASAP7_75t_SL g168 ( 
.A(n_127),
.B(n_131),
.CI(n_134),
.CON(n_168),
.SN(n_168)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_42),
.B1(n_28),
.B2(n_40),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_18),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_58),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_90),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_98),
.A2(n_40),
.B1(n_41),
.B2(n_55),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_98),
.B(n_16),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_16),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_111),
.A2(n_25),
.B1(n_20),
.B2(n_27),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_108),
.A2(n_111),
.B1(n_88),
.B2(n_86),
.Y(n_140)
);

OAI32xp33_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_86),
.A3(n_90),
.B1(n_20),
.B2(n_31),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_141),
.B(n_159),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_109),
.B(n_22),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_139),
.B(n_121),
.Y(n_172)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_146),
.B(n_156),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_120),
.A2(n_85),
.B1(n_137),
.B2(n_138),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_84),
.B1(n_63),
.B2(n_78),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_155),
.Y(n_191)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_128),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_16),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_160),
.B(n_161),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_130),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_16),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_169),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_127),
.B1(n_134),
.B2(n_106),
.Y(n_175)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_164),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_106),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_165),
.B(n_166),
.Y(n_194)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_30),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_96),
.C(n_93),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_96),
.C(n_78),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_30),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_172),
.A2(n_187),
.B1(n_190),
.B2(n_141),
.Y(n_203)
);

FAx1_ASAP7_75t_SL g173 ( 
.A(n_169),
.B(n_131),
.CI(n_154),
.CON(n_173),
.SN(n_173)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_179),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_167),
.B(n_127),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_175),
.A2(n_177),
.B1(n_183),
.B2(n_184),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_119),
.B1(n_85),
.B2(n_94),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_178),
.B(n_195),
.Y(n_221)
);

AOI32xp33_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_79),
.A3(n_78),
.B1(n_30),
.B2(n_57),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_182),
.A2(n_199),
.B1(n_147),
.B2(n_160),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_145),
.A2(n_30),
.B1(n_21),
.B2(n_24),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_41),
.B1(n_63),
.B2(n_10),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_157),
.A2(n_30),
.B(n_10),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_165),
.B(n_143),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_192),
.B(n_1),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_41),
.C(n_18),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_156),
.B(n_30),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_200),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_21),
.B1(n_24),
.B2(n_18),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_198),
.A2(n_153),
.B1(n_148),
.B2(n_168),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_142),
.A2(n_24),
.B1(n_21),
.B2(n_18),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_146),
.B(n_18),
.C(n_15),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_18),
.C(n_21),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_170),
.Y(n_205)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_217),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_203),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_186),
.C(n_195),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_185),
.A2(n_159),
.B1(n_149),
.B2(n_142),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_206),
.A2(n_213),
.B1(n_13),
.B2(n_12),
.Y(n_239)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

XOR2x1_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_168),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_208),
.A2(n_209),
.B1(n_223),
.B2(n_172),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_178),
.A2(n_158),
.B1(n_168),
.B2(n_149),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_196),
.Y(n_233)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

NAND3xp33_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_148),
.C(n_153),
.Y(n_216)
);

OA21x2_ASAP7_75t_SL g230 ( 
.A1(n_216),
.A2(n_192),
.B(n_187),
.Y(n_230)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_219),
.Y(n_241)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_222),
.Y(n_240)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_218),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_234),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_186),
.C(n_173),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_231),
.C(n_238),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_204),
.B1(n_13),
.B2(n_12),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_173),
.C(n_193),
.Y(n_231)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_214),
.A2(n_199),
.B1(n_177),
.B2(n_175),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_235),
.A2(n_236),
.B1(n_213),
.B2(n_209),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_197),
.B1(n_193),
.B2(n_184),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_200),
.C(n_201),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_12),
.B1(n_10),
.B2(n_3),
.Y(n_252)
);

FAx1_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_208),
.CI(n_218),
.CON(n_244),
.SN(n_244)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_245),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_240),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_249),
.B1(n_228),
.B2(n_225),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_203),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_253),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_235),
.A2(n_204),
.B1(n_223),
.B2(n_3),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_251),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_13),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_252),
.A2(n_256),
.B1(n_9),
.B2(n_6),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_226),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_1),
.C(n_2),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_237),
.C(n_228),
.Y(n_258)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_254),
.A2(n_229),
.B1(n_241),
.B2(n_232),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_255),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_243),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_242),
.A2(n_233),
.B1(n_232),
.B2(n_234),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_249),
.B1(n_255),
.B2(n_252),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_263),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_2),
.C(n_4),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_265),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g265 ( 
.A(n_244),
.B(n_2),
.CI(n_4),
.CON(n_265),
.SN(n_265)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_267),
.B(n_5),
.Y(n_274)
);

OAI21x1_ASAP7_75t_SL g269 ( 
.A1(n_259),
.A2(n_244),
.B(n_251),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_270),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_266),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_9),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_260),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_273),
.B(n_263),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_265),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_243),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_275),
.A2(n_268),
.B(n_261),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_6),
.C(n_7),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_260),
.C(n_258),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_280),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_281),
.B(n_282),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_285),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_275),
.A2(n_265),
.B(n_264),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_284),
.A2(n_278),
.B(n_276),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_286),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_288),
.A2(n_274),
.B(n_8),
.Y(n_292)
);

AO21x1_ASAP7_75t_L g296 ( 
.A1(n_292),
.A2(n_293),
.B(n_7),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_9),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_289),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_296),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_287),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_298),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_7),
.C(n_8),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_8),
.Y(n_301)
);


endmodule