module fake_jpeg_783_n_543 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_543);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_543;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_417;
wire n_362;
wire n_142;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_9),
.B(n_5),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_50),
.Y(n_155)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_53),
.Y(n_171)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_57),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g119 ( 
.A(n_59),
.Y(n_119)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx9p33_ASAP7_75t_R g114 ( 
.A(n_60),
.Y(n_114)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_67),
.B(n_70),
.Y(n_143)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_68),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_40),
.B(n_13),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_13),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_95),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_31),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_80),
.B(n_86),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_85),
.Y(n_167)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_31),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_88),
.B(n_92),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_89),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_17),
.Y(n_90)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_90),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_93),
.Y(n_150)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_94),
.B(n_100),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_15),
.B(n_12),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_14),
.Y(n_98)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

BUFx16f_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_103),
.B(n_27),
.Y(n_166)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_105),
.Y(n_131)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_18),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_103),
.B(n_47),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_112),
.B(n_120),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_50),
.B(n_47),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_51),
.B(n_46),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_121),
.B(n_122),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_65),
.B(n_46),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_128),
.B(n_135),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_78),
.A2(n_19),
.B1(n_38),
.B2(n_18),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_130),
.A2(n_149),
.B1(n_153),
.B2(n_22),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_98),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_49),
.B(n_38),
.C(n_45),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_156),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_68),
.A2(n_26),
.B1(n_45),
.B2(n_15),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_77),
.A2(n_26),
.B1(n_35),
.B2(n_48),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_72),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_62),
.B(n_35),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_159),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_52),
.B(n_27),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_90),
.B(n_21),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_165),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_55),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_56),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_207),
.Y(n_221)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_125),
.Y(n_173)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_173),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_174),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_84),
.B1(n_58),
.B2(n_74),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_179),
.A2(n_199),
.B1(n_215),
.B2(n_144),
.Y(n_257)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_181),
.Y(n_225)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_114),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_114),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_183),
.Y(n_229)
);

HAxp5_ASAP7_75t_SL g250 ( 
.A(n_184),
.B(n_219),
.CON(n_250),
.SN(n_250)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_64),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_188),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

CKINVDCx12_ASAP7_75t_R g190 ( 
.A(n_119),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_190),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_191),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_129),
.Y(n_192)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_193),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_147),
.B(n_59),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_194),
.B(n_162),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_64),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_195),
.Y(n_251)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_196),
.Y(n_247)
);

CKINVDCx12_ASAP7_75t_R g197 ( 
.A(n_133),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_197),
.Y(n_239)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_131),
.A2(n_82),
.B1(n_69),
.B2(n_76),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_115),
.A2(n_21),
.B1(n_89),
.B2(n_85),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_200),
.A2(n_204),
.B1(n_206),
.B2(n_211),
.Y(n_222)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_202),
.Y(n_241)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_117),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_205),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_131),
.A2(n_97),
.B1(n_101),
.B2(n_53),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_117),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_158),
.A2(n_105),
.B1(n_104),
.B2(n_60),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

NAND2x1_ASAP7_75t_SL g208 ( 
.A(n_133),
.B(n_93),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_208),
.A2(n_130),
.B(n_149),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_107),
.B(n_14),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_212),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_136),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_136),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_213),
.A2(n_163),
.B1(n_141),
.B2(n_168),
.Y(n_224)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_123),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_216),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_137),
.A2(n_96),
.B1(n_91),
.B2(n_83),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_161),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_123),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_163),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_109),
.B(n_111),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_111),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_110),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_180),
.A2(n_150),
.B1(n_148),
.B2(n_168),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_258),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_224),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_203),
.A2(n_158),
.B1(n_118),
.B2(n_110),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_231),
.A2(n_244),
.B1(n_183),
.B2(n_153),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_178),
.B(n_113),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_236),
.B(n_249),
.C(n_256),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_179),
.A2(n_138),
.B1(n_154),
.B2(n_146),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_178),
.B(n_108),
.C(n_124),
.Y(n_249)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_255),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_205),
.B(n_132),
.C(n_118),
.Y(n_256)
);

OA22x2_ASAP7_75t_L g288 ( 
.A1(n_257),
.A2(n_140),
.B1(n_127),
.B2(n_145),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_175),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_259),
.B(n_261),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_216),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_260),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_176),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_257),
.A2(n_199),
.B1(n_215),
.B2(n_210),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_264),
.A2(n_288),
.B1(n_144),
.B2(n_241),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_236),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_270),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_194),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_266),
.B(n_239),
.C(n_221),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_230),
.Y(n_267)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_267),
.Y(n_292)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_269),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_194),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_271),
.A2(n_237),
.B1(n_229),
.B2(n_234),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_177),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_272),
.B(n_273),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_227),
.B(n_220),
.Y(n_273)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_238),
.Y(n_275)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_276),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_254),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_282),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_255),
.A2(n_181),
.B(n_208),
.C(n_172),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_278),
.B(n_280),
.Y(n_306)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_238),
.Y(n_279)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_279),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_227),
.B(n_193),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_223),
.B(n_208),
.Y(n_282)
);

O2A1O1Ixp33_ASAP7_75t_L g283 ( 
.A1(n_258),
.A2(n_182),
.B(n_191),
.C(n_155),
.Y(n_283)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_283),
.Y(n_312)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_228),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_285),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_221),
.B(n_227),
.Y(n_285)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_238),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_229),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_295),
.A2(n_315),
.B1(n_270),
.B2(n_288),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_260),
.B(n_239),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_298),
.B(n_316),
.Y(n_324)
);

OAI32xp33_ASAP7_75t_L g299 ( 
.A1(n_268),
.A2(n_250),
.A3(n_225),
.B1(n_253),
.B2(n_256),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_300),
.Y(n_335)
);

XNOR2x1_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_225),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_300),
.B(n_308),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_263),
.A2(n_222),
.B1(n_225),
.B2(n_145),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_301),
.A2(n_303),
.B1(n_310),
.B2(n_309),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_304),
.C(n_307),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_243),
.C(n_230),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_235),
.C(n_241),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_266),
.B(n_243),
.C(n_235),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_309),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_263),
.A2(n_229),
.B1(n_234),
.B2(n_242),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_232),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_318),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_264),
.A2(n_277),
.B1(n_268),
.B2(n_263),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_261),
.B(n_232),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_259),
.B(n_138),
.C(n_154),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_276),
.B(n_247),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_319),
.B(n_228),
.Y(n_343)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_320),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_290),
.A2(n_278),
.B(n_282),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_321),
.B(n_331),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_290),
.Y(n_322)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_322),
.Y(n_360)
);

INVx13_ASAP7_75t_L g323 ( 
.A(n_317),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_323),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_269),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_325),
.B(n_338),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_312),
.A2(n_306),
.B(n_283),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_326),
.A2(n_328),
.B(n_332),
.Y(n_353)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_289),
.Y(n_327)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_327),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_306),
.A2(n_282),
.B(n_273),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_313),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_329),
.B(n_341),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_315),
.A2(n_286),
.B(n_280),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_312),
.A2(n_291),
.B(n_305),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_333),
.B(n_337),
.Y(n_357)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_292),
.Y(n_334)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_334),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_335),
.B(n_340),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_293),
.B(n_286),
.Y(n_336)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_336),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_291),
.A2(n_272),
.B(n_274),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_296),
.B(n_262),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_292),
.B(n_284),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_294),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_293),
.B(n_287),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_348),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_343),
.B(n_347),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_345),
.A2(n_349),
.B1(n_301),
.B2(n_318),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_296),
.B(n_288),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_294),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_303),
.A2(n_288),
.B1(n_274),
.B2(n_275),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_314),
.B(n_288),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_350),
.B(n_307),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_297),
.B(n_242),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_351),
.B(n_317),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_325),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_355),
.B(n_358),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_356),
.B(n_328),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_324),
.B(n_297),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_338),
.B(n_299),
.Y(n_363)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_363),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_364),
.A2(n_366),
.B1(n_367),
.B2(n_340),
.Y(n_399)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_345),
.A2(n_302),
.B1(n_304),
.B2(n_308),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_331),
.A2(n_347),
.B1(n_350),
.B2(n_349),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_324),
.B(n_289),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_369),
.B(n_371),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_329),
.B(n_242),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_346),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_372),
.B(n_374),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_339),
.B(n_307),
.C(n_311),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_330),
.C(n_344),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_337),
.B(n_247),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_333),
.B(n_336),
.Y(n_375)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_375),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_320),
.B(n_311),
.Y(n_377)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_377),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_339),
.B(n_218),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_380),
.B(n_198),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_339),
.B(n_214),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_382),
.B(n_380),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_364),
.A2(n_326),
.B1(n_332),
.B2(n_335),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_383),
.A2(n_394),
.B1(n_400),
.B2(n_411),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_385),
.B(n_407),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_366),
.B(n_330),
.C(n_344),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_386),
.B(n_404),
.C(n_372),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_363),
.B(n_351),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_387),
.B(n_393),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_353),
.A2(n_328),
.B(n_321),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_390),
.A2(n_395),
.B(n_375),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_391),
.B(n_401),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_367),
.A2(n_346),
.B1(n_342),
.B2(n_334),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_353),
.A2(n_330),
.B(n_343),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_376),
.A2(n_344),
.B1(n_348),
.B2(n_341),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_397),
.A2(n_399),
.B1(n_403),
.B2(n_355),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_381),
.Y(n_398)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_398),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_376),
.A2(n_327),
.B1(n_274),
.B2(n_279),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_376),
.A2(n_327),
.B1(n_274),
.B2(n_323),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_SL g404 ( 
.A(n_373),
.B(n_274),
.C(n_323),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_357),
.B(n_279),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_370),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_382),
.B(n_217),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_406),
.B(n_352),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_354),
.B(n_196),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_370),
.Y(n_409)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_409),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_354),
.B(n_356),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_410),
.B(n_359),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_362),
.A2(n_233),
.B1(n_226),
.B2(n_240),
.Y(n_411)
);

MAJx2_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_435),
.C(n_427),
.Y(n_447)
);

AOI21xp33_ASAP7_75t_SL g457 ( 
.A1(n_414),
.A2(n_201),
.B(n_185),
.Y(n_457)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_415),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_417),
.B(n_419),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_396),
.B(n_384),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_418),
.B(n_202),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_402),
.A2(n_362),
.B1(n_379),
.B2(n_359),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_389),
.B(n_377),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_421),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_430),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_388),
.B(n_360),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_424),
.B(n_431),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_423),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_385),
.B(n_386),
.C(n_395),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_436),
.C(n_406),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_392),
.A2(n_379),
.B1(n_360),
.B2(n_352),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_428),
.B(n_432),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_408),
.A2(n_378),
.B1(n_368),
.B2(n_365),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_429),
.A2(n_397),
.B1(n_393),
.B2(n_407),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_383),
.B(n_378),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_368),
.Y(n_431)
);

INVxp33_ASAP7_75t_L g432 ( 
.A(n_394),
.Y(n_432)
);

INVxp33_ASAP7_75t_L g433 ( 
.A(n_411),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_433),
.B(n_186),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_390),
.B(n_361),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_404),
.B(n_361),
.C(n_381),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_437),
.A2(n_438),
.B1(n_448),
.B2(n_449),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_434),
.A2(n_403),
.B1(n_398),
.B2(n_381),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_439),
.B(n_450),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_416),
.A2(n_400),
.B1(n_401),
.B2(n_391),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_440),
.Y(n_465)
);

AOI322xp5_ASAP7_75t_L g441 ( 
.A1(n_413),
.A2(n_186),
.A3(n_213),
.B1(n_211),
.B2(n_192),
.C1(n_189),
.C2(n_174),
.Y(n_441)
);

BUFx24_ASAP7_75t_SL g469 ( 
.A(n_441),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_414),
.A2(n_416),
.B(n_432),
.Y(n_444)
);

MAJx2_ASAP7_75t_L g463 ( 
.A(n_444),
.B(n_447),
.C(n_453),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_430),
.A2(n_233),
.B1(n_226),
.B2(n_240),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_425),
.A2(n_240),
.B1(n_234),
.B2(n_213),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_422),
.B(n_173),
.C(n_212),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_420),
.B(n_170),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_454),
.B(n_457),
.Y(n_460)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_455),
.Y(n_467)
);

FAx1_ASAP7_75t_SL g456 ( 
.A(n_419),
.B(n_126),
.CI(n_211),
.CON(n_456),
.SN(n_456)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_456),
.B(n_428),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_436),
.A2(n_174),
.B1(n_192),
.B2(n_189),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_458),
.B(n_433),
.Y(n_470)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_459),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_461),
.B(n_456),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_446),
.B(n_422),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_462),
.B(n_464),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_447),
.B(n_412),
.C(n_435),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_471),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_439),
.B(n_426),
.C(n_420),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_451),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_472),
.B(n_476),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_452),
.B(n_207),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_473),
.B(n_479),
.Y(n_490)
);

INVx13_ASAP7_75t_L g475 ( 
.A(n_455),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_475),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_443),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_443),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_477),
.B(n_478),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_445),
.B(n_151),
.C(n_171),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_453),
.B(n_151),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_445),
.C(n_444),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_481),
.B(n_484),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_472),
.A2(n_451),
.B(n_440),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_482),
.A2(n_0),
.B(n_1),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_463),
.B(n_442),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_483),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_463),
.B(n_442),
.C(n_450),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_479),
.B(n_454),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_485),
.B(n_493),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_459),
.C(n_457),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_486),
.B(n_478),
.C(n_460),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_465),
.A2(n_456),
.B1(n_140),
.B2(n_142),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_488),
.A2(n_496),
.B1(n_33),
.B2(n_42),
.Y(n_509)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_489),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_467),
.B(n_142),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_491),
.B(n_0),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_471),
.B(n_79),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_469),
.B(n_162),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_494),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_466),
.A2(n_127),
.B1(n_152),
.B2(n_14),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_492),
.A2(n_466),
.B1(n_475),
.B2(n_474),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_499),
.B(n_501),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_482),
.A2(n_460),
.B1(n_152),
.B2(n_32),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_504),
.B(n_505),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_481),
.B(n_152),
.C(n_126),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_495),
.A2(n_42),
.B1(n_66),
.B2(n_81),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_506),
.B(n_508),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_509),
.B(n_512),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_480),
.A2(n_42),
.B(n_33),
.Y(n_510)
);

AOI21x1_ASAP7_75t_L g523 ( 
.A1(n_510),
.A2(n_1),
.B(n_3),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_511),
.A2(n_497),
.B(n_486),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_487),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_512)
);

AOI21x1_ASAP7_75t_SL g529 ( 
.A1(n_513),
.A2(n_518),
.B(n_522),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_483),
.C(n_484),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_515),
.B(n_516),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_503),
.B(n_502),
.C(n_501),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_502),
.A2(n_490),
.B(n_488),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_505),
.B(n_493),
.C(n_485),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_519),
.A2(n_512),
.B(n_506),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_507),
.A2(n_496),
.B(n_2),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_523),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_521),
.B(n_511),
.C(n_504),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_524),
.B(n_525),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_514),
.A2(n_509),
.B(n_498),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_526),
.B(n_530),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_514),
.A2(n_1),
.B(n_3),
.Y(n_530)
);

AOI322xp5_ASAP7_75t_L g532 ( 
.A1(n_528),
.A2(n_520),
.A3(n_517),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_4),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_532),
.B(n_533),
.C(n_535),
.Y(n_536)
);

AOI322xp5_ASAP7_75t_L g533 ( 
.A1(n_529),
.A2(n_517),
.A3(n_5),
.B1(n_7),
.B2(n_8),
.C1(n_4),
.C2(n_10),
.Y(n_533)
);

AOI322xp5_ASAP7_75t_L g535 ( 
.A1(n_527),
.A2(n_4),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_528),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_531),
.A2(n_4),
.B(n_9),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_537),
.B(n_538),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_534),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_536),
.Y(n_539)
);

INVxp33_ASAP7_75t_L g541 ( 
.A(n_539),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_540),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_542),
.B(n_10),
.Y(n_543)
);


endmodule