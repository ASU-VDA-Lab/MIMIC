module fake_netlist_5_225_n_1838 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1838);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1838;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1644;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1731;
wire n_1453;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g171 ( 
.A(n_42),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_125),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_29),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_37),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_159),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_119),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_74),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_53),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_99),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_62),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_123),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_69),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_106),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_117),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_68),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_49),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_2),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_48),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_102),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_103),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_98),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_5),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_75),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_59),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_66),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_43),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_31),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_27),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_115),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_16),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_67),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_51),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_145),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_70),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_94),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_25),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g213 ( 
.A(n_107),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_45),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_52),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_136),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_25),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_28),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g219 ( 
.A(n_81),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_52),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_54),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_110),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_18),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_54),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_170),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_35),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_10),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_40),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_131),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_87),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_128),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_21),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_113),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_8),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_55),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_36),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_30),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_77),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_160),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_32),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_23),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_8),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_53),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_112),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_33),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_7),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_50),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_83),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_10),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_108),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_97),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_3),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_73),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_63),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_33),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_126),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_40),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_32),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_38),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_161),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_155),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_24),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_60),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_12),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_64),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_121),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_140),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_78),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_22),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_17),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_50),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_26),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_56),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_137),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_65),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_45),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_157),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_5),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_162),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_127),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_147),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_138),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_163),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_41),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_36),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_72),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_80),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_3),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_167),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_79),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_149),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_19),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_82),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_38),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_42),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_88),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_114),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_55),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_109),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_92),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_135),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_93),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_101),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_0),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_19),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_71),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_116),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_56),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_39),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_164),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_27),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_142),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_96),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_46),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_58),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g316 ( 
.A(n_15),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_124),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_13),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_156),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_41),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_34),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_151),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_76),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_95),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_30),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_12),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_144),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_100),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_20),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_130),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_29),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_133),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_17),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_129),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_49),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_285),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_316),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_281),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_183),
.B(n_0),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_239),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_316),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g342 ( 
.A(n_171),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_316),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_269),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_220),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_316),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_228),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_316),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_221),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_175),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_316),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_316),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_175),
.B(n_1),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_316),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_228),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_195),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_223),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_224),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_195),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_310),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_180),
.B(n_4),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_214),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_319),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_189),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_174),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_189),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_207),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_324),
.Y(n_368)
);

INVxp33_ASAP7_75t_SL g369 ( 
.A(n_173),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_289),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_207),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_252),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_225),
.Y(n_373)
);

INVxp33_ASAP7_75t_SL g374 ( 
.A(n_173),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_199),
.B(n_6),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_231),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_214),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_226),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_199),
.B(n_229),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_215),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_199),
.B(n_6),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_252),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_273),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_273),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_227),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_304),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_304),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_229),
.B(n_7),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_228),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_234),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_190),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_191),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_215),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_201),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_202),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_236),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_218),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_242),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_181),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_246),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_186),
.B(n_9),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_237),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_247),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_249),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_262),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_190),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_262),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_255),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_257),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_244),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_253),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_240),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_271),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_203),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_276),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_305),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_181),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_362),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_200),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_337),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_417),
.B(n_200),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_373),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_362),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_376),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_337),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_377),
.Y(n_427)
);

NOR2xp67_ASAP7_75t_L g428 ( 
.A(n_348),
.B(n_179),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_365),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_365),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_340),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_377),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_380),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_360),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_380),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_348),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_351),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_352),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_339),
.A2(n_205),
.B1(n_212),
.B2(n_235),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_338),
.B(n_254),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_375),
.B(n_280),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_410),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_341),
.Y(n_444)
);

OA21x2_ASAP7_75t_L g445 ( 
.A1(n_352),
.A2(n_266),
.B(n_233),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_350),
.B(n_280),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_354),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_354),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_344),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_363),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_365),
.Y(n_451)
);

AND2x6_ASAP7_75t_L g452 ( 
.A(n_379),
.B(n_174),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_343),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_346),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_350),
.B(n_197),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_411),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_365),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_370),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_368),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_344),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_336),
.A2(n_292),
.B1(n_333),
.B2(n_326),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_356),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_388),
.B(n_233),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_408),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_345),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_364),
.B(n_266),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_356),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_353),
.B(n_197),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_345),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_359),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_366),
.B(n_286),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_408),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_353),
.B(n_213),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_409),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_349),
.B(n_185),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_409),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_357),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_357),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_359),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_381),
.B(n_286),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_393),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_358),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_393),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_405),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_358),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_378),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_420),
.Y(n_487)
);

OR2x6_ASAP7_75t_L g488 ( 
.A(n_468),
.B(n_361),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_451),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_451),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_420),
.Y(n_491)
);

OAI221xp5_ASAP7_75t_L g492 ( 
.A1(n_463),
.A2(n_401),
.B1(n_361),
.B2(n_404),
.C(n_320),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_436),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_442),
.B(n_385),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_436),
.Y(n_495)
);

AND2x6_ASAP7_75t_L g496 ( 
.A(n_480),
.B(n_174),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_452),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_431),
.Y(n_498)
);

AND2x2_ASAP7_75t_SL g499 ( 
.A(n_480),
.B(n_174),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_442),
.B(n_392),
.Y(n_500)
);

AO21x2_ASAP7_75t_L g501 ( 
.A1(n_428),
.A2(n_184),
.B(n_182),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_437),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_420),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_480),
.A2(n_369),
.B1(n_374),
.B2(n_329),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_419),
.B(n_367),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_475),
.B(n_385),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_419),
.B(n_371),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_425),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_438),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_425),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_441),
.B(n_369),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_480),
.A2(n_374),
.B1(n_314),
.B2(n_331),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_477),
.Y(n_513)
);

OR2x6_ASAP7_75t_L g514 ( 
.A(n_468),
.B(n_372),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_439),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_451),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_442),
.B(n_394),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_421),
.B(n_390),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_455),
.B(n_390),
.Y(n_519)
);

AND2x2_ASAP7_75t_SL g520 ( 
.A(n_473),
.B(n_174),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_446),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_483),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_483),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_483),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_473),
.B(n_391),
.Y(n_525)
);

OAI22xp33_ASAP7_75t_L g526 ( 
.A1(n_440),
.A2(n_217),
.B1(n_278),
.B2(n_259),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_446),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_439),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_455),
.B(n_406),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_465),
.B(n_396),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_452),
.A2(n_308),
.B1(n_414),
.B2(n_415),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_482),
.B(n_402),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_451),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_449),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_447),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_452),
.A2(n_416),
.B1(n_413),
.B2(n_395),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_451),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_447),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_442),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_483),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_483),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_485),
.B(n_402),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_483),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_444),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_479),
.B(n_484),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_448),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_444),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_451),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_462),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_486),
.B(n_412),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_469),
.B(n_347),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_457),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_453),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_479),
.B(n_382),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_460),
.Y(n_555)
);

AND2x6_ASAP7_75t_L g556 ( 
.A(n_454),
.B(n_293),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_461),
.B(n_355),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_445),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_478),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_462),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_457),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_452),
.B(n_230),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_464),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_466),
.B(n_389),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_484),
.B(n_383),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_434),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_464),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_472),
.B(n_397),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_457),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_472),
.B(n_384),
.Y(n_570)
);

INVx5_ASAP7_75t_L g571 ( 
.A(n_452),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_457),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_457),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_462),
.Y(n_574)
);

AND2x2_ASAP7_75t_SL g575 ( 
.A(n_440),
.B(n_293),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_474),
.B(n_398),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_462),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_467),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_474),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_476),
.B(n_400),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_445),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_452),
.B(n_267),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_476),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_452),
.B(n_260),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_467),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_422),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_445),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_418),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_467),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_418),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_428),
.B(n_261),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_423),
.B(n_403),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_471),
.B(n_386),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_423),
.B(n_342),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_427),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_445),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_458),
.B(n_387),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_427),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_432),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_432),
.Y(n_600)
);

AND3x2_ASAP7_75t_L g601 ( 
.A(n_433),
.B(n_192),
.C(n_188),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_433),
.B(n_172),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_426),
.B(n_263),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_435),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_426),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_426),
.B(n_265),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_429),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_424),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_435),
.B(n_405),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_470),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_470),
.B(n_407),
.Y(n_611)
);

NAND3xp33_ASAP7_75t_L g612 ( 
.A(n_470),
.B(n_243),
.C(n_241),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_481),
.B(n_172),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_481),
.B(n_407),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_481),
.A2(n_293),
.B1(n_300),
.B2(n_334),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_429),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_429),
.B(n_198),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_430),
.B(n_176),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_430),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_430),
.B(n_268),
.Y(n_620)
);

AND2x6_ASAP7_75t_L g621 ( 
.A(n_458),
.B(n_293),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_443),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_450),
.B(n_206),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_456),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_459),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_521),
.B(n_210),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_563),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_597),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_508),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_497),
.B(n_293),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_525),
.B(n_284),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_521),
.B(n_216),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_508),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_510),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_558),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_518),
.B(n_176),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_497),
.B(n_300),
.Y(n_637)
);

OAI221xp5_ASAP7_75t_L g638 ( 
.A1(n_492),
.A2(n_512),
.B1(n_504),
.B2(n_527),
.C(n_593),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_597),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_563),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_497),
.B(n_300),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_527),
.B(n_222),
.Y(n_642)
);

INVxp33_ASAP7_75t_L g643 ( 
.A(n_564),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_510),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_506),
.B(n_511),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_520),
.B(n_238),
.Y(n_646)
);

AND2x6_ASAP7_75t_L g647 ( 
.A(n_558),
.B(n_300),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_611),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_611),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_614),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_614),
.Y(n_651)
);

BUFx8_ASAP7_75t_L g652 ( 
.A(n_608),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_497),
.B(n_300),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_502),
.Y(n_654)
);

BUFx6f_ASAP7_75t_SL g655 ( 
.A(n_575),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_583),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_502),
.Y(n_657)
);

NOR3xp33_ASAP7_75t_L g658 ( 
.A(n_526),
.B(n_272),
.C(n_258),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_499),
.B(n_250),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_499),
.B(n_256),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_583),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_575),
.A2(n_275),
.B1(n_277),
.B2(n_282),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_509),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_539),
.B(n_274),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_571),
.B(n_279),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_509),
.A2(n_546),
.B1(n_515),
.B2(n_495),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_571),
.B(n_283),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_515),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_545),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_539),
.A2(n_196),
.B1(n_332),
.B2(n_330),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_546),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_553),
.B(n_302),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_SL g673 ( 
.A(n_586),
.B(n_530),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_600),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_525),
.B(n_335),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_600),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_571),
.B(n_306),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_553),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_487),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_607),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_545),
.Y(n_681)
);

BUFx2_ASAP7_75t_L g682 ( 
.A(n_498),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_607),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_493),
.B(n_315),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_528),
.A2(n_328),
.B1(n_317),
.B2(n_213),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_567),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_594),
.B(n_232),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_551),
.B(n_177),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_571),
.B(n_177),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_535),
.B(n_178),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_538),
.B(n_178),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_505),
.B(n_245),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_579),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_554),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_487),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_554),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_531),
.B(n_187),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_496),
.A2(n_213),
.B1(n_219),
.B2(n_326),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_587),
.B(n_187),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_494),
.B(n_193),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_587),
.B(n_193),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_SL g702 ( 
.A(n_586),
.B(n_219),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_488),
.A2(n_296),
.B1(n_196),
.B2(n_332),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_529),
.B(n_488),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_500),
.B(n_194),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_500),
.B(n_194),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_565),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_562),
.B(n_204),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_517),
.B(n_204),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_491),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_519),
.B(n_208),
.Y(n_711)
);

NAND3xp33_ASAP7_75t_L g712 ( 
.A(n_529),
.B(n_507),
.C(n_505),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_607),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_517),
.B(n_208),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_604),
.B(n_581),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_581),
.B(n_209),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_581),
.B(n_211),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_596),
.B(n_211),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_513),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_532),
.B(n_248),
.Y(n_720)
);

NOR3xp33_ASAP7_75t_L g721 ( 
.A(n_542),
.B(n_270),
.C(n_264),
.Y(n_721)
);

OAI22xp33_ASAP7_75t_L g722 ( 
.A1(n_488),
.A2(n_335),
.B1(n_333),
.B2(n_309),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_596),
.B(n_248),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_491),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_503),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_596),
.B(n_251),
.Y(n_726)
);

AND2x6_ASAP7_75t_SL g727 ( 
.A(n_625),
.B(n_284),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_607),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_503),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_514),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_507),
.B(n_251),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_565),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_568),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_613),
.B(n_287),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_582),
.B(n_287),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_578),
.Y(n_736)
);

BUFx6f_ASAP7_75t_SL g737 ( 
.A(n_621),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_568),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_618),
.B(n_290),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_616),
.B(n_290),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_616),
.B(n_291),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_607),
.Y(n_742)
);

INVx1_ASAP7_75t_SL g743 ( 
.A(n_559),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_592),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_593),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_536),
.B(n_291),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_578),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_619),
.B(n_296),
.Y(n_748)
);

O2A1O1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_570),
.A2(n_330),
.B(n_327),
.C(n_297),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_623),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_550),
.B(n_557),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_549),
.B(n_299),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_568),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_557),
.B(n_299),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_592),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_585),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_585),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_592),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_619),
.B(n_301),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_623),
.B(n_301),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_623),
.B(n_303),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_570),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_549),
.B(n_303),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_621),
.A2(n_612),
.B1(n_580),
.B2(n_576),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_589),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_609),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_609),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_560),
.B(n_327),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_588),
.B(n_590),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_576),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_555),
.B(n_307),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_534),
.B(n_307),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_576),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_589),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_560),
.B(n_323),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_610),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_574),
.B(n_577),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_574),
.B(n_323),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_595),
.B(n_322),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_577),
.B(n_544),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_643),
.B(n_566),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_645),
.A2(n_584),
.B1(n_615),
.B2(n_622),
.Y(n_782)
);

O2A1O1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_646),
.A2(n_599),
.B(n_598),
.C(n_602),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_636),
.A2(n_580),
.B(n_617),
.C(n_603),
.Y(n_784)
);

OAI21xp5_ASAP7_75t_L g785 ( 
.A1(n_715),
.A2(n_544),
.B(n_547),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_643),
.B(n_745),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_648),
.A2(n_650),
.B(n_649),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_674),
.Y(n_788)
);

AOI21x1_ASAP7_75t_L g789 ( 
.A1(n_780),
.A2(n_606),
.B(n_620),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_674),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_648),
.A2(n_547),
.B(n_541),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_716),
.A2(n_540),
.B(n_522),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_649),
.A2(n_543),
.B(n_541),
.Y(n_793)
);

OAI321xp33_ASAP7_75t_L g794 ( 
.A1(n_754),
.A2(n_688),
.A3(n_638),
.B1(n_722),
.B2(n_720),
.C(n_751),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_682),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_717),
.A2(n_522),
.B(n_523),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_718),
.A2(n_540),
.B(n_523),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_652),
.Y(n_798)
);

BUFx4f_ASAP7_75t_L g799 ( 
.A(n_704),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_650),
.B(n_621),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_651),
.A2(n_524),
.B(n_543),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_687),
.B(n_624),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_651),
.A2(n_524),
.B(n_591),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_R g804 ( 
.A(n_673),
.B(n_498),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_733),
.B(n_608),
.Y(n_805)
);

OAI21xp33_ASAP7_75t_L g806 ( 
.A1(n_771),
.A2(n_580),
.B(n_318),
.Y(n_806)
);

BUFx12f_ASAP7_75t_L g807 ( 
.A(n_652),
.Y(n_807)
);

CKINVDCx6p67_ASAP7_75t_R g808 ( 
.A(n_719),
.Y(n_808)
);

AOI21x1_ASAP7_75t_L g809 ( 
.A1(n_780),
.A2(n_777),
.B(n_726),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_711),
.A2(n_617),
.B(n_610),
.C(n_625),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_628),
.B(n_621),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_692),
.B(n_501),
.Y(n_812)
);

BUFx8_ASAP7_75t_L g813 ( 
.A(n_655),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_635),
.Y(n_814)
);

AO21x1_ASAP7_75t_L g815 ( 
.A1(n_659),
.A2(n_660),
.B(n_708),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_627),
.B(n_496),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_639),
.B(n_312),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_635),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_640),
.B(n_496),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_733),
.B(n_313),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_723),
.A2(n_777),
.B(n_664),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_773),
.A2(n_490),
.B(n_537),
.C(n_569),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_769),
.A2(n_533),
.B(n_489),
.Y(n_823)
);

AOI21x1_ASAP7_75t_L g824 ( 
.A1(n_699),
.A2(n_533),
.B(n_573),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_701),
.A2(n_496),
.B(n_490),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_669),
.B(n_501),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_672),
.A2(n_533),
.B(n_572),
.Y(n_827)
);

NOR2xp67_ASAP7_75t_L g828 ( 
.A(n_712),
.B(n_490),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_656),
.B(n_496),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_661),
.B(n_537),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_626),
.A2(n_573),
.B(n_572),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_632),
.A2(n_572),
.B(n_537),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_743),
.Y(n_833)
);

NOR2xp67_ASAP7_75t_L g834 ( 
.A(n_662),
.B(n_561),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_642),
.A2(n_569),
.B(n_561),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_678),
.B(n_601),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_752),
.A2(n_768),
.B(n_763),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_763),
.A2(n_569),
.B(n_501),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_655),
.A2(n_556),
.B1(n_552),
.B2(n_548),
.Y(n_839)
);

O2A1O1Ixp5_ASAP7_75t_L g840 ( 
.A1(n_708),
.A2(n_556),
.B(n_219),
.C(n_552),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_666),
.B(n_552),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_680),
.A2(n_552),
.B(n_548),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_681),
.B(n_552),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_654),
.B(n_548),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_676),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_654),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_680),
.A2(n_548),
.B(n_516),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_772),
.B(n_288),
.Y(n_848)
);

NAND2x1p5_ASAP7_75t_L g849 ( 
.A(n_738),
.B(n_548),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_655),
.A2(n_516),
.B1(n_294),
.B2(n_318),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_657),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_764),
.A2(n_516),
.B1(n_294),
.B2(n_311),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_700),
.B(n_295),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_663),
.A2(n_556),
.B(n_605),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_760),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_680),
.A2(n_516),
.B(n_605),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_766),
.B(n_295),
.Y(n_857)
);

CKINVDCx11_ASAP7_75t_R g858 ( 
.A(n_727),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_738),
.B(n_325),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_680),
.A2(n_605),
.B(n_556),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_767),
.B(n_298),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_768),
.A2(n_605),
.B(n_325),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_697),
.A2(n_298),
.B(n_309),
.C(n_321),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_683),
.A2(n_605),
.B(n_556),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_652),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_697),
.A2(n_694),
.B1(n_696),
.B2(n_707),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_668),
.B(n_556),
.Y(n_867)
);

NOR2xp67_ASAP7_75t_L g868 ( 
.A(n_750),
.B(n_61),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_671),
.B(n_321),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_700),
.B(n_9),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_775),
.A2(n_84),
.B(n_166),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_671),
.A2(n_169),
.B(n_165),
.Y(n_872)
);

INVx1_ASAP7_75t_SL g873 ( 
.A(n_631),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_686),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_675),
.B(n_761),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_753),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_770),
.A2(n_154),
.B1(n_152),
.B2(n_150),
.Y(n_877)
);

AND2x4_ASAP7_75t_SL g878 ( 
.A(n_730),
.B(n_146),
.Y(n_878)
);

INVx4_ASAP7_75t_L g879 ( 
.A(n_753),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_775),
.A2(n_141),
.B(n_139),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_744),
.A2(n_134),
.B1(n_132),
.B2(n_120),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_693),
.B(n_734),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_732),
.B(n_11),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_755),
.A2(n_118),
.B1(n_111),
.B2(n_105),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_778),
.A2(n_104),
.B(n_91),
.Y(n_885)
);

BUFx12f_ASAP7_75t_L g886 ( 
.A(n_647),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_762),
.B(n_90),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_629),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_702),
.B(n_89),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_731),
.B(n_13),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_683),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_739),
.B(n_14),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_758),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_629),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_683),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_778),
.A2(n_86),
.B(n_85),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_684),
.B(n_15),
.Y(n_897)
);

AOI21xp33_ASAP7_75t_L g898 ( 
.A1(n_735),
.A2(n_16),
.B(n_18),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_647),
.A2(n_20),
.B(n_21),
.Y(n_899)
);

O2A1O1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_735),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_900)
);

BUFx4f_ASAP7_75t_L g901 ( 
.A(n_647),
.Y(n_901)
);

NOR2xp67_ASAP7_75t_L g902 ( 
.A(n_705),
.B(n_26),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_633),
.Y(n_903)
);

OAI21xp33_ASAP7_75t_L g904 ( 
.A1(n_658),
.A2(n_34),
.B(n_43),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_633),
.A2(n_44),
.B(n_46),
.Y(n_905)
);

AOI21x1_ASAP7_75t_L g906 ( 
.A1(n_665),
.A2(n_677),
.B(n_667),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_647),
.A2(n_44),
.B(n_47),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_634),
.A2(n_47),
.B(n_48),
.Y(n_908)
);

AOI21x1_ASAP7_75t_L g909 ( 
.A1(n_665),
.A2(n_57),
.B(n_677),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_634),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_644),
.A2(n_57),
.B(n_736),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_742),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_746),
.A2(n_647),
.B1(n_698),
.B2(n_644),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_736),
.A2(n_747),
.B(n_776),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_756),
.A2(n_776),
.B(n_774),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_703),
.B(n_691),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_756),
.A2(n_774),
.B(n_765),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_757),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_757),
.B(n_765),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_706),
.B(n_709),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_679),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_779),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_737),
.A2(n_714),
.B1(n_670),
.B2(n_740),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_690),
.B(n_759),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_741),
.B(n_748),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_SL g926 ( 
.A(n_737),
.B(n_749),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_683),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_713),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_679),
.B(n_710),
.Y(n_929)
);

AOI21xp33_ASAP7_75t_L g930 ( 
.A1(n_685),
.A2(n_689),
.B(n_729),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_695),
.A2(n_729),
.B(n_725),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_689),
.A2(n_721),
.B1(n_737),
.B2(n_667),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_695),
.A2(n_710),
.B(n_725),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_724),
.B(n_742),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_724),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_742),
.A2(n_713),
.B1(n_728),
.B2(n_641),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_713),
.A2(n_728),
.B1(n_637),
.B2(n_641),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_728),
.B(n_653),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_630),
.Y(n_939)
);

NOR3xp33_ASAP7_75t_L g940 ( 
.A(n_630),
.B(n_637),
.C(n_653),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_636),
.B(n_645),
.Y(n_941)
);

NAND2x1p5_ASAP7_75t_L g942 ( 
.A(n_635),
.B(n_733),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_678),
.B(n_733),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_643),
.B(n_645),
.Y(n_944)
);

AOI21x1_ASAP7_75t_L g945 ( 
.A1(n_780),
.A2(n_587),
.B(n_715),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_635),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_715),
.A2(n_558),
.B(n_587),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_636),
.B(n_645),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_833),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_794),
.B(n_941),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_948),
.B(n_944),
.Y(n_951)
);

AO31x2_ASAP7_75t_L g952 ( 
.A1(n_815),
.A2(n_810),
.A3(n_784),
.B(n_822),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_947),
.A2(n_901),
.B(n_821),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_786),
.B(n_875),
.Y(n_954)
);

OAI21x1_ASAP7_75t_L g955 ( 
.A1(n_793),
.A2(n_801),
.B(n_809),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_947),
.A2(n_901),
.B(n_821),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_793),
.A2(n_801),
.B(n_945),
.Y(n_957)
);

OAI21x1_ASAP7_75t_L g958 ( 
.A1(n_791),
.A2(n_803),
.B(n_914),
.Y(n_958)
);

OAI21x1_ASAP7_75t_L g959 ( 
.A1(n_791),
.A2(n_803),
.B(n_914),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_924),
.B(n_925),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_802),
.B(n_855),
.Y(n_961)
);

OAI21x1_ASAP7_75t_L g962 ( 
.A1(n_915),
.A2(n_933),
.B(n_917),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_812),
.B(n_787),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_781),
.B(n_848),
.Y(n_964)
);

AO31x2_ASAP7_75t_L g965 ( 
.A1(n_838),
.A2(n_782),
.A3(n_911),
.B(n_837),
.Y(n_965)
);

AOI21xp33_ASAP7_75t_L g966 ( 
.A1(n_916),
.A2(n_870),
.B(n_853),
.Y(n_966)
);

OR2x6_ASAP7_75t_L g967 ( 
.A(n_807),
.B(n_795),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_787),
.A2(n_838),
.B(n_837),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_882),
.B(n_890),
.Y(n_969)
);

INVx1_ASAP7_75t_SL g970 ( 
.A(n_808),
.Y(n_970)
);

O2A1O1Ixp5_ASAP7_75t_L g971 ( 
.A1(n_892),
.A2(n_920),
.B(n_840),
.C(n_923),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_922),
.B(n_866),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_836),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_818),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_827),
.A2(n_823),
.B(n_825),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_876),
.B(n_943),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_863),
.A2(n_806),
.B(n_783),
.C(n_904),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_876),
.B(n_943),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_851),
.B(n_790),
.Y(n_979)
);

BUFx4_ASAP7_75t_SL g980 ( 
.A(n_798),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_792),
.A2(n_796),
.B(n_797),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_835),
.A2(n_931),
.B(n_824),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_930),
.A2(n_902),
.B(n_898),
.C(n_874),
.Y(n_983)
);

OA21x2_ASAP7_75t_L g984 ( 
.A1(n_785),
.A2(n_800),
.B(n_835),
.Y(n_984)
);

NAND2x1p5_ASAP7_75t_L g985 ( 
.A(n_818),
.B(n_946),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_789),
.A2(n_832),
.B(n_842),
.Y(n_986)
);

AO31x2_ASAP7_75t_L g987 ( 
.A1(n_911),
.A2(n_936),
.A3(n_937),
.B(n_908),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_913),
.A2(n_826),
.B(n_841),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_818),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_893),
.B(n_879),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_845),
.Y(n_991)
);

AOI21x1_ASAP7_75t_L g992 ( 
.A1(n_831),
.A2(n_844),
.B(n_827),
.Y(n_992)
);

AOI221xp5_ASAP7_75t_L g993 ( 
.A1(n_873),
.A2(n_861),
.B1(n_857),
.B2(n_900),
.C(n_817),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_832),
.A2(n_847),
.B(n_934),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_804),
.Y(n_995)
);

INVx4_ASAP7_75t_L g996 ( 
.A(n_946),
.Y(n_996)
);

INVxp67_ASAP7_75t_SL g997 ( 
.A(n_946),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_938),
.A2(n_929),
.B(n_919),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_846),
.B(n_814),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_SL g1000 ( 
.A1(n_881),
.A2(n_897),
.B(n_896),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_799),
.B(n_869),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_811),
.A2(n_883),
.B(n_932),
.C(n_834),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_935),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_SL g1004 ( 
.A1(n_942),
.A2(n_928),
.B(n_927),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_816),
.A2(n_829),
.B(n_819),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_856),
.A2(n_912),
.B(n_906),
.Y(n_1006)
);

NOR2x1_ASAP7_75t_SL g1007 ( 
.A(n_886),
.B(n_891),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_828),
.A2(n_896),
.B(n_871),
.C(n_885),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_912),
.A2(n_830),
.B(n_843),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_849),
.A2(n_918),
.B(n_921),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_849),
.A2(n_888),
.B(n_910),
.Y(n_1011)
);

O2A1O1Ixp5_ASAP7_75t_L g1012 ( 
.A1(n_887),
.A2(n_854),
.B(n_820),
.C(n_862),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_876),
.B(n_903),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_942),
.A2(n_839),
.B1(n_799),
.B2(n_939),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_880),
.A2(n_885),
.B(n_862),
.C(n_868),
.Y(n_1015)
);

NAND3xp33_ASAP7_75t_L g1016 ( 
.A(n_859),
.B(n_850),
.C(n_805),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_852),
.B(n_836),
.Y(n_1017)
);

BUFx12f_ASAP7_75t_L g1018 ( 
.A(n_813),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_894),
.A2(n_867),
.B(n_940),
.Y(n_1019)
);

O2A1O1Ixp5_ASAP7_75t_L g1020 ( 
.A1(n_909),
.A2(n_889),
.B(n_880),
.C(n_908),
.Y(n_1020)
);

NOR2xp67_ASAP7_75t_L g1021 ( 
.A(n_865),
.B(n_905),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_926),
.B(n_813),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_891),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_860),
.A2(n_864),
.B(n_877),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_884),
.A2(n_905),
.B(n_891),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_895),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_895),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_927),
.B(n_928),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_878),
.B(n_858),
.Y(n_1029)
);

NAND2x1_ASAP7_75t_L g1030 ( 
.A(n_818),
.B(n_635),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_SL g1031 ( 
.A1(n_899),
.A2(n_907),
.B(n_872),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_784),
.A2(n_539),
.B(n_497),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_793),
.A2(n_801),
.B(n_809),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_947),
.A2(n_821),
.B(n_941),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_851),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_818),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_941),
.B(n_948),
.Y(n_1037)
);

AOI21xp33_ASAP7_75t_L g1038 ( 
.A1(n_941),
.A2(n_948),
.B(n_794),
.Y(n_1038)
);

INVxp67_ASAP7_75t_L g1039 ( 
.A(n_786),
.Y(n_1039)
);

OAI21xp33_ASAP7_75t_L g1040 ( 
.A1(n_848),
.A2(n_645),
.B(n_941),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_784),
.A2(n_539),
.B(n_497),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_944),
.B(n_941),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_833),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_784),
.A2(n_539),
.B(n_497),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_941),
.A2(n_948),
.B(n_794),
.C(n_645),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_941),
.B(n_948),
.Y(n_1046)
);

AOI21xp33_ASAP7_75t_L g1047 ( 
.A1(n_941),
.A2(n_948),
.B(n_794),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_784),
.A2(n_539),
.B(n_497),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_947),
.A2(n_821),
.B(n_941),
.Y(n_1049)
);

CKINVDCx11_ASAP7_75t_R g1050 ( 
.A(n_807),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_941),
.B(n_948),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_941),
.B(n_948),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_941),
.B(n_948),
.Y(n_1053)
);

INVx1_ASAP7_75t_SL g1054 ( 
.A(n_833),
.Y(n_1054)
);

NOR3xp33_ASAP7_75t_L g1055 ( 
.A(n_794),
.B(n_458),
.C(n_941),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_943),
.B(n_678),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_793),
.A2(n_801),
.B(n_809),
.Y(n_1057)
);

AO31x2_ASAP7_75t_L g1058 ( 
.A1(n_815),
.A2(n_810),
.A3(n_784),
.B(n_822),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_818),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_944),
.B(n_643),
.Y(n_1060)
);

OAI21xp33_ASAP7_75t_L g1061 ( 
.A1(n_848),
.A2(n_645),
.B(n_941),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_794),
.B(n_941),
.Y(n_1062)
);

AO31x2_ASAP7_75t_L g1063 ( 
.A1(n_815),
.A2(n_810),
.A3(n_784),
.B(n_822),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_SL g1064 ( 
.A(n_899),
.B(n_655),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_794),
.B(n_941),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_941),
.B(n_948),
.Y(n_1066)
);

AND2x6_ASAP7_75t_L g1067 ( 
.A(n_818),
.B(n_635),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_947),
.A2(n_821),
.B(n_941),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_804),
.Y(n_1069)
);

NAND2x1p5_ASAP7_75t_L g1070 ( 
.A(n_818),
.B(n_946),
.Y(n_1070)
);

AO31x2_ASAP7_75t_L g1071 ( 
.A1(n_815),
.A2(n_810),
.A3(n_784),
.B(n_822),
.Y(n_1071)
);

AOI21xp33_ASAP7_75t_L g1072 ( 
.A1(n_941),
.A2(n_948),
.B(n_794),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_941),
.B(n_948),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_851),
.Y(n_1074)
);

INVxp67_ASAP7_75t_SL g1075 ( 
.A(n_818),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_SL g1076 ( 
.A1(n_899),
.A2(n_907),
.B(n_872),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_941),
.B(n_948),
.Y(n_1077)
);

NAND2x1_ASAP7_75t_L g1078 ( 
.A(n_818),
.B(n_635),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_793),
.A2(n_801),
.B(n_809),
.Y(n_1079)
);

AOI21xp33_ASAP7_75t_L g1080 ( 
.A1(n_941),
.A2(n_948),
.B(n_794),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_851),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_944),
.B(n_941),
.Y(n_1082)
);

A2O1A1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_941),
.A2(n_948),
.B(n_794),
.C(n_645),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_943),
.B(n_678),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_793),
.A2(n_801),
.B(n_809),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_794),
.B(n_941),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_947),
.A2(n_821),
.B(n_941),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_793),
.A2(n_801),
.B(n_809),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_788),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_960),
.A2(n_1045),
.B1(n_1083),
.B2(n_1051),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1060),
.B(n_954),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_1043),
.Y(n_1092)
);

AOI21x1_ASAP7_75t_L g1093 ( 
.A1(n_953),
.A2(n_956),
.B(n_992),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_949),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1046),
.A2(n_1066),
.B1(n_1073),
.B2(n_964),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1042),
.B(n_1082),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_1054),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_1054),
.Y(n_1098)
);

BUFx8_ASAP7_75t_L g1099 ( 
.A(n_1018),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_1067),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_974),
.Y(n_1101)
);

BUFx4f_ASAP7_75t_L g1102 ( 
.A(n_967),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_1050),
.Y(n_1103)
);

CKINVDCx11_ASAP7_75t_R g1104 ( 
.A(n_967),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_951),
.B(n_1052),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1035),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1074),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1037),
.B(n_1055),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1052),
.B(n_1053),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_966),
.B(n_1040),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_1067),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_957),
.A2(n_1033),
.B(n_955),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_974),
.Y(n_1113)
);

INVx5_ASAP7_75t_L g1114 ( 
.A(n_1067),
.Y(n_1114)
);

OA21x2_ASAP7_75t_L g1115 ( 
.A1(n_981),
.A2(n_968),
.B(n_1034),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1056),
.B(n_1084),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1081),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1053),
.B(n_1077),
.Y(n_1118)
);

INVx5_ASAP7_75t_L g1119 ( 
.A(n_1067),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_979),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_966),
.A2(n_1061),
.B(n_1080),
.C(n_1047),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_970),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_974),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_1036),
.Y(n_1124)
);

NAND2x1p5_ASAP7_75t_L g1125 ( 
.A(n_996),
.B(n_1030),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_1036),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_979),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_1056),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_1078),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_950),
.A2(n_1062),
.B1(n_1086),
.B2(n_1065),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_991),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_958),
.Y(n_1132)
);

INVx5_ASAP7_75t_L g1133 ( 
.A(n_1036),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1077),
.B(n_969),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_1084),
.B(n_990),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1001),
.B(n_1039),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1003),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_996),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_959),
.Y(n_1139)
);

BUFx10_ASAP7_75t_L g1140 ( 
.A(n_1022),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_970),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_973),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_967),
.Y(n_1143)
);

BUFx12f_ASAP7_75t_L g1144 ( 
.A(n_1069),
.Y(n_1144)
);

INVx5_ASAP7_75t_L g1145 ( 
.A(n_1023),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1089),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1038),
.A2(n_1047),
.B1(n_1080),
.B2(n_1072),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_980),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1034),
.A2(n_1068),
.B(n_1087),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_999),
.Y(n_1150)
);

BUFx12f_ASAP7_75t_L g1151 ( 
.A(n_1029),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_961),
.B(n_993),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_990),
.B(n_976),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_972),
.B(n_963),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1064),
.A2(n_1031),
.B1(n_1076),
.B2(n_1016),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_995),
.B(n_1017),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1064),
.A2(n_988),
.B(n_977),
.C(n_1000),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_985),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_995),
.B(n_978),
.Y(n_1159)
);

INVx1_ASAP7_75t_SL g1160 ( 
.A(n_1013),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1002),
.A2(n_963),
.B1(n_983),
.B2(n_1014),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_989),
.Y(n_1162)
);

OAI21xp33_ASAP7_75t_L g1163 ( 
.A1(n_988),
.A2(n_1049),
.B(n_1087),
.Y(n_1163)
);

NOR2x1_ASAP7_75t_L g1164 ( 
.A(n_1004),
.B(n_1059),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_989),
.Y(n_1165)
);

NOR2xp67_ASAP7_75t_L g1166 ( 
.A(n_1021),
.B(n_1059),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_985),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1026),
.B(n_1027),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_1028),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_999),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1070),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_1007),
.B(n_1023),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_1070),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1049),
.A2(n_1068),
.B1(n_968),
.B2(n_1014),
.Y(n_1174)
);

INVx3_ASAP7_75t_SL g1175 ( 
.A(n_984),
.Y(n_1175)
);

INVx2_ASAP7_75t_SL g1176 ( 
.A(n_1010),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_1011),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_997),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1075),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_SL g1180 ( 
.A1(n_1008),
.A2(n_1015),
.B(n_1005),
.C(n_1019),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1019),
.A2(n_998),
.B1(n_1005),
.B2(n_984),
.Y(n_1181)
);

INVx4_ASAP7_75t_L g1182 ( 
.A(n_1025),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_965),
.B(n_971),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1057),
.A2(n_1088),
.B1(n_1085),
.B2(n_1079),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_987),
.B(n_952),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_987),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_952),
.B(n_1071),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1009),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1006),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1024),
.Y(n_1190)
);

CKINVDCx16_ASAP7_75t_R g1191 ( 
.A(n_1012),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_952),
.Y(n_1192)
);

AND2x2_ASAP7_75t_SL g1193 ( 
.A(n_1058),
.B(n_1071),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1058),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1058),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1063),
.B(n_1071),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1063),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1020),
.A2(n_1041),
.B(n_1048),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1032),
.A2(n_1044),
.B1(n_994),
.B2(n_982),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_986),
.B(n_1063),
.Y(n_1200)
);

NAND2xp33_ASAP7_75t_L g1201 ( 
.A(n_960),
.B(n_1045),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1067),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_960),
.B(n_1042),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1067),
.Y(n_1204)
);

INVxp67_ASAP7_75t_SL g1205 ( 
.A(n_960),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_1054),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_1050),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_1054),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_966),
.B(n_1042),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1056),
.B(n_1084),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1060),
.B(n_954),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_960),
.B(n_1042),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_960),
.B(n_1042),
.Y(n_1213)
);

NOR2x1_ASAP7_75t_L g1214 ( 
.A(n_949),
.B(n_624),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_981),
.A2(n_975),
.B(n_956),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_949),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1067),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1043),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_1043),
.Y(n_1219)
);

CKINVDCx11_ASAP7_75t_R g1220 ( 
.A(n_1050),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_949),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_960),
.B(n_1042),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_960),
.B(n_1042),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_966),
.B(n_794),
.Y(n_1224)
);

BUFx4f_ASAP7_75t_SL g1225 ( 
.A(n_1018),
.Y(n_1225)
);

INVxp67_ASAP7_75t_L g1226 ( 
.A(n_1043),
.Y(n_1226)
);

INVx5_ASAP7_75t_L g1227 ( 
.A(n_1067),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_981),
.A2(n_975),
.B(n_956),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1067),
.Y(n_1229)
);

OR2x6_ASAP7_75t_L g1230 ( 
.A(n_967),
.B(n_1004),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_974),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_1043),
.Y(n_1232)
);

OAI21xp33_ASAP7_75t_L g1233 ( 
.A1(n_964),
.A2(n_960),
.B(n_1040),
.Y(n_1233)
);

BUFx12f_ASAP7_75t_L g1234 ( 
.A(n_1050),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_960),
.B(n_1042),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_949),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_962),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1106),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_SL g1239 ( 
.A1(n_1209),
.A2(n_1096),
.B1(n_1110),
.B2(n_1095),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1107),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1117),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1209),
.A2(n_1224),
.B1(n_1110),
.B2(n_1233),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1224),
.A2(n_1201),
.B1(n_1090),
.B2(n_1108),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1098),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1216),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1220),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1201),
.A2(n_1152),
.B1(n_1205),
.B2(n_1130),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1150),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_1207),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1203),
.B(n_1212),
.Y(n_1250)
);

CKINVDCx11_ASAP7_75t_R g1251 ( 
.A(n_1220),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1205),
.A2(n_1130),
.B1(n_1213),
.B2(n_1235),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1216),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1222),
.A2(n_1223),
.B1(n_1118),
.B2(n_1109),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1163),
.A2(n_1134),
.B1(n_1147),
.B2(n_1161),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1206),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1131),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1137),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1105),
.B(n_1091),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_1208),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_1236),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1146),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1147),
.A2(n_1174),
.B1(n_1155),
.B2(n_1156),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1221),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1133),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1114),
.Y(n_1266)
);

AO21x2_ASAP7_75t_L g1267 ( 
.A1(n_1198),
.A2(n_1228),
.B(n_1215),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_SL g1268 ( 
.A1(n_1156),
.A2(n_1102),
.B1(n_1191),
.B2(n_1140),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1153),
.B(n_1230),
.Y(n_1269)
);

INVx4_ASAP7_75t_L g1270 ( 
.A(n_1114),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1133),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1168),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1097),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1211),
.B(n_1136),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1170),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1133),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1120),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1154),
.B(n_1160),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1094),
.Y(n_1279)
);

CKINVDCx11_ASAP7_75t_R g1280 ( 
.A(n_1207),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1133),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1112),
.A2(n_1184),
.B(n_1199),
.Y(n_1282)
);

CKINVDCx11_ASAP7_75t_R g1283 ( 
.A(n_1234),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1127),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_SL g1285 ( 
.A1(n_1102),
.A2(n_1140),
.B1(n_1159),
.B2(n_1221),
.Y(n_1285)
);

CKINVDCx11_ASAP7_75t_R g1286 ( 
.A(n_1234),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1169),
.B(n_1121),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1174),
.A2(n_1155),
.B1(n_1149),
.B2(n_1115),
.Y(n_1288)
);

AO21x1_ASAP7_75t_L g1289 ( 
.A1(n_1194),
.A2(n_1195),
.B(n_1197),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1121),
.B(n_1092),
.Y(n_1290)
);

INVx2_ASAP7_75t_SL g1291 ( 
.A(n_1145),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1157),
.A2(n_1219),
.B1(n_1226),
.B2(n_1141),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1218),
.B(n_1232),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1171),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1167),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1119),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_SL g1297 ( 
.A1(n_1157),
.A2(n_1214),
.B(n_1122),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1210),
.B(n_1135),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1153),
.A2(n_1144),
.B1(n_1151),
.B2(n_1116),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1167),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1227),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1135),
.B(n_1116),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_SL g1303 ( 
.A1(n_1143),
.A2(n_1153),
.B(n_1226),
.Y(n_1303)
);

OAI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1230),
.A2(n_1219),
.B1(n_1196),
.B2(n_1185),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1179),
.Y(n_1305)
);

CKINVDCx11_ASAP7_75t_R g1306 ( 
.A(n_1104),
.Y(n_1306)
);

BUFx8_ASAP7_75t_L g1307 ( 
.A(n_1148),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1115),
.A2(n_1104),
.B1(n_1186),
.B2(n_1193),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1184),
.A2(n_1199),
.B(n_1188),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1128),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1178),
.Y(n_1311)
);

NAND2x1p5_ASAP7_75t_L g1312 ( 
.A(n_1227),
.B(n_1164),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1144),
.A2(n_1151),
.B1(n_1230),
.B2(n_1142),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1165),
.Y(n_1314)
);

INVx6_ASAP7_75t_L g1315 ( 
.A(n_1227),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1188),
.A2(n_1139),
.B(n_1132),
.Y(n_1316)
);

BUFx12f_ASAP7_75t_L g1317 ( 
.A(n_1103),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1178),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1115),
.A2(n_1193),
.B1(n_1187),
.B2(n_1183),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1162),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1128),
.B(n_1165),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1103),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1158),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1158),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1172),
.B(n_1173),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1192),
.A2(n_1181),
.B1(n_1200),
.B2(n_1172),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1173),
.Y(n_1327)
);

AO21x2_ASAP7_75t_L g1328 ( 
.A1(n_1132),
.A2(n_1139),
.B(n_1237),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1101),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1145),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1181),
.A2(n_1200),
.B1(n_1172),
.B2(n_1166),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1101),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1101),
.Y(n_1333)
);

BUFx2_ASAP7_75t_SL g1334 ( 
.A(n_1101),
.Y(n_1334)
);

CKINVDCx11_ASAP7_75t_R g1335 ( 
.A(n_1113),
.Y(n_1335)
);

NOR2x1_ASAP7_75t_R g1336 ( 
.A(n_1225),
.B(n_1231),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1113),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1113),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1180),
.B(n_1138),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1113),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1100),
.B(n_1202),
.Y(n_1341)
);

BUFx2_ASAP7_75t_R g1342 ( 
.A(n_1177),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_1099),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1225),
.A2(n_1099),
.B1(n_1100),
.B2(n_1111),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1111),
.A2(n_1202),
.B(n_1229),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1189),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1123),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1123),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1123),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1123),
.Y(n_1350)
);

BUFx2_ASAP7_75t_R g1351 ( 
.A(n_1177),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1124),
.Y(n_1352)
);

AO21x1_ASAP7_75t_SL g1353 ( 
.A1(n_1180),
.A2(n_1175),
.B(n_1229),
.Y(n_1353)
);

CKINVDCx6p67_ASAP7_75t_R g1354 ( 
.A(n_1145),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1124),
.B(n_1231),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1204),
.A2(n_1217),
.B(n_1129),
.Y(n_1356)
);

CKINVDCx8_ASAP7_75t_R g1357 ( 
.A(n_1124),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_1182),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1176),
.A2(n_1182),
.B(n_1190),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1190),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1126),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1126),
.Y(n_1362)
);

CKINVDCx6p67_ASAP7_75t_R g1363 ( 
.A(n_1145),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1126),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1231),
.Y(n_1365)
);

NOR2x1_ASAP7_75t_R g1366 ( 
.A(n_1129),
.B(n_1190),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1125),
.A2(n_966),
.B1(n_1209),
.B2(n_1055),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1125),
.A2(n_1093),
.B(n_1112),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1319),
.B(n_1243),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1319),
.B(n_1243),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1289),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1346),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1288),
.B(n_1242),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1269),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1288),
.B(n_1242),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1328),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1308),
.B(n_1239),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1308),
.B(n_1326),
.Y(n_1378)
);

AO21x2_ASAP7_75t_L g1379 ( 
.A1(n_1309),
.A2(n_1282),
.B(n_1267),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1252),
.B(n_1254),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1328),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1318),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1346),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1326),
.B(n_1255),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1269),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1316),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1255),
.B(n_1263),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1368),
.A2(n_1356),
.B(n_1358),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1252),
.B(n_1247),
.Y(n_1389)
);

INVx4_ASAP7_75t_L g1390 ( 
.A(n_1301),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1263),
.B(n_1248),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1248),
.B(n_1275),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1353),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1359),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1277),
.B(n_1284),
.Y(n_1395)
);

OA21x2_ASAP7_75t_L g1396 ( 
.A1(n_1331),
.A2(n_1367),
.B(n_1247),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1359),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1359),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1238),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1240),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1267),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1331),
.B(n_1241),
.Y(n_1402)
);

AO21x2_ASAP7_75t_L g1403 ( 
.A1(n_1339),
.A2(n_1360),
.B(n_1290),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1269),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1356),
.B(n_1345),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1366),
.A2(n_1287),
.B(n_1312),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1311),
.B(n_1259),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1367),
.A2(n_1345),
.B(n_1257),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1258),
.Y(n_1409)
);

AO21x1_ASAP7_75t_SL g1410 ( 
.A1(n_1313),
.A2(n_1323),
.B(n_1324),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1315),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1262),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_1280),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1272),
.B(n_1274),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1305),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1325),
.B(n_1295),
.Y(n_1416)
);

BUFx2_ASAP7_75t_L g1417 ( 
.A(n_1300),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1294),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1250),
.B(n_1278),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1304),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1268),
.B(n_1285),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1320),
.B(n_1355),
.Y(n_1422)
);

INVxp67_ASAP7_75t_L g1423 ( 
.A(n_1244),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1297),
.A2(n_1303),
.B(n_1292),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1266),
.B(n_1296),
.Y(n_1425)
);

INVxp67_ASAP7_75t_L g1426 ( 
.A(n_1256),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1270),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1273),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1291),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1327),
.A2(n_1352),
.B(n_1365),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1332),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1330),
.Y(n_1432)
);

INVxp67_ASAP7_75t_L g1433 ( 
.A(n_1348),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1261),
.B(n_1260),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1245),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1329),
.B(n_1364),
.Y(n_1436)
);

INVx8_ASAP7_75t_L g1437 ( 
.A(n_1301),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1354),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1333),
.B(n_1349),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1354),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1350),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1245),
.B(n_1264),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1337),
.B(n_1338),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1363),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1340),
.B(n_1361),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1363),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1341),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1341),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1347),
.B(n_1362),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1341),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1253),
.B(n_1264),
.Y(n_1451)
);

NAND2x1_ASAP7_75t_L g1452 ( 
.A(n_1315),
.B(n_1301),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1301),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1315),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1253),
.Y(n_1455)
);

INVx5_ASAP7_75t_L g1456 ( 
.A(n_1265),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1428),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1420),
.B(n_1321),
.Y(n_1458)
);

AOI211xp5_ASAP7_75t_L g1459 ( 
.A1(n_1421),
.A2(n_1336),
.B(n_1302),
.C(n_1279),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1420),
.B(n_1314),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1401),
.B(n_1351),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1401),
.B(n_1342),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1430),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1397),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1386),
.B(n_1403),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1403),
.B(n_1299),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_SL g1467 ( 
.A(n_1387),
.B(n_1357),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1403),
.B(n_1310),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_1435),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1403),
.B(n_1310),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1398),
.B(n_1334),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1430),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1380),
.B(n_1293),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1371),
.B(n_1298),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_1413),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1380),
.B(n_1344),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1398),
.B(n_1281),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1391),
.B(n_1271),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1369),
.B(n_1357),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1399),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1399),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1369),
.B(n_1335),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1400),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1370),
.B(n_1335),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1400),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1371),
.B(n_1271),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1370),
.B(n_1265),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1430),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1382),
.B(n_1271),
.Y(n_1489)
);

INVx3_ASAP7_75t_L g1490 ( 
.A(n_1405),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1391),
.B(n_1271),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1405),
.B(n_1276),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1389),
.A2(n_1246),
.B1(n_1249),
.B2(n_1343),
.Y(n_1493)
);

CKINVDCx6p67_ASAP7_75t_R g1494 ( 
.A(n_1456),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1430),
.Y(n_1495)
);

INVx2_ASAP7_75t_SL g1496 ( 
.A(n_1405),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1394),
.B(n_1265),
.Y(n_1497)
);

AOI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1376),
.A2(n_1276),
.B(n_1306),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1435),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1430),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1405),
.B(n_1388),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1394),
.B(n_1306),
.Y(n_1502)
);

AOI221xp5_ASAP7_75t_L g1503 ( 
.A1(n_1387),
.A2(n_1246),
.B1(n_1249),
.B2(n_1322),
.C(n_1343),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1372),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1480),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1468),
.B(n_1378),
.Y(n_1506)
);

NAND3xp33_ASAP7_75t_L g1507 ( 
.A(n_1459),
.B(n_1406),
.C(n_1377),
.Y(n_1507)
);

OAI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1459),
.A2(n_1419),
.B1(n_1389),
.B2(n_1377),
.C(n_1406),
.Y(n_1508)
);

OAI221xp5_ASAP7_75t_SL g1509 ( 
.A1(n_1503),
.A2(n_1384),
.B1(n_1373),
.B2(n_1375),
.C(n_1378),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1472),
.A2(n_1388),
.B(n_1381),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1468),
.B(n_1408),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1476),
.A2(n_1396),
.B1(n_1424),
.B2(n_1384),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1473),
.B(n_1458),
.Y(n_1513)
);

NOR3xp33_ASAP7_75t_L g1514 ( 
.A(n_1493),
.B(n_1419),
.C(n_1438),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1473),
.B(n_1402),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1458),
.B(n_1402),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1468),
.B(n_1408),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1457),
.B(n_1423),
.Y(n_1518)
);

OAI221xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1503),
.A2(n_1373),
.B1(n_1375),
.B2(n_1426),
.C(n_1423),
.Y(n_1519)
);

OAI221xp5_ASAP7_75t_SL g1520 ( 
.A1(n_1476),
.A2(n_1426),
.B1(n_1434),
.B2(n_1407),
.C(n_1428),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1470),
.B(n_1408),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1457),
.B(n_1407),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1502),
.A2(n_1396),
.B1(n_1424),
.B2(n_1404),
.Y(n_1523)
);

NAND3xp33_ASAP7_75t_L g1524 ( 
.A(n_1460),
.B(n_1424),
.C(n_1396),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1496),
.B(n_1379),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1474),
.B(n_1415),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1474),
.B(n_1415),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1470),
.B(n_1408),
.Y(n_1528)
);

OAI21xp5_ASAP7_75t_SL g1529 ( 
.A1(n_1482),
.A2(n_1438),
.B(n_1440),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1460),
.B(n_1417),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1502),
.B(n_1414),
.Y(n_1531)
);

NAND3xp33_ASAP7_75t_L g1532 ( 
.A(n_1466),
.B(n_1424),
.C(n_1396),
.Y(n_1532)
);

NAND3xp33_ASAP7_75t_L g1533 ( 
.A(n_1466),
.B(n_1424),
.C(n_1396),
.Y(n_1533)
);

AOI211xp5_ASAP7_75t_L g1534 ( 
.A1(n_1482),
.A2(n_1484),
.B(n_1502),
.C(n_1466),
.Y(n_1534)
);

NAND3xp33_ASAP7_75t_L g1535 ( 
.A(n_1486),
.B(n_1450),
.C(n_1448),
.Y(n_1535)
);

NAND4xp25_ASAP7_75t_L g1536 ( 
.A(n_1482),
.B(n_1434),
.C(n_1414),
.D(n_1484),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1487),
.B(n_1409),
.Y(n_1537)
);

OAI221xp5_ASAP7_75t_L g1538 ( 
.A1(n_1467),
.A2(n_1451),
.B1(n_1442),
.B2(n_1446),
.C(n_1440),
.Y(n_1538)
);

NAND3xp33_ASAP7_75t_L g1539 ( 
.A(n_1486),
.B(n_1448),
.C(n_1450),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1470),
.B(n_1408),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1487),
.B(n_1409),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1487),
.B(n_1412),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1467),
.B(n_1425),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1477),
.B(n_1372),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1478),
.B(n_1412),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1478),
.B(n_1418),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1477),
.B(n_1383),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1461),
.B(n_1425),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1461),
.B(n_1425),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1491),
.B(n_1418),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1491),
.B(n_1418),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1464),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1504),
.B(n_1416),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1504),
.B(n_1416),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1489),
.B(n_1480),
.Y(n_1555)
);

OAI211xp5_ASAP7_75t_SL g1556 ( 
.A1(n_1489),
.A2(n_1251),
.B(n_1451),
.C(n_1442),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1481),
.B(n_1392),
.Y(n_1557)
);

NAND4xp25_ASAP7_75t_L g1558 ( 
.A(n_1484),
.B(n_1449),
.C(n_1422),
.D(n_1395),
.Y(n_1558)
);

OAI21xp33_ASAP7_75t_L g1559 ( 
.A1(n_1479),
.A2(n_1447),
.B(n_1422),
.Y(n_1559)
);

OAI221xp5_ASAP7_75t_L g1560 ( 
.A1(n_1498),
.A2(n_1444),
.B1(n_1446),
.B2(n_1454),
.C(n_1455),
.Y(n_1560)
);

NAND4xp25_ASAP7_75t_L g1561 ( 
.A(n_1479),
.B(n_1449),
.C(n_1395),
.D(n_1445),
.Y(n_1561)
);

NAND4xp25_ASAP7_75t_L g1562 ( 
.A(n_1479),
.B(n_1439),
.C(n_1443),
.D(n_1445),
.Y(n_1562)
);

AOI221xp5_ASAP7_75t_L g1563 ( 
.A1(n_1465),
.A2(n_1433),
.B1(n_1447),
.B2(n_1431),
.C(n_1441),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1530),
.B(n_1496),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1506),
.B(n_1496),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1506),
.B(n_1490),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1544),
.B(n_1490),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1552),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1513),
.B(n_1477),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1505),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1505),
.Y(n_1571)
);

INVxp67_ASAP7_75t_L g1572 ( 
.A(n_1518),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1515),
.B(n_1481),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1525),
.B(n_1490),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1516),
.B(n_1465),
.Y(n_1575)
);

NOR2x1_ASAP7_75t_L g1576 ( 
.A(n_1524),
.B(n_1469),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1552),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1555),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1547),
.B(n_1501),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1547),
.B(n_1501),
.Y(n_1580)
);

NAND2x1p5_ASAP7_75t_L g1581 ( 
.A(n_1543),
.B(n_1469),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1553),
.B(n_1465),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1510),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1522),
.B(n_1483),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1511),
.B(n_1501),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1526),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1511),
.B(n_1501),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1525),
.B(n_1501),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1560),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1510),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1507),
.B(n_1455),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1527),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1545),
.B(n_1483),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1557),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1509),
.A2(n_1519),
.B1(n_1508),
.B2(n_1520),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1546),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1517),
.B(n_1497),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1554),
.B(n_1463),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1537),
.B(n_1488),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1541),
.B(n_1495),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1510),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1542),
.B(n_1495),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1517),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1550),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1521),
.B(n_1492),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1531),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1551),
.B(n_1485),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1535),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1521),
.B(n_1500),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1512),
.B(n_1485),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1528),
.B(n_1497),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1610),
.B(n_1532),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1570),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1570),
.Y(n_1614)
);

AOI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1595),
.A2(n_1589),
.B1(n_1591),
.B2(n_1608),
.C(n_1514),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1571),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1575),
.B(n_1533),
.Y(n_1617)
);

OR2x6_ASAP7_75t_L g1618 ( 
.A(n_1576),
.B(n_1543),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1605),
.B(n_1534),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1575),
.B(n_1528),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1605),
.B(n_1540),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1605),
.B(n_1539),
.Y(n_1622)
);

NOR2x1_ASAP7_75t_L g1623 ( 
.A(n_1589),
.B(n_1576),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1605),
.B(n_1540),
.Y(n_1624)
);

INVxp67_ASAP7_75t_SL g1625 ( 
.A(n_1608),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1564),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1571),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1568),
.Y(n_1628)
);

NOR2x1_ASAP7_75t_R g1629 ( 
.A(n_1589),
.B(n_1251),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1586),
.B(n_1592),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1586),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1585),
.B(n_1548),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1588),
.B(n_1548),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1598),
.B(n_1561),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1585),
.B(n_1549),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1587),
.B(n_1549),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1572),
.A2(n_1556),
.B1(n_1529),
.B2(n_1536),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1568),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1592),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1598),
.B(n_1558),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1587),
.B(n_1566),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1566),
.B(n_1492),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1564),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1584),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1578),
.Y(n_1645)
);

INVxp67_ASAP7_75t_SL g1646 ( 
.A(n_1581),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1578),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1597),
.B(n_1611),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1577),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1588),
.B(n_1492),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_SL g1651 ( 
.A(n_1581),
.B(n_1538),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1629),
.B(n_1475),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1619),
.B(n_1588),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1634),
.B(n_1606),
.Y(n_1654)
);

NAND3xp33_ASAP7_75t_L g1655 ( 
.A(n_1615),
.B(n_1563),
.C(n_1523),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1627),
.Y(n_1656)
);

INVxp67_ASAP7_75t_SL g1657 ( 
.A(n_1623),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1625),
.B(n_1596),
.Y(n_1658)
);

NOR2x1p5_ASAP7_75t_L g1659 ( 
.A(n_1640),
.B(n_1317),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1634),
.B(n_1582),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1627),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1613),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1614),
.Y(n_1663)
);

OAI22xp33_ASAP7_75t_SL g1664 ( 
.A1(n_1651),
.A2(n_1581),
.B1(n_1609),
.B2(n_1602),
.Y(n_1664)
);

INVx2_ASAP7_75t_SL g1665 ( 
.A(n_1622),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1640),
.B(n_1612),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1616),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1631),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1639),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1637),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1619),
.B(n_1588),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1645),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1647),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1648),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1633),
.B(n_1579),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1633),
.B(n_1579),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1630),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1626),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1643),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1633),
.B(n_1580),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1644),
.B(n_1596),
.Y(n_1681)
);

INVx4_ASAP7_75t_L g1682 ( 
.A(n_1618),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1628),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1612),
.B(n_1617),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1617),
.B(n_1604),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1632),
.B(n_1604),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1628),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1632),
.B(n_1280),
.Y(n_1688)
);

OR2x6_ASAP7_75t_L g1689 ( 
.A(n_1618),
.B(n_1498),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1638),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1622),
.B(n_1580),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1620),
.B(n_1582),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1638),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1649),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1678),
.B(n_1594),
.Y(n_1695)
);

NAND3xp33_ASAP7_75t_L g1696 ( 
.A(n_1670),
.B(n_1618),
.C(n_1283),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1678),
.B(n_1594),
.Y(n_1697)
);

INVxp67_ASAP7_75t_SL g1698 ( 
.A(n_1657),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1661),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1675),
.B(n_1618),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1675),
.B(n_1646),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1661),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1666),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1655),
.A2(n_1622),
.B1(n_1562),
.B2(n_1650),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1664),
.B(n_1650),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1676),
.B(n_1650),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1659),
.A2(n_1461),
.B1(n_1462),
.B2(n_1385),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1656),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1677),
.B(n_1620),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1688),
.Y(n_1710)
);

BUFx3_ASAP7_75t_L g1711 ( 
.A(n_1652),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1676),
.B(n_1621),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1662),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1680),
.B(n_1621),
.Y(n_1714)
);

NAND2x1p5_ASAP7_75t_L g1715 ( 
.A(n_1682),
.B(n_1456),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1684),
.B(n_1609),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1674),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1679),
.B(n_1648),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1668),
.B(n_1603),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1663),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1688),
.A2(n_1462),
.B1(n_1635),
.B2(n_1636),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1658),
.B(n_1635),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1652),
.B(n_1283),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1660),
.B(n_1600),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1674),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1654),
.A2(n_1462),
.B1(n_1374),
.B2(n_1385),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1682),
.B(n_1286),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1667),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_1682),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1680),
.B(n_1624),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1703),
.B(n_1669),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1702),
.Y(n_1732)
);

OAI21xp5_ASAP7_75t_SL g1733 ( 
.A1(n_1696),
.A2(n_1665),
.B(n_1653),
.Y(n_1733)
);

O2A1O1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1698),
.A2(n_1689),
.B(n_1665),
.C(n_1685),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1706),
.B(n_1653),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1703),
.B(n_1681),
.Y(n_1736)
);

OAI311xp33_ASAP7_75t_L g1737 ( 
.A1(n_1696),
.A2(n_1686),
.A3(n_1671),
.B1(n_1692),
.C1(n_1673),
.Y(n_1737)
);

OAI32xp33_ASAP7_75t_L g1738 ( 
.A1(n_1705),
.A2(n_1671),
.A3(n_1672),
.B1(n_1590),
.B2(n_1690),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1710),
.B(n_1691),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1718),
.B(n_1694),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1702),
.Y(n_1741)
);

OAI21xp5_ASAP7_75t_SL g1742 ( 
.A1(n_1727),
.A2(n_1691),
.B(n_1636),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1702),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1704),
.A2(n_1689),
.B1(n_1472),
.B2(n_1500),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1722),
.B(n_1683),
.Y(n_1745)
);

OAI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1711),
.A2(n_1689),
.B1(n_1693),
.B2(n_1687),
.C(n_1573),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1711),
.A2(n_1689),
.B1(n_1559),
.B2(n_1444),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1729),
.B(n_1641),
.Y(n_1748)
);

NOR2xp67_ASAP7_75t_SL g1749 ( 
.A(n_1711),
.B(n_1317),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1706),
.B(n_1624),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1729),
.B(n_1641),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1721),
.A2(n_1590),
.B1(n_1603),
.B2(n_1494),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1723),
.B(n_1286),
.Y(n_1753)
);

BUFx2_ASAP7_75t_L g1754 ( 
.A(n_1700),
.Y(n_1754)
);

XOR2x2_ASAP7_75t_L g1755 ( 
.A(n_1721),
.B(n_1322),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1716),
.B(n_1307),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1700),
.A2(n_1492),
.B1(n_1574),
.B2(n_1404),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1754),
.B(n_1739),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1753),
.B(n_1701),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1744),
.A2(n_1701),
.B1(n_1716),
.B2(n_1709),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1735),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1733),
.B(n_1712),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1750),
.B(n_1712),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1732),
.Y(n_1764)
);

CKINVDCx16_ASAP7_75t_R g1765 ( 
.A(n_1756),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1741),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1743),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1736),
.B(n_1695),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1731),
.B(n_1714),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1731),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1734),
.B(n_1715),
.Y(n_1771)
);

NAND2x1_ASAP7_75t_SL g1772 ( 
.A(n_1747),
.B(n_1699),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1744),
.A2(n_1709),
.B1(n_1724),
.B2(n_1717),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1742),
.B(n_1714),
.Y(n_1774)
);

INVx2_ASAP7_75t_SL g1775 ( 
.A(n_1748),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1751),
.B(n_1695),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1740),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1749),
.B(n_1730),
.Y(n_1778)
);

NAND3xp33_ASAP7_75t_SL g1779 ( 
.A(n_1771),
.B(n_1737),
.C(n_1715),
.Y(n_1779)
);

AOI21xp33_ASAP7_75t_L g1780 ( 
.A1(n_1759),
.A2(n_1738),
.B(n_1746),
.Y(n_1780)
);

NOR3xp33_ASAP7_75t_L g1781 ( 
.A(n_1765),
.B(n_1745),
.C(n_1752),
.Y(n_1781)
);

AOI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1771),
.A2(n_1755),
.B(n_1697),
.Y(n_1782)
);

OAI221xp5_ASAP7_75t_L g1783 ( 
.A1(n_1772),
.A2(n_1707),
.B1(n_1715),
.B2(n_1752),
.C(n_1757),
.Y(n_1783)
);

AOI322xp5_ASAP7_75t_L g1784 ( 
.A1(n_1762),
.A2(n_1699),
.A3(n_1720),
.B1(n_1728),
.B2(n_1713),
.C1(n_1708),
.C2(n_1697),
.Y(n_1784)
);

NAND4xp25_ASAP7_75t_SL g1785 ( 
.A(n_1760),
.B(n_1726),
.C(n_1730),
.D(n_1717),
.Y(n_1785)
);

OAI221xp5_ASAP7_75t_L g1786 ( 
.A1(n_1774),
.A2(n_1758),
.B1(n_1773),
.B2(n_1769),
.C(n_1777),
.Y(n_1786)
);

AOI221xp5_ASAP7_75t_L g1787 ( 
.A1(n_1770),
.A2(n_1775),
.B1(n_1761),
.B2(n_1768),
.C(n_1767),
.Y(n_1787)
);

AOI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1778),
.A2(n_1720),
.B(n_1713),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1761),
.A2(n_1725),
.B1(n_1717),
.B2(n_1724),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1778),
.A2(n_1728),
.B(n_1725),
.Y(n_1790)
);

AOI221xp5_ASAP7_75t_L g1791 ( 
.A1(n_1775),
.A2(n_1725),
.B1(n_1708),
.B2(n_1719),
.C(n_1590),
.Y(n_1791)
);

CKINVDCx20_ASAP7_75t_R g1792 ( 
.A(n_1768),
.Y(n_1792)
);

NAND5xp2_ASAP7_75t_L g1793 ( 
.A(n_1781),
.B(n_1763),
.C(n_1764),
.D(n_1776),
.E(n_1766),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1782),
.B(n_1763),
.Y(n_1794)
);

AO22x2_ASAP7_75t_L g1795 ( 
.A1(n_1779),
.A2(n_1764),
.B1(n_1766),
.B2(n_1776),
.Y(n_1795)
);

BUFx2_ASAP7_75t_L g1796 ( 
.A(n_1792),
.Y(n_1796)
);

NOR2x1_ASAP7_75t_L g1797 ( 
.A(n_1786),
.B(n_1719),
.Y(n_1797)
);

NOR3xp33_ASAP7_75t_L g1798 ( 
.A(n_1780),
.B(n_1787),
.C(n_1785),
.Y(n_1798)
);

NOR4xp75_ASAP7_75t_L g1799 ( 
.A(n_1783),
.B(n_1590),
.C(n_1452),
.D(n_1307),
.Y(n_1799)
);

NOR2x1_ASAP7_75t_L g1800 ( 
.A(n_1790),
.B(n_1307),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1788),
.Y(n_1801)
);

NOR3xp33_ASAP7_75t_SL g1802 ( 
.A(n_1791),
.B(n_1569),
.C(n_1454),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1789),
.Y(n_1803)
);

NOR3x1_ASAP7_75t_L g1804 ( 
.A(n_1784),
.B(n_1452),
.C(n_1600),
.Y(n_1804)
);

NAND4xp75_ASAP7_75t_L g1805 ( 
.A(n_1797),
.B(n_1411),
.C(n_1601),
.D(n_1642),
.Y(n_1805)
);

NOR3xp33_ASAP7_75t_L g1806 ( 
.A(n_1796),
.B(n_1601),
.C(n_1583),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1803),
.B(n_1642),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1800),
.B(n_1565),
.Y(n_1808)
);

AOI211xp5_ASAP7_75t_SL g1809 ( 
.A1(n_1798),
.A2(n_1433),
.B(n_1601),
.C(n_1427),
.Y(n_1809)
);

AOI221x1_ASAP7_75t_L g1810 ( 
.A1(n_1795),
.A2(n_1583),
.B1(n_1574),
.B2(n_1593),
.C(n_1607),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1807),
.Y(n_1811)
);

AOI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1808),
.A2(n_1795),
.B1(n_1794),
.B2(n_1801),
.Y(n_1812)
);

AOI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1805),
.A2(n_1802),
.B1(n_1793),
.B2(n_1799),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1806),
.B(n_1804),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1810),
.Y(n_1815)
);

AO22x2_ASAP7_75t_L g1816 ( 
.A1(n_1809),
.A2(n_1603),
.B1(n_1574),
.B2(n_1602),
.Y(n_1816)
);

NOR3xp33_ASAP7_75t_SL g1817 ( 
.A(n_1809),
.B(n_1429),
.C(n_1432),
.Y(n_1817)
);

NAND4xp75_ASAP7_75t_L g1818 ( 
.A(n_1812),
.B(n_1411),
.C(n_1565),
.D(n_1443),
.Y(n_1818)
);

NAND3xp33_ASAP7_75t_L g1819 ( 
.A(n_1815),
.B(n_1811),
.C(n_1813),
.Y(n_1819)
);

AOI221x1_ASAP7_75t_L g1820 ( 
.A1(n_1816),
.A2(n_1574),
.B1(n_1577),
.B2(n_1429),
.C(n_1432),
.Y(n_1820)
);

NOR3xp33_ASAP7_75t_L g1821 ( 
.A(n_1814),
.B(n_1390),
.C(n_1411),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1817),
.Y(n_1822)
);

AOI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1813),
.A2(n_1494),
.B1(n_1492),
.B2(n_1439),
.Y(n_1823)
);

NAND4xp75_ASAP7_75t_L g1824 ( 
.A(n_1822),
.B(n_1611),
.C(n_1597),
.D(n_1471),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1818),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1821),
.B(n_1567),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1825),
.Y(n_1827)
);

NAND5xp2_ASAP7_75t_L g1828 ( 
.A(n_1827),
.B(n_1823),
.C(n_1819),
.D(n_1824),
.E(n_1826),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1828),
.A2(n_1824),
.B1(n_1820),
.B2(n_1410),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1828),
.A2(n_1410),
.B1(n_1390),
.B2(n_1437),
.Y(n_1830)
);

OAI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1829),
.A2(n_1599),
.B(n_1436),
.Y(n_1831)
);

OAI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1830),
.A2(n_1599),
.B1(n_1456),
.B2(n_1494),
.Y(n_1832)
);

AO221x1_ASAP7_75t_L g1833 ( 
.A1(n_1832),
.A2(n_1831),
.B1(n_1393),
.B2(n_1427),
.C(n_1453),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1832),
.A2(n_1437),
.B(n_1436),
.Y(n_1834)
);

NOR2x1_ASAP7_75t_L g1835 ( 
.A(n_1834),
.B(n_1390),
.Y(n_1835)
);

AOI22xp5_ASAP7_75t_SL g1836 ( 
.A1(n_1835),
.A2(n_1833),
.B1(n_1390),
.B2(n_1427),
.Y(n_1836)
);

OAI221xp5_ASAP7_75t_R g1837 ( 
.A1(n_1836),
.A2(n_1437),
.B1(n_1456),
.B2(n_1469),
.C(n_1499),
.Y(n_1837)
);

AOI211xp5_ASAP7_75t_L g1838 ( 
.A1(n_1837),
.A2(n_1453),
.B(n_1393),
.C(n_1427),
.Y(n_1838)
);


endmodule