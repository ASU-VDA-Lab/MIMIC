module fake_netlist_6_1849_n_1794 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1794);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1794;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_1214;
wire n_835;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_130),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_97),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_19),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_55),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_77),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_38),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_80),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_134),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_18),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_157),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_106),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_57),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_132),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_42),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_83),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_173),
.Y(n_191)
);

INVxp67_ASAP7_75t_SL g192 ( 
.A(n_22),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_138),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_24),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_85),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_136),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_8),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_119),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_166),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_92),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_87),
.Y(n_202)
);

INVxp67_ASAP7_75t_SL g203 ( 
.A(n_143),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_90),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_145),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_146),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_144),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_58),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_76),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_108),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_127),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_161),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_46),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_61),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_86),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_55),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_5),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_40),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_150),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_114),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_69),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_135),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_58),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_79),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_109),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_9),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_162),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_54),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_53),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_28),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_12),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_24),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_74),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_158),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_13),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_96),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_7),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_152),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_43),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_103),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_88),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_153),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_128),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_154),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_169),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_67),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_68),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_51),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_29),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_71),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_93),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_41),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_72),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_33),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_131),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_160),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_40),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_34),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_147),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_174),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_8),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_149),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_142),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_29),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_156),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_39),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_7),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_141),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_49),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_3),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_101),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_12),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_155),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_139),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_82),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_38),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_148),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_129),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_37),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_120),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_94),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_4),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_75),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_57),
.Y(n_284)
);

BUFx8_ASAP7_75t_SL g285 ( 
.A(n_28),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_104),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_14),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_50),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_100),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_2),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_56),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_124),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_122),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_105),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_95),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_89),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_32),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_13),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_123),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_111),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_98),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_22),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_5),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_60),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_60),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_43),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_14),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_102),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_30),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_65),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_6),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_20),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_112),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_140),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_78),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_118),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_4),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_64),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_84),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_36),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_20),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_51),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_23),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_117),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_165),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_27),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_3),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_107),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_23),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_2),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_56),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_63),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_171),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_113),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_121),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_62),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_25),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_59),
.Y(n_338)
);

BUFx10_ASAP7_75t_L g339 ( 
.A(n_50),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_151),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_116),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_15),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_21),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_34),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_168),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_49),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_0),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_32),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_167),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_81),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_17),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_27),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_39),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_133),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_30),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_53),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_187),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_312),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_187),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_190),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_285),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_235),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_262),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_217),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_199),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_201),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_235),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_218),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_327),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_327),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_229),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_339),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_276),
.B(n_0),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_230),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_237),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_206),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_194),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_233),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_276),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_344),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_208),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_176),
.B(n_1),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_216),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_262),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_241),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_226),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_248),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_252),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_207),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_257),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_258),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_316),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_268),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_264),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_339),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_178),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_228),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_231),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_259),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_313),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_232),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_266),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_268),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_249),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_267),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_270),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_281),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_234),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_254),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_220),
.B(n_341),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_178),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_288),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_302),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_304),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_305),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_317),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_272),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_322),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_323),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_281),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_279),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_220),
.B(n_1),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_330),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_282),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_284),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_286),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_346),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_205),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_347),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_224),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_225),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_236),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_353),
.B(n_6),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_222),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_283),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_180),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_240),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_242),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_202),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_179),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_287),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_341),
.B(n_9),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_204),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_243),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_244),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_245),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_290),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_291),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_246),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_261),
.B(n_10),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_363),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_431),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_411),
.B(n_289),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_432),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_433),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_358),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_363),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_438),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_364),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_383),
.B(n_437),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_364),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_423),
.B(n_318),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_436),
.Y(n_464)
);

AND2x2_ASAP7_75t_SL g465 ( 
.A(n_383),
.B(n_283),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_360),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_436),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_439),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_365),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_404),
.B(n_325),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_366),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_445),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_385),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_412),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_394),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_440),
.B(n_325),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_394),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_382),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_444),
.B(n_210),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_385),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_376),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_382),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_R g483 ( 
.A(n_368),
.B(n_247),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_379),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_446),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_384),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_384),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_379),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_368),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_447),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_443),
.B(n_408),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_450),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_380),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_361),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_420),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_361),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_380),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_381),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_371),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_441),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_408),
.B(n_177),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_371),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_374),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_381),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_421),
.B(n_215),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_409),
.B(n_427),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_377),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_387),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_398),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_374),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_397),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_399),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_402),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_429),
.B(n_349),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_405),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_378),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_410),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_397),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_451),
.A2(n_356),
.B1(n_269),
.B2(n_239),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_393),
.B(n_375),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_413),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_414),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_375),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_415),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_416),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_386),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_417),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_388),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_419),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_461),
.B(n_388),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_452),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_458),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_465),
.A2(n_434),
.B1(n_373),
.B2(n_421),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_465),
.A2(n_434),
.B1(n_424),
.B2(n_430),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_475),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_463),
.A2(n_390),
.B1(n_400),
.B2(n_401),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_507),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_507),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_452),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_524),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_463),
.A2(n_418),
.B1(n_449),
.B2(n_448),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_452),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_465),
.A2(n_451),
.B1(n_449),
.B2(n_448),
.Y(n_543)
);

INVx5_ASAP7_75t_L g544 ( 
.A(n_452),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_454),
.B(n_389),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_461),
.B(n_389),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_508),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_458),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_508),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_470),
.B(n_357),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_480),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_R g552 ( 
.A(n_460),
.B(n_462),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_470),
.B(n_359),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_458),
.Y(n_554)
);

NAND2xp33_ASAP7_75t_L g555 ( 
.A(n_491),
.B(n_197),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_511),
.B(n_372),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_524),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_454),
.B(n_391),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_511),
.B(n_396),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_473),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_514),
.B(n_197),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_475),
.B(n_428),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_480),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_475),
.B(n_362),
.Y(n_564)
);

BUFx8_ASAP7_75t_SL g565 ( 
.A(n_466),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_L g566 ( 
.A(n_491),
.B(n_197),
.Y(n_566)
);

BUFx8_ASAP7_75t_SL g567 ( 
.A(n_469),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_477),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_524),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_473),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_461),
.B(n_470),
.Y(n_571)
);

NAND3xp33_ASAP7_75t_L g572 ( 
.A(n_518),
.B(n_392),
.C(n_391),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_453),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_520),
.B(n_392),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_473),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_520),
.B(n_395),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_498),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_480),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_471),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_498),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_524),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_498),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_512),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_505),
.B(n_197),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_513),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_513),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_474),
.A2(n_442),
.B1(n_395),
.B2(n_426),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_521),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_476),
.B(n_367),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_521),
.Y(n_590)
);

INVxp33_ASAP7_75t_L g591 ( 
.A(n_457),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_498),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_501),
.B(n_403),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_524),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_498),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_498),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_477),
.B(n_369),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_476),
.B(n_479),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_484),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_484),
.Y(n_600)
);

OAI22xp33_ASAP7_75t_L g601 ( 
.A1(n_518),
.A2(n_342),
.B1(n_307),
.B2(n_306),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_525),
.Y(n_602)
);

AND2x2_ASAP7_75t_SL g603 ( 
.A(n_460),
.B(n_197),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_529),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_457),
.B(n_435),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_479),
.B(n_403),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_479),
.B(n_406),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_462),
.B(n_370),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_529),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_478),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_484),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_505),
.B(n_406),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_505),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_474),
.B(n_407),
.Y(n_614)
);

BUFx8_ASAP7_75t_SL g615 ( 
.A(n_481),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_478),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_482),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_500),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_484),
.Y(n_619)
);

AND2x6_ASAP7_75t_L g620 ( 
.A(n_476),
.B(n_280),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_482),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_488),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_505),
.A2(n_295),
.B1(n_280),
.B2(n_192),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_517),
.B(n_407),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_486),
.B(n_219),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_487),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_488),
.Y(n_627)
);

XOR2xp5_ASAP7_75t_L g628 ( 
.A(n_516),
.B(n_418),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_526),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_488),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_455),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_517),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_502),
.B(n_422),
.Y(n_633)
);

BUFx8_ASAP7_75t_SL g634 ( 
.A(n_456),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_483),
.B(n_280),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_464),
.B(n_435),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_493),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_493),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_500),
.B(n_422),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_495),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_509),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_464),
.B(n_425),
.Y(n_642)
);

AND2x6_ASAP7_75t_L g643 ( 
.A(n_467),
.B(n_280),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_493),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_467),
.B(n_425),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_509),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_493),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_509),
.B(n_515),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_497),
.Y(n_649)
);

AND2x6_ASAP7_75t_L g650 ( 
.A(n_515),
.B(n_280),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_515),
.A2(n_295),
.B1(n_350),
.B2(n_335),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_522),
.A2(n_295),
.B1(n_333),
.B2(n_319),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_489),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_522),
.A2(n_295),
.B1(n_296),
.B2(n_221),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_522),
.Y(n_655)
);

BUFx10_ASAP7_75t_L g656 ( 
.A(n_494),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_497),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_483),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_527),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_504),
.B(n_426),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_527),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_497),
.Y(n_662)
);

INVx4_ASAP7_75t_L g663 ( 
.A(n_504),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_503),
.B(n_295),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_545),
.B(n_558),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_605),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_618),
.B(n_489),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_603),
.A2(n_528),
.B1(n_523),
.B2(n_510),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_537),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_603),
.B(n_499),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_614),
.Y(n_671)
);

AND2x2_ASAP7_75t_SL g672 ( 
.A(n_555),
.B(n_499),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_571),
.B(n_203),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_598),
.A2(n_561),
.B1(n_625),
.B2(n_663),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_532),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_593),
.B(n_506),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_619),
.B(n_262),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_574),
.B(n_177),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_538),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_532),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_598),
.B(n_227),
.Y(n_681)
);

BUFx6f_ASAP7_75t_SL g682 ( 
.A(n_656),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_576),
.B(n_182),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_548),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_645),
.B(n_182),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_655),
.B(n_238),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_606),
.B(n_183),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_547),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_605),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_655),
.B(n_253),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_549),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_607),
.B(n_183),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_619),
.B(n_256),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_619),
.B(n_260),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_543),
.B(n_185),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_533),
.A2(n_265),
.B1(n_263),
.B2(n_274),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_647),
.B(n_262),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_647),
.B(n_275),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_647),
.B(n_292),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_L g700 ( 
.A(n_624),
.B(n_262),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_610),
.B(n_294),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_561),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_616),
.B(n_315),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_583),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_554),
.Y(n_705)
);

INVxp33_ASAP7_75t_L g706 ( 
.A(n_591),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_618),
.B(n_519),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_554),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_625),
.A2(n_519),
.B1(n_262),
.B2(n_222),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_613),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_572),
.B(n_468),
.C(n_492),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_638),
.B(n_530),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_552),
.Y(n_713)
);

CKINVDCx11_ASAP7_75t_R g714 ( 
.A(n_656),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_617),
.B(n_250),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_621),
.B(n_251),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_626),
.B(n_255),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_546),
.B(n_185),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_585),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_568),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_560),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_586),
.Y(n_722)
);

AND2x6_ASAP7_75t_SL g723 ( 
.A(n_633),
.B(n_213),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_556),
.B(n_459),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_640),
.B(n_632),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_556),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_560),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_570),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_632),
.B(n_271),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_R g730 ( 
.A(n_573),
.B(n_472),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_570),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_613),
.B(n_66),
.Y(n_732)
);

OAI221xp5_ASAP7_75t_L g733 ( 
.A1(n_534),
.A2(n_309),
.B1(n_298),
.B2(n_297),
.C(n_348),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_535),
.B(n_273),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_642),
.B(n_485),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_588),
.B(n_590),
.Y(n_736)
);

OR2x6_ASAP7_75t_L g737 ( 
.A(n_608),
.B(n_490),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_638),
.B(n_599),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_541),
.B(n_186),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_602),
.B(n_277),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_575),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_638),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_604),
.B(n_278),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_609),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_562),
.Y(n_745)
);

OAI22xp33_ASAP7_75t_L g746 ( 
.A1(n_559),
.A2(n_329),
.B1(n_303),
.B2(n_223),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_550),
.A2(n_179),
.B1(n_355),
.B2(n_184),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_636),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_575),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_638),
.B(n_293),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_642),
.B(n_496),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_562),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_559),
.B(n_639),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_553),
.B(n_531),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_568),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_660),
.B(n_188),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_649),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_660),
.B(n_188),
.Y(n_758)
);

OAI22xp33_ASAP7_75t_L g759 ( 
.A1(n_612),
.A2(n_181),
.B1(n_352),
.B2(n_351),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_649),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_564),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_564),
.A2(n_310),
.B1(n_308),
.B2(n_345),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_623),
.A2(n_321),
.B1(n_352),
.B2(n_351),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_597),
.Y(n_764)
);

NAND3xp33_ASAP7_75t_L g765 ( 
.A(n_587),
.B(n_664),
.C(n_639),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_664),
.B(n_191),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_658),
.B(n_191),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_599),
.B(n_600),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_539),
.B(n_193),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_653),
.B(n_184),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_591),
.B(n_608),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_597),
.Y(n_772)
);

NOR3xp33_ASAP7_75t_L g773 ( 
.A(n_601),
.B(n_321),
.C(n_343),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_539),
.B(n_193),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_539),
.B(n_195),
.Y(n_775)
);

INVx8_ASAP7_75t_L g776 ( 
.A(n_608),
.Y(n_776)
);

NOR2xp67_ASAP7_75t_L g777 ( 
.A(n_536),
.B(n_195),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_611),
.B(n_622),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_551),
.B(n_563),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_597),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_551),
.B(n_196),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_622),
.B(n_196),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_551),
.B(n_200),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_SL g784 ( 
.A(n_573),
.B(n_200),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_589),
.B(n_339),
.Y(n_785)
);

NOR2xp67_ASAP7_75t_SL g786 ( 
.A(n_635),
.B(n_209),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_563),
.B(n_209),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_563),
.B(n_211),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_578),
.B(n_211),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_555),
.A2(n_189),
.B1(n_343),
.B2(n_198),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_589),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_635),
.A2(n_608),
.B1(n_566),
.B2(n_584),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_566),
.A2(n_354),
.B(n_340),
.C(n_212),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_648),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_578),
.B(n_340),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_620),
.A2(n_189),
.B1(n_337),
.B2(n_198),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_641),
.B(n_212),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_646),
.B(n_91),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_R g799 ( 
.A(n_631),
.B(n_338),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_710),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_665),
.B(n_629),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_678),
.A2(n_644),
.B(n_627),
.C(n_630),
.Y(n_802)
);

OAI21x1_ASAP7_75t_L g803 ( 
.A1(n_779),
.A2(n_630),
.B(n_637),
.Y(n_803)
);

NOR2xp67_ASAP7_75t_L g804 ( 
.A(n_668),
.B(n_659),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_794),
.A2(n_627),
.B(n_637),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_754),
.A2(n_644),
.B(n_577),
.Y(n_806)
);

BUFx8_ASAP7_75t_L g807 ( 
.A(n_682),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_667),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_707),
.B(n_656),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_730),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_673),
.A2(n_577),
.B(n_580),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_751),
.B(n_628),
.Y(n_812)
);

AOI21x1_ASAP7_75t_L g813 ( 
.A1(n_712),
.A2(n_580),
.B(n_661),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_670),
.A2(n_657),
.B(n_654),
.C(n_652),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_735),
.B(n_579),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_671),
.B(n_579),
.Y(n_816)
);

OAI321xp33_ASAP7_75t_L g817 ( 
.A1(n_695),
.A2(n_683),
.A3(n_678),
.B1(n_709),
.B2(n_739),
.C(n_733),
.Y(n_817)
);

O2A1O1Ixp5_ASAP7_75t_L g818 ( 
.A1(n_683),
.A2(n_592),
.B(n_582),
.C(n_569),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_666),
.Y(n_819)
);

OAI21xp33_ASAP7_75t_L g820 ( 
.A1(n_739),
.A2(n_338),
.B(n_311),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_670),
.A2(n_657),
.B(n_651),
.C(n_592),
.Y(n_821)
);

AOI21x1_ASAP7_75t_L g822 ( 
.A1(n_738),
.A2(n_581),
.B(n_596),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_685),
.B(n_662),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_685),
.B(n_662),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_687),
.B(n_692),
.Y(n_825)
);

NOR2xp67_ASAP7_75t_L g826 ( 
.A(n_713),
.B(n_582),
.Y(n_826)
);

AND2x6_ASAP7_75t_L g827 ( 
.A(n_732),
.B(n_540),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_687),
.B(n_620),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_692),
.B(n_620),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_718),
.B(n_595),
.Y(n_830)
);

A2O1A1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_766),
.A2(n_214),
.B(n_336),
.C(n_314),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_771),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_674),
.A2(n_326),
.B1(n_337),
.B2(n_320),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_676),
.A2(n_732),
.B1(n_718),
.B2(n_765),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_756),
.B(n_540),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_710),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_780),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_681),
.B(n_540),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_689),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_785),
.B(n_311),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_756),
.B(n_557),
.Y(n_841)
);

OA21x2_ASAP7_75t_L g842 ( 
.A1(n_693),
.A2(n_334),
.B(n_314),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_706),
.B(n_565),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_758),
.B(n_320),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_758),
.B(n_326),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_768),
.A2(n_643),
.B(n_650),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_766),
.A2(n_695),
.B(n_792),
.C(n_748),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_737),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_706),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_672),
.A2(n_331),
.B1(n_324),
.B2(n_328),
.Y(n_850)
);

NAND2xp33_ASAP7_75t_L g851 ( 
.A(n_725),
.B(n_557),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_726),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_791),
.A2(n_214),
.B(n_324),
.C(n_328),
.Y(n_853)
);

A2O1A1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_669),
.A2(n_332),
.B(n_334),
.C(n_336),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_679),
.Y(n_855)
);

INVx1_ASAP7_75t_SL g856 ( 
.A(n_753),
.Y(n_856)
);

NOR2x1p5_ASAP7_75t_SL g857 ( 
.A(n_757),
.B(n_594),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_720),
.B(n_542),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_780),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_720),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_688),
.B(n_544),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_675),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_672),
.B(n_761),
.Y(n_863)
);

CKINVDCx10_ASAP7_75t_R g864 ( 
.A(n_682),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_755),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_680),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_691),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_767),
.B(n_565),
.Y(n_868)
);

AND2x6_ASAP7_75t_L g869 ( 
.A(n_732),
.B(n_643),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_696),
.A2(n_331),
.B1(n_332),
.B2(n_542),
.Y(n_870)
);

NOR2x1_ASAP7_75t_L g871 ( 
.A(n_755),
.B(n_634),
.Y(n_871)
);

O2A1O1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_782),
.A2(n_10),
.B(n_11),
.C(n_15),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_704),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_729),
.A2(n_542),
.B(n_650),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_719),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_798),
.Y(n_876)
);

NOR3xp33_ASAP7_75t_L g877 ( 
.A(n_746),
.B(n_567),
.C(n_615),
.Y(n_877)
);

CKINVDCx11_ASAP7_75t_R g878 ( 
.A(n_714),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_764),
.B(n_73),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_736),
.A2(n_650),
.B(n_643),
.Y(n_880)
);

AO22x1_ASAP7_75t_L g881 ( 
.A1(n_773),
.A2(n_643),
.B1(n_650),
.B2(n_634),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_702),
.A2(n_11),
.B1(n_16),
.B2(n_17),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_722),
.A2(n_643),
.B1(n_650),
.B2(n_615),
.Y(n_883)
);

AOI21x1_ASAP7_75t_L g884 ( 
.A1(n_768),
.A2(n_70),
.B(n_175),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_770),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_714),
.Y(n_886)
);

BUFx12f_ASAP7_75t_L g887 ( 
.A(n_737),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_684),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_767),
.B(n_567),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_778),
.A2(n_172),
.B(n_170),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_778),
.A2(n_164),
.B(n_163),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_734),
.A2(n_159),
.B(n_137),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_677),
.A2(n_126),
.B(n_125),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_744),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_730),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_742),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_742),
.Y(n_897)
);

NOR2xp67_ASAP7_75t_L g898 ( 
.A(n_724),
.B(n_115),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_763),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_784),
.B(n_99),
.Y(n_900)
);

O2A1O1Ixp5_ASAP7_75t_L g901 ( 
.A1(n_750),
.A2(n_25),
.B(n_26),
.C(n_31),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_745),
.A2(n_31),
.B(n_33),
.C(n_35),
.Y(n_902)
);

AO21x1_ASAP7_75t_L g903 ( 
.A1(n_700),
.A2(n_35),
.B(n_36),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_769),
.A2(n_37),
.B(n_41),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_677),
.A2(n_42),
.B(n_44),
.Y(n_905)
);

O2A1O1Ixp5_ASAP7_75t_L g906 ( 
.A1(n_786),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_697),
.A2(n_45),
.B(n_47),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_782),
.A2(n_47),
.B(n_48),
.C(n_52),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_757),
.B(n_48),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_752),
.B(n_52),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_772),
.B(n_59),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_797),
.B(n_701),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_797),
.A2(n_793),
.B(n_694),
.C(n_698),
.Y(n_913)
);

AO22x1_ASAP7_75t_L g914 ( 
.A1(n_711),
.A2(n_798),
.B1(n_781),
.B2(n_795),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_699),
.A2(n_703),
.B(n_762),
.C(n_686),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_774),
.A2(n_775),
.B(n_789),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_759),
.B(n_740),
.Y(n_917)
);

NOR2xp67_ASAP7_75t_L g918 ( 
.A(n_783),
.B(n_787),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_747),
.B(n_777),
.Y(n_919)
);

CKINVDCx10_ASAP7_75t_R g920 ( 
.A(n_737),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_743),
.B(n_715),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_788),
.A2(n_690),
.B(n_716),
.Y(n_922)
);

AND2x6_ASAP7_75t_L g923 ( 
.A(n_798),
.B(n_760),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_796),
.A2(n_790),
.B1(n_776),
.B2(n_708),
.Y(n_924)
);

INVx6_ASAP7_75t_L g925 ( 
.A(n_776),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_717),
.B(n_705),
.Y(n_926)
);

AOI21xp33_ASAP7_75t_L g927 ( 
.A1(n_799),
.A2(n_705),
.B(n_708),
.Y(n_927)
);

BUFx4f_ASAP7_75t_L g928 ( 
.A(n_776),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_723),
.B(n_721),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_727),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_728),
.B(n_731),
.Y(n_931)
);

CKINVDCx6p67_ASAP7_75t_R g932 ( 
.A(n_799),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_741),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_749),
.B(n_665),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_665),
.B(n_794),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_665),
.A2(n_533),
.B1(n_709),
.B2(n_603),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_665),
.B(n_678),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_665),
.B(n_603),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_667),
.B(n_707),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_665),
.B(n_678),
.Y(n_940)
);

OR2x6_ASAP7_75t_L g941 ( 
.A(n_925),
.B(n_887),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_849),
.Y(n_942)
);

OAI22x1_ASAP7_75t_L g943 ( 
.A1(n_834),
.A2(n_940),
.B1(n_937),
.B2(n_801),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_935),
.B(n_825),
.Y(n_944)
);

OA22x2_ASAP7_75t_L g945 ( 
.A1(n_936),
.A2(n_820),
.B1(n_856),
.B2(n_899),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_808),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_939),
.B(n_809),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_935),
.B(n_817),
.Y(n_948)
);

NAND2x1_ASAP7_75t_SL g949 ( 
.A(n_919),
.B(n_871),
.Y(n_949)
);

NAND2xp33_ASAP7_75t_L g950 ( 
.A(n_876),
.B(n_827),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_936),
.A2(n_847),
.B1(n_938),
.B2(n_934),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_865),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_876),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_921),
.B(n_912),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_852),
.B(n_816),
.Y(n_955)
);

AND2x2_ASAP7_75t_SL g956 ( 
.A(n_877),
.B(n_928),
.Y(n_956)
);

AOI221x1_ASAP7_75t_L g957 ( 
.A1(n_913),
.A2(n_916),
.B1(n_835),
.B2(n_841),
.C(n_823),
.Y(n_957)
);

AO22x1_ASAP7_75t_L g958 ( 
.A1(n_899),
.A2(n_812),
.B1(n_905),
.B2(n_907),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_838),
.A2(n_824),
.B(n_830),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_837),
.B(n_917),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_844),
.B(n_845),
.Y(n_961)
);

INVx1_ASAP7_75t_SL g962 ( 
.A(n_832),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_855),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_840),
.B(n_885),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_838),
.A2(n_922),
.B(n_851),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_806),
.A2(n_818),
.B(n_802),
.Y(n_966)
);

AO31x2_ASAP7_75t_L g967 ( 
.A1(n_903),
.A2(n_915),
.A3(n_828),
.B(n_829),
.Y(n_967)
);

AO21x1_ASAP7_75t_L g968 ( 
.A1(n_905),
.A2(n_907),
.B(n_908),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_839),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_867),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_815),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_932),
.B(n_889),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_876),
.A2(n_873),
.B1(n_875),
.B2(n_894),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_819),
.B(n_868),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_918),
.A2(n_804),
.B(n_814),
.C(n_831),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_811),
.A2(n_805),
.B(n_821),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_860),
.B(n_865),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_865),
.Y(n_978)
);

BUFx2_ASAP7_75t_SL g979 ( 
.A(n_886),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_923),
.B(n_926),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_SL g981 ( 
.A1(n_882),
.A2(n_872),
.B(n_893),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_923),
.B(n_926),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_927),
.A2(n_909),
.B(n_924),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_837),
.B(n_898),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_800),
.A2(n_836),
.B(n_863),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_810),
.Y(n_986)
);

BUFx2_ASAP7_75t_L g987 ( 
.A(n_848),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_929),
.B(n_895),
.Y(n_988)
);

OAI22xp33_ASAP7_75t_L g989 ( 
.A1(n_910),
.A2(n_911),
.B1(n_859),
.B2(n_837),
.Y(n_989)
);

OAI21x1_ASAP7_75t_L g990 ( 
.A1(n_896),
.A2(n_897),
.B(n_884),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_896),
.A2(n_897),
.B(n_874),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_853),
.A2(n_924),
.B(n_893),
.C(n_854),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_923),
.B(n_827),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_858),
.Y(n_994)
);

AO31x2_ASAP7_75t_L g995 ( 
.A1(n_909),
.A2(n_902),
.A3(n_904),
.B(n_880),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_864),
.Y(n_996)
);

NAND2x1p5_ASAP7_75t_L g997 ( 
.A(n_859),
.B(n_928),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_862),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_923),
.B(n_827),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_866),
.Y(n_1000)
);

AOI21x1_ASAP7_75t_L g1001 ( 
.A1(n_861),
.A2(n_826),
.B(n_888),
.Y(n_1001)
);

BUFx4_ASAP7_75t_SL g1002 ( 
.A(n_920),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_827),
.B(n_933),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_858),
.B(n_879),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_930),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_879),
.B(n_827),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_930),
.Y(n_1007)
);

BUFx2_ASAP7_75t_R g1008 ( 
.A(n_900),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_933),
.B(n_869),
.Y(n_1009)
);

AOI21x1_ASAP7_75t_L g1010 ( 
.A1(n_892),
.A2(n_891),
.B(n_890),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_869),
.B(n_857),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_901),
.A2(n_846),
.B(n_906),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_925),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_869),
.B(n_850),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_883),
.A2(n_842),
.B(n_870),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_869),
.B(n_843),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_850),
.B(n_833),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_842),
.A2(n_870),
.B(n_833),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_925),
.Y(n_1019)
);

AOI21x1_ASAP7_75t_L g1020 ( 
.A1(n_881),
.A2(n_869),
.B(n_807),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_807),
.B(n_878),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_931),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_937),
.B(n_940),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_838),
.A2(n_824),
.B(n_823),
.Y(n_1024)
);

NAND2x1p5_ASAP7_75t_L g1025 ( 
.A(n_876),
.B(n_859),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_855),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_937),
.A2(n_665),
.B1(n_940),
.B2(n_825),
.Y(n_1027)
);

NAND2x1_ASAP7_75t_L g1028 ( 
.A(n_827),
.B(n_923),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_SL g1029 ( 
.A1(n_905),
.A2(n_907),
.B(n_893),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_SL g1030 ( 
.A1(n_905),
.A2(n_907),
.B(n_893),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_803),
.A2(n_822),
.B(n_813),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_939),
.B(n_809),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_865),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_937),
.A2(n_940),
.B(n_817),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_937),
.A2(n_665),
.B(n_940),
.C(n_817),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_937),
.A2(n_665),
.B(n_940),
.C(n_817),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_SL g1037 ( 
.A1(n_905),
.A2(n_907),
.B(n_893),
.Y(n_1037)
);

AND3x4_ASAP7_75t_L g1038 ( 
.A(n_877),
.B(n_711),
.C(n_871),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_937),
.B(n_940),
.Y(n_1039)
);

NAND2x1p5_ASAP7_75t_L g1040 ( 
.A(n_876),
.B(n_859),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_849),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_SL g1042 ( 
.A1(n_905),
.A2(n_907),
.B(n_893),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_810),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_939),
.B(n_809),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_803),
.A2(n_822),
.B(n_813),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_937),
.B(n_940),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_803),
.A2(n_822),
.B(n_813),
.Y(n_1047)
);

AOI21x1_ASAP7_75t_L g1048 ( 
.A1(n_914),
.A2(n_841),
.B(n_835),
.Y(n_1048)
);

NAND3xp33_ASAP7_75t_L g1049 ( 
.A(n_937),
.B(n_665),
.C(n_678),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_931),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_860),
.B(n_865),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_SL g1052 ( 
.A(n_936),
.B(n_665),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_803),
.A2(n_822),
.B(n_813),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_937),
.A2(n_940),
.B1(n_665),
.B2(n_935),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_937),
.B(n_940),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_937),
.A2(n_665),
.B(n_940),
.C(n_817),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_803),
.A2(n_822),
.B(n_813),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_SL g1058 ( 
.A1(n_905),
.A2(n_907),
.B(n_893),
.Y(n_1058)
);

OR2x6_ASAP7_75t_L g1059 ( 
.A(n_925),
.B(n_776),
.Y(n_1059)
);

AND2x6_ASAP7_75t_L g1060 ( 
.A(n_876),
.B(n_834),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_937),
.B(n_940),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_839),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_937),
.B(n_665),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_939),
.B(n_809),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_937),
.B(n_940),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_937),
.B(n_940),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_856),
.B(n_753),
.Y(n_1067)
);

AOI21x1_ASAP7_75t_L g1068 ( 
.A1(n_914),
.A2(n_841),
.B(n_835),
.Y(n_1068)
);

O2A1O1Ixp5_ASAP7_75t_L g1069 ( 
.A1(n_825),
.A2(n_665),
.B(n_940),
.C(n_937),
.Y(n_1069)
);

AO31x2_ASAP7_75t_L g1070 ( 
.A1(n_913),
.A2(n_847),
.A3(n_802),
.B(n_903),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_970),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_1063),
.B(n_954),
.Y(n_1072)
);

NOR2x1_ASAP7_75t_SL g1073 ( 
.A(n_984),
.B(n_1059),
.Y(n_1073)
);

OR2x2_ASAP7_75t_SL g1074 ( 
.A(n_1049),
.B(n_1067),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1026),
.Y(n_1075)
);

BUFx12f_ASAP7_75t_L g1076 ( 
.A(n_996),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_942),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_1041),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1039),
.B(n_1046),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_1062),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_1059),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_942),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_1059),
.B(n_1004),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_969),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_1004),
.B(n_977),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_947),
.B(n_1032),
.Y(n_1086)
);

INVx5_ASAP7_75t_L g1087 ( 
.A(n_952),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_1006),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_977),
.B(n_1051),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1044),
.B(n_1064),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_998),
.Y(n_1091)
);

NAND2x1_ASAP7_75t_L g1092 ( 
.A(n_953),
.B(n_1006),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1000),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_954),
.B(n_1027),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_971),
.B(n_1039),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_946),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1023),
.B(n_1066),
.Y(n_1097)
);

OA21x2_ASAP7_75t_L g1098 ( 
.A1(n_966),
.A2(n_957),
.B(n_976),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_1052),
.A2(n_1017),
.B1(n_948),
.B2(n_958),
.Y(n_1099)
);

NOR2x1_ASAP7_75t_L g1100 ( 
.A(n_1043),
.B(n_1019),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_987),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_1051),
.B(n_1019),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1022),
.Y(n_1103)
);

INVxp67_ASAP7_75t_L g1104 ( 
.A(n_964),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1035),
.A2(n_1036),
.B1(n_1055),
.B2(n_1061),
.Y(n_1105)
);

OR2x2_ASAP7_75t_SL g1106 ( 
.A(n_1046),
.B(n_1055),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1061),
.B(n_1065),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_1013),
.B(n_941),
.Y(n_1108)
);

INVxp67_ASAP7_75t_L g1109 ( 
.A(n_955),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_1056),
.A2(n_1054),
.B(n_1034),
.C(n_1065),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1050),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1052),
.A2(n_945),
.B1(n_1034),
.B2(n_1029),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_945),
.A2(n_1058),
.B1(n_1042),
.B2(n_1037),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_951),
.A2(n_966),
.B(n_975),
.Y(n_1114)
);

CKINVDCx9p33_ASAP7_75t_R g1115 ( 
.A(n_974),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_952),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1054),
.B(n_944),
.Y(n_1117)
);

INVxp67_ASAP7_75t_SL g1118 ( 
.A(n_950),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_952),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_961),
.B(n_971),
.Y(n_1120)
);

INVx1_ASAP7_75t_SL g1121 ( 
.A(n_962),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_944),
.B(n_962),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_988),
.B(n_986),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_943),
.B(n_972),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_981),
.A2(n_992),
.B1(n_1014),
.B2(n_1018),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_981),
.A2(n_1018),
.B1(n_1008),
.B2(n_973),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_941),
.B(n_978),
.Y(n_1127)
);

BUFx4_ASAP7_75t_SL g1128 ( 
.A(n_941),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_1028),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_978),
.B(n_1033),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_960),
.B(n_949),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_978),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_1016),
.B(n_994),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_1033),
.B(n_994),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_1005),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_1007),
.Y(n_1136)
);

CKINVDCx6p67_ASAP7_75t_R g1137 ( 
.A(n_979),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_997),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1016),
.B(n_953),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1069),
.B(n_956),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_1025),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_1002),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_983),
.B(n_1060),
.Y(n_1143)
);

CKINVDCx8_ASAP7_75t_R g1144 ( 
.A(n_1060),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_989),
.B(n_982),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_980),
.B(n_982),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_997),
.B(n_1040),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1060),
.B(n_1030),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_SL g1149 ( 
.A1(n_1012),
.A2(n_1011),
.B(n_993),
.C(n_999),
.Y(n_1149)
);

O2A1O1Ixp5_ASAP7_75t_L g1150 ( 
.A1(n_968),
.A2(n_1048),
.B(n_1068),
.C(n_1010),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_1021),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1060),
.A2(n_1038),
.B1(n_980),
.B2(n_1015),
.Y(n_1152)
);

INVx5_ASAP7_75t_L g1153 ( 
.A(n_1025),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_1009),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1040),
.B(n_1070),
.Y(n_1155)
);

AND2x6_ASAP7_75t_L g1156 ( 
.A(n_1009),
.B(n_1003),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_985),
.B(n_1003),
.Y(n_1157)
);

OR2x2_ASAP7_75t_SL g1158 ( 
.A(n_1011),
.B(n_1020),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1070),
.B(n_995),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1001),
.B(n_990),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_995),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1070),
.Y(n_1162)
);

INVxp67_ASAP7_75t_SL g1163 ( 
.A(n_991),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_967),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_967),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_967),
.B(n_1057),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1031),
.B(n_1045),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1047),
.B(n_1053),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1017),
.A2(n_665),
.B1(n_940),
.B2(n_937),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_963),
.Y(n_1170)
);

NAND2x1p5_ASAP7_75t_L g1171 ( 
.A(n_1028),
.B(n_1006),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_1059),
.B(n_1004),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1067),
.B(n_856),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1059),
.B(n_1004),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_947),
.B(n_939),
.Y(n_1175)
);

OAI211xp5_ASAP7_75t_L g1176 ( 
.A1(n_1017),
.A2(n_665),
.B(n_820),
.C(n_739),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1059),
.B(n_1004),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1052),
.A2(n_665),
.B1(n_1017),
.B2(n_940),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_942),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1052),
.A2(n_665),
.B1(n_1017),
.B2(n_940),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_1006),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_952),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1063),
.B(n_954),
.Y(n_1183)
);

NOR2x1_ASAP7_75t_SL g1184 ( 
.A(n_984),
.B(n_1059),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_1041),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1035),
.A2(n_665),
.B(n_940),
.C(n_937),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_1062),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_963),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1062),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1067),
.B(n_856),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_965),
.A2(n_959),
.B(n_1024),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1062),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1041),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_963),
.Y(n_1194)
);

INVxp67_ASAP7_75t_L g1195 ( 
.A(n_1041),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1035),
.A2(n_1036),
.B(n_940),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_947),
.B(n_939),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_963),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_965),
.A2(n_959),
.B(n_1024),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_942),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1063),
.B(n_954),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_952),
.Y(n_1202)
);

OR2x6_ASAP7_75t_L g1203 ( 
.A(n_1059),
.B(n_941),
.Y(n_1203)
);

INVxp67_ASAP7_75t_L g1204 ( 
.A(n_1041),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_947),
.B(n_939),
.Y(n_1205)
);

BUFx12f_ASAP7_75t_L g1206 ( 
.A(n_996),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1006),
.Y(n_1207)
);

O2A1O1Ixp5_ASAP7_75t_L g1208 ( 
.A1(n_1034),
.A2(n_665),
.B(n_825),
.C(n_940),
.Y(n_1208)
);

INVx3_ASAP7_75t_SL g1209 ( 
.A(n_986),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_965),
.A2(n_959),
.B(n_1024),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1063),
.A2(n_937),
.B1(n_940),
.B2(n_1027),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_963),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1126),
.A2(n_1180),
.B1(n_1178),
.B2(n_1169),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1155),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_1077),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1144),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1212),
.Y(n_1217)
);

INVxp67_ASAP7_75t_SL g1218 ( 
.A(n_1078),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_1087),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1080),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1071),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1178),
.A2(n_1180),
.B1(n_1072),
.B2(n_1176),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_1142),
.Y(n_1223)
);

INVx4_ASAP7_75t_SL g1224 ( 
.A(n_1156),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1126),
.A2(n_1099),
.B1(n_1211),
.B2(n_1125),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1099),
.B(n_1079),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1107),
.B(n_1183),
.Y(n_1227)
);

OAI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1201),
.A2(n_1097),
.B1(n_1211),
.B2(n_1094),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1079),
.B(n_1154),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1109),
.B(n_1086),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1075),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1125),
.A2(n_1140),
.B1(n_1124),
.B2(n_1112),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1170),
.Y(n_1233)
);

BUFx2_ASAP7_75t_R g1234 ( 
.A(n_1209),
.Y(n_1234)
);

CKINVDCx11_ASAP7_75t_R g1235 ( 
.A(n_1076),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1188),
.Y(n_1236)
);

INVx3_ASAP7_75t_SL g1237 ( 
.A(n_1137),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_1143),
.B(n_1117),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1194),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1077),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_1115),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1196),
.A2(n_1131),
.B1(n_1175),
.B2(n_1197),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1091),
.Y(n_1243)
);

BUFx2_ASAP7_75t_R g1244 ( 
.A(n_1151),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1196),
.A2(n_1205),
.B1(n_1090),
.B2(n_1145),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1148),
.A2(n_1120),
.B1(n_1146),
.B2(n_1114),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1103),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1111),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1123),
.A2(n_1100),
.B1(n_1122),
.B2(n_1104),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1095),
.A2(n_1173),
.B1(n_1190),
.B2(n_1152),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1189),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1093),
.Y(n_1252)
);

AO21x2_ASAP7_75t_L g1253 ( 
.A1(n_1191),
.A2(n_1210),
.B(n_1199),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1135),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1135),
.Y(n_1255)
);

OR2x6_ASAP7_75t_L g1256 ( 
.A(n_1203),
.B(n_1161),
.Y(n_1256)
);

INVx4_ASAP7_75t_L g1257 ( 
.A(n_1087),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1192),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1096),
.B(n_1195),
.Y(n_1259)
);

CKINVDCx9p33_ASAP7_75t_R g1260 ( 
.A(n_1185),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1150),
.Y(n_1261)
);

NAND2x1_ASAP7_75t_L g1262 ( 
.A(n_1129),
.B(n_1167),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1105),
.A2(n_1113),
.B1(n_1152),
.B2(n_1156),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1084),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1136),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1159),
.B(n_1105),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1156),
.A2(n_1193),
.B1(n_1101),
.B2(n_1139),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1082),
.Y(n_1268)
);

CKINVDCx11_ASAP7_75t_R g1269 ( 
.A(n_1206),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1162),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1129),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1157),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1163),
.A2(n_1168),
.B(n_1166),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1106),
.B(n_1098),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1082),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_1074),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1179),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1156),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1179),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1200),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1200),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1204),
.A2(n_1085),
.B1(n_1121),
.B2(n_1083),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1171),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1208),
.B(n_1186),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1141),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1088),
.B(n_1207),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1085),
.A2(n_1121),
.B1(n_1177),
.B2(n_1172),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1160),
.A2(n_1164),
.B(n_1165),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1118),
.Y(n_1289)
);

BUFx2_ASAP7_75t_SL g1290 ( 
.A(n_1087),
.Y(n_1290)
);

CKINVDCx11_ASAP7_75t_R g1291 ( 
.A(n_1089),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1172),
.A2(n_1174),
.B1(n_1177),
.B2(n_1133),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1134),
.Y(n_1293)
);

BUFx12f_ASAP7_75t_L g1294 ( 
.A(n_1187),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1181),
.B(n_1110),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1203),
.A2(n_1081),
.B1(n_1158),
.B2(n_1108),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1102),
.B(n_1127),
.Y(n_1297)
);

BUFx12f_ASAP7_75t_L g1298 ( 
.A(n_1102),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1147),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1171),
.A2(n_1092),
.B(n_1149),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1138),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1138),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1153),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1127),
.B(n_1132),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1116),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1119),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1153),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1081),
.B(n_1073),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_SL g1309 ( 
.A1(n_1184),
.A2(n_1203),
.B1(n_1153),
.B2(n_1128),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1182),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1130),
.A2(n_665),
.B1(n_1017),
.B2(n_1052),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1202),
.B(n_665),
.Y(n_1312)
);

BUFx2_ASAP7_75t_SL g1313 ( 
.A(n_1202),
.Y(n_1313)
);

BUFx12f_ASAP7_75t_L g1314 ( 
.A(n_1142),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1169),
.A2(n_665),
.B1(n_940),
.B2(n_937),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1099),
.B(n_1178),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1142),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1176),
.A2(n_665),
.B1(n_1063),
.B2(n_816),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1072),
.B(n_1063),
.Y(n_1319)
);

INVx4_ASAP7_75t_L g1320 ( 
.A(n_1087),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1139),
.B(n_1088),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1099),
.B(n_1178),
.Y(n_1322)
);

CKINVDCx11_ASAP7_75t_R g1323 ( 
.A(n_1076),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_1099),
.B(n_1143),
.Y(n_1324)
);

NAND2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1145),
.B(n_1161),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1144),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_SL g1327 ( 
.A1(n_1176),
.A2(n_665),
.B(n_536),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1176),
.A2(n_665),
.B1(n_1052),
.B2(n_1017),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1126),
.A2(n_665),
.B1(n_1017),
.B2(n_1052),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1173),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1155),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1176),
.A2(n_665),
.B1(n_1052),
.B2(n_1017),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1072),
.B(n_1063),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1198),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1198),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1214),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1220),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1329),
.A2(n_1225),
.B1(n_1332),
.B2(n_1328),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1318),
.A2(n_1315),
.B(n_1327),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1270),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1266),
.B(n_1316),
.Y(n_1341)
);

OR2x6_ASAP7_75t_L g1342 ( 
.A(n_1256),
.B(n_1325),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1262),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1322),
.B(n_1226),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1288),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1322),
.B(n_1226),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1274),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_1262),
.Y(n_1348)
);

AO21x2_ASAP7_75t_L g1349 ( 
.A1(n_1253),
.A2(n_1261),
.B(n_1284),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1220),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1274),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1272),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1254),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1224),
.B(n_1256),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1251),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1324),
.B(n_1238),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1276),
.A2(n_1222),
.B1(n_1241),
.B2(n_1319),
.Y(n_1357)
);

NAND2xp33_ASAP7_75t_R g1358 ( 
.A(n_1223),
.B(n_1317),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1215),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1251),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1324),
.B(n_1238),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1223),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1214),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1240),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1268),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1331),
.B(n_1232),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1258),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1273),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1284),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1277),
.Y(n_1370)
);

BUFx5_ASAP7_75t_L g1371 ( 
.A(n_1295),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1300),
.A2(n_1271),
.B(n_1325),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1276),
.A2(n_1241),
.B1(n_1333),
.B2(n_1296),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1221),
.Y(n_1374)
);

INVx4_ASAP7_75t_L g1375 ( 
.A(n_1257),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1231),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1233),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1256),
.B(n_1250),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1258),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1229),
.B(n_1295),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1236),
.Y(n_1381)
);

AOI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1213),
.A2(n_1228),
.B1(n_1249),
.B2(n_1242),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1263),
.B(n_1278),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1278),
.B(n_1246),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1239),
.Y(n_1385)
);

AO21x2_ASAP7_75t_L g1386 ( 
.A1(n_1253),
.A2(n_1243),
.B(n_1289),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1264),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1253),
.A2(n_1308),
.B(n_1252),
.Y(n_1388)
);

INVxp67_ASAP7_75t_L g1389 ( 
.A(n_1281),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1217),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1264),
.Y(n_1391)
);

INVx11_ASAP7_75t_L g1392 ( 
.A(n_1314),
.Y(n_1392)
);

NAND2x1_ASAP7_75t_L g1393 ( 
.A(n_1256),
.B(n_1283),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1325),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1224),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1298),
.Y(n_1396)
);

AO21x2_ASAP7_75t_L g1397 ( 
.A1(n_1247),
.A2(n_1248),
.B(n_1334),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1224),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1330),
.B(n_1275),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1335),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1311),
.A2(n_1245),
.B(n_1267),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1255),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_1260),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1227),
.B(n_1279),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1299),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1280),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1218),
.B(n_1312),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1283),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1283),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1286),
.B(n_1321),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1286),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_1235),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1285),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1265),
.Y(n_1414)
);

INVxp67_ASAP7_75t_L g1415 ( 
.A(n_1230),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1309),
.A2(n_1259),
.B(n_1282),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1303),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1293),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1307),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1307),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1301),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1369),
.B(n_1302),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1347),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1347),
.B(n_1321),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1351),
.B(n_1304),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1340),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1349),
.B(n_1305),
.Y(n_1427)
);

INVx5_ASAP7_75t_SL g1428 ( 
.A(n_1342),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1393),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1386),
.Y(n_1430)
);

NOR2x1_ASAP7_75t_SL g1431 ( 
.A(n_1342),
.B(n_1290),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1349),
.B(n_1310),
.Y(n_1432)
);

AND2x4_ASAP7_75t_SL g1433 ( 
.A(n_1354),
.B(n_1216),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1368),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1386),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1386),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1339),
.B(n_1326),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1388),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1368),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1382),
.B(n_1216),
.Y(n_1440)
);

OAI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1366),
.A2(n_1216),
.B1(n_1326),
.B2(n_1297),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1356),
.B(n_1216),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1371),
.B(n_1292),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1388),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1388),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1356),
.B(n_1216),
.Y(n_1446)
);

OR2x6_ASAP7_75t_L g1447 ( 
.A(n_1342),
.B(n_1290),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1393),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1371),
.B(n_1345),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1397),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1338),
.A2(n_1291),
.B1(n_1326),
.B2(n_1287),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1397),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1397),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1361),
.B(n_1306),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1361),
.B(n_1219),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1359),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1336),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1336),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1363),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1357),
.A2(n_1244),
.B1(n_1234),
.B2(n_1237),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1341),
.B(n_1313),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1352),
.B(n_1219),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1363),
.Y(n_1463)
);

NAND2x1p5_ASAP7_75t_L g1464 ( 
.A(n_1372),
.B(n_1257),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1343),
.B(n_1257),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1416),
.A2(n_1320),
.B(n_1317),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1460),
.A2(n_1373),
.B1(n_1403),
.B2(n_1366),
.Y(n_1467)
);

NAND3xp33_ASAP7_75t_L g1468 ( 
.A(n_1466),
.B(n_1437),
.C(n_1440),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_SL g1469 ( 
.A(n_1466),
.B(n_1378),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1437),
.B(n_1407),
.Y(n_1470)
);

NAND3xp33_ASAP7_75t_L g1471 ( 
.A(n_1440),
.B(n_1394),
.C(n_1378),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1454),
.B(n_1442),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1460),
.A2(n_1415),
.B1(n_1401),
.B2(n_1346),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_SL g1474 ( 
.A(n_1454),
.B(n_1362),
.Y(n_1474)
);

NOR3xp33_ASAP7_75t_L g1475 ( 
.A(n_1441),
.B(n_1404),
.C(n_1389),
.Y(n_1475)
);

NAND3xp33_ASAP7_75t_L g1476 ( 
.A(n_1451),
.B(n_1456),
.C(n_1444),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1451),
.A2(n_1401),
.B1(n_1384),
.B2(n_1383),
.Y(n_1477)
);

OAI21xp33_ASAP7_75t_L g1478 ( 
.A1(n_1442),
.A2(n_1384),
.B(n_1446),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1454),
.B(n_1364),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1441),
.A2(n_1383),
.B(n_1346),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1446),
.B(n_1365),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1456),
.B(n_1370),
.Y(n_1482)
);

NOR3xp33_ASAP7_75t_L g1483 ( 
.A(n_1462),
.B(n_1375),
.C(n_1291),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1425),
.B(n_1455),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1455),
.B(n_1380),
.Y(n_1485)
);

OAI21xp5_ASAP7_75t_SL g1486 ( 
.A1(n_1433),
.A2(n_1344),
.B(n_1398),
.Y(n_1486)
);

OAI221xp5_ASAP7_75t_L g1487 ( 
.A1(n_1447),
.A2(n_1237),
.B1(n_1399),
.B2(n_1396),
.C(n_1367),
.Y(n_1487)
);

NAND3xp33_ASAP7_75t_L g1488 ( 
.A(n_1438),
.B(n_1418),
.C(n_1408),
.Y(n_1488)
);

NAND4xp25_ASAP7_75t_L g1489 ( 
.A(n_1462),
.B(n_1399),
.C(n_1414),
.D(n_1406),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1457),
.B(n_1344),
.Y(n_1490)
);

OAI221xp5_ASAP7_75t_SL g1491 ( 
.A1(n_1447),
.A2(n_1414),
.B1(n_1406),
.B2(n_1396),
.C(n_1402),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1457),
.B(n_1353),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1449),
.B(n_1374),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1458),
.B(n_1353),
.Y(n_1494)
);

OAI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1447),
.A2(n_1401),
.B1(n_1350),
.B2(n_1367),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1464),
.A2(n_1372),
.B(n_1417),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1443),
.A2(n_1401),
.B1(n_1410),
.B2(n_1413),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1458),
.B(n_1413),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1465),
.B(n_1410),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1443),
.A2(n_1410),
.B1(n_1402),
.B2(n_1298),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_SL g1501 ( 
.A(n_1465),
.B(n_1410),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_L g1502 ( 
.A(n_1438),
.B(n_1408),
.C(n_1409),
.Y(n_1502)
);

NAND3xp33_ASAP7_75t_L g1503 ( 
.A(n_1444),
.B(n_1409),
.C(n_1419),
.Y(n_1503)
);

NAND2xp33_ASAP7_75t_SL g1504 ( 
.A(n_1461),
.B(n_1412),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1459),
.B(n_1374),
.Y(n_1505)
);

NAND3xp33_ASAP7_75t_L g1506 ( 
.A(n_1445),
.B(n_1435),
.C(n_1430),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1459),
.B(n_1463),
.Y(n_1507)
);

AOI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1427),
.A2(n_1411),
.B1(n_1405),
.B2(n_1400),
.C(n_1376),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1443),
.A2(n_1411),
.B1(n_1405),
.B2(n_1390),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1447),
.A2(n_1360),
.B1(n_1350),
.B2(n_1337),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1463),
.B(n_1422),
.Y(n_1511)
);

NAND3xp33_ASAP7_75t_L g1512 ( 
.A(n_1445),
.B(n_1435),
.C(n_1430),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1464),
.A2(n_1419),
.B(n_1417),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1429),
.B(n_1348),
.Y(n_1514)
);

NOR3xp33_ASAP7_75t_L g1515 ( 
.A(n_1450),
.B(n_1375),
.C(n_1395),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1447),
.A2(n_1355),
.B1(n_1360),
.B2(n_1379),
.Y(n_1516)
);

NAND3xp33_ASAP7_75t_L g1517 ( 
.A(n_1436),
.B(n_1420),
.C(n_1377),
.Y(n_1517)
);

AOI221x1_ASAP7_75t_SL g1518 ( 
.A1(n_1426),
.A2(n_1377),
.B1(n_1376),
.B2(n_1385),
.C(n_1381),
.Y(n_1518)
);

OAI221xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1447),
.A2(n_1337),
.B1(n_1355),
.B2(n_1379),
.C(n_1400),
.Y(n_1519)
);

AND2x4_ASAP7_75t_SL g1520 ( 
.A(n_1514),
.B(n_1447),
.Y(n_1520)
);

NAND2x1_ASAP7_75t_L g1521 ( 
.A(n_1514),
.B(n_1434),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1493),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1507),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1514),
.B(n_1429),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1505),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1484),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1517),
.Y(n_1527)
);

INVxp67_ASAP7_75t_SL g1528 ( 
.A(n_1503),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1498),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1511),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1518),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1492),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1499),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1499),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1468),
.B(n_1429),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1494),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1501),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1479),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1490),
.B(n_1434),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1502),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1472),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1501),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1485),
.B(n_1423),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1506),
.B(n_1434),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1482),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1497),
.B(n_1439),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1497),
.B(n_1439),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1512),
.Y(n_1548)
);

INVxp67_ASAP7_75t_L g1549 ( 
.A(n_1488),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_L g1550 ( 
.A(n_1469),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1481),
.B(n_1423),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1513),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1489),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1478),
.B(n_1423),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1508),
.B(n_1427),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1474),
.B(n_1429),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1496),
.B(n_1432),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1510),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1516),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1471),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1515),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1509),
.B(n_1432),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1509),
.B(n_1432),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1553),
.B(n_1470),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1560),
.B(n_1450),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1520),
.B(n_1448),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1522),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1524),
.B(n_1428),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1522),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1553),
.B(n_1470),
.Y(n_1570)
);

NAND2xp33_ASAP7_75t_SL g1571 ( 
.A(n_1556),
.B(n_1467),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1522),
.Y(n_1572)
);

INVxp33_ASAP7_75t_SL g1573 ( 
.A(n_1556),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1524),
.B(n_1428),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1560),
.B(n_1452),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_SL g1576 ( 
.A(n_1550),
.B(n_1519),
.Y(n_1576)
);

INVxp67_ASAP7_75t_SL g1577 ( 
.A(n_1540),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1539),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1520),
.B(n_1448),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1539),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1538),
.B(n_1475),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1539),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1529),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1538),
.B(n_1424),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1551),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1524),
.B(n_1428),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1524),
.B(n_1428),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1544),
.Y(n_1588)
);

OAI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1549),
.A2(n_1476),
.B(n_1477),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1544),
.Y(n_1590)
);

INVxp67_ASAP7_75t_SL g1591 ( 
.A(n_1540),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1529),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1544),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1551),
.Y(n_1594)
);

OAI21xp33_ASAP7_75t_L g1595 ( 
.A1(n_1555),
.A2(n_1552),
.B(n_1535),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1524),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1533),
.B(n_1428),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1533),
.B(n_1428),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1560),
.B(n_1452),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1533),
.B(n_1431),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1545),
.B(n_1424),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_1552),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1534),
.B(n_1431),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1554),
.B(n_1453),
.Y(n_1604)
);

NOR2x1_ASAP7_75t_L g1605 ( 
.A(n_1535),
.B(n_1487),
.Y(n_1605)
);

NOR2x1_ASAP7_75t_L g1606 ( 
.A(n_1548),
.B(n_1448),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1581),
.B(n_1531),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1594),
.B(n_1548),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1583),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1564),
.B(n_1392),
.Y(n_1610)
);

INVxp67_ASAP7_75t_SL g1611 ( 
.A(n_1606),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1596),
.B(n_1600),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1570),
.B(n_1531),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1567),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1589),
.B(n_1595),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1596),
.B(n_1557),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1583),
.Y(n_1617)
);

NOR2xp67_ASAP7_75t_L g1618 ( 
.A(n_1602),
.B(n_1549),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1592),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1577),
.B(n_1561),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1594),
.B(n_1528),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1567),
.Y(n_1622)
);

NAND2x1_ASAP7_75t_L g1623 ( 
.A(n_1566),
.B(n_1550),
.Y(n_1623)
);

AND2x2_ASAP7_75t_SL g1624 ( 
.A(n_1576),
.B(n_1550),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1600),
.B(n_1557),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1592),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1603),
.B(n_1557),
.Y(n_1627)
);

AOI32xp33_ASAP7_75t_L g1628 ( 
.A1(n_1571),
.A2(n_1528),
.A3(n_1555),
.B1(n_1563),
.B2(n_1562),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1578),
.B(n_1527),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1578),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1603),
.B(n_1534),
.Y(n_1631)
);

NOR2x1p5_ASAP7_75t_L g1632 ( 
.A(n_1591),
.B(n_1550),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1566),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1605),
.B(n_1561),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1573),
.A2(n_1473),
.B1(n_1550),
.B2(n_1469),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1573),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1585),
.B(n_1545),
.Y(n_1637)
);

INVxp67_ASAP7_75t_SL g1638 ( 
.A(n_1565),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1568),
.B(n_1534),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1580),
.Y(n_1640)
);

INVx2_ASAP7_75t_SL g1641 ( 
.A(n_1566),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1568),
.B(n_1537),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1574),
.B(n_1537),
.Y(n_1643)
);

INVx2_ASAP7_75t_SL g1644 ( 
.A(n_1579),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1580),
.Y(n_1645)
);

XNOR2xp5_ASAP7_75t_L g1646 ( 
.A(n_1574),
.B(n_1362),
.Y(n_1646)
);

OAI21xp33_ASAP7_75t_L g1647 ( 
.A1(n_1582),
.A2(n_1480),
.B(n_1550),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1569),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1588),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1582),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1601),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1584),
.B(n_1523),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1636),
.B(n_1607),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1609),
.Y(n_1654)
);

NAND3xp33_ASAP7_75t_L g1655 ( 
.A(n_1628),
.B(n_1550),
.C(n_1527),
.Y(n_1655)
);

AND3x2_ASAP7_75t_L g1656 ( 
.A(n_1611),
.B(n_1558),
.C(n_1483),
.Y(n_1656)
);

INVx5_ASAP7_75t_L g1657 ( 
.A(n_1633),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1609),
.Y(n_1658)
);

AOI21xp33_ASAP7_75t_SL g1659 ( 
.A1(n_1624),
.A2(n_1358),
.B(n_1558),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1618),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1617),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1633),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1615),
.B(n_1235),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1624),
.B(n_1588),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1632),
.B(n_1590),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1634),
.A2(n_1559),
.B1(n_1537),
.B2(n_1542),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1617),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1621),
.B(n_1590),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1623),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1646),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1641),
.B(n_1579),
.Y(n_1671)
);

CKINVDCx16_ASAP7_75t_R g1672 ( 
.A(n_1646),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1612),
.B(n_1593),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1621),
.B(n_1593),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1619),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1619),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1626),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1623),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1626),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1612),
.B(n_1586),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1608),
.B(n_1565),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1608),
.B(n_1575),
.Y(n_1682)
);

NOR2xp67_ASAP7_75t_L g1683 ( 
.A(n_1641),
.B(n_1579),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1639),
.B(n_1586),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1629),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1630),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1639),
.B(n_1587),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1630),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1635),
.A2(n_1559),
.B1(n_1542),
.B2(n_1491),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1660),
.B(n_1644),
.Y(n_1690)
);

OA21x2_ASAP7_75t_L g1691 ( 
.A1(n_1655),
.A2(n_1620),
.B(n_1640),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1670),
.B(n_1613),
.Y(n_1692)
);

AOI22x1_ASAP7_75t_L g1693 ( 
.A1(n_1672),
.A2(n_1629),
.B1(n_1649),
.B2(n_1644),
.Y(n_1693)
);

AOI21xp33_ASAP7_75t_SL g1694 ( 
.A1(n_1663),
.A2(n_1647),
.B(n_1610),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1657),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1657),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1659),
.A2(n_1645),
.B1(n_1650),
.B2(n_1640),
.C(n_1638),
.Y(n_1697)
);

OAI322xp33_ASAP7_75t_SL g1698 ( 
.A1(n_1653),
.A2(n_1651),
.A3(n_1637),
.B1(n_1652),
.B2(n_1614),
.C1(n_1622),
.C2(n_1648),
.Y(n_1698)
);

A2O1A1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1663),
.A2(n_1504),
.B(n_1616),
.C(n_1547),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1656),
.A2(n_1504),
.B1(n_1643),
.B2(n_1642),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1657),
.Y(n_1701)
);

AOI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1689),
.A2(n_1666),
.B1(n_1685),
.B2(n_1662),
.C(n_1664),
.Y(n_1702)
);

OAI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1683),
.A2(n_1616),
.B1(n_1643),
.B2(n_1642),
.C(n_1521),
.Y(n_1703)
);

AOI21xp33_ASAP7_75t_L g1704 ( 
.A1(n_1678),
.A2(n_1599),
.B(n_1575),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1680),
.B(n_1631),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1680),
.B(n_1631),
.Y(n_1706)
);

INVxp67_ASAP7_75t_L g1707 ( 
.A(n_1664),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1654),
.Y(n_1708)
);

OAI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1678),
.A2(n_1599),
.B(n_1598),
.Y(n_1709)
);

AOI21xp33_ASAP7_75t_SL g1710 ( 
.A1(n_1669),
.A2(n_1323),
.B(n_1269),
.Y(n_1710)
);

OAI21xp33_ASAP7_75t_L g1711 ( 
.A1(n_1665),
.A2(n_1627),
.B(n_1625),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1673),
.B(n_1625),
.Y(n_1712)
);

AOI21xp33_ASAP7_75t_L g1713 ( 
.A1(n_1668),
.A2(n_1622),
.B(n_1614),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_1657),
.Y(n_1714)
);

OAI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1665),
.A2(n_1598),
.B(n_1597),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1657),
.B(n_1627),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1707),
.B(n_1673),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1708),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1690),
.B(n_1684),
.Y(n_1719)
);

NOR2x1_ASAP7_75t_L g1720 ( 
.A(n_1695),
.B(n_1669),
.Y(n_1720)
);

INVx2_ASAP7_75t_SL g1721 ( 
.A(n_1690),
.Y(n_1721)
);

NAND2xp33_ASAP7_75t_SL g1722 ( 
.A(n_1716),
.B(n_1714),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1710),
.B(n_1269),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1714),
.B(n_1695),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1692),
.B(n_1684),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1702),
.A2(n_1687),
.B1(n_1671),
.B2(n_1669),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1712),
.B(n_1668),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1694),
.B(n_1323),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1700),
.B(n_1314),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1705),
.B(n_1687),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1696),
.Y(n_1731)
);

NOR3xp33_ASAP7_75t_L g1732 ( 
.A(n_1716),
.B(n_1661),
.C(n_1658),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1696),
.Y(n_1733)
);

INVxp33_ASAP7_75t_L g1734 ( 
.A(n_1693),
.Y(n_1734)
);

INVxp33_ASAP7_75t_L g1735 ( 
.A(n_1705),
.Y(n_1735)
);

NAND2x1_ASAP7_75t_L g1736 ( 
.A(n_1701),
.B(n_1671),
.Y(n_1736)
);

OAI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1691),
.A2(n_1674),
.B1(n_1521),
.B2(n_1559),
.Y(n_1737)
);

OAI221xp5_ASAP7_75t_L g1738 ( 
.A1(n_1726),
.A2(n_1699),
.B1(n_1697),
.B2(n_1691),
.C(n_1715),
.Y(n_1738)
);

NAND3xp33_ASAP7_75t_SL g1739 ( 
.A(n_1734),
.B(n_1699),
.C(n_1701),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1731),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1723),
.B(n_1711),
.Y(n_1741)
);

OAI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1722),
.A2(n_1691),
.B1(n_1703),
.B2(n_1709),
.C(n_1698),
.Y(n_1742)
);

NAND4xp25_ASAP7_75t_SL g1743 ( 
.A(n_1732),
.B(n_1706),
.C(n_1704),
.D(n_1713),
.Y(n_1743)
);

AOI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1728),
.A2(n_1706),
.B(n_1688),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1735),
.A2(n_1671),
.B1(n_1674),
.B2(n_1686),
.Y(n_1745)
);

OAI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1737),
.A2(n_1675),
.B(n_1667),
.Y(n_1746)
);

OAI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1721),
.A2(n_1542),
.B1(n_1681),
.B2(n_1682),
.Y(n_1747)
);

OAI211xp5_ASAP7_75t_SL g1748 ( 
.A1(n_1725),
.A2(n_1679),
.B(n_1677),
.C(n_1676),
.Y(n_1748)
);

NAND4xp25_ASAP7_75t_SL g1749 ( 
.A(n_1719),
.B(n_1682),
.C(n_1681),
.D(n_1597),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1729),
.B(n_1392),
.Y(n_1750)
);

NAND5xp2_ASAP7_75t_L g1751 ( 
.A(n_1738),
.B(n_1717),
.C(n_1733),
.D(n_1730),
.E(n_1718),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_SL g1752 ( 
.A(n_1747),
.B(n_1745),
.Y(n_1752)
);

NAND3xp33_ASAP7_75t_SL g1753 ( 
.A(n_1742),
.B(n_1736),
.C(n_1717),
.Y(n_1753)
);

NAND3xp33_ASAP7_75t_SL g1754 ( 
.A(n_1744),
.B(n_1727),
.C(n_1720),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1741),
.B(n_1724),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1740),
.Y(n_1756)
);

NAND4xp25_ASAP7_75t_L g1757 ( 
.A(n_1739),
.B(n_1724),
.C(n_1391),
.D(n_1387),
.Y(n_1757)
);

NOR3x1_ASAP7_75t_L g1758 ( 
.A(n_1746),
.B(n_1604),
.C(n_1554),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1750),
.B(n_1587),
.Y(n_1759)
);

NAND4xp25_ASAP7_75t_L g1760 ( 
.A(n_1748),
.B(n_1391),
.C(n_1500),
.D(n_1546),
.Y(n_1760)
);

NOR3xp33_ASAP7_75t_L g1761 ( 
.A(n_1743),
.B(n_1495),
.C(n_1648),
.Y(n_1761)
);

NOR3xp33_ASAP7_75t_L g1762 ( 
.A(n_1751),
.B(n_1749),
.C(n_1320),
.Y(n_1762)
);

OAI221xp5_ASAP7_75t_L g1763 ( 
.A1(n_1761),
.A2(n_1554),
.B1(n_1604),
.B2(n_1523),
.C(n_1536),
.Y(n_1763)
);

AOI211x1_ASAP7_75t_SL g1764 ( 
.A1(n_1754),
.A2(n_1543),
.B(n_1530),
.C(n_1421),
.Y(n_1764)
);

XOR2xp5_ASAP7_75t_L g1765 ( 
.A(n_1753),
.B(n_1500),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1755),
.Y(n_1766)
);

OAI211xp5_ASAP7_75t_SL g1767 ( 
.A1(n_1752),
.A2(n_1536),
.B(n_1532),
.C(n_1526),
.Y(n_1767)
);

A2O1A1Ixp33_ASAP7_75t_L g1768 ( 
.A1(n_1760),
.A2(n_1547),
.B(n_1546),
.C(n_1563),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1766),
.Y(n_1769)
);

INVxp67_ASAP7_75t_SL g1770 ( 
.A(n_1762),
.Y(n_1770)
);

NOR2x1_ASAP7_75t_L g1771 ( 
.A(n_1765),
.B(n_1756),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1763),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1764),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1768),
.B(n_1757),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1769),
.B(n_1767),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1771),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1774),
.Y(n_1777)
);

NOR4xp75_ASAP7_75t_SL g1778 ( 
.A(n_1770),
.B(n_1758),
.C(n_1759),
.D(n_1294),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1772),
.B(n_1569),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1776),
.Y(n_1780)
);

INVx3_ASAP7_75t_L g1781 ( 
.A(n_1779),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1775),
.B(n_1773),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1780),
.A2(n_1777),
.B1(n_1779),
.B2(n_1778),
.Y(n_1783)
);

XNOR2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1783),
.B(n_1781),
.Y(n_1784)
);

AOI21xp33_ASAP7_75t_L g1785 ( 
.A1(n_1784),
.A2(n_1782),
.B(n_1781),
.Y(n_1785)
);

AO21x2_ASAP7_75t_L g1786 ( 
.A1(n_1784),
.A2(n_1294),
.B(n_1572),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1785),
.A2(n_1572),
.B(n_1320),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1786),
.Y(n_1788)
);

AOI21xp33_ASAP7_75t_L g1789 ( 
.A1(n_1788),
.A2(n_1532),
.B(n_1525),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1787),
.B(n_1541),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1790),
.A2(n_1541),
.B1(n_1526),
.B2(n_1525),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1791),
.Y(n_1792)
);

OAI221xp5_ASAP7_75t_R g1793 ( 
.A1(n_1792),
.A2(n_1789),
.B1(n_1520),
.B2(n_1551),
.C(n_1530),
.Y(n_1793)
);

AOI211xp5_ASAP7_75t_L g1794 ( 
.A1(n_1793),
.A2(n_1486),
.B(n_1398),
.C(n_1395),
.Y(n_1794)
);


endmodule