module real_jpeg_13890_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_258, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_258;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_105;
wire n_40;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_44),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_2),
.A2(n_44),
.B1(n_61),
.B2(n_62),
.Y(n_121)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_4),
.A2(n_55),
.B1(n_57),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_67),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_4),
.A2(n_41),
.B1(n_42),
.B2(n_67),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_67),
.Y(n_177)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_22)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_7),
.A2(n_27),
.B1(n_41),
.B2(n_42),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_7),
.A2(n_27),
.B1(n_61),
.B2(n_62),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_7),
.A2(n_27),
.B1(n_55),
.B2(n_57),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_10),
.A2(n_33),
.B1(n_55),
.B2(n_57),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_10),
.A2(n_33),
.B1(n_61),
.B2(n_62),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_10),
.A2(n_33),
.B1(n_41),
.B2(n_42),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_10),
.B(n_99),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_10),
.B(n_24),
.C(n_38),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_10),
.B(n_34),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_10),
.B(n_37),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_10),
.A2(n_62),
.B(n_73),
.C(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_10),
.B(n_58),
.Y(n_197)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_125),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_124),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_105),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_16),
.B(n_105),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_81),
.C(n_88),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_17),
.A2(n_18),
.B1(n_81),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_49),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_19),
.B(n_50),
.C(n_69),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_20),
.B(n_35),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_30),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_21),
.B(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_21),
.A2(n_29),
.B(n_91),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_22),
.B(n_29),
.Y(n_93)
);

AO22x1_ASAP7_75t_L g37 ( 
.A1(n_23),
.A2(n_24),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_24),
.B(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_28),
.A2(n_29),
.B(n_32),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_28),
.A2(n_91),
.B(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_28),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_28),
.B(n_32),
.Y(n_159)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_29),
.B(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_30),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_33),
.A2(n_41),
.B(n_74),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_33),
.B(n_59),
.C(n_62),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_40),
.B(n_45),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_36),
.A2(n_85),
.B(n_97),
.Y(n_222)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_37),
.B(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_37),
.B(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_37),
.B(n_141),
.Y(n_151)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_40),
.A2(n_85),
.B(n_86),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_42),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_42),
.B(n_149),
.Y(n_148)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_45),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_45),
.B(n_151),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_46),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_46),
.B(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_68),
.B2(n_69),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_63),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_54),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_54),
.B(n_114),
.Y(n_216)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_55),
.B(n_209),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_66),
.Y(n_102)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_58),
.B(n_104),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_62),
.B1(n_73),
.B2(n_74),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_63),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_64),
.B(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_75),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_70),
.B(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_71),
.B(n_78),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_76),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_80),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_78),
.B(n_194),
.Y(n_193)
);

NAND2x1_ASAP7_75t_SL g230 ( 
.A(n_80),
.B(n_99),
.Y(n_230)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_81),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_87),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_83),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_82),
.A2(n_83),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_84),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_83),
.B(n_180),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_84),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_86),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_88),
.B(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_98),
.C(n_100),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_89),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_90),
.B(n_94),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_93),
.B(n_135),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_93),
.B(n_159),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_95),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_98),
.A2(n_100),
.B1(n_101),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_98),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_99),
.B(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_102),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_116),
.B2(n_117),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_120),
.B(n_123),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_120),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_119),
.B(n_140),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_122),
.B(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_250),
.B(n_255),
.Y(n_125)
);

AOI321xp33_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_224),
.A3(n_243),
.B1(n_248),
.B2(n_249),
.C(n_258),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_200),
.B(n_223),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_184),
.B(n_199),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_171),
.B(n_183),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_152),
.B(n_170),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_146),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_146),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_137),
.B1(n_138),
.B2(n_145),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_133),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_139),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_143),
.C(n_145),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_164),
.B(n_169),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_160),
.B(n_163),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_162),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_167),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_173),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_179),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_178),
.C(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_180),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_198),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_198),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_191),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_189),
.C(n_191),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_196),
.C(n_197),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_202),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_212),
.B2(n_213),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_206),
.C(n_212),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_211),
.Y(n_232)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_219),
.C(n_221),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_238),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_238),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_233),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_234),
.C(n_237),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.C(n_232),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_227),
.B(n_229),
.CI(n_232),
.CON(n_240),
.SN(n_240)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.C(n_242),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_240),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g256 ( 
.A(n_240),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_242),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_247),
.Y(n_248)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);


endmodule