module fake_jpeg_10591_n_170 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_170);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_38),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_20),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_35),
.A2(n_28),
.B1(n_19),
.B2(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_1),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_24),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_18),
.B(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_25),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_40),
.Y(n_60)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_2),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_57),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_20),
.B1(n_16),
.B2(n_17),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_62),
.B1(n_23),
.B2(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_5),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_25),
.Y(n_56)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_25),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_19),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_58),
.B(n_54),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_65),
.A2(n_47),
.B(n_59),
.Y(n_96)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_76),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_74),
.Y(n_90)
);

AND2x6_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_4),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_79),
.C(n_82),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_78),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_72),
.B(n_73),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_18),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_26),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_53),
.B(n_23),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_22),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_4),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_84),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_27),
.B1(n_26),
.B2(n_21),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_81),
.A2(n_60),
.B1(n_42),
.B2(n_5),
.Y(n_105)
);

AND2x6_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_4),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_51),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_85),
.B(n_5),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_44),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_89),
.B(n_96),
.Y(n_117)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_101),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_46),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_9),
.Y(n_121)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_52),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_48),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_103),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_45),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_68),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_76),
.B1(n_75),
.B2(n_86),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_42),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_80),
.Y(n_115)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_114),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_77),
.B1(n_73),
.B2(n_65),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_66),
.C(n_71),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_118),
.C(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_121),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_82),
.B1(n_70),
.B2(n_83),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_80),
.C(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_106),
.B1(n_95),
.B2(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_32),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_112),
.Y(n_136)
);

A2O1A1O1Ixp25_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_93),
.B(n_88),
.C(n_89),
.D(n_96),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_118),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_129),
.C(n_110),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_109),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_130),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_104),
.C(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_133),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_120),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_145),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_142),
.C(n_144),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_107),
.Y(n_139)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_134),
.A2(n_107),
.B1(n_121),
.B2(n_115),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_135),
.B1(n_131),
.B2(n_132),
.Y(n_151)
);

BUFx12_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_125),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_113),
.C(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_91),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_130),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_148),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_141),
.B(n_129),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_151),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_131),
.Y(n_155)
);

AOI31xp67_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_135),
.A3(n_124),
.B(n_144),
.Y(n_154)
);

OAI31xp33_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_121),
.A3(n_153),
.B(n_32),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_155),
.B(n_156),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_141),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_99),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_157),
.B(n_10),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_142),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_60),
.C(n_11),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_159),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_154),
.C(n_153),
.Y(n_165)
);

BUFx24_ASAP7_75t_SL g167 ( 
.A(n_164),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

AOI32xp33_ASAP7_75t_L g169 ( 
.A1(n_167),
.A2(n_168),
.A3(n_161),
.B1(n_166),
.B2(n_162),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_13),
.Y(n_170)
);


endmodule