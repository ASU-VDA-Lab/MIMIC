module fake_netlist_5_589_n_1919 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1919);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1919;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_174;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_177;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx2_ASAP7_75t_L g158 ( 
.A(n_53),
.Y(n_158)
);

BUFx2_ASAP7_75t_SL g159 ( 
.A(n_39),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_17),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_46),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_90),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_24),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_0),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_17),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_0),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_125),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_21),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_35),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_5),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_118),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_41),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_102),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_25),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_59),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_119),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_116),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_50),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_64),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_96),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_24),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_40),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_106),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_5),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_1),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_94),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_123),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_137),
.Y(n_191)
);

BUFx2_ASAP7_75t_SL g192 ( 
.A(n_113),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_86),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_33),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_99),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_107),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_42),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_141),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_89),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_39),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_33),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_124),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_84),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_15),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_41),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_95),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_72),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_55),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_70),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_31),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_87),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_47),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_121),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_93),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_54),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_77),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_9),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_4),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_126),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_34),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_144),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_73),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_16),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_35),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_138),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_12),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_79),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_40),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_26),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_91),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_74),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_156),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_14),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_75),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_7),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_139),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_150),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_25),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_27),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_85),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_20),
.Y(n_244)
);

BUFx2_ASAP7_75t_SL g245 ( 
.A(n_154),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_20),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_134),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_30),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_92),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_1),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_63),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_56),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_2),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_44),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_32),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_36),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_112),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_83),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_8),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_136),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_2),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_37),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_14),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_109),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_133),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_140),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_45),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_120),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_81),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_131),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_31),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_32),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_62),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_65),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_29),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_22),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_115),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_28),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_80),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_66),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_98),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_67),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_28),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_23),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_12),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_157),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_37),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_6),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_10),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_4),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_15),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_88),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_30),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_61),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_51),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_58),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_153),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_130),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_143),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_18),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_21),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_105),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_8),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_18),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_76),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_101),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_114),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_22),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_129),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_11),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_29),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_34),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_60),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_177),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_188),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_188),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_203),
.Y(n_317)
);

INVxp33_ASAP7_75t_SL g318 ( 
.A(n_163),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_189),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_203),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_172),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_253),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_293),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_187),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_196),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_284),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_163),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_256),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_293),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_247),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_173),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_279),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_293),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_234),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_209),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_190),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_293),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_194),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_256),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_293),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_209),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_160),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_165),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_199),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_174),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_183),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_202),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_184),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_221),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_258),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_226),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_313),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_227),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_206),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_238),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_207),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_241),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_258),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_242),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_191),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_313),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_256),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_248),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_213),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_195),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_250),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_254),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_272),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_285),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_165),
.Y(n_370)
);

BUFx2_ASAP7_75t_SL g371 ( 
.A(n_170),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_170),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_223),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_287),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_291),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_308),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_159),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_311),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_167),
.Y(n_379)
);

INVxp33_ASAP7_75t_SL g380 ( 
.A(n_164),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_167),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_236),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_197),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_236),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_229),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_231),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_158),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_161),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_312),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_332),
.B(n_267),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_338),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_323),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_338),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_338),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_388),
.B(n_158),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_336),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_323),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_329),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_338),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_338),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_329),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_314),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_333),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_333),
.Y(n_404)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_387),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_362),
.B(n_170),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_337),
.B(n_181),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_337),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_340),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_335),
.B(n_341),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_360),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_350),
.B(n_273),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_343),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_352),
.B(n_181),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_358),
.B(n_193),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_343),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_365),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_370),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_370),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_379),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_379),
.Y(n_422)
);

NAND2x1_ASAP7_75t_L g423 ( 
.A(n_381),
.B(n_194),
.Y(n_423)
);

NOR2xp67_ASAP7_75t_L g424 ( 
.A(n_377),
.B(n_166),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_381),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_382),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_382),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_384),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_383),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_384),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_342),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_345),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_346),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_324),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_371),
.Y(n_435)
);

BUFx12f_ASAP7_75t_L g436 ( 
.A(n_324),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_361),
.B(n_162),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_325),
.B(n_162),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_372),
.B(n_168),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_372),
.B(n_168),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_348),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_349),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_351),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_353),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_319),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_325),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_315),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_355),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_344),
.B(n_175),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_357),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_330),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_316),
.B(n_317),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_359),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_320),
.B(n_193),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_344),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_363),
.B(n_180),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_331),
.A2(n_255),
.B1(n_310),
.B2(n_283),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_366),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_390),
.B(n_347),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_409),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_409),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_443),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_409),
.Y(n_463)
);

AO21x2_ASAP7_75t_L g464 ( 
.A1(n_415),
.A2(n_185),
.B(n_182),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_435),
.B(n_318),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_443),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_402),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_421),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_421),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_391),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_443),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_443),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_413),
.B(n_347),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_392),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_392),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_413),
.B(n_354),
.Y(n_476)
);

OR2x2_ASAP7_75t_SL g477 ( 
.A(n_455),
.B(n_327),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_396),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_421),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_410),
.B(n_354),
.Y(n_480)
);

AO21x2_ASAP7_75t_L g481 ( 
.A1(n_416),
.A2(n_201),
.B(n_186),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_421),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_R g483 ( 
.A(n_411),
.B(n_356),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_410),
.A2(n_322),
.B1(n_326),
.B2(n_321),
.Y(n_484)
);

NAND3xp33_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_456),
.C(n_410),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_421),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_397),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_410),
.B(n_371),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_437),
.B(n_356),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_447),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_397),
.Y(n_491)
);

BUFx10_ASAP7_75t_L g492 ( 
.A(n_434),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_418),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_398),
.Y(n_494)
);

AND3x2_ASAP7_75t_L g495 ( 
.A(n_439),
.B(n_322),
.C(n_328),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_421),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_391),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_437),
.B(n_364),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_398),
.Y(n_499)
);

OR2x6_ASAP7_75t_L g500 ( 
.A(n_436),
.B(n_192),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_401),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_447),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_391),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_404),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_401),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_404),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_391),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_408),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_456),
.A2(n_380),
.B1(n_318),
.B2(n_245),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_L g510 ( 
.A1(n_456),
.A2(n_380),
.B1(n_368),
.B2(n_375),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_401),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_401),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_391),
.Y(n_513)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_391),
.Y(n_514)
);

BUFx10_ASAP7_75t_L g515 ( 
.A(n_446),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_440),
.B(n_364),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_438),
.B(n_373),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_408),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_405),
.B(n_373),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_401),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_449),
.B(n_385),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_441),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_441),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_405),
.B(n_385),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_441),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_441),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_441),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_406),
.B(n_386),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_401),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_403),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_447),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_405),
.B(n_386),
.Y(n_532)
);

BUFx10_ASAP7_75t_L g533 ( 
.A(n_429),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_441),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_L g535 ( 
.A(n_452),
.B(n_194),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_405),
.B(n_198),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_394),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_403),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_403),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_403),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_407),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_445),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_456),
.B(n_200),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_424),
.B(n_389),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_403),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_403),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_394),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_394),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_393),
.B(n_204),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_407),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_407),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_419),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_395),
.Y(n_553)
);

INVx6_ASAP7_75t_L g554 ( 
.A(n_395),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_412),
.B(n_367),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_407),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_419),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_393),
.B(n_210),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_394),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_393),
.B(n_211),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_451),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_395),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_424),
.B(n_334),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_394),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_395),
.A2(n_378),
.B1(n_376),
.B2(n_374),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_394),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_423),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_419),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_419),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_399),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_431),
.A2(n_369),
.B1(n_194),
.B2(n_266),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_444),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_431),
.A2(n_266),
.B1(n_194),
.B2(n_205),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_444),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_444),
.B(n_208),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_436),
.B(n_339),
.Y(n_576)
);

BUFx10_ASAP7_75t_L g577 ( 
.A(n_432),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_432),
.B(n_266),
.Y(n_578)
);

OAI22xp33_ASAP7_75t_L g579 ( 
.A1(n_436),
.A2(n_275),
.B1(n_220),
.B2(n_232),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_433),
.A2(n_266),
.B1(n_252),
.B2(n_309),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_423),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_399),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_457),
.B(n_175),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_448),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_433),
.B(n_244),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_417),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_417),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_417),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_442),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_442),
.B(n_178),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_448),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_448),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_458),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_450),
.B(n_246),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_399),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_458),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_450),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_400),
.B(n_212),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_420),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_453),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_400),
.B(n_214),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_420),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_400),
.B(n_215),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_453),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_420),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_458),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_414),
.B(n_178),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_412),
.B(n_179),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_460),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_597),
.Y(n_610)
);

INVx8_ASAP7_75t_L g611 ( 
.A(n_500),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_478),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_460),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_489),
.B(n_179),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_460),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_597),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_461),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_541),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_490),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_541),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_550),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_550),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_490),
.B(n_414),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_490),
.B(n_430),
.Y(n_624)
);

NAND2x1p5_ASAP7_75t_L g625 ( 
.A(n_581),
.B(n_218),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_551),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_488),
.B(n_422),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_597),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_502),
.B(n_426),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_461),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_585),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_551),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_581),
.Y(n_633)
);

OAI22xp33_ASAP7_75t_L g634 ( 
.A1(n_498),
.A2(n_283),
.B1(n_169),
.B2(n_164),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_585),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_488),
.B(n_426),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_556),
.Y(n_637)
);

INVxp67_ASAP7_75t_SL g638 ( 
.A(n_556),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_502),
.B(n_430),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_555),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_581),
.Y(n_641)
);

BUFx2_ASAP7_75t_L g642 ( 
.A(n_542),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_555),
.Y(n_643)
);

NAND3xp33_ASAP7_75t_L g644 ( 
.A(n_465),
.B(n_261),
.C(n_262),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_483),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_461),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_500),
.B(n_240),
.Y(n_647)
);

AO22x2_ASAP7_75t_L g648 ( 
.A1(n_583),
.A2(n_274),
.B1(n_296),
.B2(n_295),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_554),
.Y(n_649)
);

A2O1A1Ixp33_ASAP7_75t_L g650 ( 
.A1(n_485),
.A2(n_286),
.B(n_269),
.C(n_270),
.Y(n_650)
);

NAND2x1p5_ASAP7_75t_L g651 ( 
.A(n_553),
.B(n_249),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_462),
.B(n_422),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_553),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_493),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_606),
.B(n_428),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_562),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_561),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_462),
.B(n_422),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_484),
.B(n_428),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_562),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_474),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_477),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_474),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_463),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_466),
.B(n_425),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_475),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_475),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_463),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_531),
.B(n_425),
.Y(n_669)
);

AND2x4_ASAP7_75t_SL g670 ( 
.A(n_533),
.B(n_266),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_487),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_533),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_554),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_594),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_464),
.A2(n_216),
.B1(n_169),
.B2(n_312),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_487),
.Y(n_676)
);

AO22x2_ASAP7_75t_L g677 ( 
.A1(n_485),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_463),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_509),
.A2(n_517),
.B1(n_510),
.B2(n_528),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_467),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_491),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_473),
.B(n_228),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_466),
.B(n_425),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_531),
.B(n_427),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_491),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_586),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_554),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_476),
.B(n_228),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_586),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_587),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_587),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_494),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_608),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_494),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_533),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_589),
.B(n_427),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_499),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_471),
.B(n_427),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_471),
.B(n_216),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_499),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_589),
.B(n_259),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_600),
.B(n_277),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_554),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_504),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_600),
.B(n_277),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_519),
.B(n_280),
.Y(n_706)
);

INVx4_ASAP7_75t_L g707 ( 
.A(n_582),
.Y(n_707)
);

NAND2x1p5_ASAP7_75t_L g708 ( 
.A(n_567),
.B(n_48),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_588),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_504),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_533),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_582),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_472),
.B(n_552),
.Y(n_713)
);

BUFx4f_ASAP7_75t_L g714 ( 
.A(n_500),
.Y(n_714)
);

NAND2x1p5_ASAP7_75t_L g715 ( 
.A(n_567),
.B(n_49),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_604),
.B(n_280),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_492),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_506),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_594),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_506),
.Y(n_720)
);

AO22x2_ASAP7_75t_L g721 ( 
.A1(n_459),
.A2(n_3),
.B1(n_9),
.B2(n_10),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_508),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_472),
.B(n_216),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_508),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_575),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_477),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_552),
.B(n_216),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_604),
.B(n_577),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_582),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_557),
.B(n_216),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_588),
.Y(n_731)
);

AND2x6_ASAP7_75t_L g732 ( 
.A(n_568),
.B(n_216),
.Y(n_732)
);

OAI221xp5_ASAP7_75t_L g733 ( 
.A1(n_565),
.A2(n_310),
.B1(n_171),
.B2(n_176),
.C(n_271),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_500),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_518),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_518),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_500),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_480),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_577),
.B(n_216),
.Y(n_739)
);

BUFx4f_ASAP7_75t_L g740 ( 
.A(n_575),
.Y(n_740)
);

OAI22xp33_ASAP7_75t_L g741 ( 
.A1(n_524),
.A2(n_532),
.B1(n_300),
.B2(n_290),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_599),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_575),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_599),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_557),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_568),
.Y(n_746)
);

AO21x2_ASAP7_75t_L g747 ( 
.A1(n_464),
.A2(n_216),
.B(n_307),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_568),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_582),
.Y(n_749)
);

OR2x2_ASAP7_75t_SL g750 ( 
.A(n_579),
.B(n_171),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_577),
.B(n_217),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_577),
.B(n_306),
.Y(n_752)
);

AND2x6_ASAP7_75t_L g753 ( 
.A(n_569),
.B(n_468),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_464),
.A2(n_289),
.B1(n_271),
.B2(n_276),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_602),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_575),
.B(n_281),
.Y(n_756)
);

AO22x2_ASAP7_75t_L g757 ( 
.A1(n_521),
.A2(n_11),
.B1(n_13),
.B2(n_16),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_569),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_569),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_572),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_492),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_543),
.A2(n_219),
.B1(n_302),
.B2(n_298),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_572),
.B(n_222),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_544),
.B(n_281),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_574),
.B(n_224),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_492),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_590),
.B(n_282),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_574),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_564),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_481),
.A2(n_176),
.B1(n_276),
.B2(n_278),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_492),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_584),
.B(n_305),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_495),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_516),
.B(n_292),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_584),
.B(n_268),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_563),
.B(n_292),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_591),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_591),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_592),
.B(n_282),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_592),
.B(n_294),
.Y(n_780)
);

INVx8_ASAP7_75t_L g781 ( 
.A(n_470),
.Y(n_781)
);

CKINVDCx8_ASAP7_75t_R g782 ( 
.A(n_612),
.Y(n_782)
);

NOR2x1p5_ASAP7_75t_L g783 ( 
.A(n_695),
.B(n_278),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_669),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_636),
.B(n_481),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_654),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_693),
.B(n_481),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_693),
.B(n_679),
.Y(n_788)
);

INVx5_ASAP7_75t_L g789 ( 
.A(n_611),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_627),
.B(n_593),
.Y(n_790)
);

OR2x6_ASAP7_75t_L g791 ( 
.A(n_611),
.B(n_576),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_679),
.A2(n_593),
.B1(n_596),
.B2(n_580),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_669),
.Y(n_793)
);

NOR2x1p5_ASAP7_75t_L g794 ( 
.A(n_711),
.B(n_288),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_680),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_728),
.B(n_515),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_680),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_633),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_633),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_729),
.A2(n_558),
.B(n_603),
.Y(n_800)
);

AO22x1_ASAP7_75t_L g801 ( 
.A1(n_774),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_801)
);

AO22x1_ASAP7_75t_L g802 ( 
.A1(n_774),
.A2(n_300),
.B1(n_303),
.B2(n_301),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_627),
.B(n_596),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_640),
.B(n_607),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_638),
.B(n_602),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_633),
.Y(n_806)
);

AND2x6_ASAP7_75t_SL g807 ( 
.A(n_682),
.B(n_515),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_638),
.B(n_605),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_754),
.A2(n_573),
.B1(n_571),
.B2(n_263),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_618),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_620),
.Y(n_811)
);

NAND2x1p5_ASAP7_75t_L g812 ( 
.A(n_641),
.B(n_522),
.Y(n_812)
);

NAND2xp33_ASAP7_75t_SL g813 ( 
.A(n_717),
.B(n_294),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_741),
.A2(n_536),
.B(n_535),
.C(n_598),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_641),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_621),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_622),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_675),
.A2(n_527),
.B1(n_522),
.B2(n_523),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_SL g819 ( 
.A1(n_682),
.A2(n_515),
.B1(n_297),
.B2(n_299),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_R g820 ( 
.A(n_657),
.B(n_672),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_655),
.B(n_515),
.Y(n_821)
);

NOR2xp67_ASAP7_75t_L g822 ( 
.A(n_644),
.B(n_549),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_696),
.B(n_560),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_706),
.B(n_601),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_706),
.B(n_523),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_642),
.Y(n_826)
);

OAI21xp33_ASAP7_75t_SL g827 ( 
.A1(n_661),
.A2(n_526),
.B(n_525),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_629),
.B(n_525),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_641),
.B(n_297),
.Y(n_829)
);

INVx6_ASAP7_75t_L g830 ( 
.A(n_761),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_675),
.A2(n_526),
.B1(n_527),
.B2(n_534),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_631),
.B(n_299),
.Y(n_832)
);

OR2x6_ASAP7_75t_L g833 ( 
.A(n_611),
.B(n_468),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_729),
.Y(n_834)
);

CKINVDCx8_ASAP7_75t_R g835 ( 
.A(n_773),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_663),
.B(n_605),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_674),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_749),
.A2(n_534),
.B(n_529),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_626),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_632),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_674),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_684),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_684),
.Y(n_843)
);

NOR3xp33_ASAP7_75t_SL g844 ( 
.A(n_634),
.B(n_304),
.C(n_243),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_629),
.B(n_470),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_639),
.B(n_470),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_639),
.B(n_470),
.Y(n_847)
);

NAND2x1p5_ASAP7_75t_L g848 ( 
.A(n_740),
.B(n_468),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_662),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_666),
.B(n_497),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_610),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_635),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_719),
.B(n_497),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_667),
.B(n_497),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_671),
.B(n_497),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_719),
.A2(n_482),
.B1(n_486),
.B2(n_469),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_676),
.B(n_681),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_685),
.B(n_503),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_779),
.Y(n_859)
);

NAND2x1p5_ASAP7_75t_L g860 ( 
.A(n_740),
.B(n_469),
.Y(n_860)
);

AND2x6_ASAP7_75t_L g861 ( 
.A(n_643),
.B(n_564),
.Y(n_861)
);

INVx4_ASAP7_75t_L g862 ( 
.A(n_610),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_637),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_735),
.Y(n_864)
);

INVx5_ASAP7_75t_L g865 ( 
.A(n_753),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_692),
.B(n_479),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_694),
.B(n_479),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_610),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_741),
.A2(n_482),
.B1(n_486),
.B2(n_496),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_736),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_713),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_616),
.B(n_628),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_697),
.B(n_496),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_713),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_616),
.B(n_225),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_700),
.B(n_501),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_766),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_704),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_710),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_616),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_648),
.A2(n_538),
.B1(n_529),
.B2(n_530),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_745),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_718),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_726),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_738),
.B(n_503),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_720),
.B(n_501),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_628),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_779),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_701),
.B(n_570),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_722),
.B(n_501),
.Y(n_890)
);

INVx1_ASAP7_75t_SL g891 ( 
.A(n_738),
.Y(n_891)
);

BUFx5_ASAP7_75t_L g892 ( 
.A(n_753),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_724),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_628),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_760),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_768),
.Y(n_896)
);

OR2x6_ASAP7_75t_L g897 ( 
.A(n_771),
.B(n_505),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_777),
.Y(n_898)
);

AND2x6_ASAP7_75t_SL g899 ( 
.A(n_688),
.B(n_13),
.Y(n_899)
);

AND2x4_ASAP7_75t_SL g900 ( 
.A(n_647),
.B(n_530),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_614),
.A2(n_656),
.B1(n_653),
.B2(n_660),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_778),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_746),
.Y(n_903)
);

BUFx8_ASAP7_75t_L g904 ( 
.A(n_734),
.Y(n_904)
);

NOR2x1p5_ASAP7_75t_L g905 ( 
.A(n_767),
.B(n_230),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_749),
.B(n_520),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_614),
.B(n_623),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_748),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_758),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_645),
.Y(n_910)
);

OAI21xp33_ASAP7_75t_L g911 ( 
.A1(n_688),
.A2(n_233),
.B(n_265),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_623),
.B(n_547),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_759),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_756),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_624),
.B(n_547),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_609),
.Y(n_916)
);

OAI22xp33_ASAP7_75t_L g917 ( 
.A1(n_714),
.A2(n_235),
.B1(n_264),
.B2(n_237),
.Y(n_917)
);

INVx5_ASAP7_75t_L g918 ( 
.A(n_753),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_SL g919 ( 
.A1(n_750),
.A2(n_733),
.B1(n_645),
.B2(n_770),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_634),
.A2(n_578),
.B(n_595),
.C(n_570),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_780),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_714),
.B(n_239),
.Y(n_922)
);

INVxp33_ASAP7_75t_SL g923 ( 
.A(n_776),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_613),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_702),
.B(n_251),
.Y(n_925)
);

INVx5_ASAP7_75t_L g926 ( 
.A(n_753),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_702),
.B(n_705),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_615),
.Y(n_928)
);

NOR2x2_ASAP7_75t_L g929 ( 
.A(n_647),
.B(n_564),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_776),
.B(n_513),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_650),
.A2(n_595),
.B(n_570),
.C(n_538),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_624),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_725),
.B(n_539),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_780),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_617),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_769),
.Y(n_936)
);

AND2x2_ASAP7_75t_SL g937 ( 
.A(n_754),
.B(n_770),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_659),
.B(n_520),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_743),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_705),
.B(n_507),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_648),
.A2(n_539),
.B1(n_545),
.B2(n_546),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_677),
.A2(n_595),
.B1(n_257),
.B2(n_260),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_716),
.B(n_546),
.Y(n_943)
);

AO22x1_ASAP7_75t_L g944 ( 
.A1(n_767),
.A2(n_545),
.B1(n_540),
.B2(n_511),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_652),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_716),
.B(n_566),
.Y(n_946)
);

NAND2x1p5_ASAP7_75t_L g947 ( 
.A(n_619),
.B(n_566),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_630),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_652),
.A2(n_540),
.B(n_511),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_658),
.B(n_505),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_646),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_756),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_764),
.B(n_505),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_619),
.B(n_566),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_764),
.B(n_649),
.Y(n_955)
);

NAND2x1p5_ASAP7_75t_L g956 ( 
.A(n_707),
.B(n_566),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_772),
.A2(n_511),
.B1(n_512),
.B2(n_520),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_664),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_658),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_649),
.B(n_673),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_665),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_737),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_665),
.B(n_512),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_683),
.B(n_512),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_668),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_678),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_649),
.B(n_559),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_673),
.B(n_559),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_751),
.B(n_559),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_673),
.B(n_687),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_683),
.B(n_559),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_698),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_686),
.Y(n_973)
);

INVxp67_ASAP7_75t_SL g974 ( 
.A(n_687),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_903),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_795),
.Y(n_976)
);

INVx2_ASAP7_75t_SL g977 ( 
.A(n_797),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_788),
.A2(n_751),
.B(n_752),
.C(n_733),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_799),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_810),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_871),
.B(n_752),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_799),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_821),
.B(n_670),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_811),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_923),
.B(n_625),
.Y(n_985)
);

AOI22x1_ASAP7_75t_L g986 ( 
.A1(n_945),
.A2(n_648),
.B1(n_625),
.B2(n_677),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_799),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_816),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_806),
.Y(n_989)
);

AND3x1_ASAP7_75t_L g990 ( 
.A(n_844),
.B(n_762),
.C(n_757),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_782),
.Y(n_991)
);

INVxp67_ASAP7_75t_SL g992 ( 
.A(n_834),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_916),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_817),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_874),
.B(n_763),
.Y(n_995)
);

OR2x6_ASAP7_75t_L g996 ( 
.A(n_830),
.B(n_791),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_924),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_797),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_839),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_959),
.B(n_763),
.Y(n_1000)
);

BUFx12f_ASAP7_75t_L g1001 ( 
.A(n_826),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_SL g1002 ( 
.A1(n_937),
.A2(n_647),
.B1(n_715),
.B2(n_708),
.Y(n_1002)
);

AND3x1_ASAP7_75t_SL g1003 ( 
.A(n_905),
.B(n_721),
.C(n_757),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_961),
.B(n_765),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_891),
.B(n_910),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_806),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_928),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_935),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_837),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_840),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_838),
.A2(n_698),
.B(n_699),
.Y(n_1011)
);

AO21x2_ASAP7_75t_L g1012 ( 
.A1(n_949),
.A2(n_747),
.B(n_739),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_863),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_878),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_891),
.B(n_841),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_806),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_914),
.B(n_757),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_972),
.B(n_765),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_849),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_907),
.B(n_775),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_948),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_952),
.B(n_721),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_951),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_786),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_958),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_852),
.B(n_721),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_789),
.B(n_784),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_865),
.B(n_707),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_789),
.B(n_687),
.Y(n_1029)
);

CKINVDCx11_ASAP7_75t_R g1030 ( 
.A(n_835),
.Y(n_1030)
);

AO22x1_ASAP7_75t_L g1031 ( 
.A1(n_962),
.A2(n_677),
.B1(n_753),
.B2(n_732),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_880),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_884),
.Y(n_1033)
);

INVxp67_ASAP7_75t_L g1034 ( 
.A(n_927),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_965),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_879),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_787),
.B(n_775),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_857),
.B(n_651),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_824),
.B(n_651),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_901),
.A2(n_712),
.B1(n_703),
.B2(n_708),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_793),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_804),
.B(n_859),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_820),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_919),
.B(n_842),
.Y(n_1044)
);

AO22x1_ASAP7_75t_L g1045 ( 
.A1(n_904),
.A2(n_732),
.B1(n_723),
.B2(n_699),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_904),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_843),
.Y(n_1047)
);

NOR2x1_ASAP7_75t_L g1048 ( 
.A(n_862),
.B(n_739),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_883),
.B(n_712),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_893),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_880),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_938),
.B(n_703),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_938),
.B(n_772),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_SL g1054 ( 
.A1(n_819),
.A2(n_715),
.B1(n_723),
.B2(n_730),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_880),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_804),
.B(n_709),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_888),
.A2(n_747),
.B1(n_690),
.B2(n_755),
.Y(n_1057)
);

CKINVDCx20_ASAP7_75t_R g1058 ( 
.A(n_877),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_921),
.B(n_730),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_895),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_889),
.B(n_691),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_789),
.B(n_769),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_823),
.B(n_689),
.Y(n_1063)
);

OR2x2_ASAP7_75t_SL g1064 ( 
.A(n_830),
.B(n_727),
.Y(n_1064)
);

INVx4_ASAP7_75t_L g1065 ( 
.A(n_887),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_934),
.B(n_769),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_955),
.B(n_744),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_887),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_943),
.B(n_742),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_932),
.B(n_802),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_939),
.B(n_731),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_896),
.B(n_781),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_942),
.A2(n_727),
.B(n_507),
.C(n_513),
.Y(n_1073)
);

NAND2x1p5_ASAP7_75t_L g1074 ( 
.A(n_865),
.B(n_537),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_833),
.B(n_503),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_785),
.A2(n_732),
.B(n_537),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_801),
.B(n_732),
.Y(n_1077)
);

INVx5_ASAP7_75t_L g1078 ( 
.A(n_865),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_966),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_898),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_929),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_908),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_833),
.B(n_503),
.Y(n_1083)
);

INVx2_ASAP7_75t_SL g1084 ( 
.A(n_783),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_902),
.Y(n_1085)
);

AND2x6_ASAP7_75t_L g1086 ( 
.A(n_969),
.B(n_548),
.Y(n_1086)
);

NAND2xp33_ASAP7_75t_SL g1087 ( 
.A(n_887),
.B(n_548),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_836),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_909),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_853),
.B(n_781),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_885),
.B(n_781),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_833),
.B(n_732),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_913),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_790),
.B(n_548),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_894),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_894),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_894),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_836),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_866),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_973),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_866),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_882),
.Y(n_1102)
);

NOR2x2_ASAP7_75t_L g1103 ( 
.A(n_791),
.B(n_19),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_897),
.Y(n_1104)
);

INVx2_ASAP7_75t_SL g1105 ( 
.A(n_794),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_790),
.B(n_548),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_930),
.A2(n_547),
.B1(n_537),
.B2(n_513),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_892),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_897),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_803),
.B(n_547),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_803),
.B(n_537),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_832),
.B(n_19),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_805),
.B(n_507),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_892),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_805),
.B(n_808),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_892),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_808),
.B(n_507),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_825),
.B(n_513),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_950),
.B(n_23),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_892),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_829),
.A2(n_514),
.B1(n_100),
.B2(n_103),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_867),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_892),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_867),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_900),
.B(n_97),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_873),
.Y(n_1126)
);

INVx5_ASAP7_75t_L g1127 ( 
.A(n_918),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_918),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_950),
.B(n_26),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1044),
.A2(n_911),
.B1(n_809),
.B2(n_925),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_1128),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_SL g1132 ( 
.A1(n_986),
.A2(n_942),
.B1(n_809),
.B2(n_899),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_1104),
.B(n_791),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_976),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1082),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_998),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_SL g1137 ( 
.A1(n_981),
.A2(n_946),
.B(n_940),
.Y(n_1137)
);

OR2x6_ASAP7_75t_L g1138 ( 
.A(n_996),
.B(n_862),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_980),
.Y(n_1139)
);

INVx4_ASAP7_75t_L g1140 ( 
.A(n_1078),
.Y(n_1140)
);

AOI221xp5_ASAP7_75t_L g1141 ( 
.A1(n_978),
.A2(n_813),
.B1(n_917),
.B2(n_814),
.C(n_870),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_977),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_976),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1082),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1088),
.B(n_963),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_1128),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_1005),
.B(n_918),
.Y(n_1147)
);

INVx5_ASAP7_75t_L g1148 ( 
.A(n_1128),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1115),
.A2(n_792),
.B1(n_926),
.B2(n_818),
.Y(n_1149)
);

INVx4_ASAP7_75t_L g1150 ( 
.A(n_1078),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_979),
.Y(n_1151)
);

INVxp67_ASAP7_75t_L g1152 ( 
.A(n_1015),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_1058),
.Y(n_1153)
);

OR2x6_ASAP7_75t_L g1154 ( 
.A(n_996),
.B(n_868),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1089),
.Y(n_1155)
);

AOI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1045),
.A2(n_944),
.B(n_800),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_979),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1128),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1044),
.A2(n_926),
.B1(n_831),
.B2(n_828),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1098),
.B(n_963),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_984),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_988),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1089),
.Y(n_1163)
);

BUFx4_ASAP7_75t_SL g1164 ( 
.A(n_1046),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1099),
.B(n_964),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_994),
.Y(n_1166)
);

BUFx12f_ASAP7_75t_L g1167 ( 
.A(n_1030),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_1009),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_1019),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_1033),
.B(n_953),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_1058),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_992),
.A2(n_926),
.B1(n_864),
.B2(n_964),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1024),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1078),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_985),
.A2(n_922),
.B1(n_796),
.B2(n_875),
.Y(n_1175)
);

AOI221xp5_ASAP7_75t_L g1176 ( 
.A1(n_990),
.A2(n_920),
.B1(n_827),
.B2(n_869),
.C(n_873),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1104),
.B(n_868),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_991),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1034),
.B(n_995),
.Y(n_1179)
);

AND2x2_ASAP7_75t_SL g1180 ( 
.A(n_1017),
.B(n_807),
.Y(n_1180)
);

INVx5_ASAP7_75t_L g1181 ( 
.A(n_1078),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_1001),
.Y(n_1182)
);

AOI221xp5_ASAP7_75t_L g1183 ( 
.A1(n_1112),
.A2(n_886),
.B1(n_890),
.B2(n_876),
.C(n_881),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1127),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1093),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1101),
.B(n_1122),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_991),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1037),
.A2(n_906),
.B(n_971),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1093),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_983),
.B(n_1042),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_1001),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_979),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_979),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1039),
.A2(n_822),
.B(n_856),
.C(n_845),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_SL g1195 ( 
.A1(n_1002),
.A2(n_861),
.B1(n_815),
.B2(n_798),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_975),
.Y(n_1196)
);

NAND2x1_ASAP7_75t_SL g1197 ( 
.A(n_1029),
.B(n_798),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_975),
.Y(n_1198)
);

INVxp67_ASAP7_75t_L g1199 ( 
.A(n_1081),
.Y(n_1199)
);

BUFx12f_ASAP7_75t_L g1200 ( 
.A(n_1030),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_999),
.Y(n_1201)
);

INVx5_ASAP7_75t_L g1202 ( 
.A(n_1127),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1020),
.A2(n_906),
.B(n_971),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1102),
.Y(n_1204)
);

BUFx12f_ASAP7_75t_L g1205 ( 
.A(n_1024),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1000),
.A2(n_847),
.B(n_846),
.C(n_886),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1124),
.B(n_876),
.Y(n_1207)
);

NOR2x1p5_ASAP7_75t_L g1208 ( 
.A(n_1043),
.B(n_974),
.Y(n_1208)
);

OAI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1034),
.A2(n_897),
.B1(n_912),
.B2(n_915),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1043),
.B(n_1004),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_982),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1126),
.B(n_890),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_1022),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1046),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_985),
.A2(n_1070),
.B1(n_1084),
.B2(n_1105),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1018),
.A2(n_933),
.B1(n_872),
.B2(n_815),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_996),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_982),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_992),
.A2(n_941),
.B1(n_851),
.B2(n_848),
.Y(n_1219)
);

INVxp67_ASAP7_75t_L g1220 ( 
.A(n_1041),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1064),
.A2(n_1010),
.B1(n_1060),
.B2(n_1050),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1053),
.B(n_851),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1026),
.B(n_933),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_1097),
.Y(n_1224)
);

INVxp67_ASAP7_75t_SL g1225 ( 
.A(n_1041),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1056),
.A2(n_861),
.B1(n_960),
.B2(n_970),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1047),
.A2(n_861),
.B1(n_936),
.B2(n_854),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1102),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1056),
.A2(n_861),
.B1(n_968),
.B2(n_967),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1013),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1097),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_993),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_982),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1011),
.A2(n_931),
.B(n_949),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1059),
.B(n_936),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1014),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1127),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1036),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1080),
.Y(n_1239)
);

INVxp67_ASAP7_75t_L g1240 ( 
.A(n_1047),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1109),
.B(n_858),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_993),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_982),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_997),
.Y(n_1244)
);

INVxp67_ASAP7_75t_SL g1245 ( 
.A(n_1096),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1016),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_997),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1127),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_1092),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1063),
.B(n_855),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1096),
.Y(n_1251)
);

AND2x2_ASAP7_75t_SL g1252 ( 
.A(n_1125),
.B(n_954),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1007),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1016),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1085),
.A2(n_848),
.B1(n_860),
.B2(n_812),
.Y(n_1255)
);

AOI221xp5_ASAP7_75t_L g1256 ( 
.A1(n_1119),
.A2(n_850),
.B1(n_957),
.B2(n_860),
.C(n_812),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_1016),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1109),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1038),
.A2(n_1067),
.B(n_1129),
.C(n_1057),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1125),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1007),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1067),
.A2(n_956),
.B(n_947),
.C(n_38),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1077),
.A2(n_1071),
.B1(n_1054),
.B2(n_1100),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1016),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1071),
.A2(n_947),
.B1(n_956),
.B2(n_514),
.Y(n_1265)
);

NAND3xp33_ASAP7_75t_L g1266 ( 
.A(n_1121),
.B(n_514),
.C(n_36),
.Y(n_1266)
);

INVxp67_ASAP7_75t_SL g1267 ( 
.A(n_1051),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1051),
.Y(n_1268)
);

NAND2x1p5_ASAP7_75t_L g1269 ( 
.A(n_1062),
.B(n_514),
.Y(n_1269)
);

INVx5_ASAP7_75t_L g1270 ( 
.A(n_1051),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1051),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1049),
.A2(n_27),
.B1(n_38),
.B2(n_42),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1076),
.A2(n_514),
.B(n_110),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1055),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1061),
.B(n_514),
.Y(n_1275)
);

OR2x6_ASAP7_75t_L g1276 ( 
.A(n_1092),
.B(n_1029),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1052),
.B(n_43),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1066),
.B(n_43),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1069),
.B(n_44),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1055),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1055),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1008),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1021),
.Y(n_1283)
);

NAND3xp33_ASAP7_75t_L g1284 ( 
.A(n_1130),
.B(n_1031),
.C(n_1040),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1234),
.A2(n_1118),
.B(n_1113),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1234),
.A2(n_1073),
.B(n_1117),
.Y(n_1286)
);

AO21x2_ASAP7_75t_L g1287 ( 
.A1(n_1273),
.A2(n_1156),
.B(n_1259),
.Y(n_1287)
);

AOI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1273),
.A2(n_1091),
.B(n_1107),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1135),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1188),
.A2(n_1110),
.B(n_1106),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1181),
.B(n_1062),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1139),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_1134),
.Y(n_1293)
);

O2A1O1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1221),
.A2(n_1072),
.B(n_1100),
.C(n_1023),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1161),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1260),
.B(n_1027),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1179),
.B(n_1066),
.Y(n_1297)
);

INVx4_ASAP7_75t_L g1298 ( 
.A(n_1148),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1215),
.A2(n_1090),
.B1(n_1027),
.B2(n_1048),
.Y(n_1299)
);

BUFx12f_ASAP7_75t_L g1300 ( 
.A(n_1167),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1223),
.B(n_1025),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1188),
.A2(n_1111),
.B(n_1094),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1162),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1203),
.A2(n_1123),
.B(n_1120),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1190),
.B(n_1023),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1166),
.Y(n_1306)
);

INVxp33_ASAP7_75t_SL g1307 ( 
.A(n_1164),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1266),
.A2(n_1090),
.B(n_1028),
.Y(n_1308)
);

INVx5_ASAP7_75t_L g1309 ( 
.A(n_1181),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1203),
.A2(n_1123),
.B(n_1120),
.Y(n_1310)
);

OA21x2_ASAP7_75t_L g1311 ( 
.A1(n_1176),
.A2(n_1116),
.B(n_1114),
.Y(n_1311)
);

O2A1O1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1221),
.A2(n_1021),
.B(n_1025),
.C(n_1079),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1132),
.A2(n_1035),
.B1(n_1079),
.B2(n_1003),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1169),
.Y(n_1314)
);

OA21x2_ASAP7_75t_L g1315 ( 
.A1(n_1176),
.A2(n_1116),
.B(n_1114),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1270),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1201),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1276),
.B(n_1027),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1144),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1137),
.A2(n_1108),
.B(n_1028),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1255),
.A2(n_1108),
.B(n_1074),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1213),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1148),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1255),
.A2(n_1074),
.B(n_1035),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1155),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1252),
.A2(n_1029),
.B1(n_1062),
.B2(n_1092),
.Y(n_1326)
);

AOI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1172),
.A2(n_1083),
.B(n_1075),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1163),
.Y(n_1328)
);

AO21x2_ASAP7_75t_L g1329 ( 
.A1(n_1172),
.A2(n_1209),
.B(n_1262),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1266),
.A2(n_1003),
.B(n_1087),
.C(n_1075),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1222),
.A2(n_987),
.B(n_1095),
.Y(n_1331)
);

AOI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1219),
.A2(n_1083),
.B(n_1012),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1230),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1141),
.A2(n_1012),
.B(n_1086),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1132),
.A2(n_1086),
.B1(n_1103),
.B2(n_987),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1213),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1148),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1173),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1185),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1187),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1222),
.A2(n_989),
.B(n_1095),
.Y(n_1341)
);

AO21x1_ASAP7_75t_L g1342 ( 
.A1(n_1272),
.A2(n_1277),
.B(n_1149),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1219),
.A2(n_989),
.B(n_1006),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1275),
.A2(n_1006),
.B(n_1032),
.Y(n_1344)
);

INVxp67_ASAP7_75t_SL g1345 ( 
.A(n_1186),
.Y(n_1345)
);

INVxp67_ASAP7_75t_L g1346 ( 
.A(n_1136),
.Y(n_1346)
);

O2A1O1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1272),
.A2(n_1210),
.B(n_1159),
.C(n_1186),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1270),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1275),
.A2(n_1263),
.B(n_1256),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1189),
.Y(n_1350)
);

INVxp67_ASAP7_75t_SL g1351 ( 
.A(n_1145),
.Y(n_1351)
);

A2O1A1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1149),
.A2(n_1087),
.B(n_1103),
.C(n_1032),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1256),
.A2(n_1086),
.B(n_1068),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1169),
.A2(n_1065),
.B1(n_1068),
.B2(n_1055),
.Y(n_1354)
);

A2O1A1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1141),
.A2(n_1086),
.B(n_1068),
.C(n_68),
.Y(n_1355)
);

O2A1O1Ixp33_ASAP7_75t_SL g1356 ( 
.A1(n_1194),
.A2(n_1086),
.B(n_1068),
.C(n_69),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1236),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1276),
.B(n_1065),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1232),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_SL g1360 ( 
.A1(n_1159),
.A2(n_52),
.B(n_57),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1206),
.A2(n_71),
.B(n_78),
.Y(n_1361)
);

A2O1A1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1183),
.A2(n_82),
.B(n_104),
.C(n_108),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1276),
.B(n_111),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1180),
.A2(n_155),
.B1(n_122),
.B2(n_127),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1277),
.A2(n_117),
.B(n_128),
.Y(n_1365)
);

OAI21xp33_ASAP7_75t_L g1366 ( 
.A1(n_1175),
.A2(n_132),
.B(n_135),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1238),
.Y(n_1367)
);

A2O1A1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1183),
.A2(n_146),
.B(n_152),
.C(n_1145),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1225),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1196),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1152),
.B(n_1235),
.Y(n_1371)
);

BUFx12f_ASAP7_75t_L g1372 ( 
.A(n_1200),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1250),
.A2(n_1165),
.B(n_1160),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1242),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1148),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1250),
.A2(n_1160),
.B(n_1165),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1199),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1220),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1207),
.A2(n_1212),
.B(n_1283),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1240),
.B(n_1220),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1279),
.A2(n_1226),
.B(n_1216),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1239),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1174),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_SL g1384 ( 
.A1(n_1279),
.A2(n_1212),
.B(n_1207),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1261),
.A2(n_1265),
.B(n_1237),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1198),
.Y(n_1386)
);

OA21x2_ASAP7_75t_L g1387 ( 
.A1(n_1227),
.A2(n_1229),
.B(n_1228),
.Y(n_1387)
);

OR2x6_ASAP7_75t_L g1388 ( 
.A(n_1138),
.B(n_1154),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1204),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1231),
.Y(n_1390)
);

OAI222xp33_ASAP7_75t_L g1391 ( 
.A1(n_1195),
.A2(n_1147),
.B1(n_1138),
.B2(n_1154),
.C1(n_1217),
.C2(n_1170),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1195),
.A2(n_1154),
.B1(n_1138),
.B2(n_1208),
.Y(n_1392)
);

BUFx2_ASAP7_75t_R g1393 ( 
.A(n_1214),
.Y(n_1393)
);

O2A1O1Ixp33_ASAP7_75t_SL g1394 ( 
.A1(n_1280),
.A2(n_1267),
.B(n_1244),
.C(n_1282),
.Y(n_1394)
);

INVx1_ASAP7_75t_SL g1395 ( 
.A(n_1142),
.Y(n_1395)
);

AO21x1_ASAP7_75t_L g1396 ( 
.A1(n_1241),
.A2(n_1245),
.B(n_1140),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1174),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1247),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1181),
.A2(n_1202),
.B(n_1140),
.Y(n_1399)
);

AO31x2_ASAP7_75t_L g1400 ( 
.A1(n_1253),
.A2(n_1248),
.A3(n_1150),
.B(n_1254),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1184),
.A2(n_1249),
.B(n_1131),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1181),
.A2(n_1202),
.B(n_1248),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_1153),
.Y(n_1403)
);

AO22x1_ASAP7_75t_L g1404 ( 
.A1(n_1258),
.A2(n_1133),
.B1(n_1177),
.B2(n_1178),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1251),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1249),
.A2(n_1131),
.B(n_1158),
.Y(n_1406)
);

AOI221xp5_ASAP7_75t_L g1407 ( 
.A1(n_1278),
.A2(n_1133),
.B1(n_1168),
.B2(n_1143),
.C(n_1171),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1205),
.A2(n_1182),
.B1(n_1191),
.B2(n_1202),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1264),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1241),
.B(n_1177),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1257),
.Y(n_1411)
);

OA21x2_ASAP7_75t_L g1412 ( 
.A1(n_1197),
.A2(n_1274),
.B(n_1271),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1270),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1233),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1224),
.B(n_1146),
.Y(n_1415)
);

AO31x2_ASAP7_75t_L g1416 ( 
.A1(n_1150),
.A2(n_1202),
.A3(n_1270),
.B(n_1269),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1146),
.A2(n_1158),
.B(n_1269),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1268),
.Y(n_1418)
);

AO21x1_ASAP7_75t_L g1419 ( 
.A1(n_1151),
.A2(n_1157),
.B(n_1192),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1151),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1151),
.B(n_1157),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1157),
.Y(n_1422)
);

O2A1O1Ixp33_ASAP7_75t_SL g1423 ( 
.A1(n_1192),
.A2(n_1193),
.B(n_1211),
.C(n_1218),
.Y(n_1423)
);

OAI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1192),
.A2(n_1193),
.B1(n_1211),
.B2(n_1218),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1193),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1211),
.B(n_1218),
.Y(n_1426)
);

INVx4_ASAP7_75t_L g1427 ( 
.A(n_1243),
.Y(n_1427)
);

AOI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1243),
.A2(n_1246),
.B(n_1281),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1243),
.Y(n_1429)
);

O2A1O1Ixp33_ASAP7_75t_SL g1430 ( 
.A1(n_1246),
.A2(n_978),
.B(n_1262),
.C(n_1259),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1338),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1345),
.B(n_1246),
.Y(n_1432)
);

AOI221xp5_ASAP7_75t_L g1433 ( 
.A1(n_1347),
.A2(n_1281),
.B1(n_1368),
.B2(n_1430),
.C(n_1342),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1284),
.A2(n_1281),
.B1(n_1297),
.B2(n_1361),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1335),
.A2(n_1366),
.B1(n_1364),
.B2(n_1381),
.Y(n_1435)
);

BUFx8_ASAP7_75t_L g1436 ( 
.A(n_1300),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_SL g1437 ( 
.A(n_1308),
.B(n_1355),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1307),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1289),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1301),
.B(n_1305),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1322),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1335),
.A2(n_1364),
.B1(n_1384),
.B2(n_1329),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1319),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1371),
.B(n_1322),
.Y(n_1444)
);

AOI21xp33_ASAP7_75t_L g1445 ( 
.A1(n_1347),
.A2(n_1329),
.B(n_1299),
.Y(n_1445)
);

CKINVDCx8_ASAP7_75t_R g1446 ( 
.A(n_1409),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1336),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1336),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1345),
.B(n_1351),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1369),
.B(n_1405),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1355),
.A2(n_1313),
.B1(n_1352),
.B2(n_1407),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1292),
.Y(n_1452)
);

INVx4_ASAP7_75t_SL g1453 ( 
.A(n_1416),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1313),
.A2(n_1377),
.B1(n_1378),
.B2(n_1403),
.Y(n_1454)
);

A2O1A1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1368),
.A2(n_1362),
.B(n_1330),
.C(n_1352),
.Y(n_1455)
);

AOI221xp5_ASAP7_75t_L g1456 ( 
.A1(n_1430),
.A2(n_1362),
.B1(n_1360),
.B2(n_1346),
.C(n_1356),
.Y(n_1456)
);

AOI221xp5_ASAP7_75t_L g1457 ( 
.A1(n_1346),
.A2(n_1356),
.B1(n_1395),
.B2(n_1314),
.C(n_1330),
.Y(n_1457)
);

BUFx12f_ASAP7_75t_L g1458 ( 
.A(n_1372),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1378),
.A2(n_1351),
.B1(n_1392),
.B2(n_1388),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1318),
.B(n_1410),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1369),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1388),
.A2(n_1363),
.B1(n_1287),
.B2(n_1357),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1318),
.B(n_1411),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1390),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1339),
.Y(n_1465)
);

AOI221xp5_ASAP7_75t_L g1466 ( 
.A1(n_1380),
.A2(n_1391),
.B1(n_1294),
.B2(n_1312),
.C(n_1367),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1388),
.B(n_1358),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1332),
.Y(n_1468)
);

INVx1_ASAP7_75t_SL g1469 ( 
.A(n_1340),
.Y(n_1469)
);

OAI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1295),
.A2(n_1303),
.B1(n_1382),
.B2(n_1306),
.Y(n_1470)
);

INVx4_ASAP7_75t_L g1471 ( 
.A(n_1316),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1363),
.A2(n_1287),
.B1(n_1333),
.B2(n_1317),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1350),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1370),
.B(n_1386),
.Y(n_1474)
);

AO21x2_ASAP7_75t_L g1475 ( 
.A1(n_1288),
.A2(n_1286),
.B(n_1327),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1408),
.A2(n_1326),
.B1(n_1340),
.B2(n_1414),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_1390),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1373),
.B(n_1376),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1408),
.A2(n_1296),
.B1(n_1293),
.B2(n_1415),
.Y(n_1479)
);

AO22x1_ASAP7_75t_L g1480 ( 
.A1(n_1293),
.A2(n_1309),
.B1(n_1296),
.B2(n_1358),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1389),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1418),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1373),
.B(n_1398),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1316),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1325),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1373),
.A2(n_1312),
.B(n_1394),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1425),
.B(n_1328),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1331),
.Y(n_1488)
);

AOI221xp5_ASAP7_75t_L g1489 ( 
.A1(n_1391),
.A2(n_1294),
.B1(n_1404),
.B2(n_1394),
.C(n_1415),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1341),
.Y(n_1490)
);

INVx1_ASAP7_75t_SL g1491 ( 
.A(n_1393),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1425),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1359),
.Y(n_1493)
);

BUFx8_ASAP7_75t_L g1494 ( 
.A(n_1420),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1291),
.A2(n_1354),
.B1(n_1417),
.B2(n_1424),
.Y(n_1495)
);

AOI22x1_ASAP7_75t_L g1496 ( 
.A1(n_1399),
.A2(n_1402),
.B1(n_1291),
.B2(n_1413),
.Y(n_1496)
);

INVx2_ASAP7_75t_SL g1497 ( 
.A(n_1422),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1396),
.B(n_1397),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1359),
.B(n_1374),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1374),
.Y(n_1500)
);

BUFx12f_ASAP7_75t_L g1501 ( 
.A(n_1422),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1426),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1379),
.B(n_1383),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1344),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1316),
.Y(n_1505)
);

CKINVDCx8_ASAP7_75t_R g1506 ( 
.A(n_1426),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1383),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1290),
.A2(n_1302),
.B(n_1320),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1424),
.A2(n_1309),
.B1(n_1412),
.B2(n_1413),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1349),
.B(n_1400),
.Y(n_1510)
);

OR2x6_ASAP7_75t_L g1511 ( 
.A(n_1353),
.B(n_1343),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_1316),
.Y(n_1512)
);

NAND2x1p5_ASAP7_75t_L g1513 ( 
.A(n_1309),
.B(n_1337),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1365),
.A2(n_1387),
.B1(n_1334),
.B2(n_1311),
.Y(n_1514)
);

BUFx10_ASAP7_75t_L g1515 ( 
.A(n_1421),
.Y(n_1515)
);

NAND3xp33_ASAP7_75t_SL g1516 ( 
.A(n_1419),
.B(n_1421),
.C(n_1298),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1397),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1406),
.B(n_1401),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1311),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1348),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1365),
.A2(n_1387),
.B1(n_1334),
.B2(n_1315),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1400),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1315),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1323),
.B(n_1375),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1387),
.A2(n_1285),
.B1(n_1412),
.B2(n_1385),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_SL g1526 ( 
.A1(n_1309),
.A2(n_1348),
.B1(n_1298),
.B2(n_1337),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1422),
.Y(n_1527)
);

AOI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1428),
.A2(n_1324),
.B(n_1321),
.Y(n_1528)
);

OAI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1348),
.A2(n_1285),
.B1(n_1427),
.B2(n_1429),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1400),
.B(n_1427),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1429),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1304),
.Y(n_1532)
);

O2A1O1Ixp5_ASAP7_75t_SL g1533 ( 
.A1(n_1285),
.A2(n_1310),
.B(n_1423),
.C(n_1416),
.Y(n_1533)
);

AOI21xp33_ASAP7_75t_L g1534 ( 
.A1(n_1348),
.A2(n_1429),
.B(n_1416),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1429),
.B(n_1416),
.Y(n_1535)
);

AND2x4_ASAP7_75t_SL g1536 ( 
.A(n_1305),
.B(n_1058),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1338),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1342),
.A2(n_937),
.B1(n_679),
.B2(n_788),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1342),
.A2(n_937),
.B1(n_679),
.B2(n_788),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1342),
.A2(n_937),
.B1(n_679),
.B2(n_788),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1335),
.A2(n_923),
.B1(n_1132),
.B2(n_937),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1388),
.B(n_1318),
.Y(n_1542)
);

CKINVDCx20_ASAP7_75t_R g1543 ( 
.A(n_1338),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1342),
.A2(n_937),
.B1(n_679),
.B2(n_788),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1342),
.A2(n_937),
.B1(n_679),
.B2(n_788),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1338),
.Y(n_1546)
);

OAI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1344),
.A2(n_1302),
.B(n_1290),
.Y(n_1547)
);

INVx5_ASAP7_75t_L g1548 ( 
.A(n_1511),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1461),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1444),
.B(n_1441),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1464),
.Y(n_1551)
);

AO31x2_ASAP7_75t_L g1552 ( 
.A1(n_1486),
.A2(n_1455),
.A3(n_1523),
.B(n_1519),
.Y(n_1552)
);

NOR3xp33_ASAP7_75t_SL g1553 ( 
.A(n_1541),
.B(n_1451),
.C(n_1438),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1460),
.B(n_1440),
.Y(n_1554)
);

CKINVDCx16_ASAP7_75t_R g1555 ( 
.A(n_1431),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1463),
.B(n_1536),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1461),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1482),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1447),
.B(n_1448),
.Y(n_1559)
);

OR2x6_ASAP7_75t_L g1560 ( 
.A(n_1480),
.B(n_1511),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1449),
.B(n_1450),
.Y(n_1561)
);

OAI21xp5_ASAP7_75t_SL g1562 ( 
.A1(n_1435),
.A2(n_1545),
.B(n_1544),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_R g1563 ( 
.A(n_1537),
.B(n_1546),
.Y(n_1563)
);

NAND2xp33_ASAP7_75t_R g1564 ( 
.A(n_1498),
.B(n_1467),
.Y(n_1564)
);

INVxp33_ASAP7_75t_L g1565 ( 
.A(n_1487),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1452),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1542),
.B(n_1502),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1470),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_R g1569 ( 
.A(n_1506),
.B(n_1543),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1481),
.Y(n_1570)
);

BUFx12f_ASAP7_75t_L g1571 ( 
.A(n_1436),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1474),
.B(n_1432),
.Y(n_1572)
);

BUFx12f_ASAP7_75t_L g1573 ( 
.A(n_1436),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1470),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1483),
.Y(n_1575)
);

NAND2xp33_ASAP7_75t_SL g1576 ( 
.A(n_1437),
.B(n_1435),
.Y(n_1576)
);

OAI21xp33_ASAP7_75t_L g1577 ( 
.A1(n_1437),
.A2(n_1538),
.B(n_1539),
.Y(n_1577)
);

OR2x6_ASAP7_75t_L g1578 ( 
.A(n_1511),
.B(n_1510),
.Y(n_1578)
);

BUFx4f_ASAP7_75t_SL g1579 ( 
.A(n_1458),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1538),
.B(n_1539),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1540),
.B(n_1544),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1493),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1478),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1455),
.A2(n_1434),
.B(n_1456),
.Y(n_1584)
);

INVx4_ASAP7_75t_L g1585 ( 
.A(n_1512),
.Y(n_1585)
);

NAND2xp33_ASAP7_75t_SL g1586 ( 
.A(n_1454),
.B(n_1476),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1446),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1485),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1515),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1540),
.B(n_1545),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1503),
.B(n_1459),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1530),
.B(n_1467),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1459),
.B(n_1535),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1542),
.B(n_1492),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1491),
.Y(n_1595)
);

BUFx6f_ASAP7_75t_L g1596 ( 
.A(n_1515),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1498),
.B(n_1499),
.Y(n_1597)
);

INVxp67_ASAP7_75t_L g1598 ( 
.A(n_1488),
.Y(n_1598)
);

INVx3_ASAP7_75t_SL g1599 ( 
.A(n_1469),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1439),
.B(n_1473),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1530),
.B(n_1517),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1434),
.B(n_1479),
.Y(n_1602)
);

NAND3xp33_ASAP7_75t_L g1603 ( 
.A(n_1457),
.B(n_1433),
.C(n_1445),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1500),
.Y(n_1604)
);

NAND2xp33_ASAP7_75t_SL g1605 ( 
.A(n_1454),
.B(n_1477),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1507),
.B(n_1462),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1494),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1527),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1443),
.B(n_1465),
.Y(n_1609)
);

INVxp67_ASAP7_75t_L g1610 ( 
.A(n_1488),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_R g1611 ( 
.A(n_1516),
.B(n_1484),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1522),
.B(n_1490),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1490),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_R g1614 ( 
.A(n_1516),
.B(n_1484),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1462),
.B(n_1472),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1472),
.B(n_1524),
.Y(n_1616)
);

AND2x2_ASAP7_75t_SL g1617 ( 
.A(n_1442),
.B(n_1514),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1504),
.B(n_1475),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1532),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1552),
.B(n_1514),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1599),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1552),
.B(n_1521),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1613),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1584),
.A2(n_1442),
.B1(n_1521),
.B2(n_1489),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1613),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1552),
.Y(n_1626)
);

NOR2x1_ASAP7_75t_L g1627 ( 
.A(n_1560),
.B(n_1618),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1619),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1597),
.B(n_1583),
.Y(n_1629)
);

INVx3_ASAP7_75t_SL g1630 ( 
.A(n_1607),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1589),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1557),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1566),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1583),
.B(n_1468),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1548),
.B(n_1453),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1549),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1549),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1575),
.B(n_1565),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1561),
.B(n_1532),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1576),
.A2(n_1466),
.B1(n_1495),
.B2(n_1496),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1548),
.B(n_1518),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1560),
.B(n_1518),
.Y(n_1642)
);

INVx2_ASAP7_75t_SL g1643 ( 
.A(n_1551),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1552),
.B(n_1525),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1578),
.B(n_1525),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1570),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1568),
.B(n_1529),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1578),
.B(n_1475),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1565),
.B(n_1547),
.Y(n_1649)
);

INVx5_ASAP7_75t_L g1650 ( 
.A(n_1560),
.Y(n_1650)
);

INVx1_ASAP7_75t_SL g1651 ( 
.A(n_1599),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1563),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1582),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1588),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1619),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1574),
.B(n_1509),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1616),
.B(n_1508),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1559),
.B(n_1550),
.Y(n_1658)
);

NOR2x1_ASAP7_75t_L g1659 ( 
.A(n_1551),
.B(n_1527),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1598),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1629),
.B(n_1578),
.Y(n_1661)
);

OAI221xp5_ASAP7_75t_L g1662 ( 
.A1(n_1640),
.A2(n_1586),
.B1(n_1562),
.B2(n_1553),
.C(n_1577),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1629),
.B(n_1617),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1657),
.B(n_1617),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1638),
.B(n_1572),
.Y(n_1665)
);

OAI21xp33_ASAP7_75t_L g1666 ( 
.A1(n_1624),
.A2(n_1553),
.B(n_1602),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1638),
.B(n_1591),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1621),
.B(n_1603),
.Y(n_1668)
);

NAND3xp33_ASAP7_75t_L g1669 ( 
.A(n_1624),
.B(n_1602),
.C(n_1605),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1621),
.A2(n_1580),
.B1(n_1590),
.B2(n_1581),
.Y(n_1670)
);

OAI21xp33_ASAP7_75t_SL g1671 ( 
.A1(n_1659),
.A2(n_1615),
.B(n_1606),
.Y(n_1671)
);

NAND4xp25_ASAP7_75t_L g1672 ( 
.A(n_1656),
.B(n_1593),
.C(n_1564),
.D(n_1610),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1658),
.B(n_1554),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1643),
.B(n_1657),
.Y(n_1674)
);

NAND3xp33_ASAP7_75t_L g1675 ( 
.A(n_1647),
.B(n_1564),
.C(n_1598),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1658),
.B(n_1594),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1639),
.B(n_1601),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_SL g1678 ( 
.A(n_1659),
.B(n_1589),
.Y(n_1678)
);

NAND3xp33_ASAP7_75t_L g1679 ( 
.A(n_1647),
.B(n_1610),
.C(n_1609),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1651),
.A2(n_1526),
.B1(n_1558),
.B2(n_1589),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1651),
.B(n_1596),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1639),
.B(n_1604),
.Y(n_1682)
);

OA21x2_ASAP7_75t_L g1683 ( 
.A1(n_1626),
.A2(n_1612),
.B(n_1534),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1656),
.B(n_1567),
.Y(n_1684)
);

NAND3xp33_ASAP7_75t_L g1685 ( 
.A(n_1627),
.B(n_1634),
.C(n_1648),
.Y(n_1685)
);

NAND4xp25_ASAP7_75t_L g1686 ( 
.A(n_1627),
.B(n_1600),
.C(n_1556),
.D(n_1526),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1634),
.B(n_1592),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1645),
.B(n_1592),
.Y(n_1688)
);

NAND4xp25_ASAP7_75t_L g1689 ( 
.A(n_1644),
.B(n_1531),
.C(n_1585),
.D(n_1608),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1631),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1643),
.B(n_1596),
.Y(n_1691)
);

NAND3xp33_ASAP7_75t_L g1692 ( 
.A(n_1648),
.B(n_1596),
.C(n_1589),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1633),
.B(n_1596),
.Y(n_1693)
);

OA21x2_ASAP7_75t_L g1694 ( 
.A1(n_1626),
.A2(n_1528),
.B(n_1524),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1650),
.A2(n_1513),
.B1(n_1471),
.B2(n_1595),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1633),
.B(n_1608),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1620),
.A2(n_1622),
.B1(n_1644),
.B2(n_1649),
.C(n_1632),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1620),
.A2(n_1571),
.B1(n_1573),
.B2(n_1579),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1646),
.B(n_1611),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1645),
.B(n_1614),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1646),
.B(n_1611),
.Y(n_1701)
);

NAND3xp33_ASAP7_75t_SL g1702 ( 
.A(n_1652),
.B(n_1569),
.C(n_1614),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1632),
.B(n_1585),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1654),
.B(n_1533),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1667),
.B(n_1636),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1700),
.B(n_1642),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1679),
.B(n_1685),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1699),
.B(n_1649),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1694),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1692),
.B(n_1650),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1682),
.B(n_1637),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1694),
.Y(n_1712)
);

INVx2_ASAP7_75t_SL g1713 ( 
.A(n_1690),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1700),
.B(n_1642),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1663),
.B(n_1642),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1697),
.B(n_1660),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1678),
.B(n_1650),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1704),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1696),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1694),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1701),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1663),
.B(n_1642),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1688),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1677),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1688),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1703),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1678),
.Y(n_1727)
);

NAND4xp25_ASAP7_75t_L g1728 ( 
.A(n_1662),
.B(n_1620),
.C(n_1622),
.D(n_1644),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1693),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1665),
.B(n_1637),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1664),
.B(n_1660),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1674),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1664),
.B(n_1636),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1661),
.B(n_1650),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1673),
.B(n_1655),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1661),
.B(n_1650),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1691),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1671),
.B(n_1650),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1687),
.B(n_1650),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1676),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1681),
.B(n_1645),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1709),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1721),
.B(n_1668),
.Y(n_1743)
);

NAND2x1p5_ASAP7_75t_L g1744 ( 
.A(n_1710),
.B(n_1683),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1721),
.B(n_1630),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1711),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1727),
.Y(n_1747)
);

AOI211xp5_ASAP7_75t_L g1748 ( 
.A1(n_1728),
.A2(n_1666),
.B(n_1669),
.C(n_1670),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1728),
.B(n_1630),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1726),
.B(n_1668),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1718),
.B(n_1684),
.Y(n_1751)
);

INVx2_ASAP7_75t_SL g1752 ( 
.A(n_1717),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1711),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1734),
.B(n_1698),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_SL g1755 ( 
.A(n_1710),
.B(n_1675),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1726),
.B(n_1681),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1707),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1734),
.B(n_1698),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1730),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1718),
.B(n_1672),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1709),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1738),
.B(n_1648),
.Y(n_1762)
);

INVxp67_ASAP7_75t_SL g1763 ( 
.A(n_1707),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1717),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1719),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1719),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1730),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1716),
.B(n_1625),
.Y(n_1768)
);

INVx5_ASAP7_75t_L g1769 ( 
.A(n_1710),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1738),
.B(n_1643),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1736),
.B(n_1631),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1736),
.B(n_1631),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1705),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1723),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1736),
.B(n_1631),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1705),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1729),
.B(n_1686),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1736),
.B(n_1631),
.Y(n_1778)
);

NOR2xp67_ASAP7_75t_L g1779 ( 
.A(n_1717),
.B(n_1702),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1716),
.B(n_1623),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1733),
.B(n_1623),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1723),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1715),
.B(n_1631),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1744),
.Y(n_1784)
);

AOI322xp5_ASAP7_75t_L g1785 ( 
.A1(n_1763),
.A2(n_1710),
.A3(n_1740),
.B1(n_1724),
.B2(n_1741),
.C1(n_1717),
.C2(n_1731),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1754),
.B(n_1722),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1782),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1779),
.B(n_1680),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1748),
.B(n_1725),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1754),
.B(n_1722),
.Y(n_1790)
);

AOI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1757),
.A2(n_1755),
.B1(n_1749),
.B2(n_1758),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1758),
.B(n_1715),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1771),
.B(n_1714),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1782),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1746),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1746),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1753),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1744),
.Y(n_1798)
);

BUFx2_ASAP7_75t_L g1799 ( 
.A(n_1752),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1771),
.B(n_1714),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1760),
.B(n_1731),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1772),
.B(n_1775),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1774),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1760),
.A2(n_1739),
.B1(n_1706),
.B2(n_1708),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1772),
.B(n_1706),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1765),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1766),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1753),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1773),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1773),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1743),
.B(n_1725),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1768),
.B(n_1733),
.Y(n_1812)
);

OAI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1777),
.A2(n_1737),
.B1(n_1741),
.B2(n_1732),
.Y(n_1813)
);

O2A1O1Ixp33_ASAP7_75t_L g1814 ( 
.A1(n_1750),
.A2(n_1713),
.B(n_1630),
.C(n_1712),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1768),
.B(n_1735),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1776),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1756),
.B(n_1729),
.Y(n_1817)
);

NOR2xp67_ASAP7_75t_L g1818 ( 
.A(n_1769),
.B(n_1713),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1787),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1818),
.B(n_1799),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1803),
.B(n_1747),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1808),
.B(n_1751),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1786),
.B(n_1745),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1788),
.B(n_1579),
.Y(n_1824)
);

NAND2x1_ASAP7_75t_L g1825 ( 
.A(n_1799),
.B(n_1764),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1794),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1786),
.B(n_1751),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1795),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1802),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1791),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1802),
.B(n_1769),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1801),
.B(n_1767),
.Y(n_1832)
);

NOR2x1_ASAP7_75t_L g1833 ( 
.A(n_1814),
.B(n_1761),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1790),
.B(n_1776),
.Y(n_1834)
);

OAI221xp5_ASAP7_75t_L g1835 ( 
.A1(n_1804),
.A2(n_1752),
.B1(n_1764),
.B2(n_1769),
.C(n_1744),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1810),
.B(n_1759),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1816),
.B(n_1759),
.Y(n_1837)
);

BUFx2_ASAP7_75t_L g1838 ( 
.A(n_1790),
.Y(n_1838)
);

NOR2xp67_ASAP7_75t_SL g1839 ( 
.A(n_1801),
.B(n_1555),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1792),
.B(n_1778),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1789),
.B(n_1780),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1792),
.B(n_1780),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1793),
.B(n_1778),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1838),
.Y(n_1844)
);

O2A1O1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1833),
.A2(n_1813),
.B(n_1798),
.C(n_1784),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1830),
.B(n_1785),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1820),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1829),
.B(n_1800),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1828),
.Y(n_1849)
);

A2O1A1Ixp33_ASAP7_75t_L g1850 ( 
.A1(n_1835),
.A2(n_1769),
.B(n_1817),
.C(n_1784),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1824),
.B(n_1793),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1840),
.B(n_1839),
.Y(n_1852)
);

AOI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1831),
.A2(n_1775),
.B1(n_1800),
.B2(n_1805),
.Y(n_1853)
);

OAI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1841),
.A2(n_1769),
.B1(n_1811),
.B2(n_1805),
.Y(n_1854)
);

OAI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1825),
.A2(n_1823),
.B1(n_1842),
.B2(n_1827),
.Y(n_1855)
);

O2A1O1Ixp33_ASAP7_75t_L g1856 ( 
.A1(n_1821),
.A2(n_1798),
.B(n_1807),
.C(n_1806),
.Y(n_1856)
);

AOI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1821),
.A2(n_1795),
.B(n_1809),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1819),
.Y(n_1858)
);

AOI221x1_ASAP7_75t_L g1859 ( 
.A1(n_1820),
.A2(n_1809),
.B1(n_1797),
.B2(n_1796),
.C(n_1742),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1843),
.B(n_1797),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1831),
.Y(n_1861)
);

OAI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1834),
.A2(n_1796),
.B(n_1812),
.Y(n_1862)
);

AO21x1_ASAP7_75t_L g1863 ( 
.A1(n_1845),
.A2(n_1826),
.B(n_1836),
.Y(n_1863)
);

OAI22xp5_ASAP7_75t_L g1864 ( 
.A1(n_1846),
.A2(n_1832),
.B1(n_1822),
.B2(n_1812),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1844),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1847),
.B(n_1861),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1860),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1848),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1855),
.B(n_1822),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1849),
.Y(n_1870)
);

AOI21xp33_ASAP7_75t_SL g1871 ( 
.A1(n_1845),
.A2(n_1587),
.B(n_1837),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1852),
.Y(n_1872)
);

NAND3xp33_ASAP7_75t_L g1873 ( 
.A(n_1856),
.B(n_1837),
.C(n_1836),
.Y(n_1873)
);

OAI221xp5_ASAP7_75t_SL g1874 ( 
.A1(n_1869),
.A2(n_1850),
.B1(n_1853),
.B2(n_1857),
.C(n_1851),
.Y(n_1874)
);

XOR2xp5_ASAP7_75t_L g1875 ( 
.A(n_1864),
.B(n_1854),
.Y(n_1875)
);

AOI22xp33_ASAP7_75t_L g1876 ( 
.A1(n_1863),
.A2(n_1862),
.B1(n_1857),
.B2(n_1858),
.Y(n_1876)
);

NAND2xp33_ASAP7_75t_SL g1877 ( 
.A(n_1866),
.B(n_1563),
.Y(n_1877)
);

AOI22xp33_ASAP7_75t_SL g1878 ( 
.A1(n_1873),
.A2(n_1859),
.B1(n_1569),
.B2(n_1762),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1872),
.B(n_1815),
.Y(n_1879)
);

NAND4xp75_ASAP7_75t_L g1880 ( 
.A(n_1865),
.B(n_1762),
.C(n_1770),
.D(n_1742),
.Y(n_1880)
);

O2A1O1Ixp33_ASAP7_75t_L g1881 ( 
.A1(n_1871),
.A2(n_1815),
.B(n_1761),
.C(n_1720),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1870),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1868),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1874),
.B(n_1867),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1876),
.B(n_1873),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1879),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1875),
.B(n_1883),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1882),
.Y(n_1888)
);

AOI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1877),
.A2(n_1770),
.B1(n_1783),
.B2(n_1695),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_SL g1890 ( 
.A1(n_1881),
.A2(n_1783),
.B(n_1720),
.Y(n_1890)
);

AOI211xp5_ASAP7_75t_L g1891 ( 
.A1(n_1885),
.A2(n_1884),
.B(n_1887),
.C(n_1886),
.Y(n_1891)
);

NOR2x1_ASAP7_75t_L g1892 ( 
.A(n_1888),
.B(n_1890),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1889),
.B(n_1878),
.Y(n_1893)
);

NAND5xp2_ASAP7_75t_L g1894 ( 
.A(n_1887),
.B(n_1880),
.C(n_1739),
.D(n_1513),
.E(n_1732),
.Y(n_1894)
);

NOR4xp25_ASAP7_75t_L g1895 ( 
.A(n_1885),
.B(n_1712),
.C(n_1720),
.D(n_1709),
.Y(n_1895)
);

NAND4xp25_ASAP7_75t_L g1896 ( 
.A(n_1887),
.B(n_1689),
.C(n_1781),
.D(n_1735),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1892),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1893),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1891),
.Y(n_1899)
);

NAND4xp75_ASAP7_75t_L g1900 ( 
.A(n_1894),
.B(n_1712),
.C(n_1737),
.D(n_1683),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1896),
.A2(n_1494),
.B1(n_1781),
.B2(n_1635),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1897),
.Y(n_1902)
);

HB1xp67_ASAP7_75t_L g1903 ( 
.A(n_1898),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_SL g1904 ( 
.A(n_1899),
.B(n_1501),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1903),
.B(n_1901),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_1905),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1906),
.B(n_1902),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1906),
.Y(n_1908)
);

XOR2xp5_ASAP7_75t_L g1909 ( 
.A(n_1908),
.B(n_1900),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1907),
.Y(n_1910)
);

OAI221xp5_ASAP7_75t_SL g1911 ( 
.A1(n_1909),
.A2(n_1895),
.B1(n_1904),
.B2(n_1625),
.C(n_1655),
.Y(n_1911)
);

CKINVDCx20_ASAP7_75t_R g1912 ( 
.A(n_1910),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1912),
.B(n_1641),
.Y(n_1913)
);

AOI221xp5_ASAP7_75t_L g1914 ( 
.A1(n_1913),
.A2(n_1911),
.B1(n_1628),
.B2(n_1653),
.C(n_1471),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1914),
.Y(n_1915)
);

OAI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1915),
.A2(n_1505),
.B(n_1497),
.Y(n_1916)
);

OAI21x1_ASAP7_75t_SL g1917 ( 
.A1(n_1916),
.A2(n_1683),
.B(n_1653),
.Y(n_1917)
);

AOI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1917),
.A2(n_1520),
.B1(n_1512),
.B2(n_1635),
.Y(n_1918)
);

AOI211xp5_ASAP7_75t_L g1919 ( 
.A1(n_1918),
.A2(n_1512),
.B(n_1520),
.C(n_1505),
.Y(n_1919)
);


endmodule