module real_jpeg_2036_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_286;
wire n_288;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_1),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_53),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_1),
.A2(n_53),
.B1(n_59),
.B2(n_60),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_2),
.Y(n_93)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_3),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_41),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_41),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_4),
.A2(n_41),
.B1(n_59),
.B2(n_60),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_4),
.A2(n_41),
.B1(n_48),
.B2(n_49),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_5),
.A2(n_38),
.B1(n_48),
.B2(n_49),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_5),
.A2(n_38),
.B1(n_59),
.B2(n_60),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_5),
.B(n_29),
.C(n_34),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_5),
.B(n_32),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_5),
.B(n_45),
.C(n_49),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_5),
.B(n_93),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_5),
.B(n_57),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_5),
.B(n_58),
.C(n_60),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_5),
.B(n_51),
.Y(n_233)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_22)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_8),
.A2(n_27),
.B1(n_48),
.B2(n_49),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_8),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_8),
.A2(n_27),
.B1(n_59),
.B2(n_60),
.Y(n_158)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_15),
.B(n_290),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_12),
.B(n_291),
.Y(n_290)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_78),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_76),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_73),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_18),
.B(n_73),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_67),
.C(n_69),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_19),
.B(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.C(n_54),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_20),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_20),
.A2(n_104),
.B1(n_142),
.B2(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_20),
.B(n_142),
.C(n_152),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_20),
.A2(n_104),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_28),
.B1(n_32),
.B2(n_37),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g126 ( 
.A1(n_22),
.A2(n_70),
.B(n_72),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_29),
.B(n_31),
.C(n_32),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_29),
.Y(n_31)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_24),
.B(n_155),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_28),
.B(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

AO22x1_ASAP7_75t_SL g32 ( 
.A1(n_29),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_34),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_34),
.B(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_37),
.B(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_39),
.A2(n_54),
.B1(n_264),
.B2(n_279),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_39),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_42),
.B1(n_51),
.B2(n_52),
.Y(n_39)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_40),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_42),
.A2(n_51),
.B1(n_100),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_43),
.B(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_43),
.B(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_43),
.A2(n_47),
.B(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

AOI22x1_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_47),
.A2(n_266),
.B(n_267),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_49),
.B1(n_58),
.B2(n_63),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_49),
.B(n_226),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AO21x1_ASAP7_75t_L g99 ( 
.A1(n_51),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_54),
.A2(n_264),
.B1(n_265),
.B2(n_268),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_54),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_54),
.B(n_126),
.C(n_265),
.Y(n_280)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_66),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_64),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_64),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_56),
.A2(n_111),
.B(n_112),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_56),
.A2(n_64),
.B1(n_88),
.B2(n_89),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_56),
.A2(n_64),
.B(n_89),
.Y(n_168)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_57),
.A2(n_66),
.B1(n_114),
.B2(n_141),
.Y(n_140)
);

AO22x1_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_57)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_60),
.B(n_219),
.Y(n_218)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_67),
.B(n_69),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B(n_72),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_70),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_70),
.B(n_74),
.Y(n_136)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21x1_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_285),
.B(n_289),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_256),
.B(n_282),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_146),
.B(n_255),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_127),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_82),
.B(n_127),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_105),
.C(n_116),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_83),
.B(n_105),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_97),
.B2(n_98),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_84),
.B(n_99),
.C(n_104),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_86),
.A2(n_87),
.B1(n_90),
.B2(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_86),
.A2(n_87),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_86),
.A2(n_87),
.B1(n_206),
.B2(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_87),
.B(n_201),
.C(n_206),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_87),
.B(n_157),
.C(n_233),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_90),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_92),
.A2(n_93),
.B1(n_121),
.B2(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_95),
.B(n_120),
.Y(n_119)
);

OA21x2_ASAP7_75t_L g177 ( 
.A1(n_95),
.A2(n_120),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_99),
.B(n_125),
.C(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_99),
.A2(n_103),
.B1(n_168),
.B2(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_99),
.A2(n_103),
.B1(n_122),
.B2(n_123),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_99),
.B(n_122),
.C(n_241),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_101),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_115),
.Y(n_105)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_110),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_115),
.B1(n_135),
.B2(n_137),
.Y(n_134)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_108),
.B(n_121),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_115),
.A2(n_131),
.B(n_137),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_116),
.B(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_124),
.C(n_125),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_117),
.A2(n_118),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_119),
.A2(n_122),
.B1(n_123),
.B2(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_119),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_122),
.A2(n_123),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_122),
.B(n_227),
.Y(n_235)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_125),
.A2(n_126),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_125),
.A2(n_126),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_125),
.A2(n_126),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_126),
.B(n_276),
.C(n_280),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_145),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_138),
.B2(n_139),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_130),
.B(n_138),
.C(n_145),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_135),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_142),
.B(n_144),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_142),
.Y(n_144)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_176),
.C(n_177),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_142),
.A2(n_160),
.B1(n_202),
.B2(n_205),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_144),
.A2(n_260),
.B1(n_261),
.B2(n_269),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_144),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_250),
.B(n_254),
.Y(n_146)
);

OAI211xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_179),
.B(n_193),
.C(n_194),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_169),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_169),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_161),
.B2(n_162),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_164),
.C(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_159),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_154),
.B1(n_156),
.B2(n_157),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_156),
.A2(n_157),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_157),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_157),
.B(n_221),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.C(n_175),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_175),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_177),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_176),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND3xp33_ASAP7_75t_SL g194 ( 
.A(n_180),
.B(n_195),
.C(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_182),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_183),
.B(n_185),
.C(n_191),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_190),
.B2(n_191),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI21x1_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_212),
.B(n_249),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_198),
.B(n_200),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_201),
.B(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

NOR2xp67_ASAP7_75t_SL g223 ( 
.A(n_204),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_224),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_207),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_243),
.B(n_248),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_237),
.B(n_242),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_229),
.B(n_236),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_223),
.B(n_228),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_220),
.B(n_222),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_225),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_235),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_235),
.Y(n_236)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_239),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_247),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_252),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_272),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_271),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_271),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_270),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_269),
.C(n_270),
.Y(n_281)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_265),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_281),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_281),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_280),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_288),
.Y(n_289)
);


endmodule