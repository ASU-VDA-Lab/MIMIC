module fake_jpeg_24625_n_328 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_46),
.Y(n_52)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx6p67_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_48),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_49),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_9),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_19),
.B(n_0),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_59),
.Y(n_95)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_62),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_18),
.B1(n_24),
.B2(n_37),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_63),
.A2(n_37),
.B1(n_48),
.B2(n_36),
.Y(n_96)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_64),
.B(n_69),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_18),
.B1(n_29),
.B2(n_21),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_67),
.A2(n_72),
.B1(n_74),
.B2(n_60),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_68),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_29),
.B1(n_30),
.B2(n_21),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_29),
.B1(n_30),
.B2(n_21),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_20),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_77),
.Y(n_120)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_25),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_20),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_82),
.Y(n_116)
);

AO22x1_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_23),
.B1(n_22),
.B2(n_40),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_83),
.A2(n_88),
.B1(n_94),
.B2(n_66),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_48),
.B1(n_43),
.B2(n_30),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_84),
.A2(n_98),
.B1(n_101),
.B2(n_102),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_78),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_87),
.A2(n_89),
.B(n_90),
.C(n_105),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_23),
.B1(n_22),
.B2(n_30),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_40),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_40),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_37),
.B1(n_22),
.B2(n_43),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_96),
.B1(n_97),
.B2(n_115),
.Y(n_130)
);

AO22x2_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_23),
.B1(n_38),
.B2(n_47),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_97),
.B(n_33),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_70),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_99),
.A2(n_118),
.B1(n_35),
.B2(n_33),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_52),
.A2(n_19),
.B1(n_26),
.B2(n_31),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_58),
.A2(n_38),
.B1(n_23),
.B2(n_34),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_23),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_54),
.B(n_17),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_25),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_58),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_32),
.B(n_28),
.C(n_79),
.Y(n_140)
);

AND2x4_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_38),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_94),
.C(n_104),
.Y(n_144)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_75),
.A2(n_26),
.B1(n_28),
.B2(n_27),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_64),
.A2(n_33),
.B(n_25),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_2),
.Y(n_150)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_126),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_75),
.B1(n_71),
.B2(n_80),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_141),
.B1(n_146),
.B2(n_106),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_128),
.B1(n_129),
.B2(n_133),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_71),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_73),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_134),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_83),
.A2(n_96),
.B1(n_90),
.B2(n_119),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_83),
.A2(n_81),
.B1(n_76),
.B2(n_55),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_130),
.A2(n_145),
.B1(n_148),
.B2(n_151),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_132),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_87),
.A2(n_55),
.B1(n_79),
.B2(n_57),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_35),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_136),
.Y(n_182)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_35),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_137),
.B(n_139),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_147),
.B1(n_149),
.B2(n_91),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_87),
.A2(n_25),
.B1(n_33),
.B2(n_17),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_68),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_142),
.B(n_143),
.Y(n_187)
);

AOI32xp33_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_55),
.A3(n_47),
.B1(n_59),
.B2(n_53),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_144),
.A2(n_150),
.B(n_104),
.Y(n_157)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_94),
.A2(n_17),
.B1(n_47),
.B2(n_33),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_89),
.A2(n_33),
.B1(n_2),
.B2(n_5),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_157),
.B(n_6),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_106),
.B(n_91),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_160),
.A2(n_144),
.B(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_161),
.B(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_121),
.A2(n_120),
.B1(n_88),
.B2(n_92),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_168),
.B1(n_113),
.B2(n_136),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_166),
.B(n_170),
.Y(n_213)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_169),
.B(n_177),
.Y(n_200)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_125),
.B(n_120),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_173),
.B(n_176),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_88),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_180),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_142),
.A2(n_116),
.B(n_88),
.C(n_86),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_179),
.B(n_181),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_4),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_183),
.B(n_7),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_128),
.A2(n_113),
.B1(n_117),
.B2(n_108),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_184),
.A2(n_155),
.B1(n_145),
.B2(n_143),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_140),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_186),
.Y(n_207)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_188),
.Y(n_208)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_198),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_191),
.A2(n_195),
.B(n_206),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_150),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_211),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_196),
.B1(n_215),
.B2(n_218),
.Y(n_231)
);

XNOR2x1_ASAP7_75t_SL g195 ( 
.A(n_175),
.B(n_124),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_149),
.B(n_154),
.C(n_117),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_219),
.B1(n_186),
.B2(n_166),
.Y(n_225)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_100),
.Y(n_202)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_107),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_203),
.B(n_205),
.Y(n_235)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_160),
.A2(n_95),
.B(n_5),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_4),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_187),
.Y(n_230)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_217),
.B(n_15),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_16),
.B1(n_7),
.B2(n_8),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_170),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_216),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_164),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_181),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_218)
);

AND2x4_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_200),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_236),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_214),
.A2(n_159),
.B1(n_169),
.B2(n_177),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_224),
.B1(n_237),
.B2(n_242),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_214),
.A2(n_159),
.B1(n_179),
.B2(n_178),
.Y(n_224)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_225),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_201),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_187),
.C(n_156),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_234),
.C(n_206),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_172),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_156),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_212),
.A2(n_178),
.B1(n_172),
.B2(n_176),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_161),
.B1(n_163),
.B2(n_171),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_213),
.A2(n_163),
.B1(n_188),
.B2(n_180),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_194),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_200),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_197),
.A2(n_15),
.B1(n_12),
.B2(n_13),
.Y(n_244)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_228),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_226),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_246),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_247),
.B(n_249),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_233),
.C(n_229),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_205),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_220),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_256),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_230),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_207),
.B1(n_219),
.B2(n_198),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_260),
.B1(n_263),
.B2(n_218),
.Y(n_279)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_220),
.Y(n_259)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_221),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_231),
.A2(n_207),
.B1(n_221),
.B2(n_241),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_208),
.B1(n_244),
.B2(n_242),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_267),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_258),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_236),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_256),
.A2(n_221),
.B1(n_232),
.B2(n_203),
.Y(n_271)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_234),
.C(n_229),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_274),
.C(n_277),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_243),
.C(n_223),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_237),
.B1(n_196),
.B2(n_215),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_275),
.A2(n_276),
.B1(n_279),
.B2(n_253),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_202),
.C(n_190),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_262),
.C(n_190),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_250),
.C(n_254),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_274),
.B1(n_280),
.B2(n_273),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_266),
.B(n_189),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_208),
.Y(n_285)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_291),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_259),
.B(n_252),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_296),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_281),
.B(n_254),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_294),
.C(n_295),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_216),
.C(n_252),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_199),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_277),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_297),
.B(n_298),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_295),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_192),
.B(n_12),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_286),
.A2(n_275),
.B1(n_292),
.B2(n_287),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_192),
.C(n_267),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_296),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_10),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_290),
.C(n_288),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_307),
.A2(n_309),
.B(n_311),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_299),
.A2(n_268),
.B1(n_210),
.B2(n_199),
.Y(n_308)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_308),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_290),
.C(n_272),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_306),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_303),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_301),
.A2(n_14),
.B1(n_305),
.B2(n_303),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_313),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_309),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_319),
.B(n_307),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_321),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_323),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_314),
.C(n_324),
.Y(n_326)
);

A2O1A1Ixp33_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_318),
.B(n_300),
.C(n_315),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_14),
.Y(n_328)
);


endmodule