module fake_ariane_2017_n_110 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_10, n_110);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_110;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_40;
wire n_106;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_109;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_58;
wire n_37;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_108;
wire n_102;
wire n_22;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVxp67_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVxp67_ASAP7_75t_SL g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

AOI21x1_ASAP7_75t_L g37 ( 
.A1(n_20),
.A2(n_0),
.B(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_21),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_39),
.Y(n_51)
);

AND2x4_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_31),
.Y(n_52)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

AND2x6_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_25),
.B(n_23),
.C(n_47),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_33),
.B(n_30),
.C(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_57),
.B(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_42),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_57),
.B2(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_40),
.Y(n_65)
);

AO31x2_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_56),
.A3(n_54),
.B(n_50),
.Y(n_66)
);

BUFx2_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_52),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_58),
.Y(n_69)
);

AO21x2_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_37),
.B(n_53),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_41),
.Y(n_73)
);

OR2x6_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_74),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

OR2x6_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_76),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_82),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_78),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_53),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_45),
.B1(n_46),
.B2(n_76),
.Y(n_89)
);

OAI32xp33_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_45),
.A3(n_85),
.B1(n_87),
.B2(n_86),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_69),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_0),
.B(n_1),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_84),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_4),
.Y(n_97)
);

OAI211xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_76),
.B(n_5),
.C(n_7),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_94),
.B(n_93),
.C(n_96),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_52),
.B(n_53),
.C(n_70),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_100),
.B(n_76),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_72),
.B1(n_24),
.B2(n_68),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_102),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_SL g105 ( 
.A(n_103),
.B(n_101),
.C(n_99),
.Y(n_105)
);

AOI222xp33_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_42),
.B1(n_55),
.B2(n_56),
.C1(n_54),
.C2(n_4),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_104),
.B1(n_70),
.B2(n_42),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_50),
.B1(n_55),
.B2(n_42),
.Y(n_108)
);

AOI222xp33_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_55),
.B1(n_13),
.B2(n_17),
.C1(n_19),
.C2(n_11),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_55),
.B(n_107),
.Y(n_110)
);


endmodule