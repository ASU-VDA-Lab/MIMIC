module fake_jpeg_2677_n_168 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_29),
.B(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_9),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_31),
.B(n_35),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_33),
.Y(n_69)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_39),
.Y(n_66)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_55),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_8),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_51),
.Y(n_63)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_53),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_26),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_54),
.B(n_5),
.Y(n_74)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_7),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_26),
.C(n_23),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_61),
.B(n_86),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_23),
.B1(n_21),
.B2(n_3),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_68),
.B1(n_76),
.B2(n_57),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_32),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_46),
.B1(n_48),
.B2(n_63),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_79),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_7),
.B1(n_8),
.B2(n_38),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_52),
.B(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_83),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_53),
.Y(n_83)
);

HAxp5_ASAP7_75t_SL g86 ( 
.A(n_43),
.B(n_46),
.CON(n_86),
.SN(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_59),
.B(n_63),
.C(n_66),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_58),
.B(n_49),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_103),
.Y(n_109)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_90),
.Y(n_121)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_36),
.B1(n_41),
.B2(n_50),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_100),
.B1(n_85),
.B2(n_103),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_62),
.B1(n_75),
.B2(n_72),
.Y(n_112)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_71),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_99),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_80),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_67),
.A2(n_68),
.B1(n_81),
.B2(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_77),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_73),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_73),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_101),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_120),
.B1(n_102),
.B2(n_85),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_75),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_109),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_117),
.A2(n_91),
.B1(n_89),
.B2(n_105),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_85),
.B1(n_87),
.B2(n_100),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_90),
.B(n_104),
.C(n_88),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_126),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_130),
.B1(n_131),
.B2(n_112),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_116),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_132),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_96),
.B1(n_97),
.B2(n_89),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_109),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_133),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_136),
.Y(n_145)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_113),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_123),
.C(n_121),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_147),
.C(n_148),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_137),
.B(n_132),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_149),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_137),
.B(n_138),
.Y(n_146)
);

XNOR2x1_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_131),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_115),
.C(n_111),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_114),
.C(n_107),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_145),
.A2(n_127),
.B1(n_134),
.B2(n_120),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_150),
.A2(n_140),
.B1(n_128),
.B2(n_116),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_149),
.B(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_158),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_152),
.A2(n_130),
.B1(n_142),
.B2(n_140),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_156),
.A2(n_157),
.B1(n_153),
.B2(n_155),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_159),
.B(n_108),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_154),
.Y(n_161)
);

AOI31xp33_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_154),
.A3(n_160),
.B(n_159),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_163),
.Y(n_164)
);

AOI221xp5_ASAP7_75t_L g165 ( 
.A1(n_163),
.A2(n_161),
.B1(n_160),
.B2(n_110),
.C(n_119),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_164),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);


endmodule