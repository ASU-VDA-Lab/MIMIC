module fake_jpeg_19961_n_316 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_48),
.Y(n_50)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_21),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_37),
.C(n_34),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_9),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_28),
.B1(n_25),
.B2(n_17),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_51),
.A2(n_63),
.B1(n_69),
.B2(n_72),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_36),
.B(n_17),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_53),
.B(n_61),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_55),
.Y(n_98)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_31),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_70),
.Y(n_85)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_24),
.B1(n_35),
.B2(n_19),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_38),
.B(n_31),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_19),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_74),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_22),
.B1(n_35),
.B2(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_43),
.B(n_32),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_24),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_37),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_23),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_91),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_42),
.B1(n_40),
.B2(n_17),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_78),
.A2(n_96),
.B1(n_100),
.B2(n_107),
.Y(n_118)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_80),
.B(n_82),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_63),
.A2(n_23),
.B1(n_29),
.B2(n_28),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_83),
.A2(n_15),
.B(n_8),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_84),
.Y(n_121)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_89),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_75),
.B1(n_74),
.B2(n_61),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_90),
.B1(n_109),
.B2(n_113),
.Y(n_117)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_50),
.A2(n_45),
.B1(n_26),
.B2(n_25),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_21),
.C(n_37),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_69),
.A2(n_28),
.B(n_25),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_93),
.A2(n_104),
.B(n_20),
.Y(n_135)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_102),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_56),
.A2(n_26),
.B1(n_47),
.B2(n_29),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_51),
.A2(n_47),
.B1(n_37),
.B2(n_34),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_70),
.B(n_67),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_101),
.B(n_103),
.Y(n_140)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_SL g104 ( 
.A1(n_73),
.A2(n_18),
.B(n_34),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_114),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_66),
.A2(n_27),
.B1(n_30),
.B2(n_34),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_56),
.A2(n_30),
.B1(n_27),
.B2(n_18),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_67),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_20),
.B1(n_55),
.B2(n_54),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_58),
.A2(n_30),
.B1(n_18),
.B2(n_20),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_62),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_68),
.Y(n_115)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_73),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_119),
.B(n_120),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_30),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_122),
.A2(n_135),
.B(n_106),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_92),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_123),
.A2(n_128),
.B1(n_98),
.B2(n_79),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_81),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_0),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_131),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_93),
.B1(n_91),
.B2(n_99),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_81),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_83),
.B(n_0),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_0),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_144),
.Y(n_153)
);

INVxp33_ASAP7_75t_SL g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_137),
.B(n_123),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_96),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_139),
.A2(n_118),
.B1(n_125),
.B2(n_140),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_1),
.B(n_2),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_4),
.B(n_6),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_76),
.B(n_1),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_84),
.B(n_1),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_146),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_2),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_4),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_106),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_150),
.Y(n_151)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_159),
.A2(n_166),
.B(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_162),
.B(n_177),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_164),
.B1(n_168),
.B2(n_121),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_128),
.A2(n_82),
.B1(n_102),
.B2(n_95),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_138),
.A2(n_108),
.B1(n_94),
.B2(n_86),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_108),
.C(n_7),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_176),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_6),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_135),
.A2(n_8),
.B(n_10),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_137),
.B(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_141),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_175),
.A2(n_179),
.B1(n_182),
.B2(n_139),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_12),
.C(n_13),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_122),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_141),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_116),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_149),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_181),
.A2(n_117),
.B1(n_146),
.B2(n_144),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_149),
.A2(n_124),
.B1(n_147),
.B2(n_122),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_183),
.A2(n_196),
.B(n_177),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_152),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_192),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_197),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_172),
.B(n_120),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_178),
.Y(n_194)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_122),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_158),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_199),
.A2(n_210),
.B1(n_151),
.B2(n_154),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_160),
.Y(n_201)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_155),
.B(n_119),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_202),
.B(n_156),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_209),
.Y(n_227)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_161),
.B(n_166),
.Y(n_215)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_181),
.A2(n_117),
.B1(n_127),
.B2(n_145),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_163),
.A2(n_148),
.B1(n_132),
.B2(n_142),
.Y(n_210)
);

NAND3xp33_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_159),
.C(n_176),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_164),
.B(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_215),
.A2(n_229),
.B1(n_204),
.B2(n_186),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_161),
.C(n_170),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_218),
.C(n_221),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_197),
.C(n_209),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_220),
.A2(n_233),
.B(n_215),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_153),
.Y(n_221)
);

A2O1A1O1Ixp25_ASAP7_75t_L g222 ( 
.A1(n_193),
.A2(n_156),
.B(n_171),
.C(n_157),
.D(n_168),
.Y(n_222)
);

NOR3xp33_ASAP7_75t_SL g251 ( 
.A(n_222),
.B(n_229),
.C(n_235),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_231),
.C(n_187),
.Y(n_248)
);

AOI22x1_ASAP7_75t_SL g229 ( 
.A1(n_193),
.A2(n_171),
.B1(n_157),
.B2(n_151),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_230),
.A2(n_234),
.B1(n_196),
.B2(n_191),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_154),
.C(n_210),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_183),
.A2(n_188),
.B(n_196),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_199),
.A2(n_206),
.B1(n_190),
.B2(n_189),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_198),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_239),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_189),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_252),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_214),
.B(n_208),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_244),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_248),
.Y(n_257)
);

NOR3xp33_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_186),
.C(n_187),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_255),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_234),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_200),
.Y(n_246)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_246),
.Y(n_258)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_200),
.Y(n_249)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_205),
.B1(n_207),
.B2(n_227),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_213),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_252),
.A2(n_227),
.B1(n_231),
.B2(n_220),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_253),
.B1(n_233),
.B2(n_245),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_239),
.Y(n_261)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

INVxp67_ASAP7_75t_SL g265 ( 
.A(n_255),
.Y(n_265)
);

INVx11_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_270),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_218),
.C(n_221),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_238),
.C(n_248),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_240),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_242),
.Y(n_277)
);

O2A1O1Ixp33_ASAP7_75t_SL g290 ( 
.A1(n_277),
.A2(n_269),
.B(n_272),
.C(n_273),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_266),
.B(n_247),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_280),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_271),
.C(n_263),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_257),
.B(n_260),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_284),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_259),
.A2(n_250),
.B1(n_251),
.B2(n_222),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_254),
.B1(n_216),
.B2(n_228),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_286),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_226),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_258),
.B(n_225),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_267),
.Y(n_292)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_290),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_292),
.B(n_293),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_277),
.A2(n_269),
.B(n_256),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_274),
.B(n_273),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_281),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_296),
.B(n_288),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_279),
.C(n_284),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_297),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_294),
.A2(n_262),
.B1(n_286),
.B2(n_275),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_298),
.A2(n_302),
.B1(n_274),
.B2(n_289),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_294),
.A2(n_268),
.B(n_275),
.Y(n_299)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_299),
.Y(n_303)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_290),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_306),
.A2(n_307),
.B1(n_300),
.B2(n_296),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_308),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_305),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_310),
.A2(n_306),
.B(n_303),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_312),
.B(n_309),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_224),
.C(n_297),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_314),
.A2(n_276),
.B1(n_311),
.B2(n_305),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_315),
.Y(n_316)
);


endmodule