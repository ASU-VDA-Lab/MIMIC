module fake_jpeg_12194_n_69 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_69);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_69;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

INVx2_ASAP7_75t_SL g22 ( 
.A(n_21),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_31),
.Y(n_40)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_0),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_26),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_41),
.B(n_6),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_22),
.B1(n_24),
.B2(n_30),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_43),
.B1(n_3),
.B2(n_5),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_27),
.B1(n_28),
.B2(n_13),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_28),
.C(n_27),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_1),
.B(n_2),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_52),
.C(n_53),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_51),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_3),
.B1(n_7),
.B2(n_9),
.Y(n_60)
);

HAxp5_ASAP7_75t_SL g63 ( 
.A(n_60),
.B(n_11),
.CON(n_63),
.SN(n_63)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_56),
.B(n_51),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_63),
.C(n_58),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_65),
.B(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_66),
.B(n_62),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_61),
.B(n_59),
.C(n_57),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_17),
.Y(n_69)
);


endmodule