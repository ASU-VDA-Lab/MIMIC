module fake_jpeg_9528_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_1),
.B(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_19),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_57),
.Y(n_93)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_49),
.B(n_65),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_55),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_24),
.B1(n_31),
.B2(n_16),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_66),
.B1(n_30),
.B2(n_23),
.Y(n_88)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_16),
.B1(n_24),
.B2(n_18),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_42),
.B1(n_39),
.B2(n_36),
.Y(n_85)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_41),
.Y(n_82)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_36),
.A2(n_31),
.B1(n_27),
.B2(n_28),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_42),
.B1(n_41),
.B2(n_40),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_72),
.A2(n_78),
.B1(n_84),
.B2(n_86),
.Y(n_99)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_75),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_42),
.B1(n_41),
.B2(n_40),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_57),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_42),
.B1(n_41),
.B2(n_36),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_18),
.B1(n_43),
.B2(n_26),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_70),
.A2(n_20),
.B1(n_30),
.B2(n_26),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g114 ( 
.A(n_87),
.B(n_15),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_88),
.A2(n_96),
.B1(n_64),
.B2(n_52),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_47),
.A2(n_27),
.B(n_33),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_66),
.Y(n_100)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_94),
.Y(n_124)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_33),
.B1(n_28),
.B2(n_43),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_54),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_100),
.B(n_112),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_101),
.A2(n_119),
.B(n_123),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_63),
.Y(n_103)
);

BUFx24_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_77),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_110),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_109),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_70),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_60),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_117),
.B1(n_83),
.B2(n_95),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_77),
.B1(n_80),
.B2(n_33),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_82),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_43),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_71),
.B(n_79),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_79),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_64),
.B1(n_52),
.B2(n_43),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_86),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_35),
.C(n_60),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_35),
.C(n_62),
.Y(n_146)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

AO22x1_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_43),
.B1(n_35),
.B2(n_62),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_121),
.B1(n_119),
.B2(n_110),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_129),
.B1(n_138),
.B2(n_151),
.Y(n_156)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_133),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_102),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_134),
.B(n_136),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_11),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_75),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_137),
.B(n_140),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_83),
.B1(n_45),
.B2(n_68),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_117),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_76),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_142),
.B(n_147),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_111),
.A2(n_91),
.B1(n_77),
.B2(n_94),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_104),
.B(n_50),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_90),
.B1(n_123),
.B2(n_28),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_106),
.C(n_124),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_80),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_97),
.B(n_35),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_149),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_67),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_67),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_101),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_99),
.A2(n_45),
.B1(n_90),
.B2(n_35),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_119),
.B1(n_100),
.B2(n_99),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_163),
.B1(n_130),
.B2(n_140),
.Y(n_186)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_164),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_167),
.C(n_172),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_129),
.B1(n_135),
.B2(n_138),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_101),
.Y(n_164)
);

AO22x1_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_123),
.B1(n_113),
.B2(n_50),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_174),
.B(n_141),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_118),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_127),
.Y(n_169)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

NAND2xp33_ASAP7_75t_SL g194 ( 
.A(n_170),
.B(n_143),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_171),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_104),
.C(n_118),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_177),
.B(n_179),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_0),
.Y(n_174)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_127),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_176),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_128),
.A2(n_0),
.B(n_1),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_104),
.Y(n_178)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_125),
.A2(n_17),
.B1(n_25),
.B2(n_13),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_148),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_184),
.C(n_206),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_183),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_150),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_186),
.A2(n_201),
.B(n_202),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_191),
.B(n_192),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_195),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_194),
.A2(n_173),
.B1(n_170),
.B2(n_163),
.Y(n_213)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_156),
.A2(n_130),
.B1(n_129),
.B2(n_147),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_179),
.B1(n_151),
.B2(n_161),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_142),
.B(n_141),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_152),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_160),
.A2(n_139),
.B(n_136),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_205),
.A2(n_152),
.B(n_160),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_167),
.B(n_146),
.C(n_151),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_210),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_229),
.B(n_231),
.Y(n_248)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_200),
.Y(n_210)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_157),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_204),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_182),
.Y(n_233)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_218),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_184),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_222),
.C(n_212),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_155),
.Y(n_217)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_217),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_198),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_156),
.B1(n_153),
.B2(n_165),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_219),
.A2(n_227),
.B1(n_185),
.B2(n_165),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_155),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_220),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_174),
.B(n_176),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_197),
.B(n_190),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_164),
.C(n_153),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_228),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_144),
.B1(n_165),
.B2(n_169),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_189),
.B(n_177),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_230),
.Y(n_240)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_233),
.B(n_224),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_206),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_239),
.C(n_242),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_182),
.Y(n_235)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_236),
.A2(n_223),
.B(n_221),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_185),
.B1(n_190),
.B2(n_188),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_238),
.A2(n_223),
.B1(n_210),
.B2(n_208),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_205),
.Y(n_239)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_174),
.C(n_133),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_246),
.C(n_247),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_174),
.C(n_131),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_159),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_231),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_228),
.C(n_209),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_175),
.Y(n_253)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_253),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_255),
.B(n_270),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_264),
.C(n_268),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_259),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_215),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_260),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_217),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_234),
.Y(n_264)
);

BUFx4f_ASAP7_75t_SL g265 ( 
.A(n_236),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_265),
.A2(n_251),
.B1(n_235),
.B2(n_248),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_271),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_244),
.A2(n_213),
.B1(n_219),
.B2(n_227),
.Y(n_268)
);

NAND4xp25_ASAP7_75t_SL g269 ( 
.A(n_238),
.B(n_183),
.C(n_131),
.D(n_107),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_269),
.B(n_237),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_220),
.C(n_230),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_243),
.C(n_246),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_242),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_276),
.C(n_279),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_275),
.A2(n_277),
.B1(n_0),
.B2(n_1),
.Y(n_297)
);

A2O1A1Ixp33_ASAP7_75t_SL g277 ( 
.A1(n_265),
.A2(n_241),
.B(n_211),
.C(n_245),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_283),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_239),
.C(n_233),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_13),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_286),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_11),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_281),
.A2(n_265),
.B(n_262),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_287),
.A2(n_293),
.B(n_2),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_282),
.B(n_266),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_291),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_270),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_263),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_295),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_284),
.A2(n_258),
.B(n_257),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_257),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_256),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_296),
.B(n_298),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_299),
.B(n_0),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_11),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_280),
.C(n_277),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_306),
.B(n_3),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_277),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_303),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_280),
.A3(n_17),
.B1(n_25),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_305),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_297),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_2),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_307),
.B(n_3),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_308),
.A2(n_2),
.B(n_3),
.Y(n_310)
);

OAI321xp33_ASAP7_75t_L g318 ( 
.A1(n_310),
.A2(n_311),
.A3(n_4),
.B1(n_5),
.B2(n_7),
.C(n_8),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_3),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_315),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_4),
.B(n_7),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_305),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_8),
.C(n_9),
.Y(n_322)
);

A2O1A1O1Ixp25_ASAP7_75t_L g324 ( 
.A1(n_318),
.A2(n_322),
.B(n_8),
.C(n_9),
.D(n_313),
.Y(n_324)
);

NAND4xp25_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_302),
.C(n_7),
.D(n_8),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_321),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_9),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_320),
.B(n_316),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_323),
.Y(n_327)
);


endmodule