module fake_jpeg_13814_n_185 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_185);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_51),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx6p67_ASAP7_75t_R g79 ( 
.A(n_41),
.Y(n_79)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_47),
.Y(n_83)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx4f_ASAP7_75t_SL g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_57),
.Y(n_62)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_52),
.B(n_54),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_0),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_56),
.Y(n_58)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_54),
.A2(n_22),
.B1(n_27),
.B2(n_18),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_74),
.B1(n_70),
.B2(n_84),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_16),
.B1(n_28),
.B2(n_19),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_63),
.A2(n_72),
.B(n_75),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_16),
.B1(n_28),
.B2(n_19),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_65),
.A2(n_80),
.B1(n_63),
.B2(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_30),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_86),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_24),
.B1(n_14),
.B2(n_23),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_30),
.B1(n_29),
.B2(n_4),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_32),
.A2(n_29),
.B1(n_3),
.B2(n_4),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_34),
.B(n_1),
.C(n_3),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_70),
.B(n_62),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_38),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_5),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_35),
.B(n_36),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_89),
.B(n_41),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_94),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_6),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_95),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_41),
.B1(n_7),
.B2(n_53),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_58),
.A2(n_63),
.B1(n_72),
.B2(n_59),
.Y(n_97)
);

OAI22x1_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_99),
.B1(n_101),
.B2(n_111),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_102),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_100),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_71),
.B1(n_66),
.B2(n_88),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_SL g102 ( 
.A(n_61),
.B(n_81),
.C(n_73),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_84),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_107),
.B(n_108),
.C(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_105),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_79),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_113),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_83),
.B(n_90),
.C(n_77),
.Y(n_107)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_64),
.A2(n_68),
.B1(n_77),
.B2(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_99),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_123),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g146 ( 
.A(n_116),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_93),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_118),
.Y(n_143)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

OR2x4_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_102),
.Y(n_132)
);

A2O1A1O1Ixp25_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_107),
.B(n_95),
.C(n_113),
.D(n_112),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_96),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_96),
.C(n_105),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_141),
.C(n_117),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_126),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_137),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_124),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_128),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_125),
.A2(n_104),
.B1(n_109),
.B2(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_145),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_117),
.C(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_143),
.B(n_132),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_147),
.Y(n_155)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_131),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_134),
.C(n_136),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_147),
.B(n_131),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_129),
.B1(n_130),
.B2(n_122),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_156),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_157),
.A2(n_136),
.B(n_138),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_141),
.C(n_146),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_160),
.C(n_163),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_157),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_140),
.C(n_145),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_144),
.C(n_121),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_153),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_171),
.Y(n_175)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_161),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_170),
.Y(n_173)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_158),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_166),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_155),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_176),
.B(n_177),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_174),
.A2(n_153),
.B1(n_154),
.B2(n_168),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_178),
.A2(n_172),
.B1(n_175),
.B2(n_150),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_180),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_178),
.B1(n_175),
.B2(n_142),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_181),
.A2(n_179),
.B(n_121),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_182),
.B(n_120),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_128),
.Y(n_185)
);


endmodule