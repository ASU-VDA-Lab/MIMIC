module real_aes_5118_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_599;
wire n_887;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_592;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_400;
wire n_1160;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_417;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_552;
wire n_590;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1250;
wire n_1095;
wire n_859;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1161;
wire n_686;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_837;
wire n_829;
wire n_1030;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1129;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_807;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1163;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1162;
wire n_762;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_459;
wire n_1172;
wire n_998;
wire n_836;
wire n_1184;
wire n_583;
wire n_414;
wire n_776;
wire n_1138;
wire n_890;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_1102;
wire n_661;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_577;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_937;
wire n_773;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_816;
wire n_625;
wire n_953;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_609;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1050;
wire n_426;
wire n_1134;
wire n_616;
wire n_880;
wire n_1103;
wire n_832;
wire n_1060;
wire n_1154;
wire n_632;
wire n_714;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1033;
wire n_1028;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1240;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_974;
wire n_857;
wire n_376;
wire n_491;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_408;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1198;
wire n_993;
wire n_819;
wire n_737;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_449;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_986;
wire n_451;
wire n_1037;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1057;
wire n_907;
wire n_1005;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_698;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_483;
wire n_394;
wire n_729;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_603;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g1257 ( .A1(n_0), .A2(n_265), .B1(n_831), .B2(n_835), .Y(n_1257) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_1), .A2(n_360), .B1(n_622), .B2(n_623), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_2), .A2(n_82), .B1(n_591), .B2(n_592), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g1256 ( .A1(n_3), .A2(n_199), .B1(n_619), .B2(n_620), .Y(n_1256) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_4), .A2(n_206), .B1(n_674), .B2(n_757), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_5), .A2(n_153), .B1(n_622), .B2(n_623), .Y(n_773) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_6), .A2(n_261), .B1(n_435), .B2(n_507), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_7), .A2(n_166), .B1(n_508), .B2(n_588), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_8), .A2(n_325), .B1(n_619), .B2(n_620), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_9), .A2(n_170), .B1(n_412), .B2(n_510), .Y(n_724) );
INVx1_ASAP7_75t_L g632 ( .A(n_10), .Y(n_632) );
INVx1_ASAP7_75t_SL g973 ( .A(n_11), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_12), .A2(n_340), .B1(n_550), .B2(n_588), .Y(n_781) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_13), .A2(n_309), .B1(n_535), .B2(n_567), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_14), .A2(n_29), .B1(n_419), .B2(n_424), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_15), .A2(n_109), .B1(n_439), .B2(n_757), .Y(n_888) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_16), .B(n_394), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_17), .A2(n_203), .B1(n_535), .B2(n_597), .Y(n_891) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_18), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_19), .A2(n_250), .B1(n_622), .B2(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_20), .B(n_474), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g907 ( .A1(n_21), .A2(n_213), .B1(n_775), .B2(n_776), .Y(n_907) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_22), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g987 ( .A1(n_23), .A2(n_100), .B1(n_988), .B2(n_990), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_24), .A2(n_343), .B1(n_562), .B2(n_743), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_25), .A2(n_73), .B1(n_468), .B2(n_471), .Y(n_467) );
INVx1_ASAP7_75t_L g1223 ( .A(n_26), .Y(n_1223) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_27), .A2(n_151), .B1(n_446), .B2(n_503), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_28), .A2(n_599), .B(n_602), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_30), .A2(n_144), .B1(n_584), .B2(n_585), .Y(n_583) );
INVx1_ASAP7_75t_L g384 ( .A(n_31), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_32), .A2(n_216), .B1(n_634), .B2(n_640), .Y(n_864) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_33), .A2(n_519), .B(n_522), .Y(n_518) );
INVx1_ASAP7_75t_L g523 ( .A(n_34), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_35), .A2(n_240), .B1(n_978), .B2(n_980), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_36), .A2(n_101), .B1(n_776), .B2(n_835), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_37), .A2(n_121), .B1(n_443), .B2(n_546), .Y(n_1217) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_38), .A2(n_372), .B1(n_775), .B2(n_776), .Y(n_774) );
XOR2x2_ASAP7_75t_L g898 ( .A(n_39), .B(n_899), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g1228 ( .A1(n_40), .A2(n_54), .B1(n_595), .B2(n_812), .Y(n_1228) );
AOI22xp33_ASAP7_75t_SL g1253 ( .A1(n_41), .A2(n_363), .B1(n_562), .B2(n_634), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_42), .A2(n_50), .B1(n_424), .B2(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_43), .A2(n_149), .B1(n_552), .B2(n_588), .Y(n_695) );
INVx1_ASAP7_75t_L g1001 ( .A(n_44), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_45), .A2(n_108), .B1(n_535), .B2(n_597), .Y(n_813) );
INVx1_ASAP7_75t_L g559 ( .A(n_46), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_47), .A2(n_160), .B1(n_670), .B2(n_745), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_48), .A2(n_135), .B1(n_535), .B2(n_597), .Y(n_846) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_49), .A2(n_94), .B1(n_443), .B2(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_51), .A2(n_141), .B1(n_591), .B2(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_52), .A2(n_167), .B1(n_516), .B2(n_676), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_53), .A2(n_181), .B1(n_513), .B2(n_554), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_55), .A2(n_105), .B1(n_622), .B2(n_623), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_56), .A2(n_237), .B1(n_619), .B2(n_620), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_57), .A2(n_259), .B1(n_557), .B2(n_719), .Y(n_867) );
OA22x2_ASAP7_75t_L g400 ( .A1(n_58), .A2(n_165), .B1(n_394), .B2(n_398), .Y(n_400) );
INVx1_ASAP7_75t_L g431 ( .A(n_58), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_59), .A2(n_316), .B1(n_503), .B2(n_546), .Y(n_545) );
XNOR2x1_ASAP7_75t_L g578 ( .A(n_60), .B(n_579), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_61), .A2(n_64), .B1(n_622), .B2(n_623), .Y(n_910) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_62), .A2(n_303), .B1(n_674), .B2(n_757), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_63), .A2(n_359), .B1(n_595), .B2(n_692), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_65), .A2(n_263), .B1(n_516), .B2(n_552), .Y(n_739) );
XNOR2x2_ASAP7_75t_L g653 ( .A(n_66), .B(n_654), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_67), .A2(n_256), .B1(n_631), .B2(n_770), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_68), .A2(n_308), .B1(n_622), .B2(n_623), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_69), .A2(n_266), .B1(n_548), .B2(n_550), .Y(n_738) );
INVx1_ASAP7_75t_L g685 ( .A(n_70), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_71), .A2(n_104), .B1(n_548), .B2(n_674), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_72), .A2(n_268), .B1(n_775), .B2(n_776), .Y(n_948) );
AOI221xp5_ASAP7_75t_L g900 ( .A1(n_74), .A2(n_190), .B1(n_475), .B2(n_639), .C(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g397 ( .A(n_75), .Y(n_397) );
OAI21xp33_ASAP7_75t_L g432 ( .A1(n_75), .A2(n_165), .B(n_433), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_75), .B(n_184), .Y(n_464) );
AOI21xp33_ASAP7_75t_L g451 ( .A1(n_76), .A2(n_452), .B(n_455), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g667 ( .A1(n_77), .A2(n_152), .B1(n_668), .B2(n_670), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g894 ( .A1(n_78), .A2(n_319), .B1(n_452), .B2(n_750), .C(n_895), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g1258 ( .A1(n_79), .A2(n_355), .B1(n_622), .B2(n_623), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_80), .A2(n_305), .B1(n_631), .B2(n_634), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_81), .A2(n_279), .B1(n_435), .B2(n_438), .Y(n_434) );
INVx1_ASAP7_75t_L g946 ( .A(n_83), .Y(n_946) );
AOI22xp5_ASAP7_75t_L g852 ( .A1(n_84), .A2(n_188), .B1(n_443), .B2(n_853), .Y(n_852) );
AOI22xp33_ASAP7_75t_SL g442 ( .A1(n_85), .A2(n_220), .B1(n_443), .B2(n_446), .Y(n_442) );
INVx1_ASAP7_75t_L g748 ( .A(n_86), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g1216 ( .A1(n_87), .A2(n_91), .B1(n_508), .B2(n_588), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_88), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_89), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g972 ( .A(n_90), .Y(n_972) );
AND2x4_ASAP7_75t_L g979 ( .A(n_90), .B(n_277), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_92), .A2(n_321), .B1(n_775), .B2(n_776), .Y(n_1255) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_93), .A2(n_243), .B1(n_446), .B2(n_508), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_95), .A2(n_212), .B1(n_529), .B2(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g792 ( .A(n_96), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_97), .A2(n_225), .B1(n_588), .B2(n_589), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_98), .A2(n_99), .B1(n_388), .B2(n_412), .Y(n_387) );
XNOR2x2_ASAP7_75t_L g1213 ( .A(n_100), .B(n_1214), .Y(n_1213) );
AOI22xp33_ASAP7_75t_L g1235 ( .A1(n_100), .A2(n_1236), .B1(n_1260), .B2(n_1262), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_102), .A2(n_201), .B1(n_521), .B2(n_770), .Y(n_769) );
AOI221xp5_ASAP7_75t_L g789 ( .A1(n_103), .A2(n_107), .B1(n_700), .B2(n_764), .C(n_790), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_106), .A2(n_557), .B(n_558), .Y(n_556) );
XNOR2x1_ASAP7_75t_L g680 ( .A(n_110), .B(n_681), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g763 ( .A1(n_111), .A2(n_764), .B(n_766), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_112), .A2(n_326), .B1(n_557), .B2(n_619), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_113), .B(n_845), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_114), .A2(n_208), .B1(n_535), .B2(n_597), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_115), .A2(n_155), .B1(n_591), .B2(n_809), .Y(n_808) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_116), .A2(n_147), .B1(n_502), .B2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_117), .A2(n_183), .B1(n_634), .B2(n_770), .Y(n_943) );
INVx1_ASAP7_75t_L g791 ( .A(n_118), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_119), .A2(n_140), .B1(n_503), .B2(n_546), .Y(n_735) );
INVx1_ASAP7_75t_L g970 ( .A(n_120), .Y(n_970) );
AND2x4_ASAP7_75t_L g975 ( .A(n_120), .B(n_958), .Y(n_975) );
INVx1_ASAP7_75t_SL g989 ( .A(n_120), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_122), .A2(n_264), .B1(n_521), .B2(n_535), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_123), .A2(n_297), .B1(n_502), .B2(n_504), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_124), .A2(n_196), .B1(n_664), .B2(n_665), .Y(n_663) );
XNOR2x2_ASAP7_75t_SL g610 ( .A(n_125), .B(n_611), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_126), .A2(n_286), .B1(n_438), .B2(n_504), .Y(n_721) );
INVx1_ASAP7_75t_L g926 ( .A(n_127), .Y(n_926) );
CKINVDCx16_ASAP7_75t_R g1042 ( .A(n_128), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_129), .A2(n_154), .B1(n_968), .B2(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g818 ( .A(n_130), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_131), .B(n_750), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_132), .A2(n_270), .B1(n_552), .B2(n_591), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_133), .A2(n_346), .B1(n_510), .B2(n_513), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_134), .A2(n_357), .B1(n_557), .B2(n_631), .Y(n_942) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_136), .A2(n_366), .B1(n_637), .B2(n_639), .C(n_641), .Y(n_636) );
INVx1_ASAP7_75t_L g998 ( .A(n_137), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_138), .A2(n_150), .B1(n_588), .B2(n_674), .Y(n_673) );
XNOR2x1_ASAP7_75t_L g753 ( .A(n_139), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g761 ( .A(n_142), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_143), .A2(n_180), .B1(n_831), .B2(n_835), .Y(n_924) );
AOI22xp5_ASAP7_75t_L g920 ( .A1(n_145), .A2(n_365), .B1(n_622), .B2(n_623), .Y(n_920) );
AOI21xp5_ASAP7_75t_L g847 ( .A1(n_146), .A2(n_452), .B(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g626 ( .A(n_148), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_156), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g896 ( .A(n_157), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_158), .A2(n_234), .B1(n_843), .B2(n_893), .Y(n_892) );
AOI22xp5_ASAP7_75t_L g1237 ( .A1(n_159), .A2(n_1238), .B1(n_1239), .B2(n_1259), .Y(n_1237) );
CKINVDCx20_ASAP7_75t_R g1259 ( .A(n_159), .Y(n_1259) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_161), .A2(n_307), .B1(n_584), .B2(n_585), .Y(n_804) );
CKINVDCx6p67_ASAP7_75t_R g1041 ( .A(n_162), .Y(n_1041) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_163), .A2(n_350), .B1(n_775), .B2(n_776), .Y(n_921) );
INVx1_ASAP7_75t_L g411 ( .A(n_164), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_164), .B(n_429), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_164), .B(n_224), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_165), .B(n_289), .Y(n_463) );
INVx1_ASAP7_75t_L g456 ( .A(n_168), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_169), .A2(n_282), .B1(n_566), .B2(n_567), .Y(n_565) );
AOI21xp33_ASAP7_75t_L g1221 ( .A1(n_171), .A2(n_562), .B(n_1222), .Y(n_1221) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_172), .A2(n_185), .B1(n_700), .B2(n_701), .C(n_702), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_173), .A2(n_315), .B1(n_554), .B2(n_585), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_174), .A2(n_245), .B1(n_554), .B2(n_585), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_175), .A2(n_177), .B1(n_567), .B2(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g849 ( .A(n_176), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g1008 ( .A1(n_178), .A2(n_335), .B1(n_992), .B2(n_993), .Y(n_1008) );
AOI21xp5_ASAP7_75t_L g1246 ( .A1(n_179), .A2(n_532), .B(n_1247), .Y(n_1246) );
AOI22xp5_ASAP7_75t_L g1225 ( .A1(n_182), .A2(n_217), .B1(n_554), .B2(n_585), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_184), .B(n_404), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_186), .A2(n_218), .B1(n_516), .B2(n_552), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_187), .A2(n_262), .B1(n_831), .B2(n_835), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_189), .A2(n_373), .B1(n_554), .B2(n_585), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_191), .A2(n_374), .B1(n_388), .B2(n_585), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_192), .A2(n_232), .B1(n_446), .B2(n_676), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g991 ( .A1(n_193), .A2(n_293), .B1(n_992), .B2(n_993), .Y(n_991) );
INVx1_ASAP7_75t_L g767 ( .A(n_194), .Y(n_767) );
INVx1_ASAP7_75t_L g1219 ( .A(n_195), .Y(n_1219) );
INVx1_ASAP7_75t_L g603 ( .A(n_197), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_198), .A2(n_306), .B1(n_591), .B2(n_678), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_200), .B(n_605), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_202), .B(n_607), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_204), .A2(n_352), .B1(n_567), .B2(n_843), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_205), .A2(n_211), .B1(n_615), .B2(n_853), .Y(n_886) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_207), .A2(n_801), .B1(n_802), .B2(n_819), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_207), .Y(n_801) );
AOI21xp33_ASAP7_75t_L g746 ( .A1(n_209), .A2(n_521), .B(n_747), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_210), .A2(n_312), .B1(n_968), .B2(n_1015), .Y(n_1014) );
XNOR2x1_ASAP7_75t_L g542 ( .A(n_214), .B(n_543), .Y(n_542) );
BUFx2_ASAP7_75t_L g1249 ( .A(n_215), .Y(n_1249) );
AOI22xp5_ASAP7_75t_L g1007 ( .A1(n_219), .A2(n_349), .B1(n_988), .B2(n_990), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_221), .A2(n_287), .B1(n_980), .B2(n_1012), .Y(n_1019) );
INVx1_ASAP7_75t_L g703 ( .A(n_222), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_223), .A2(n_348), .B1(n_516), .B2(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g395 ( .A(n_224), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_226), .A2(n_339), .B1(n_513), .B2(n_737), .Y(n_736) );
XNOR2x1_ASAP7_75t_L g820 ( .A(n_227), .B(n_821), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_227), .A2(n_239), .B1(n_1012), .B2(n_1013), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_228), .A2(n_345), .B1(n_479), .B2(n_488), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_229), .A2(n_344), .B1(n_567), .B2(n_595), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_230), .A2(n_320), .B1(n_591), .B2(n_592), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g1226 ( .A1(n_231), .A2(n_332), .B1(n_591), .B2(n_678), .Y(n_1226) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_233), .A2(n_284), .B1(n_528), .B2(n_529), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g918 ( .A1(n_235), .A2(n_244), .B1(n_529), .B2(n_670), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_236), .B(n_532), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_238), .A2(n_330), .B1(n_548), .B2(n_550), .Y(n_547) );
OR2x2_ASAP7_75t_L g740 ( .A(n_241), .B(n_741), .Y(n_740) );
INVxp67_ASAP7_75t_L g752 ( .A(n_241), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_242), .A2(n_301), .B1(n_435), .B2(n_678), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g1229 ( .A1(n_246), .A2(n_358), .B1(n_670), .B2(n_743), .Y(n_1229) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_247), .A2(n_267), .B1(n_831), .B2(n_835), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_248), .A2(n_318), .B1(n_443), .B2(n_616), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_249), .A2(n_300), .B1(n_619), .B2(n_620), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_251), .A2(n_273), .B1(n_968), .B2(n_1015), .Y(n_1026) );
NAND2xp5_ASAP7_75t_SL g865 ( .A(n_252), .B(n_866), .Y(n_865) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_253), .A2(n_254), .B1(n_554), .B2(n_885), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_255), .A2(n_322), .B1(n_452), .B2(n_714), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_257), .A2(n_295), .B1(n_631), .B2(n_770), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_258), .A2(n_296), .B1(n_516), .B2(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_260), .A2(n_356), .B1(n_615), .B2(n_616), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_269), .A2(n_281), .B1(n_631), .B2(n_770), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_271), .A2(n_369), .B1(n_711), .B2(n_712), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_272), .A2(n_310), .B1(n_620), .B2(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g635 ( .A(n_274), .Y(n_635) );
AOI22x1_ASAP7_75t_L g880 ( .A1(n_275), .A2(n_881), .B1(n_882), .B2(n_897), .Y(n_880) );
INVx1_ASAP7_75t_L g897 ( .A(n_275), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_276), .A2(n_294), .B1(n_978), .B2(n_1013), .Y(n_1025) );
HB1xp67_ASAP7_75t_L g960 ( .A(n_277), .Y(n_960) );
AND2x4_ASAP7_75t_L g971 ( .A(n_277), .B(n_972), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_278), .B(n_701), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_280), .A2(n_314), .B1(n_831), .B2(n_835), .Y(n_951) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_283), .A2(n_370), .B1(n_468), .B2(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g687 ( .A(n_285), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_288), .A2(n_333), .B1(n_557), .B2(n_634), .Y(n_908) );
INVx1_ASAP7_75t_L g409 ( .A(n_289), .Y(n_409) );
INVxp67_ASAP7_75t_L g487 ( .A(n_289), .Y(n_487) );
AOI21xp33_ASAP7_75t_SL g1243 ( .A1(n_290), .A2(n_521), .B(n_1244), .Y(n_1243) );
INVx1_ASAP7_75t_L g902 ( .A(n_291), .Y(n_902) );
INVx1_ASAP7_75t_L g930 ( .A(n_292), .Y(n_930) );
INVx1_ASAP7_75t_L g860 ( .A(n_294), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_298), .A2(n_317), .B1(n_619), .B2(n_620), .Y(n_949) );
INVxp67_ASAP7_75t_R g1045 ( .A(n_299), .Y(n_1045) );
INVx2_ASAP7_75t_L g958 ( .A(n_302), .Y(n_958) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_304), .A2(n_657), .B(n_658), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_311), .A2(n_313), .B1(n_634), .B2(n_775), .Y(n_824) );
INVx1_ASAP7_75t_L g642 ( .A(n_323), .Y(n_642) );
INVx1_ASAP7_75t_L g1245 ( .A(n_324), .Y(n_1245) );
AOI21xp33_ASAP7_75t_L g826 ( .A1(n_327), .A2(n_640), .B(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g828 ( .A(n_328), .Y(n_828) );
INVx1_ASAP7_75t_L g689 ( .A(n_329), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_331), .B(n_716), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_334), .A2(n_347), .B1(n_535), .B2(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g839 ( .A(n_335), .Y(n_839) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_336), .A2(n_499), .B(n_536), .Y(n_498) );
INVx1_ASAP7_75t_L g538 ( .A(n_336), .Y(n_538) );
INVx1_ASAP7_75t_L g999 ( .A(n_337), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_338), .B(n_661), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_341), .A2(n_368), .B1(n_775), .B2(n_776), .Y(n_869) );
INVx1_ASAP7_75t_L g938 ( .A(n_342), .Y(n_938) );
INVx1_ASAP7_75t_L g931 ( .A(n_351), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_353), .B(n_866), .Y(n_941) );
BUFx2_ASAP7_75t_L g1251 ( .A(n_354), .Y(n_1251) );
AOI21xp5_ASAP7_75t_L g928 ( .A1(n_361), .A2(n_638), .B(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g976 ( .A(n_362), .Y(n_976) );
INVx1_ASAP7_75t_L g659 ( .A(n_364), .Y(n_659) );
AOI21xp33_ASAP7_75t_L g944 ( .A1(n_367), .A2(n_640), .B(n_945), .Y(n_944) );
AOI21xp33_ASAP7_75t_SL g816 ( .A1(n_371), .A2(n_668), .B(n_817), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_954), .B(n_961), .Y(n_375) );
XNOR2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_648), .Y(n_376) );
OAI21xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_573), .B(n_645), .Y(n_377) );
OAI21xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_492), .B(n_569), .Y(n_378) );
AND2x2_ASAP7_75t_L g570 ( .A(n_379), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_380), .A2(n_493), .B(n_570), .C(n_646), .Y(n_645) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
XNOR2x1_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
NOR2x1_ASAP7_75t_L g385 ( .A(n_386), .B(n_448), .Y(n_385) );
NAND4xp25_ASAP7_75t_L g386 ( .A(n_387), .B(n_418), .C(n_434), .D(n_442), .Y(n_386) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx3_ASAP7_75t_L g512 ( .A(n_389), .Y(n_512) );
BUFx12f_ASAP7_75t_L g554 ( .A(n_389), .Y(n_554) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_401), .Y(n_389) );
AND2x2_ASAP7_75t_L g415 ( .A(n_390), .B(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_L g420 ( .A(n_390), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g444 ( .A(n_390), .B(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g622 ( .A(n_390), .B(n_401), .Y(n_622) );
AND2x4_ASAP7_75t_L g623 ( .A(n_390), .B(n_416), .Y(n_623) );
AND2x4_ASAP7_75t_L g775 ( .A(n_390), .B(n_440), .Y(n_775) );
AND2x4_ASAP7_75t_L g831 ( .A(n_390), .B(n_421), .Y(n_831) );
AND2x4_ASAP7_75t_L g390 ( .A(n_391), .B(n_399), .Y(n_390) );
AND2x2_ASAP7_75t_L g454 ( .A(n_391), .B(n_400), .Y(n_454) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g437 ( .A(n_392), .B(n_400), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_396), .Y(n_392) );
NAND2xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx2_ASAP7_75t_L g398 ( .A(n_394), .Y(n_398) );
INVx3_ASAP7_75t_L g404 ( .A(n_394), .Y(n_404) );
NAND2xp33_ASAP7_75t_L g410 ( .A(n_394), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g433 ( .A(n_394), .Y(n_433) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_394), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_395), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_397), .A2(n_433), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g485 ( .A(n_400), .B(n_486), .Y(n_485) );
AND2x4_ASAP7_75t_L g453 ( .A(n_401), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g491 ( .A(n_401), .B(n_437), .Y(n_491) );
AND2x4_ASAP7_75t_L g557 ( .A(n_401), .B(n_454), .Y(n_557) );
AND2x4_ASAP7_75t_L g631 ( .A(n_401), .B(n_437), .Y(n_631) );
AND2x4_ASAP7_75t_L g401 ( .A(n_402), .B(n_406), .Y(n_401) );
INVx2_ASAP7_75t_L g417 ( .A(n_402), .Y(n_417) );
AND2x4_ASAP7_75t_L g421 ( .A(n_402), .B(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g441 ( .A(n_402), .B(n_423), .Y(n_441) );
AND2x2_ASAP7_75t_L g482 ( .A(n_402), .B(n_483), .Y(n_482) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_405), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_404), .B(n_409), .Y(n_408) );
INVxp67_ASAP7_75t_L g429 ( .A(n_404), .Y(n_429) );
NAND3xp33_ASAP7_75t_L g465 ( .A(n_405), .B(n_428), .C(n_466), .Y(n_465) );
AND2x4_ASAP7_75t_L g416 ( .A(n_406), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g423 ( .A(n_407), .Y(n_423) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx3_ASAP7_75t_L g513 ( .A(n_415), .Y(n_513) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_415), .Y(n_585) );
BUFx5_ASAP7_75t_L g885 ( .A(n_415), .Y(n_885) );
AND2x4_ASAP7_75t_L g470 ( .A(n_416), .B(n_454), .Y(n_470) );
AND2x4_ASAP7_75t_L g472 ( .A(n_416), .B(n_427), .Y(n_472) );
AND2x2_ASAP7_75t_L g477 ( .A(n_416), .B(n_437), .Y(n_477) );
AND2x4_ASAP7_75t_L g634 ( .A(n_416), .B(n_427), .Y(n_634) );
AND2x2_ASAP7_75t_L g638 ( .A(n_416), .B(n_437), .Y(n_638) );
AND2x2_ASAP7_75t_L g640 ( .A(n_416), .B(n_454), .Y(n_640) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx12f_ASAP7_75t_L g516 ( .A(n_420), .Y(n_516) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_420), .Y(n_591) );
AND2x4_ASAP7_75t_L g426 ( .A(n_421), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g436 ( .A(n_421), .B(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g549 ( .A(n_421), .B(n_437), .Y(n_549) );
AND2x4_ASAP7_75t_L g619 ( .A(n_421), .B(n_437), .Y(n_619) );
AND2x4_ASAP7_75t_L g835 ( .A(n_421), .B(n_427), .Y(n_835) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx4_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g552 ( .A(n_425), .Y(n_552) );
INVx4_ASAP7_75t_L g592 ( .A(n_425), .Y(n_592) );
INVx4_ASAP7_75t_L g678 ( .A(n_425), .Y(n_678) );
INVx1_ASAP7_75t_L g759 ( .A(n_425), .Y(n_759) );
INVx2_ASAP7_75t_L g809 ( .A(n_425), .Y(n_809) );
INVx8_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g447 ( .A(n_427), .B(n_445), .Y(n_447) );
AND2x4_ASAP7_75t_L g776 ( .A(n_427), .B(n_445), .Y(n_776) );
AND2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_432), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
BUFx8_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_436), .Y(n_588) );
AND2x4_ASAP7_75t_L g439 ( .A(n_437), .B(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g620 ( .A(n_437), .B(n_445), .Y(n_620) );
BUFx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx12f_ASAP7_75t_L g508 ( .A(n_439), .Y(n_508) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_439), .Y(n_550) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_439), .Y(n_589) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_439), .Y(n_674) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g445 ( .A(n_441), .Y(n_445) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_444), .Y(n_503) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_444), .Y(n_615) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_444), .Y(n_676) );
BUFx12f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx6_ASAP7_75t_L g505 ( .A(n_447), .Y(n_505) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_473), .C(n_478), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_467), .Y(n_450) );
INVx4_ASAP7_75t_L g690 ( .A(n_452), .Y(n_690) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx3_ASAP7_75t_L g521 ( .A(n_453), .Y(n_521) );
BUFx3_ASAP7_75t_L g595 ( .A(n_453), .Y(n_595) );
INVx1_ASAP7_75t_L g669 ( .A(n_453), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_457), .B(n_791), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g929 ( .A(n_457), .B(n_930), .Y(n_929) );
NOR2xp33_ASAP7_75t_L g1244 ( .A(n_457), .B(n_1245), .Y(n_1244) );
INVx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx4_ASAP7_75t_L g662 ( .A(n_458), .Y(n_662) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_459), .Y(n_526) );
AO21x2_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_462), .B(n_465), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_461), .B(n_484), .Y(n_483) );
HB1xp67_ASAP7_75t_L g959 ( .A(n_462), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_470), .Y(n_562) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_470), .Y(n_597) );
BUFx8_ASAP7_75t_SL g664 ( .A(n_470), .Y(n_664) );
BUFx3_ASAP7_75t_L g700 ( .A(n_470), .Y(n_700) );
BUFx3_ASAP7_75t_L g712 ( .A(n_471), .Y(n_712) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_472), .Y(n_535) );
INVx3_ASAP7_75t_L g666 ( .A(n_472), .Y(n_666) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g564 ( .A(n_476), .Y(n_564) );
INVx2_ASAP7_75t_L g750 ( .A(n_476), .Y(n_750) );
INVx2_ASAP7_75t_L g845 ( .A(n_476), .Y(n_845) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx3_ASAP7_75t_L g532 ( .A(n_477), .Y(n_532) );
INVx2_ASAP7_75t_L g601 ( .A(n_477), .Y(n_601) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx3_ASAP7_75t_L g529 ( .A(n_480), .Y(n_529) );
INVx4_ASAP7_75t_L g812 ( .A(n_480), .Y(n_812) );
INVx2_ASAP7_75t_L g843 ( .A(n_480), .Y(n_843) );
INVx5_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx2_ASAP7_75t_L g566 ( .A(n_481), .Y(n_566) );
BUFx4f_ASAP7_75t_L g692 ( .A(n_481), .Y(n_692) );
BUFx2_ASAP7_75t_L g745 ( .A(n_481), .Y(n_745) );
AND2x4_ASAP7_75t_L g481 ( .A(n_482), .B(n_485), .Y(n_481) );
AND2x4_ASAP7_75t_L g605 ( .A(n_482), .B(n_485), .Y(n_605) );
AND2x2_ASAP7_75t_L g770 ( .A(n_482), .B(n_485), .Y(n_770) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g528 ( .A(n_489), .Y(n_528) );
INVx2_ASAP7_75t_L g714 ( .A(n_489), .Y(n_714) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g893 ( .A(n_490), .Y(n_893) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx3_ASAP7_75t_L g567 ( .A(n_491), .Y(n_567) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_491), .Y(n_670) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g572 ( .A(n_496), .Y(n_572) );
OA22x2_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B1(n_540), .B2(n_568), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_517), .Y(n_499) );
INVxp67_ASAP7_75t_L g539 ( .A(n_500), .Y(n_539) );
NAND4xp25_ASAP7_75t_L g500 ( .A(n_501), .B(n_506), .C(n_509), .D(n_514), .Y(n_500) );
BUFx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx5_ASAP7_75t_L g546 ( .A(n_505), .Y(n_546) );
INVx1_ASAP7_75t_L g582 ( .A(n_505), .Y(n_582) );
INVx3_ASAP7_75t_L g616 ( .A(n_505), .Y(n_616) );
INVx2_ASAP7_75t_L g853 ( .A(n_505), .Y(n_853) );
BUFx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx4f_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g584 ( .A(n_512), .Y(n_584) );
INVx1_ASAP7_75t_L g737 ( .A(n_512), .Y(n_737) );
BUFx12f_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_516), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_517), .B(n_538), .Y(n_537) );
NAND4xp25_ASAP7_75t_L g517 ( .A(n_518), .B(n_527), .C(n_530), .D(n_533), .Y(n_517) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g1222 ( .A(n_524), .B(n_1223), .Y(n_1222) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_526), .Y(n_560) );
BUFx6f_ASAP7_75t_L g850 ( .A(n_526), .Y(n_850) );
BUFx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g717 ( .A(n_532), .Y(n_717) );
BUFx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx3_ASAP7_75t_L g686 ( .A(n_535), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OA22x2_ASAP7_75t_L g576 ( .A1(n_541), .A2(n_542), .B1(n_577), .B2(n_578), .Y(n_576) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_SL g568 ( .A(n_542), .Y(n_568) );
NOR2x1_ASAP7_75t_L g543 ( .A(n_544), .B(n_555), .Y(n_543) );
NAND4xp25_ASAP7_75t_L g544 ( .A(n_545), .B(n_547), .C(n_551), .D(n_553), .Y(n_544) );
BUFx4f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx6f_ASAP7_75t_L g757 ( .A(n_549), .Y(n_757) );
NAND4xp25_ASAP7_75t_SL g555 ( .A(n_556), .B(n_561), .C(n_563), .D(n_565), .Y(n_555) );
INVx2_ASAP7_75t_L g627 ( .A(n_557), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx1_ASAP7_75t_L g607 ( .A(n_560), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_560), .B(n_642), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_560), .B(n_748), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_560), .B(n_767), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_560), .B(n_818), .Y(n_817) );
BUFx3_ASAP7_75t_L g711 ( .A(n_562), .Y(n_711) );
INVx2_ASAP7_75t_L g762 ( .A(n_562), .Y(n_762) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
BUFx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g647 ( .A(n_575), .Y(n_647) );
OAI22x1_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_608), .B1(n_643), .B2(n_644), .Y(n_575) );
INVx2_ASAP7_75t_L g643 ( .A(n_576), .Y(n_643) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND4xp75_ASAP7_75t_L g579 ( .A(n_580), .B(n_586), .C(n_593), .D(n_598), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_590), .Y(n_586) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g657 ( .A(n_600), .Y(n_657) );
INVx2_ASAP7_75t_L g701 ( .A(n_600), .Y(n_701) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g866 ( .A(n_601), .Y(n_866) );
OAI21xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B(n_606), .Y(n_602) );
OAI21xp33_ASAP7_75t_L g658 ( .A1(n_604), .A2(n_659), .B(n_660), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g1247 ( .A1(n_604), .A2(n_1248), .B1(n_1250), .B2(n_1252), .Y(n_1247) );
INVx4_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g644 ( .A(n_610), .Y(n_644) );
NAND4xp75_ASAP7_75t_L g611 ( .A(n_612), .B(n_617), .C(n_624), .D(n_636), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_621), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_629), .Y(n_624) );
OAI21xp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B(n_628), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_632), .B1(n_633), .B2(n_635), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g1252 ( .A(n_631), .Y(n_1252) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g765 ( .A(n_638), .Y(n_765) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
XNOR2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_795), .Y(n_648) );
XNOR2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_729), .Y(n_649) );
OAI22x1_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_706), .B1(n_727), .B2(n_728), .Y(n_650) );
INVx1_ASAP7_75t_L g727 ( .A(n_651), .Y(n_727) );
OA22x2_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B1(n_679), .B2(n_705), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_671), .Y(n_654) );
NAND3xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_663), .C(n_667), .Y(n_655) );
INVx2_ASAP7_75t_L g704 ( .A(n_661), .Y(n_704) );
INVx4_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g719 ( .A(n_662), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_662), .B(n_828), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g895 ( .A(n_662), .B(n_896), .Y(n_895) );
NOR2xp33_ASAP7_75t_L g901 ( .A(n_662), .B(n_902), .Y(n_901) );
NOR2xp33_ASAP7_75t_L g945 ( .A(n_662), .B(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g927 ( .A(n_664), .Y(n_927) );
INVx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g743 ( .A(n_666), .Y(n_743) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx3_ASAP7_75t_L g684 ( .A(n_670), .Y(n_684) );
NAND4xp25_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .C(n_675), .D(n_677), .Y(n_671) );
INVx1_ASAP7_75t_L g705 ( .A(n_679), .Y(n_705) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND4xp75_ASAP7_75t_L g681 ( .A(n_682), .B(n_693), .C(n_696), .D(n_699), .Y(n_681) );
NOR2xp67_ASAP7_75t_L g682 ( .A(n_683), .B(n_688), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_685), .B1(n_686), .B2(n_687), .Y(n_683) );
OAI21xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_690), .B(n_691), .Y(n_688) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
INVx1_ASAP7_75t_L g1220 ( .A(n_701), .Y(n_1220) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g728 ( .A(n_706), .Y(n_728) );
BUFx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
XOR2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_726), .Y(n_707) );
NOR2x1_ASAP7_75t_L g708 ( .A(n_709), .B(n_720), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g709 ( .A(n_710), .B(n_713), .C(n_715), .D(n_718), .Y(n_709) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND4xp25_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .C(n_724), .D(n_725), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g1000 ( .A1(n_726), .A2(n_1001), .B1(n_1002), .B2(n_1003), .Y(n_1000) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AO22x2_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_777), .B1(n_793), .B2(n_794), .Y(n_730) );
INVx2_ASAP7_75t_L g794 ( .A(n_731), .Y(n_794) );
XNOR2x1_ASAP7_75t_L g731 ( .A(n_732), .B(n_753), .Y(n_731) );
OAI22x1_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_740), .B1(n_751), .B2(n_752), .Y(n_732) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_734), .B(n_741), .Y(n_751) );
NAND4xp25_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .C(n_738), .D(n_739), .Y(n_734) );
NAND4xp25_ASAP7_75t_L g741 ( .A(n_742), .B(n_744), .C(n_746), .D(n_749), .Y(n_741) );
NAND4xp75_ASAP7_75t_L g754 ( .A(n_755), .B(n_760), .C(n_768), .D(n_772), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_758), .Y(n_755) );
OA21x2_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_762), .B(n_763), .Y(n_760) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_771), .Y(n_768) );
AND2x2_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
BUFx3_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g793 ( .A(n_778), .Y(n_793) );
XNOR2x1_ASAP7_75t_L g778 ( .A(n_779), .B(n_792), .Y(n_778) );
NAND4xp75_ASAP7_75t_L g779 ( .A(n_780), .B(n_783), .C(n_786), .D(n_789), .Y(n_779) );
AND2x2_ASAP7_75t_L g780 ( .A(n_781), .B(n_782), .Y(n_780) );
AND2x2_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
AND2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
XNOR2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_875), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_798), .B1(n_836), .B2(n_874), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
XOR2x2_ASAP7_75t_L g799 ( .A(n_800), .B(n_820), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_801), .A2(n_1044), .B1(n_1045), .B2(n_1046), .Y(n_1043) );
INVx1_ASAP7_75t_L g819 ( .A(n_802), .Y(n_819) );
NAND4xp75_ASAP7_75t_L g802 ( .A(n_803), .B(n_806), .C(n_810), .D(n_814), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
AND2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
AND2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_813), .Y(n_810) );
AND2x2_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
OA22x2_ASAP7_75t_L g857 ( .A1(n_820), .A2(n_858), .B1(n_859), .B2(n_873), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_820), .Y(n_858) );
OR2x2_ASAP7_75t_L g821 ( .A(n_822), .B(n_829), .Y(n_821) );
NAND4xp25_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .C(n_825), .D(n_826), .Y(n_822) );
NAND4xp25_ASAP7_75t_L g829 ( .A(n_830), .B(n_832), .C(n_833), .D(n_834), .Y(n_829) );
INVx1_ASAP7_75t_L g874 ( .A(n_836), .Y(n_874) );
XOR2x2_ASAP7_75t_L g836 ( .A(n_837), .B(n_857), .Y(n_836) );
HB1xp67_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
XNOR2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
NOR2xp67_ASAP7_75t_L g840 ( .A(n_841), .B(n_851), .Y(n_840) );
NAND4xp25_ASAP7_75t_L g841 ( .A(n_842), .B(n_844), .C(n_846), .D(n_847), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_849), .B(n_850), .Y(n_848) );
NAND4xp25_ASAP7_75t_SL g851 ( .A(n_852), .B(n_854), .C(n_855), .D(n_856), .Y(n_851) );
XNOR2xp5_ASAP7_75t_L g859 ( .A(n_860), .B(n_861), .Y(n_859) );
XOR2xp5_ASAP7_75t_L g873 ( .A(n_860), .B(n_861), .Y(n_873) );
OR2x2_ASAP7_75t_L g861 ( .A(n_862), .B(n_868), .Y(n_861) );
NAND4xp25_ASAP7_75t_L g862 ( .A(n_863), .B(n_864), .C(n_865), .D(n_867), .Y(n_862) );
NAND4xp25_ASAP7_75t_L g868 ( .A(n_869), .B(n_870), .C(n_871), .D(n_872), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_935), .B1(n_936), .B2(n_952), .Y(n_875) );
OAI21xp5_ASAP7_75t_L g876 ( .A1(n_877), .A2(n_912), .B(n_932), .Y(n_876) );
AOI22x1_ASAP7_75t_SL g952 ( .A1(n_877), .A2(n_913), .B1(n_933), .B2(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx2_ASAP7_75t_L g934 ( .A(n_878), .Y(n_934) );
AO22x2_ASAP7_75t_L g878 ( .A1(n_879), .A2(n_880), .B1(n_898), .B2(n_911), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx2_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
NAND4xp75_ASAP7_75t_L g882 ( .A(n_883), .B(n_887), .C(n_890), .D(n_894), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_884), .B(n_886), .Y(n_883) );
AND2x2_ASAP7_75t_L g887 ( .A(n_888), .B(n_889), .Y(n_887) );
AND2x2_ASAP7_75t_L g890 ( .A(n_891), .B(n_892), .Y(n_890) );
INVx1_ASAP7_75t_L g911 ( .A(n_898), .Y(n_911) );
NAND3x1_ASAP7_75t_L g899 ( .A(n_900), .B(n_903), .C(n_906), .Y(n_899) );
AND2x2_ASAP7_75t_L g903 ( .A(n_904), .B(n_905), .Y(n_903) );
AND4x1_ASAP7_75t_L g906 ( .A(n_907), .B(n_908), .C(n_909), .D(n_910), .Y(n_906) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
HB1xp67_ASAP7_75t_L g933 ( .A(n_914), .Y(n_933) );
XOR2x2_ASAP7_75t_L g914 ( .A(n_915), .B(n_931), .Y(n_914) );
NOR4xp75_ASAP7_75t_L g915 ( .A(n_916), .B(n_919), .C(n_922), .D(n_925), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_917), .B(n_918), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_920), .B(n_921), .Y(n_919) );
NAND2xp5_ASAP7_75t_SL g922 ( .A(n_923), .B(n_924), .Y(n_922) );
OAI21x1_ASAP7_75t_SL g925 ( .A1(n_926), .A2(n_927), .B(n_928), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_933), .B(n_934), .Y(n_932) );
INVx2_ASAP7_75t_L g953 ( .A(n_934), .Y(n_953) );
INVx3_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
BUFx3_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
XNOR2x1_ASAP7_75t_L g937 ( .A(n_938), .B(n_939), .Y(n_937) );
OR2x2_ASAP7_75t_L g939 ( .A(n_940), .B(n_947), .Y(n_939) );
NAND4xp25_ASAP7_75t_L g940 ( .A(n_941), .B(n_942), .C(n_943), .D(n_944), .Y(n_940) );
NAND4xp25_ASAP7_75t_L g947 ( .A(n_948), .B(n_949), .C(n_950), .D(n_951), .Y(n_947) );
INVx2_ASAP7_75t_SL g954 ( .A(n_955), .Y(n_954) );
NAND3xp33_ASAP7_75t_L g955 ( .A(n_956), .B(n_959), .C(n_960), .Y(n_955) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_956), .B(n_1233), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_956), .B(n_1234), .Y(n_1261) );
INVx1_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
OA21x2_ASAP7_75t_L g1263 ( .A1(n_957), .A2(n_989), .B(n_1264), .Y(n_1263) );
HB1xp67_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
AND2x2_ASAP7_75t_L g969 ( .A(n_958), .B(n_970), .Y(n_969) );
AND3x4_ASAP7_75t_L g988 ( .A(n_958), .B(n_971), .C(n_989), .Y(n_988) );
NOR2xp33_ASAP7_75t_L g1233 ( .A(n_959), .B(n_1234), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_960), .Y(n_1234) );
OAI221xp5_ASAP7_75t_L g961 ( .A1(n_962), .A2(n_1211), .B1(n_1212), .B2(n_1230), .C(n_1235), .Y(n_961) );
AOI211xp5_ASAP7_75t_L g962 ( .A1(n_963), .A2(n_981), .B(n_1115), .C(n_1178), .Y(n_962) );
HB1xp67_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
CKINVDCx16_ASAP7_75t_R g1129 ( .A(n_964), .Y(n_1129) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_965), .B(n_1155), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1176 ( .A(n_965), .B(n_1018), .Y(n_1176) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_965), .B(n_1049), .Y(n_1196) );
BUFx3_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx2_ASAP7_75t_L g1147 ( .A(n_966), .Y(n_1147) );
OAI221xp5_ASAP7_75t_L g966 ( .A1(n_967), .A2(n_973), .B1(n_974), .B2(n_976), .C(n_977), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g1040 ( .A1(n_967), .A2(n_974), .B1(n_1041), .B2(n_1042), .Y(n_1040) );
INVx3_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
AND2x4_ASAP7_75t_L g968 ( .A(n_969), .B(n_971), .Y(n_968) );
AND2x4_ASAP7_75t_L g978 ( .A(n_969), .B(n_979), .Y(n_978) );
AND2x2_ASAP7_75t_L g992 ( .A(n_969), .B(n_979), .Y(n_992) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_969), .B(n_979), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_971), .B(n_975), .Y(n_974) );
AND2x4_ASAP7_75t_L g990 ( .A(n_971), .B(n_975), .Y(n_990) );
AND2x4_ASAP7_75t_L g1015 ( .A(n_971), .B(n_975), .Y(n_1015) );
CKINVDCx5p33_ASAP7_75t_R g1264 ( .A(n_971), .Y(n_1264) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_974), .A2(n_997), .B1(n_998), .B2(n_999), .Y(n_996) );
BUFx2_ASAP7_75t_L g1211 ( .A(n_974), .Y(n_1211) );
AND2x4_ASAP7_75t_L g980 ( .A(n_975), .B(n_979), .Y(n_980) );
AND2x2_ASAP7_75t_L g993 ( .A(n_975), .B(n_979), .Y(n_993) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_975), .B(n_979), .Y(n_1013) );
INVx3_ASAP7_75t_L g1044 ( .A(n_978), .Y(n_1044) );
INVx2_ASAP7_75t_L g1046 ( .A(n_980), .Y(n_1046) );
NAND4xp25_ASAP7_75t_L g981 ( .A(n_982), .B(n_1070), .C(n_1093), .D(n_1111), .Y(n_981) );
AOI211xp5_ASAP7_75t_SL g982 ( .A1(n_983), .A2(n_1016), .B(n_1027), .C(n_1052), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_984), .B(n_994), .Y(n_983) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_984), .B(n_1037), .Y(n_1060) );
NOR2xp33_ASAP7_75t_L g1173 ( .A(n_984), .B(n_1009), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_984), .B(n_1009), .Y(n_1188) );
INVx1_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_986), .B(n_1033), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_986), .B(n_1051), .Y(n_1050) );
CKINVDCx6p67_ASAP7_75t_R g1057 ( .A(n_986), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_986), .B(n_1137), .Y(n_1136) );
OR2x2_ASAP7_75t_L g1146 ( .A(n_986), .B(n_1006), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1166 ( .A(n_986), .B(n_1006), .Y(n_1166) );
NOR2xp33_ASAP7_75t_L g1182 ( .A(n_986), .B(n_1005), .Y(n_1182) );
AND2x2_ASAP7_75t_L g986 ( .A(n_987), .B(n_991), .Y(n_986) );
INVx1_ASAP7_75t_L g997 ( .A(n_988), .Y(n_997) );
INVx2_ASAP7_75t_SL g1022 ( .A(n_990), .Y(n_1022) );
INVx1_ASAP7_75t_L g1003 ( .A(n_992), .Y(n_1003) );
INVx1_ASAP7_75t_L g1002 ( .A(n_993), .Y(n_1002) );
AND2x2_ASAP7_75t_L g994 ( .A(n_995), .B(n_1004), .Y(n_994) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_995), .B(n_1032), .Y(n_1031) );
CKINVDCx6p67_ASAP7_75t_R g1037 ( .A(n_995), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_995), .B(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1105 ( .A(n_995), .Y(n_1105) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_995), .B(n_1110), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_995), .B(n_1068), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g1149 ( .A1(n_995), .A2(n_1086), .B1(n_1150), .B2(n_1152), .Y(n_1149) );
NOR2xp33_ASAP7_75t_L g1174 ( .A(n_995), .B(n_1039), .Y(n_1174) );
NAND4xp25_ASAP7_75t_L g1177 ( .A(n_995), .B(n_1005), .C(n_1129), .D(n_1133), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_995), .B(n_1048), .Y(n_1206) );
OR2x6_ASAP7_75t_SL g995 ( .A(n_996), .B(n_1000), .Y(n_995) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1004), .B(n_1060), .Y(n_1123) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_1004), .B(n_1037), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1004), .B(n_1069), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1009), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_1005), .B(n_1010), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_1005), .B(n_1060), .Y(n_1085) );
CKINVDCx5p33_ASAP7_75t_R g1005 ( .A(n_1006), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_1006), .B(n_1009), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1006), .B(n_1010), .Y(n_1068) );
OAI32xp33_ASAP7_75t_L g1101 ( .A1(n_1006), .A2(n_1079), .A3(n_1102), .B1(n_1106), .B2(n_1109), .Y(n_1101) );
AND2x4_ASAP7_75t_SL g1006 ( .A(n_1007), .B(n_1008), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1009), .B(n_1057), .Y(n_1110) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1009), .Y(n_1120) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1014), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1016), .B(n_1100), .Y(n_1099) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
O2A1O1Ixp33_ASAP7_75t_L g1142 ( .A1(n_1017), .A2(n_1143), .B(n_1144), .C(n_1147), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1023), .Y(n_1017) );
INVx3_ASAP7_75t_L g1049 ( .A(n_1018), .Y(n_1049) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1018), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_1018), .B(n_1024), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_1018), .B(n_1038), .Y(n_1092) );
NOR2xp33_ASAP7_75t_L g1103 ( .A(n_1018), .B(n_1104), .Y(n_1103) );
OR2x2_ASAP7_75t_L g1108 ( .A(n_1018), .B(n_1023), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1018), .B(n_1134), .Y(n_1133) );
AND2x4_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1020), .Y(n_1018) );
INVx2_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx3_ASAP7_75t_L g1029 ( .A(n_1023), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_1023), .B(n_1039), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_1023), .B(n_1049), .Y(n_1113) );
INVx2_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_1024), .B(n_1039), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1024), .B(n_1048), .Y(n_1080) );
OR2x2_ASAP7_75t_L g1088 ( .A(n_1024), .B(n_1039), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1026), .Y(n_1024) );
OAI21xp33_ASAP7_75t_L g1027 ( .A1(n_1028), .A2(n_1030), .B(n_1034), .Y(n_1027) );
AOI21xp5_ASAP7_75t_L g1180 ( .A1(n_1028), .A2(n_1135), .B(n_1181), .Y(n_1180) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
INVx3_ASAP7_75t_L g1155 ( .A(n_1029), .Y(n_1155) );
INVxp67_ASAP7_75t_SL g1030 ( .A(n_1031), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_1032), .B(n_1159), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_1033), .B(n_1060), .Y(n_1059) );
OR2x2_ASAP7_75t_L g1095 ( .A(n_1033), .B(n_1051), .Y(n_1095) );
NAND2xp5_ASAP7_75t_L g1141 ( .A(n_1033), .B(n_1104), .Y(n_1141) );
AND2x2_ASAP7_75t_SL g1151 ( .A(n_1033), .B(n_1057), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1033), .B(n_1069), .Y(n_1160) );
OAI21xp5_ASAP7_75t_L g1034 ( .A1(n_1035), .A2(n_1047), .B(n_1050), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1038), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_1037), .B(n_1057), .Y(n_1069) );
NOR2xp33_ASAP7_75t_L g1096 ( .A(n_1037), .B(n_1088), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1121 ( .A(n_1037), .B(n_1084), .Y(n_1121) );
NOR2x1p5_ASAP7_75t_L g1145 ( .A(n_1037), .B(n_1146), .Y(n_1145) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1037), .Y(n_1170) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1038), .Y(n_1131) );
INVx3_ASAP7_75t_L g1048 ( .A(n_1039), .Y(n_1048) );
INVx2_ASAP7_75t_L g1063 ( .A(n_1039), .Y(n_1063) );
OR2x2_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1043), .Y(n_1039) );
AOI322xp5_ASAP7_75t_L g1207 ( .A1(n_1047), .A2(n_1054), .A3(n_1062), .B1(n_1096), .B2(n_1182), .C1(n_1208), .C2(n_1209), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1049), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_1048), .B(n_1073), .Y(n_1072) );
NOR2xp33_ASAP7_75t_L g1107 ( .A(n_1048), .B(n_1108), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1048), .B(n_1059), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1048), .B(n_1083), .Y(n_1199) );
INVx2_ASAP7_75t_L g1083 ( .A(n_1049), .Y(n_1083) );
HB1xp67_ASAP7_75t_L g1124 ( .A(n_1049), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1050), .B(n_1104), .Y(n_1114) );
NOR2xp33_ASAP7_75t_L g1150 ( .A(n_1050), .B(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1051), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_1051), .B(n_1057), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_1051), .B(n_1091), .Y(n_1090) );
A2O1A1Ixp33_ASAP7_75t_L g1052 ( .A1(n_1053), .A2(n_1058), .B(n_1061), .C(n_1065), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
NOR2xp33_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1056), .Y(n_1054) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1056), .Y(n_1078) );
NOR2xp33_ASAP7_75t_L g1094 ( .A(n_1057), .B(n_1095), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1057), .B(n_1068), .Y(n_1098) );
NOR2xp33_ASAP7_75t_L g1127 ( .A(n_1057), .B(n_1128), .Y(n_1127) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_1060), .B(n_1068), .Y(n_1073) );
NOR2xp33_ASAP7_75t_L g1125 ( .A(n_1061), .B(n_1126), .Y(n_1125) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
NOR2xp33_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1064), .Y(n_1062) );
NOR2xp33_ASAP7_75t_L g1066 ( .A(n_1063), .B(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1063), .Y(n_1100) );
BUFx2_ASAP7_75t_L g1159 ( .A(n_1063), .Y(n_1159) );
INVxp67_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1067), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1069), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1068), .B(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1068), .Y(n_1128) );
AOI211xp5_ASAP7_75t_L g1070 ( .A1(n_1071), .A2(n_1074), .B(n_1075), .C(n_1089), .Y(n_1070) );
INVxp67_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1073), .B(n_1100), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1074), .B(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1074), .Y(n_1204) );
OAI222xp33_ASAP7_75t_L g1075 ( .A1(n_1076), .A2(n_1079), .B1(n_1081), .B2(n_1085), .C1(n_1086), .C2(n_1088), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
NOR2xp33_ASAP7_75t_L g1202 ( .A(n_1079), .B(n_1147), .Y(n_1202) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
AOI322xp5_ASAP7_75t_L g1164 ( .A1(n_1080), .A2(n_1123), .A3(n_1165), .B1(n_1167), .B2(n_1169), .C1(n_1171), .C2(n_1175), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1084), .Y(n_1081) );
INVx3_ASAP7_75t_L g1152 ( .A(n_1082), .Y(n_1152) );
INVx3_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_1084), .B(n_1104), .Y(n_1190) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1201 ( .A(n_1087), .B(n_1202), .Y(n_1201) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1088), .Y(n_1134) );
INVxp67_ASAP7_75t_SL g1089 ( .A(n_1090), .Y(n_1089) );
O2A1O1Ixp33_ASAP7_75t_L g1138 ( .A1(n_1091), .A2(n_1139), .B(n_1140), .C(n_1142), .Y(n_1138) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
AOI221xp5_ASAP7_75t_L g1093 ( .A1(n_1094), .A2(n_1096), .B1(n_1097), .B2(n_1099), .C(n_1101), .Y(n_1093) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
INVxp33_ASAP7_75t_SL g1102 ( .A(n_1103), .Y(n_1102) );
INVx3_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1108), .Y(n_1163) );
INVxp67_ASAP7_75t_SL g1111 ( .A(n_1112), .Y(n_1111) );
NOR2xp33_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1114), .Y(n_1112) );
NAND5xp2_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1148), .C(n_1156), .D(n_1164), .E(n_1177), .Y(n_1115) );
O2A1O1Ixp33_ASAP7_75t_L g1116 ( .A1(n_1117), .A2(n_1125), .B(n_1129), .C(n_1130), .Y(n_1116) );
O2A1O1Ixp33_ASAP7_75t_SL g1117 ( .A1(n_1118), .A2(n_1121), .B(n_1122), .C(n_1124), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
A2O1A1Ixp33_ASAP7_75t_L g1130 ( .A1(n_1131), .A2(n_1132), .B(n_1135), .C(n_1138), .Y(n_1130) );
AOI21xp33_ASAP7_75t_L g1183 ( .A1(n_1131), .A2(n_1169), .B(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
AOI222xp33_ASAP7_75t_L g1148 ( .A1(n_1133), .A2(n_1134), .B1(n_1149), .B2(n_1151), .C1(n_1153), .C2(n_1155), .Y(n_1148) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
OAI31xp33_ASAP7_75t_L g1156 ( .A1(n_1136), .A2(n_1157), .A3(n_1161), .B(n_1163), .Y(n_1156) );
INVxp67_ASAP7_75t_L g1192 ( .A(n_1137), .Y(n_1192) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
CKINVDCx16_ASAP7_75t_R g1185 ( .A(n_1147), .Y(n_1185) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1151), .Y(n_1184) );
INVx3_ASAP7_75t_L g1208 ( .A(n_1152), .Y(n_1208) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1160), .Y(n_1157) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1158), .Y(n_1193) );
INVx2_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
AOI211xp5_ASAP7_75t_L g1197 ( .A1(n_1160), .A2(n_1198), .B(n_1200), .C(n_1203), .Y(n_1197) );
INVxp33_ASAP7_75t_SL g1161 ( .A(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
CKINVDCx14_ASAP7_75t_R g1169 ( .A(n_1170), .Y(n_1169) );
INVxp67_ASAP7_75t_SL g1171 ( .A(n_1172), .Y(n_1171) );
NAND2xp5_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1174), .Y(n_1172) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_1174), .B(n_1182), .Y(n_1181) );
CKINVDCx14_ASAP7_75t_R g1175 ( .A(n_1176), .Y(n_1175) );
AOI21xp33_ASAP7_75t_SL g1203 ( .A1(n_1176), .A2(n_1204), .B(n_1205), .Y(n_1203) );
NAND4xp25_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1186), .C(n_1197), .D(n_1207), .Y(n_1178) );
OAI21xp5_ASAP7_75t_SL g1179 ( .A1(n_1180), .A2(n_1183), .B(n_1185), .Y(n_1179) );
A2O1A1Ixp33_ASAP7_75t_L g1191 ( .A1(n_1184), .A2(n_1192), .B(n_1193), .C(n_1194), .Y(n_1191) );
A2O1A1Ixp33_ASAP7_75t_L g1186 ( .A1(n_1187), .A2(n_1189), .B(n_1191), .C(n_1195), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1188), .B(n_1206), .Y(n_1205) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
INVxp67_ASAP7_75t_SL g1200 ( .A(n_1201), .Y(n_1200) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
HB1xp67_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
NAND4xp75_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1218), .C(n_1224), .D(n_1227), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1216), .B(n_1217), .Y(n_1215) );
OA21x2_ASAP7_75t_L g1218 ( .A1(n_1219), .A2(n_1220), .B(n_1221), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1226), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1228), .B(n_1229), .Y(n_1227) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
HB1xp67_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
INVxp33_ASAP7_75t_SL g1236 ( .A(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
HB1xp67_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
NOR2x1_ASAP7_75t_L g1241 ( .A(n_1242), .B(n_1254), .Y(n_1241) );
NAND3xp33_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1246), .C(n_1253), .Y(n_1242) );
CKINVDCx16_ASAP7_75t_R g1248 ( .A(n_1249), .Y(n_1248) );
CKINVDCx9p33_ASAP7_75t_R g1250 ( .A(n_1251), .Y(n_1250) );
NAND4xp25_ASAP7_75t_L g1254 ( .A(n_1255), .B(n_1256), .C(n_1257), .D(n_1258), .Y(n_1254) );
BUFx2_ASAP7_75t_SL g1260 ( .A(n_1261), .Y(n_1260) );
HB1xp67_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
endmodule