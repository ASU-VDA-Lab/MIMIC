module fake_jpeg_2164_n_698 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_698);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_698;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_17),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_22),
.B(n_19),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_61),
.B(n_73),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_22),
.B(n_9),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_63),
.B(n_116),
.Y(n_137)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_66),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_67),
.Y(n_192)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_68),
.Y(n_209)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_69),
.Y(n_214)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_71),
.Y(n_162)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_28),
.B(n_10),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_28),
.B(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_74),
.B(n_83),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_76),
.Y(n_187)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_78),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_79),
.Y(n_195)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_80),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_81),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_82),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_30),
.B(n_10),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_30),
.B(n_10),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_84),
.B(n_88),
.Y(n_164)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_85),
.Y(n_166)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_87),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_10),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_36),
.Y(n_89)
);

CKINVDCx6p67_ASAP7_75t_R g203 ( 
.A(n_89),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_91),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g218 ( 
.A(n_92),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

BUFx24_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

BUFx8_ASAP7_75t_L g189 ( 
.A(n_94),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_96),
.Y(n_190)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_97),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_36),
.Y(n_100)
);

INVx13_ASAP7_75t_L g221 ( 
.A(n_100),
.Y(n_221)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_102),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_59),
.B1(n_31),
.B2(n_21),
.Y(n_135)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_104),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_107),
.Y(n_227)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_109),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g200 ( 
.A(n_110),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_111),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_112),
.Y(n_230)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_29),
.Y(n_113)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_39),
.Y(n_115)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_115),
.Y(n_191)
);

AOI21xp33_ASAP7_75t_SL g116 ( 
.A1(n_39),
.A2(n_8),
.B(n_18),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_39),
.Y(n_117)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_118),
.Y(n_197)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_120),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_50),
.B(n_8),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_58),
.Y(n_140)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_122),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_43),
.Y(n_123)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_123),
.Y(n_215)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_124),
.Y(n_217)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_45),
.Y(n_125)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_125),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_43),
.Y(n_126)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_126),
.Y(n_224)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_36),
.Y(n_127)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_127),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_43),
.Y(n_128)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_36),
.Y(n_129)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_24),
.Y(n_130)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_20),
.B(n_19),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_16),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_53),
.Y(n_133)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_133),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_33),
.B1(n_34),
.B2(n_56),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_134),
.A2(n_161),
.B1(n_168),
.B2(n_182),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_135),
.A2(n_156),
.B1(n_185),
.B2(n_205),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_140),
.B(n_94),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_63),
.B(n_35),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_146),
.B(n_153),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_66),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_121),
.A2(n_34),
.B1(n_56),
.B2(n_54),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_120),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_157),
.B(n_188),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_89),
.B(n_40),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_158),
.B(n_171),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_100),
.A2(n_54),
.B1(n_49),
.B2(n_48),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g240 ( 
.A1(n_160),
.A2(n_165),
.B1(n_206),
.B2(n_228),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_21),
.B1(n_31),
.B2(n_59),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_133),
.A2(n_53),
.B1(n_44),
.B2(n_46),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_76),
.A2(n_40),
.B1(n_49),
.B2(n_48),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_72),
.B(n_33),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_174),
.B(n_175),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_35),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_67),
.B(n_20),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_181),
.B(n_186),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_126),
.A2(n_53),
.B1(n_38),
.B2(n_24),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_128),
.A2(n_38),
.B1(n_46),
.B2(n_44),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_67),
.B(n_47),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_91),
.B(n_47),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_91),
.B(n_47),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_196),
.B(n_201),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_90),
.B(n_44),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_98),
.B(n_46),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_202),
.B(n_220),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_62),
.A2(n_25),
.B1(n_7),
.B2(n_11),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_105),
.A2(n_25),
.B1(n_17),
.B2(n_16),
.Y(n_206)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_106),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_65),
.B(n_25),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_71),
.B(n_17),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_223),
.B(n_155),
.Y(n_239)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_79),
.Y(n_225)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_118),
.B(n_17),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_226),
.B(n_0),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_94),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_228)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_138),
.Y(n_232)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_232),
.Y(n_329)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_233),
.Y(n_316)
);

OAI22xp33_ASAP7_75t_L g234 ( 
.A1(n_161),
.A2(n_82),
.B1(n_112),
.B2(n_111),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_234),
.A2(n_241),
.B1(n_277),
.B2(n_300),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_236),
.Y(n_318)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_237),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_L g361 ( 
.A1(n_238),
.A2(n_262),
.B(n_263),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_239),
.B(n_276),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_L g241 ( 
.A1(n_165),
.A2(n_114),
.B1(n_110),
.B2(n_107),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_141),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_242),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_141),
.Y(n_243)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_243),
.Y(n_325)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_244),
.Y(n_378)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_245),
.Y(n_375)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_138),
.Y(n_246)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_246),
.Y(n_368)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_139),
.Y(n_248)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_248),
.Y(n_324)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_170),
.Y(n_249)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_249),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_137),
.B(n_75),
.C(n_99),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_250),
.B(n_282),
.C(n_293),
.Y(n_376)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_251),
.Y(n_327)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_152),
.Y(n_252)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_252),
.Y(n_335)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_154),
.Y(n_253)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_253),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_144),
.B(n_102),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_254),
.B(n_279),
.Y(n_341)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_150),
.Y(n_255)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_255),
.Y(n_347)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_169),
.Y(n_256)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_256),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_189),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_257),
.Y(n_328)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_145),
.Y(n_258)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_258),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_189),
.A2(n_93),
.B1(n_87),
.B2(n_81),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_259),
.Y(n_320)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_145),
.Y(n_260)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_260),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_203),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_261),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_203),
.A2(n_13),
.B(n_12),
.Y(n_262)
);

A2O1A1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_164),
.A2(n_12),
.B(n_1),
.C(n_2),
.Y(n_263)
);

INVx6_ASAP7_75t_SL g264 ( 
.A(n_203),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_264),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_185),
.A2(n_95),
.B1(n_12),
.B2(n_2),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_265),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_176),
.A2(n_214),
.B1(n_209),
.B2(n_190),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_268),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_170),
.Y(n_269)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_269),
.Y(n_369)
);

INVx3_ASAP7_75t_SL g270 ( 
.A(n_199),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_270),
.Y(n_364)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_219),
.Y(n_273)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_273),
.Y(n_373)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_275),
.B(n_280),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_L g277 ( 
.A1(n_160),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_184),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_278),
.B(n_281),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_187),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_184),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_192),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g282 ( 
.A(n_166),
.B(n_0),
.Y(n_282)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_192),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_285),
.B(n_290),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_187),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_286),
.B(n_287),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_167),
.B(n_1),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_172),
.B(n_3),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_288),
.B(n_291),
.Y(n_367)
);

INVx8_ASAP7_75t_L g289 ( 
.A(n_200),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_289),
.A2(n_297),
.B1(n_298),
.B2(n_301),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_209),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_173),
.B(n_4),
.Y(n_291)
);

AOI32xp33_ASAP7_75t_L g292 ( 
.A1(n_191),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_198),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_292),
.A2(n_305),
.B1(n_312),
.B2(n_149),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_193),
.B(n_4),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_214),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_294),
.Y(n_353)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_136),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_295),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_204),
.B(n_5),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_296),
.B(n_211),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_190),
.A2(n_5),
.B1(n_6),
.B2(n_194),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_163),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_147),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_299),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_L g300 ( 
.A1(n_206),
.A2(n_5),
.B1(n_230),
.B2(n_222),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_163),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_151),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_302),
.Y(n_372)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_179),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_303),
.A2(n_304),
.B1(n_306),
.B2(n_308),
.Y(n_357)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_222),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_182),
.A2(n_5),
.B1(n_230),
.B2(n_228),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_179),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_213),
.B(n_199),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_310),
.Y(n_317)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_194),
.Y(n_308)
);

BUFx6f_ASAP7_75t_SL g309 ( 
.A(n_221),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_309),
.A2(n_148),
.B1(n_236),
.B2(n_257),
.Y(n_370)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_143),
.Y(n_310)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_183),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_143),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_313),
.B(n_264),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_142),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_142),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_326),
.B(n_280),
.Y(n_411)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_331),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_272),
.A2(n_231),
.B1(n_210),
.B2(n_208),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_332),
.A2(n_333),
.B1(n_340),
.B2(n_354),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_283),
.A2(n_231),
.B1(n_210),
.B2(n_208),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_336),
.B(n_377),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_283),
.A2(n_227),
.B1(n_159),
.B2(n_207),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_337),
.A2(n_346),
.B1(n_351),
.B2(n_366),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_234),
.A2(n_195),
.B1(n_162),
.B2(n_183),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_282),
.B(n_227),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_342),
.B(n_365),
.Y(n_382)
);

AOI22x1_ASAP7_75t_L g344 ( 
.A1(n_240),
.A2(n_221),
.B1(n_218),
.B2(n_200),
.Y(n_344)
);

OA22x2_ASAP7_75t_L g427 ( 
.A1(n_344),
.A2(n_249),
.B1(n_269),
.B2(n_309),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_250),
.B(n_271),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_345),
.B(n_311),
.C(n_238),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_267),
.A2(n_274),
.B1(n_315),
.B2(n_284),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_282),
.A2(n_207),
.B1(n_159),
.B2(n_178),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_241),
.A2(n_195),
.B1(n_162),
.B2(n_180),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_238),
.A2(n_180),
.B1(n_212),
.B2(n_218),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_362),
.A2(n_270),
.B(n_312),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_293),
.B(n_178),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_240),
.A2(n_200),
.B1(n_212),
.B2(n_148),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_370),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_293),
.B(n_148),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_374),
.B(n_296),
.Y(n_388)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_377),
.Y(n_380)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_380),
.Y(n_438)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_347),
.Y(n_381)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_381),
.Y(n_453)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_383),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_384),
.B(n_390),
.C(n_421),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_344),
.A2(n_300),
.B(n_277),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_385),
.A2(n_387),
.B(n_415),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_344),
.A2(n_240),
.B(n_262),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_388),
.B(n_396),
.Y(n_459)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_324),
.Y(n_389)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_389),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_345),
.B(n_376),
.C(n_326),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_366),
.A2(n_240),
.B1(n_266),
.B2(n_306),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_391),
.A2(n_424),
.B(n_357),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_371),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_392),
.B(n_401),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_332),
.A2(n_333),
.B1(n_336),
.B2(n_321),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_393),
.A2(n_398),
.B1(n_413),
.B2(n_422),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_342),
.B(n_296),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_394),
.B(n_397),
.Y(n_432)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_335),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_395),
.Y(n_430)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_335),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_263),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_321),
.A2(n_310),
.B1(n_295),
.B2(n_299),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_341),
.B(n_235),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_399),
.B(n_405),
.Y(n_429)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_324),
.Y(n_400)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_400),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_371),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_320),
.A2(n_350),
.B1(n_360),
.B2(n_353),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_SL g440 ( 
.A1(n_403),
.A2(n_418),
.B1(n_318),
.B2(n_402),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_358),
.B(n_308),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_349),
.B(n_247),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_406),
.B(n_410),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_322),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_407),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_375),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_408),
.B(n_412),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_376),
.B(n_245),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_373),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_372),
.B(n_255),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_340),
.A2(n_244),
.B1(n_237),
.B2(n_251),
.Y(n_413)
);

CKINVDCx14_ASAP7_75t_R g414 ( 
.A(n_355),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_414),
.B(n_416),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_360),
.A2(n_290),
.B(n_232),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_355),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_359),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_417),
.B(n_419),
.Y(n_455)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_325),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_361),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_351),
.A2(n_317),
.B1(n_350),
.B2(n_320),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_420),
.A2(n_368),
.B1(n_329),
.B2(n_327),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_317),
.B(n_294),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_354),
.A2(n_314),
.B1(n_243),
.B2(n_242),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_359),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_423),
.B(n_426),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_365),
.A2(n_303),
.B1(n_301),
.B2(n_298),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_425),
.A2(n_331),
.B1(n_353),
.B2(n_348),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_374),
.A2(n_246),
.B1(n_281),
.B2(n_285),
.Y(n_426)
);

OA21x2_ASAP7_75t_L g444 ( 
.A1(n_427),
.A2(n_352),
.B(n_369),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_356),
.B(n_289),
.C(n_343),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_428),
.B(n_334),
.C(n_355),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_433),
.B(n_434),
.C(n_441),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_390),
.B(n_356),
.C(n_363),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_412),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_435),
.B(n_467),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_419),
.A2(n_362),
.B(n_339),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_436),
.A2(n_458),
.B(n_443),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_437),
.B(n_442),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_440),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_410),
.B(n_363),
.C(n_343),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_384),
.B(n_411),
.C(n_421),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_444),
.B(n_452),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_380),
.B(n_319),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_445),
.B(n_446),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_382),
.B(n_373),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_382),
.B(n_394),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_447),
.B(n_450),
.Y(n_484)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_448),
.Y(n_472)
);

MAJx2_ASAP7_75t_L g450 ( 
.A(n_409),
.B(n_352),
.C(n_323),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_388),
.B(n_352),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_379),
.B(n_327),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_460),
.B(n_400),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_461),
.A2(n_470),
.B1(n_444),
.B2(n_422),
.Y(n_482)
);

OAI211xp5_ASAP7_75t_SL g463 ( 
.A1(n_387),
.A2(n_316),
.B(n_330),
.C(n_378),
.Y(n_463)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_463),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_415),
.A2(n_369),
.B(n_338),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_465),
.A2(n_466),
.B(n_427),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_424),
.A2(n_338),
.B(n_368),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_406),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_391),
.A2(n_325),
.B1(n_322),
.B2(n_329),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_458),
.A2(n_409),
.B(n_401),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_471),
.A2(n_473),
.B(n_480),
.Y(n_520)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_449),
.Y(n_474)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_474),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_443),
.A2(n_386),
.B1(n_409),
.B2(n_385),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_477),
.B(n_479),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_464),
.A2(n_386),
.B1(n_420),
.B2(n_379),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_455),
.A2(n_392),
.B(n_397),
.Y(n_480)
);

INVxp33_ASAP7_75t_L g528 ( 
.A(n_482),
.Y(n_528)
);

AO22x1_ASAP7_75t_SL g483 ( 
.A1(n_438),
.A2(n_393),
.B1(n_404),
.B2(n_398),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_483),
.B(n_488),
.Y(n_516)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_430),
.Y(n_486)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_486),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_435),
.B(n_459),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_464),
.A2(n_438),
.B1(n_454),
.B2(n_432),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_489),
.B(n_490),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_454),
.A2(n_404),
.B1(n_416),
.B2(n_399),
.Y(n_490)
);

OAI32xp33_ASAP7_75t_L g491 ( 
.A1(n_432),
.A2(n_405),
.A3(n_396),
.B1(n_395),
.B2(n_423),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_491),
.B(n_492),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_451),
.B(n_417),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_439),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_493),
.B(n_494),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_439),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_470),
.A2(n_413),
.B1(n_425),
.B2(n_426),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_495),
.A2(n_482),
.B1(n_472),
.B2(n_502),
.Y(n_522)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_453),
.Y(n_496)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_496),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_455),
.A2(n_462),
.B1(n_461),
.B2(n_463),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_497),
.A2(n_500),
.B(n_509),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_429),
.B(n_408),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_498),
.B(n_499),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_462),
.A2(n_428),
.B(n_381),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_453),
.Y(n_501)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_501),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_460),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_502),
.B(n_503),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_457),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_459),
.B(n_389),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_505),
.B(n_506),
.Y(n_542)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_456),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_445),
.B(n_383),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_507),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_429),
.B(n_418),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_508),
.B(n_449),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_485),
.B(n_431),
.C(n_434),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_511),
.B(n_515),
.C(n_523),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_492),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_514),
.B(n_541),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_485),
.B(n_431),
.C(n_442),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_478),
.B(n_441),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_517),
.B(n_526),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_476),
.B(n_447),
.Y(n_518)
);

XNOR2x1_ASAP7_75t_L g568 ( 
.A(n_518),
.B(n_531),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_503),
.A2(n_444),
.B1(n_457),
.B2(n_466),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_519),
.A2(n_530),
.B1(n_536),
.B2(n_548),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_522),
.A2(n_538),
.B1(n_546),
.B2(n_479),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_478),
.B(n_452),
.C(n_446),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_476),
.B(n_433),
.C(n_437),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_525),
.B(n_540),
.C(n_523),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_484),
.B(n_450),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_475),
.A2(n_444),
.B1(n_465),
.B2(n_467),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_SL g531 ( 
.A(n_484),
.B(n_507),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_533),
.B(n_474),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_471),
.A2(n_436),
.B(n_456),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_535),
.A2(n_545),
.B(n_520),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_475),
.A2(n_468),
.B1(n_469),
.B2(n_427),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_497),
.A2(n_468),
.B1(n_469),
.B2(n_427),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_500),
.B(n_316),
.C(n_378),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_498),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_489),
.B(n_427),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_543),
.B(n_544),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_504),
.B(n_375),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_471),
.A2(n_328),
.B(n_318),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_504),
.A2(n_407),
.B1(n_328),
.B2(n_330),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_509),
.A2(n_364),
.B1(n_407),
.B2(n_493),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_534),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_549),
.B(n_560),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_520),
.A2(n_473),
.B(n_504),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_SL g584 ( 
.A1(n_552),
.A2(n_535),
.B(n_527),
.Y(n_584)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_537),
.Y(n_553)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_553),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_515),
.B(n_490),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g596 ( 
.A(n_555),
.B(n_561),
.Y(n_596)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_537),
.Y(n_557)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_557),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_545),
.B(n_477),
.Y(n_558)
);

AND2x2_ASAP7_75t_SL g597 ( 
.A(n_558),
.B(n_573),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_559),
.A2(n_527),
.B(n_530),
.Y(n_589)
);

CKINVDCx16_ASAP7_75t_R g560 ( 
.A(n_534),
.Y(n_560)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_542),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_562),
.B(n_574),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_511),
.B(n_480),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_563),
.B(n_570),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_517),
.B(n_487),
.C(n_488),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_564),
.B(n_566),
.C(n_578),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_532),
.A2(n_494),
.B1(n_481),
.B2(n_472),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_565),
.B(n_569),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_525),
.B(n_487),
.C(n_499),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_567),
.A2(n_516),
.B1(n_510),
.B2(n_543),
.Y(n_585)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_513),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_518),
.B(n_491),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_531),
.B(n_508),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_571),
.B(n_572),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_526),
.B(n_505),
.Y(n_572)
);

XNOR2x1_ASAP7_75t_L g573 ( 
.A(n_544),
.B(n_486),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_542),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_514),
.B(n_496),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_575),
.B(n_576),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_539),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_532),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_577),
.B(n_581),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_529),
.B(n_483),
.Y(n_578)
);

CKINVDCx16_ASAP7_75t_R g601 ( 
.A(n_579),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_541),
.B(n_501),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_580),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_539),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_SL g610 ( 
.A1(n_584),
.A2(n_559),
.B(n_558),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_585),
.A2(n_594),
.B1(n_569),
.B2(n_524),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_589),
.A2(n_584),
.B(n_609),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_567),
.A2(n_554),
.B1(n_516),
.B2(n_582),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_591),
.A2(n_604),
.B1(n_606),
.B2(n_579),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_550),
.B(n_540),
.C(n_512),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_592),
.B(n_593),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_550),
.B(n_561),
.C(n_555),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_582),
.A2(n_528),
.B1(n_529),
.B2(n_510),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_563),
.B(n_512),
.C(n_548),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_598),
.B(n_607),
.Y(n_630)
);

XNOR2x2_ASAP7_75t_SL g600 ( 
.A(n_552),
.B(n_519),
.Y(n_600)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_600),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_578),
.A2(n_522),
.B1(n_538),
.B2(n_536),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_558),
.A2(n_546),
.B1(n_483),
.B2(n_521),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_551),
.B(n_521),
.C(n_513),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_551),
.B(n_524),
.C(n_547),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_608),
.B(n_564),
.C(n_573),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_L g635 ( 
.A1(n_610),
.A2(n_603),
.B(n_600),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_608),
.B(n_566),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g651 ( 
.A(n_611),
.B(n_618),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_612),
.B(n_615),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_595),
.B(n_570),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_SL g637 ( 
.A(n_614),
.B(n_623),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_593),
.B(n_556),
.C(n_572),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_607),
.B(n_571),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g638 ( 
.A(n_616),
.B(n_617),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_596),
.B(n_556),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_590),
.B(n_568),
.Y(n_618)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_619),
.Y(n_648)
);

CKINVDCx16_ASAP7_75t_R g620 ( 
.A(n_587),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_620),
.B(n_583),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_SL g646 ( 
.A1(n_621),
.A2(n_599),
.B1(n_597),
.B2(n_601),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_SL g622 ( 
.A1(n_604),
.A2(n_483),
.B1(n_495),
.B2(n_547),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_622),
.B(n_628),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_SL g623 ( 
.A(n_595),
.B(n_506),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_596),
.B(n_568),
.C(n_364),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_624),
.B(n_625),
.C(n_590),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_592),
.B(n_583),
.C(n_598),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_586),
.Y(n_626)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_626),
.Y(n_640)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_586),
.Y(n_628)
);

AOI21x1_ASAP7_75t_L g634 ( 
.A1(n_629),
.A2(n_589),
.B(n_603),
.Y(n_634)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_609),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_631),
.B(n_632),
.Y(n_644)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_602),
.Y(n_632)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_633),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_634),
.B(n_636),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_SL g658 ( 
.A1(n_635),
.A2(n_610),
.B(n_591),
.Y(n_658)
);

NOR2xp67_ASAP7_75t_L g636 ( 
.A(n_628),
.B(n_605),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_SL g639 ( 
.A1(n_627),
.A2(n_600),
.B(n_606),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_639),
.B(n_643),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_613),
.B(n_605),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_645),
.B(n_616),
.Y(n_659)
);

XOR2xp5_ASAP7_75t_L g661 ( 
.A(n_646),
.B(n_621),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_629),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_647),
.B(n_649),
.Y(n_656)
);

INVx11_ASAP7_75t_L g649 ( 
.A(n_632),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_631),
.B(n_599),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_650),
.B(n_627),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_638),
.B(n_625),
.C(n_611),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_652),
.B(n_655),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_637),
.B(n_630),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_SL g673 ( 
.A(n_653),
.B(n_659),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_SL g655 ( 
.A(n_642),
.B(n_615),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_657),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_658),
.A2(n_639),
.B(n_646),
.Y(n_672)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_661),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_647),
.B(n_612),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_663),
.B(n_664),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_644),
.B(n_594),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_644),
.B(n_640),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_665),
.B(n_666),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_638),
.B(n_617),
.C(n_588),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_645),
.B(n_624),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_667),
.B(n_666),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_SL g668 ( 
.A1(n_654),
.A2(n_634),
.B(n_635),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_668),
.B(n_622),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_670),
.B(n_672),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_662),
.A2(n_648),
.B(n_640),
.Y(n_674)
);

AOI21x1_ASAP7_75t_L g682 ( 
.A1(n_674),
.A2(n_641),
.B(n_660),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_652),
.B(n_648),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_675),
.B(n_669),
.Y(n_680)
);

AND3x1_ASAP7_75t_L g677 ( 
.A(n_656),
.B(n_641),
.C(n_650),
.Y(n_677)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_677),
.Y(n_681)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_680),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_682),
.A2(n_685),
.B(n_687),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_673),
.B(n_659),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_684),
.B(n_686),
.Y(n_688)
);

A2O1A1O1Ixp25_ASAP7_75t_L g685 ( 
.A1(n_676),
.A2(n_672),
.B(n_679),
.C(n_671),
.D(n_677),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_678),
.B(n_661),
.Y(n_686)
);

MAJIxp5_ASAP7_75t_L g691 ( 
.A(n_683),
.B(n_674),
.C(n_668),
.Y(n_691)
);

A2O1A1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_691),
.A2(n_681),
.B(n_649),
.C(n_651),
.Y(n_693)
);

XOR2xp5_ASAP7_75t_L g692 ( 
.A(n_687),
.B(n_658),
.Y(n_692)
);

OAI21x1_ASAP7_75t_L g694 ( 
.A1(n_692),
.A2(n_689),
.B(n_688),
.Y(n_694)
);

AO21x1_ASAP7_75t_L g695 ( 
.A1(n_693),
.A2(n_694),
.B(n_690),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g696 ( 
.A1(n_695),
.A2(n_692),
.B(n_651),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_SL g697 ( 
.A(n_696),
.B(n_588),
.Y(n_697)
);

A2O1A1O1Ixp25_ASAP7_75t_L g698 ( 
.A1(n_697),
.A2(n_585),
.B(n_597),
.C(n_618),
.D(n_693),
.Y(n_698)
);


endmodule