module real_jpeg_35_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx2_ASAP7_75t_L g79 ( 
.A(n_0),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_1),
.B(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_1),
.B(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_1),
.B(n_27),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_1),
.B(n_39),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_1),
.B(n_77),
.Y(n_156)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_1),
.Y(n_163)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_2),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_2),
.B(n_45),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_2),
.B(n_77),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_2),
.B(n_49),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_2),
.B(n_105),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_2),
.B(n_36),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_4),
.B(n_27),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_4),
.B(n_39),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_4),
.B(n_45),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_4),
.B(n_32),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_4),
.B(n_49),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_4),
.B(n_77),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_4),
.B(n_105),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_4),
.B(n_36),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_5),
.B(n_32),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_5),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_5),
.B(n_27),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_5),
.B(n_39),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_5),
.B(n_45),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_10),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_10),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_10),
.B(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_10),
.B(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_10),
.B(n_36),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_10),
.B(n_105),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_10),
.B(n_77),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_10),
.B(n_49),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_11),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_39),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_11),
.B(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_11),
.B(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_11),
.B(n_77),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_11),
.B(n_105),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_12),
.B(n_27),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_12),
.B(n_32),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_12),
.B(n_39),
.Y(n_177)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_12),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_12),
.B(n_45),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_12),
.B(n_49),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_14),
.B(n_39),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_14),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_14),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_14),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_14),
.B(n_36),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_14),
.B(n_27),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_124),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_122),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_107),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_19),
.B(n_107),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_60),
.C(n_80),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_20),
.A2(n_21),
.B1(n_60),
.B2(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_42),
.B2(n_59),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_22),
.B(n_43),
.C(n_51),
.Y(n_109)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_25),
.B(n_31),
.C(n_34),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_25),
.A2(n_26),
.B1(n_332),
.B2(n_333),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_25),
.A2(n_26),
.B1(n_106),
.B2(n_359),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_26),
.B(n_100),
.C(n_106),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_26),
.B(n_330),
.C(n_333),
.Y(n_355)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_27),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.C(n_40),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_35),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_35),
.Y(n_97)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_36),
.Y(n_144)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_38),
.A2(n_40),
.B1(n_41),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_38),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_38),
.A2(n_96),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_38),
.B(n_296),
.C(n_300),
.Y(n_330)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_39),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_51),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.C(n_50),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_47),
.B1(n_48),
.B2(n_54),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_44),
.A2(n_54),
.B1(n_88),
.B2(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_44),
.B(n_88),
.C(n_142),
.Y(n_186)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_45),
.Y(n_297)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_SL g72 ( 
.A(n_47),
.B(n_73),
.C(n_75),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_48),
.B1(n_75),
.B2(n_76),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_47),
.A2(n_48),
.B1(n_167),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_48),
.B(n_167),
.C(n_168),
.Y(n_166)
);

INVx13_ASAP7_75t_L g191 ( 
.A(n_49),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_54),
.B(n_56),
.C(n_57),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_55),
.A2(n_56),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_55),
.A2(n_56),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_56),
.B(n_69),
.C(n_196),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_60),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.C(n_72),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_61),
.A2(n_62),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_64),
.B(n_72),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.C(n_70),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_65),
.A2(n_91),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_66),
.B(n_152),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_68),
.A2(n_69),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_74),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_75),
.A2(n_76),
.B1(n_206),
.B2(n_209),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_75),
.A2(n_76),
.B1(n_104),
.B2(n_230),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_102),
.C(n_104),
.Y(n_101)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_78),
.B(n_211),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_80),
.B(n_374),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_94),
.C(n_99),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_81),
.B(n_378),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.C(n_90),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_82),
.A2(n_83),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_86),
.B(n_90),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.C(n_89),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_87),
.B(n_89),
.Y(n_345)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_88),
.A2(n_146),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_94),
.B(n_99),
.Y(n_378)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_100),
.A2(n_101),
.B1(n_357),
.B2(n_358),
.Y(n_356)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_102),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_102),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_104),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_104),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_104),
.A2(n_134),
.B1(n_164),
.B2(n_230),
.Y(n_303)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_105),
.Y(n_162)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_106),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_121),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_119),
.A2(n_120),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_120),
.B(n_316),
.C(n_317),
.Y(n_328)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_371),
.B(n_386),
.Y(n_124)
);

OAI31xp33_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_320),
.A3(n_360),
.B(n_365),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_288),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_212),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_180),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_129),
.B(n_180),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_147),
.C(n_170),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_130),
.B(n_285),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g389 ( 
.A(n_130),
.Y(n_389)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_137),
.CI(n_141),
.CON(n_130),
.SN(n_130)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_131),
.B(n_137),
.C(n_141),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.C(n_136),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_132),
.A2(n_133),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g343 ( 
.A1(n_133),
.A2(n_164),
.B(n_230),
.C(n_304),
.Y(n_343)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_161),
.B1(n_164),
.B2(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_135),
.B(n_136),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B(n_140),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_139),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_140),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_140),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_143),
.B(n_162),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_143),
.B(n_191),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_144),
.B(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_147),
.B(n_170),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_158),
.B2(n_169),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_159),
.C(n_166),
.Y(n_182)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_150),
.B(n_155),
.C(n_157),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_154),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_165),
.B2(n_166),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.Y(n_160)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_163),
.B(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_167),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.C(n_178),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_171),
.B(n_174),
.CI(n_178),
.CON(n_275),
.SN(n_275)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.C(n_177),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_175),
.B(n_177),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_223),
.Y(n_222)
);

BUFx24_ASAP7_75t_SL g391 ( 
.A(n_180),
.Y(n_391)
);

FAx1_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_198),
.CI(n_199),
.CON(n_180),
.SN(n_180)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_181),
.B(n_198),
.C(n_199),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_182),
.B(n_185),
.C(n_192),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_192),
.B2(n_193),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_186),
.B(n_188),
.C(n_190),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_196),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_201),
.B(n_202),
.C(n_204),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_210),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_206),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_206),
.B(n_208),
.C(n_210),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_283),
.B(n_287),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_271),
.B(n_282),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_243),
.B(n_270),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_234),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_216),
.B(n_234),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_226),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_218),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.C(n_221),
.Y(n_218)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_219),
.B(n_220),
.CI(n_221),
.CON(n_235),
.SN(n_235)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_222),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_222),
.B(n_224),
.C(n_226),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_227),
.B(n_232),
.C(n_233),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.C(n_242),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_267),
.Y(n_266)
);

BUFx24_ASAP7_75t_SL g395 ( 
.A(n_235),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_236),
.A2(n_237),
.B1(n_242),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_242),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_264),
.B(n_269),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_255),
.B(n_263),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_251),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_251),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_249),
.C(n_250),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_258),
.B(n_262),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_260),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_272),
.B(n_273),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_278),
.C(n_279),
.Y(n_286)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx24_ASAP7_75t_SL g396 ( 
.A(n_275),
.Y(n_396)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_286),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_289),
.A2(n_367),
.B(n_368),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_319),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_290),
.B(n_319),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_291),
.B(n_293),
.C(n_306),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_305),
.B2(n_306),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx24_ASAP7_75t_SL g390 ( 
.A(n_294),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_301),
.CI(n_302),
.CON(n_294),
.SN(n_294)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_295),
.B(n_301),
.C(n_302),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_311),
.C(n_312),
.Y(n_335)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_317),
.B2(n_318),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g365 ( 
.A1(n_321),
.A2(n_361),
.B(n_366),
.C(n_369),
.D(n_370),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_347),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_322),
.B(n_347),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_335),
.C(n_336),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_323),
.A2(n_324),
.B1(n_336),
.B2(n_337),
.Y(n_363)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_334),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_328),
.C(n_329),
.Y(n_348)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_327),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_332),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_335),
.B(n_363),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_342),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_343),
.C(n_344),
.Y(n_354)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_339),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_345),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_348),
.B(n_350),
.C(n_353),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_353),
.Y(n_349)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_351),
.Y(n_352)
);

BUFx24_ASAP7_75t_SL g393 ( 
.A(n_353),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_355),
.CI(n_356),
.CON(n_353),
.SN(n_353)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_354),
.B(n_355),
.C(n_356),
.Y(n_382)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_364),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_362),
.B(n_364),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_383),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_372),
.A2(n_387),
.B(n_388),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_376),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_373),
.B(n_376),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_379),
.C(n_382),
.Y(n_376)
);

FAx1_ASAP7_75t_SL g384 ( 
.A(n_377),
.B(n_379),
.CI(n_382),
.CON(n_384),
.SN(n_384)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_380),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_385),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_384),
.B(n_385),
.Y(n_387)
);

BUFx24_ASAP7_75t_SL g394 ( 
.A(n_384),
.Y(n_394)
);


endmodule