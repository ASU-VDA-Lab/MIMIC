module fake_ariane_533_n_2347 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_236, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_232, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_2347);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_236;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2347;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_899;
wire n_352;
wire n_1703;
wire n_2332;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_851;
wire n_355;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_274;
wire n_337;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_2294;
wire n_2274;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_347;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_552;
wire n_348;
wire n_2312;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_2336;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_48),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_198),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_19),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_28),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_78),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_82),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_29),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_14),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_168),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_178),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_53),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_110),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_63),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_218),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_137),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_174),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_12),
.Y(n_254)
);

BUFx2_ASAP7_75t_SL g255 ( 
.A(n_24),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_8),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_6),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_195),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_10),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_64),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_40),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_139),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_200),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_134),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_155),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_98),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_62),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_150),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_25),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_33),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_235),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_76),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_30),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_213),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_17),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_84),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_109),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_38),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_94),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_54),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_180),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_183),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_113),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_175),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_133),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_166),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_189),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_31),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_78),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_86),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_234),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_81),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_22),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_69),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_35),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_225),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_77),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_32),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_17),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_89),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_227),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_32),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_128),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_184),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_63),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_96),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_64),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_104),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_203),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_136),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_52),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_27),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_40),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_199),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_25),
.Y(n_316)
);

BUFx10_ASAP7_75t_L g317 ( 
.A(n_173),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_95),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_147),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_138),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_18),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_62),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_43),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_204),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_172),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_161),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_46),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_219),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_162),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_217),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_226),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_41),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_192),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_24),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_158),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_41),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_170),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_237),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_70),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_74),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_12),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_57),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_118),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_38),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_206),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_107),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_59),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_165),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_117),
.Y(n_349)
);

BUFx5_ASAP7_75t_L g350 ( 
.A(n_181),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_152),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_169),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_21),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_11),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_2),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_222),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_5),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_61),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_69),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_72),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_119),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_61),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_22),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_39),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_127),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_211),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_126),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_132),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_20),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_79),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_221),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_229),
.Y(n_372)
);

BUFx2_ASAP7_75t_SL g373 ( 
.A(n_20),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_99),
.Y(n_374)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_66),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_45),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_11),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_72),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_231),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_34),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_56),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_97),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_45),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_51),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_46),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_146),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_71),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_43),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_35),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_185),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_232),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_18),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_3),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_190),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_33),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_236),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_210),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_10),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_39),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_34),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_135),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_75),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_156),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_103),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_93),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_102),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_108),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_116),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_197),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_55),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_124),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_160),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_149),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_106),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_5),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_21),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_80),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_58),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_67),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_191),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_153),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_23),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_57),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_105),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_66),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_111),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_55),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_74),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_123),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_59),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_194),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_121),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_145),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_16),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_85),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_75),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_125),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_7),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_115),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_122),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_193),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_51),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_14),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_53),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_48),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_26),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_29),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_212),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_224),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_2),
.Y(n_450)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_15),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_49),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_209),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_19),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_31),
.Y(n_455)
);

BUFx2_ASAP7_75t_SL g456 ( 
.A(n_52),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_216),
.Y(n_457)
);

BUFx10_ASAP7_75t_L g458 ( 
.A(n_1),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_73),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_27),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_228),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_171),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_164),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_214),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_77),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_308),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_344),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_344),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_451),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_285),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_243),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_285),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_285),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_358),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_317),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_317),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_245),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_307),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_261),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_317),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_329),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_405),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_279),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_440),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_316),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_239),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_239),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_339),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_342),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_387),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_286),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_257),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_353),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_246),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_300),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_357),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_300),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_290),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_298),
.Y(n_499)
);

CKINVDCx14_ASAP7_75t_R g500 ( 
.A(n_295),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_336),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_362),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_364),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_376),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_381),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_385),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_434),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_294),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_380),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_299),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_415),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_399),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_240),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_303),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_459),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_286),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_410),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_295),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_423),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_312),
.B(n_0),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_428),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_306),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_R g523 ( 
.A(n_291),
.B(n_83),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_313),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_445),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_314),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_246),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_247),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_447),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_271),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_271),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_360),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_300),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_391),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_360),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_247),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_363),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_391),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_448),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_251),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_363),
.Y(n_541)
);

INVxp67_ASAP7_75t_SL g542 ( 
.A(n_300),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_402),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_402),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_356),
.B(n_0),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_251),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_253),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_273),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_448),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_295),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_253),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_259),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_273),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_296),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_340),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_296),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_259),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_300),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_340),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_263),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_263),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_255),
.Y(n_562)
);

NOR2xp67_ASAP7_75t_L g563 ( 
.A(n_248),
.B(n_1),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_392),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_392),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_266),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_392),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_392),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_340),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_392),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_375),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_373),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_375),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_375),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_266),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_458),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_456),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_275),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_238),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_275),
.Y(n_580)
);

INVxp33_ASAP7_75t_SL g581 ( 
.A(n_238),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_278),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_458),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_458),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_278),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_249),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_284),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_252),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_256),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_264),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_241),
.Y(n_591)
);

INVxp33_ASAP7_75t_SL g592 ( 
.A(n_241),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_284),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_287),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_495),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_495),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_558),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_564),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_497),
.B(n_265),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_586),
.B(n_411),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_565),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_567),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_568),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_471),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_570),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_466),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_530),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_533),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_491),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_542),
.B(n_267),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_491),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_588),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_531),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_474),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_532),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_523),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_589),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_535),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_590),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g620 ( 
.A(n_492),
.B(n_499),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_537),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_541),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_543),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_467),
.B(n_411),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_544),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_477),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_479),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_483),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_485),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_468),
.B(n_272),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_488),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_489),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_493),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_496),
.Y(n_634)
);

CKINVDCx16_ASAP7_75t_R g635 ( 
.A(n_518),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_502),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_505),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_591),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_506),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_512),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_517),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_490),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_519),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_521),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_525),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_529),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_548),
.B(n_277),
.Y(n_647)
);

OA21x2_ASAP7_75t_L g648 ( 
.A1(n_553),
.A2(n_346),
.B(n_305),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_554),
.Y(n_649)
);

INVx5_ASAP7_75t_L g650 ( 
.A(n_498),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_556),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_571),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_470),
.B(n_305),
.Y(n_653)
);

INVx5_ASAP7_75t_L g654 ( 
.A(n_500),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_563),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_573),
.B(n_280),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_545),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_574),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_576),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_486),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_520),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_486),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_516),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_562),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_572),
.B(n_282),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_577),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_487),
.B(n_283),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_534),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_579),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_487),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_513),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_538),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_539),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_494),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_507),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_469),
.B(n_287),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_470),
.B(n_292),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_501),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_549),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_472),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_494),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_594),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_594),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_472),
.B(n_346),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_593),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_593),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_473),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_527),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_469),
.B(n_288),
.Y(n_689)
);

INVx4_ASAP7_75t_L g690 ( 
.A(n_527),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_528),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_473),
.B(n_288),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_475),
.B(n_293),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_651),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_680),
.B(n_528),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_681),
.B(n_536),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_601),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_601),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_650),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_661),
.B(n_475),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_597),
.Y(n_701)
);

INVx4_ASAP7_75t_L g702 ( 
.A(n_654),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_661),
.B(n_476),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_680),
.B(n_536),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_609),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_624),
.B(n_476),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_680),
.B(n_540),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_651),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_680),
.B(n_540),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_597),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_601),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_601),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_604),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_609),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_597),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_601),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_602),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_620),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_609),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_609),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_598),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_680),
.B(n_546),
.Y(n_722)
);

INVxp33_ASAP7_75t_L g723 ( 
.A(n_606),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_681),
.B(n_688),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_602),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_602),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_609),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_598),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_603),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_603),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_606),
.B(n_614),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_598),
.Y(n_732)
);

BUFx4f_ASAP7_75t_L g733 ( 
.A(n_680),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_609),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_603),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_651),
.Y(n_736)
);

NAND3xp33_ASAP7_75t_L g737 ( 
.A(n_667),
.B(n_547),
.C(n_546),
.Y(n_737)
);

AND2x6_ASAP7_75t_L g738 ( 
.A(n_680),
.B(n_687),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_SL g739 ( 
.A(n_635),
.B(n_581),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_608),
.Y(n_740)
);

INVxp33_ASAP7_75t_L g741 ( 
.A(n_614),
.Y(n_741)
);

OAI22xp33_ASAP7_75t_L g742 ( 
.A1(n_669),
.A2(n_581),
.B1(n_592),
.B2(n_480),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_609),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_598),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_680),
.B(n_547),
.Y(n_745)
);

INVx4_ASAP7_75t_L g746 ( 
.A(n_654),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_654),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_680),
.B(n_551),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_687),
.B(n_551),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_596),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_681),
.B(n_552),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_608),
.Y(n_752)
);

BUFx6f_ASAP7_75t_SL g753 ( 
.A(n_687),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_661),
.B(n_480),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_609),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_687),
.B(n_552),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_609),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_629),
.Y(n_758)
);

AO22x2_ASAP7_75t_L g759 ( 
.A1(n_657),
.A2(n_383),
.B1(n_250),
.B2(n_368),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_667),
.A2(n_592),
.B1(n_560),
.B2(n_561),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_608),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_629),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_SL g763 ( 
.A1(n_660),
.A2(n_555),
.B1(n_559),
.B2(n_550),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_596),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_654),
.Y(n_765)
);

NAND3xp33_ASAP7_75t_L g766 ( 
.A(n_666),
.B(n_560),
.C(n_557),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_612),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_596),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_664),
.B(n_557),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_624),
.B(n_681),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_650),
.Y(n_771)
);

CKINVDCx6p67_ASAP7_75t_R g772 ( 
.A(n_635),
.Y(n_772)
);

XOR2xp5_ASAP7_75t_L g773 ( 
.A(n_620),
.B(n_478),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_605),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_595),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_605),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_605),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_642),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_595),
.Y(n_779)
);

INVx4_ASAP7_75t_L g780 ( 
.A(n_654),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_612),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_657),
.A2(n_575),
.B1(n_578),
.B2(n_566),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_595),
.Y(n_783)
);

CKINVDCx6p67_ASAP7_75t_R g784 ( 
.A(n_650),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_595),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_657),
.A2(n_575),
.B1(n_578),
.B2(n_566),
.Y(n_786)
);

INVx4_ASAP7_75t_L g787 ( 
.A(n_654),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_664),
.B(n_580),
.Y(n_788)
);

NOR2x1p5_ASAP7_75t_L g789 ( 
.A(n_671),
.B(n_508),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_650),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_687),
.B(n_580),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_687),
.B(n_582),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_629),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_595),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_653),
.A2(n_585),
.B1(n_587),
.B2(n_582),
.Y(n_795)
);

AND2x6_ASAP7_75t_L g796 ( 
.A(n_687),
.B(n_269),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_607),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_612),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_687),
.B(n_585),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_664),
.B(n_587),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_624),
.A2(n_652),
.B1(n_684),
.B2(n_653),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_617),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_617),
.Y(n_803)
);

AO22x2_ASAP7_75t_L g804 ( 
.A1(n_684),
.A2(n_318),
.B1(n_309),
.B2(n_302),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_629),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_687),
.B(n_510),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_629),
.Y(n_807)
);

INVxp33_ASAP7_75t_SL g808 ( 
.A(n_678),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_617),
.Y(n_809)
);

AND2x6_ASAP7_75t_L g810 ( 
.A(n_688),
.B(n_269),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_607),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_674),
.B(n_514),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_654),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_619),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_624),
.B(n_522),
.Y(n_815)
);

OR2x2_ASAP7_75t_L g816 ( 
.A(n_642),
.B(n_675),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_619),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_654),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_688),
.B(n_524),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_624),
.A2(n_526),
.B1(n_454),
.B2(n_569),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_607),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_607),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_619),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_688),
.B(n_583),
.Y(n_824)
);

XOR2x2_ASAP7_75t_L g825 ( 
.A(n_620),
.B(n_503),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_627),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_615),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_627),
.Y(n_828)
);

NAND3xp33_ASAP7_75t_SL g829 ( 
.A(n_692),
.B(n_244),
.C(n_242),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_624),
.B(n_426),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_615),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_648),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_615),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_650),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_648),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_650),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_675),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_654),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_652),
.B(n_426),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_652),
.B(n_429),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_627),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_682),
.A2(n_322),
.B1(n_323),
.B2(n_321),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_691),
.B(n_584),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_650),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_615),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_682),
.A2(n_685),
.B1(n_686),
.B2(n_683),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_618),
.Y(n_847)
);

CKINVDCx6p67_ASAP7_75t_R g848 ( 
.A(n_650),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_629),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_691),
.B(n_481),
.Y(n_850)
);

OR2x6_ASAP7_75t_L g851 ( 
.A(n_691),
.B(n_326),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_652),
.B(n_429),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_629),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_666),
.B(n_433),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_600),
.B(n_242),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_638),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_733),
.B(n_660),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_701),
.Y(n_858)
);

NOR3xp33_ASAP7_75t_L g859 ( 
.A(n_742),
.B(n_662),
.C(n_660),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_721),
.Y(n_860)
);

INVxp67_ASAP7_75t_SL g861 ( 
.A(n_770),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_696),
.B(n_660),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_733),
.B(n_660),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_706),
.B(n_650),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_700),
.A2(n_691),
.B1(n_670),
.B2(n_662),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_837),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_701),
.Y(n_867)
);

NOR2xp67_ASAP7_75t_L g868 ( 
.A(n_760),
.B(n_678),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_837),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_728),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_710),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_733),
.B(n_770),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_751),
.B(n_662),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_819),
.B(n_662),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_724),
.B(n_662),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_731),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_770),
.B(n_670),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_731),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_728),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_706),
.B(n_670),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_804),
.A2(n_655),
.B1(n_683),
.B2(n_682),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_710),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_846),
.A2(n_685),
.B1(n_686),
.B2(n_683),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_801),
.B(n_670),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_856),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_703),
.B(n_670),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_715),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_706),
.B(n_674),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_754),
.B(n_685),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_815),
.B(n_674),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_793),
.B(n_674),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_715),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_793),
.B(n_674),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_793),
.B(n_674),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_732),
.Y(n_895)
);

OAI221xp5_ASAP7_75t_L g896 ( 
.A1(n_842),
.A2(n_665),
.B1(n_630),
.B2(n_656),
.C(n_693),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_816),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_717),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_772),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_718),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_732),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_717),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_737),
.B(n_686),
.Y(n_903)
);

NAND3xp33_ASAP7_75t_L g904 ( 
.A(n_782),
.B(n_690),
.C(n_692),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_769),
.B(n_690),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_816),
.B(n_663),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_788),
.B(n_690),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_800),
.B(n_690),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_725),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_740),
.B(n_690),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_725),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_723),
.B(n_692),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_786),
.A2(n_677),
.B1(n_693),
.B2(n_669),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_789),
.B(n_658),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_744),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_744),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_726),
.Y(n_917)
);

NOR3xp33_ASAP7_75t_SL g918 ( 
.A(n_829),
.B(n_254),
.C(n_244),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_797),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_726),
.Y(n_920)
);

NAND2xp33_ASAP7_75t_L g921 ( 
.A(n_738),
.B(n_658),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_729),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_797),
.Y(n_923)
);

O2A1O1Ixp5_ASAP7_75t_L g924 ( 
.A1(n_695),
.A2(n_677),
.B(n_628),
.C(n_634),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_811),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_752),
.B(n_666),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_772),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_723),
.B(n_741),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_811),
.Y(n_929)
);

NAND2xp33_ASAP7_75t_SL g930 ( 
.A(n_753),
.B(n_658),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_697),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_729),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_850),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_761),
.B(n_665),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_793),
.B(n_658),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_821),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_793),
.B(n_658),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_821),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_822),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_713),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_741),
.B(n_669),
.Y(n_941)
);

NAND2xp33_ASAP7_75t_L g942 ( 
.A(n_738),
.B(n_658),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_778),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_830),
.B(n_600),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_824),
.B(n_689),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_822),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_730),
.Y(n_947)
);

OR2x2_ASAP7_75t_SL g948 ( 
.A(n_825),
.B(n_671),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_827),
.Y(n_949)
);

BUFx5_ASAP7_75t_L g950 ( 
.A(n_738),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_843),
.B(n_689),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_807),
.B(n_658),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_739),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_827),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_831),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_720),
.Y(n_956)
);

BUFx6f_ASAP7_75t_SL g957 ( 
.A(n_851),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_767),
.A2(n_628),
.B(n_634),
.C(n_626),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_730),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_831),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_697),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_694),
.B(n_600),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_708),
.B(n_658),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_735),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_736),
.B(n_658),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_735),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_781),
.B(n_659),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_807),
.B(n_659),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_798),
.B(n_659),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_833),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_802),
.B(n_659),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_807),
.B(n_659),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_795),
.B(n_808),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_807),
.B(n_659),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_804),
.A2(n_655),
.B1(n_648),
.B2(n_659),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_807),
.B(n_659),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_849),
.B(n_659),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_713),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_774),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_774),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_803),
.B(n_630),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_833),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_849),
.B(n_698),
.Y(n_983)
);

NAND2xp33_ASAP7_75t_L g984 ( 
.A(n_738),
.B(n_616),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_776),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_845),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_776),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_809),
.B(n_626),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_845),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_855),
.B(n_671),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_849),
.B(n_616),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_814),
.B(n_626),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_855),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_817),
.B(n_626),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_823),
.B(n_626),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_714),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_718),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_808),
.B(n_689),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_820),
.B(n_668),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_854),
.B(n_628),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_847),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_851),
.B(n_628),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_777),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_704),
.A2(n_647),
.B(n_628),
.C(n_636),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_851),
.A2(n_676),
.B1(n_655),
.B2(n_656),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_804),
.A2(n_648),
.B1(n_629),
.B2(n_631),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_773),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_784),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_847),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_777),
.Y(n_1010)
);

OR2x6_ASAP7_75t_L g1011 ( 
.A(n_759),
.B(n_672),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_750),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_851),
.A2(n_676),
.B1(n_634),
.B2(n_637),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_698),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_812),
.B(n_839),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_750),
.Y(n_1016)
);

OR2x6_ASAP7_75t_L g1017 ( 
.A(n_804),
.B(n_672),
.Y(n_1017)
);

OR2x6_ASAP7_75t_L g1018 ( 
.A(n_759),
.B(n_672),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_766),
.B(n_634),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_849),
.B(n_616),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_849),
.B(n_616),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_759),
.B(n_668),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_806),
.B(n_676),
.Y(n_1023)
);

NAND2x1p5_ASAP7_75t_L g1024 ( 
.A(n_699),
.B(n_611),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_764),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_840),
.B(n_634),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_707),
.B(n_663),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_SL g1028 ( 
.A(n_773),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_973),
.A2(n_945),
.B1(n_951),
.B2(n_861),
.Y(n_1029)
);

AOI22x1_ASAP7_75t_L g1030 ( 
.A1(n_858),
.A2(n_711),
.B1(n_716),
.B2(n_712),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_874),
.A2(n_709),
.B1(n_745),
.B2(n_722),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_933),
.A2(n_998),
.B1(n_889),
.B2(n_912),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_867),
.B(n_826),
.Y(n_1033)
);

NOR3xp33_ASAP7_75t_L g1034 ( 
.A(n_978),
.B(n_638),
.C(n_763),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_864),
.B(n_883),
.Y(n_1035)
);

AO21x1_ASAP7_75t_L g1036 ( 
.A1(n_862),
.A2(n_749),
.B(n_748),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_871),
.B(n_828),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_869),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_882),
.B(n_841),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_887),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_875),
.A2(n_791),
.B(n_756),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_864),
.B(n_792),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_857),
.A2(n_799),
.B(n_753),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_958),
.A2(n_835),
.B(n_832),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_857),
.A2(n_753),
.B(n_746),
.Y(n_1045)
);

NAND2x1p5_ASAP7_75t_L g1046 ( 
.A(n_864),
.B(n_672),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_906),
.B(n_482),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_958),
.A2(n_835),
.B(n_832),
.Y(n_1048)
);

OAI22x1_ASAP7_75t_L g1049 ( 
.A1(n_997),
.A2(n_638),
.B1(n_825),
.B2(n_673),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_863),
.A2(n_746),
.B(n_702),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_913),
.A2(n_852),
.B(n_636),
.C(n_637),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_885),
.B(n_484),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_924),
.A2(n_719),
.B(n_705),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_863),
.A2(n_746),
.B(n_702),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_860),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_873),
.A2(n_747),
.B(n_702),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_899),
.B(n_668),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_892),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_896),
.A2(n_636),
.B(n_637),
.C(n_711),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_983),
.A2(n_780),
.B(n_747),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_876),
.B(n_668),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_878),
.B(n_673),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1004),
.A2(n_716),
.B(n_712),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_898),
.B(n_764),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_866),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_902),
.B(n_768),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_909),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_983),
.A2(n_780),
.B(n_747),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_905),
.A2(n_787),
.B(n_780),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_877),
.A2(n_848),
.B1(n_784),
.B2(n_771),
.Y(n_1070)
);

BUFx12f_ASAP7_75t_L g1071 ( 
.A(n_899),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_911),
.B(n_768),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_1026),
.A2(n_762),
.B(n_758),
.Y(n_1073)
);

AOI21xp33_ASAP7_75t_L g1074 ( 
.A1(n_881),
.A2(n_1017),
.B(n_884),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_917),
.B(n_738),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_920),
.B(n_738),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1000),
.A2(n_762),
.B(n_758),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_907),
.A2(n_787),
.B(n_699),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_908),
.A2(n_834),
.B(n_790),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_1008),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_886),
.A2(n_834),
.B(n_790),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_940),
.Y(n_1082)
);

O2A1O1Ixp5_ASAP7_75t_L g1083 ( 
.A1(n_890),
.A2(n_853),
.B(n_762),
.C(n_805),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_963),
.A2(n_805),
.B(n_758),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_927),
.B(n_673),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_903),
.A2(n_759),
.B1(n_679),
.B2(n_673),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_922),
.B(n_636),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_890),
.A2(n_844),
.B(n_836),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_897),
.B(n_679),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_910),
.A2(n_844),
.B(n_836),
.Y(n_1090)
);

INVx4_ASAP7_75t_L g1091 ( 
.A(n_927),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_932),
.B(n_636),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_928),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1015),
.A2(n_719),
.B(n_705),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_947),
.B(n_637),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_891),
.A2(n_719),
.B(n_705),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_959),
.B(n_637),
.Y(n_1097)
);

INVx4_ASAP7_75t_L g1098 ( 
.A(n_957),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_964),
.B(n_805),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_891),
.A2(n_853),
.B(n_813),
.Y(n_1100)
);

CKINVDCx6p67_ASAP7_75t_R g1101 ( 
.A(n_940),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_966),
.B(n_853),
.Y(n_1102)
);

OR2x2_ASAP7_75t_L g1103 ( 
.A(n_1007),
.B(n_679),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_893),
.A2(n_813),
.B(n_765),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_941),
.B(n_679),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_893),
.A2(n_818),
.B(n_765),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_957),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_953),
.B(n_504),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_894),
.A2(n_838),
.B(n_818),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_965),
.A2(n_779),
.B(n_775),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_943),
.Y(n_1111)
);

AO21x1_ASAP7_75t_L g1112 ( 
.A1(n_865),
.A2(n_366),
.B(n_328),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_993),
.B(n_632),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_967),
.A2(n_779),
.B(n_775),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_894),
.A2(n_838),
.B(n_727),
.Y(n_1115)
);

BUFx4f_ASAP7_75t_L g1116 ( 
.A(n_914),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_870),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_984),
.A2(n_727),
.B(n_714),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_969),
.A2(n_785),
.B(n_783),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_859),
.B(n_616),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_1027),
.B(n_509),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_984),
.A2(n_743),
.B(n_734),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_971),
.A2(n_743),
.B(n_734),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_979),
.B(n_783),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_980),
.B(n_785),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_1008),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_868),
.B(n_616),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_921),
.A2(n_942),
.B(n_988),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_985),
.A2(n_1003),
.B1(n_1010),
.B2(n_987),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_934),
.B(n_794),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_900),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_981),
.B(n_794),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_921),
.A2(n_755),
.B(n_720),
.Y(n_1133)
);

NOR2x1p5_ASAP7_75t_SL g1134 ( 
.A(n_950),
.B(n_350),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_942),
.A2(n_755),
.B(n_720),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_900),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1005),
.B(n_616),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_992),
.A2(n_796),
.B(n_648),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1013),
.A2(n_848),
.B1(n_258),
.B2(n_260),
.Y(n_1139)
);

OAI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1017),
.A2(n_904),
.B1(n_1018),
.B2(n_1011),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_956),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_944),
.A2(n_258),
.B1(n_260),
.B2(n_254),
.Y(n_1142)
);

NAND2xp33_ASAP7_75t_L g1143 ( 
.A(n_950),
.B(n_796),
.Y(n_1143)
);

NAND2x1p5_ASAP7_75t_L g1144 ( 
.A(n_1008),
.B(n_613),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_880),
.B(n_511),
.Y(n_1145)
);

AO21x1_ASAP7_75t_L g1146 ( 
.A1(n_930),
.A2(n_386),
.B(n_371),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_990),
.B(n_515),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_994),
.A2(n_757),
.B(n_720),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1023),
.A2(n_599),
.B(n_610),
.C(n_632),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_995),
.A2(n_757),
.B(n_720),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_935),
.A2(n_757),
.B(n_616),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_935),
.A2(n_757),
.B(n_616),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_962),
.A2(n_268),
.B1(n_270),
.B2(n_262),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1016),
.B(n_599),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1016),
.B(n_1019),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_870),
.Y(n_1156)
);

INVxp67_ASAP7_75t_L g1157 ( 
.A(n_999),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_937),
.A2(n_796),
.B(n_648),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_956),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_880),
.A2(n_268),
.B1(n_270),
.B2(n_262),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_888),
.A2(n_643),
.B(n_644),
.C(n_632),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_937),
.A2(n_968),
.B(n_952),
.Y(n_1162)
);

BUFx4f_ASAP7_75t_L g1163 ( 
.A(n_914),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1012),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_888),
.A2(n_274),
.B1(n_281),
.B2(n_276),
.Y(n_1165)
);

AO21x1_ASAP7_75t_L g1166 ( 
.A1(n_930),
.A2(n_401),
.B(n_390),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_914),
.Y(n_1167)
);

INVxp67_ASAP7_75t_L g1168 ( 
.A(n_1028),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_879),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_948),
.B(n_643),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1019),
.B(n_610),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_952),
.A2(n_757),
.B(n_647),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1017),
.A2(n_810),
.B1(n_796),
.B2(n_643),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_968),
.A2(n_631),
.B(n_627),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1019),
.B(n_796),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_931),
.B(n_796),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_926),
.B(n_644),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1017),
.B(n_644),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_972),
.A2(n_335),
.B(n_645),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_956),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_972),
.A2(n_646),
.B(n_645),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1025),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_974),
.A2(n_646),
.B(n_645),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_974),
.A2(n_646),
.B(n_649),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1011),
.B(n_631),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_976),
.A2(n_649),
.B(n_633),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_976),
.A2(n_649),
.B(n_633),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_879),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_977),
.A2(n_649),
.B(n_633),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1002),
.A2(n_633),
.B(n_641),
.C(n_640),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_950),
.B(n_629),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1011),
.B(n_631),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_977),
.A2(n_640),
.B(n_639),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_872),
.A2(n_640),
.B(n_639),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_872),
.A2(n_1020),
.B(n_991),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_991),
.A2(n_640),
.B(n_639),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_931),
.A2(n_961),
.B1(n_1014),
.B2(n_956),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_950),
.B(n_433),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_895),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1020),
.A2(n_641),
.B(n_639),
.Y(n_1200)
);

INVx1_ASAP7_75t_SL g1201 ( 
.A(n_1022),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1018),
.B(n_641),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_996),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1021),
.A2(n_961),
.B(n_931),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_996),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_961),
.A2(n_810),
.B(n_641),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1014),
.B(n_895),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1014),
.A2(n_810),
.B(n_625),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_918),
.A2(n_621),
.B(n_613),
.C(n_622),
.Y(n_1209)
);

BUFx24_ASAP7_75t_L g1210 ( 
.A(n_1028),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_901),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_950),
.B(n_439),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1021),
.A2(n_441),
.B(n_439),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1018),
.B(n_901),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_915),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_915),
.A2(n_810),
.B(n_625),
.Y(n_1216)
);

O2A1O1Ixp5_ASAP7_75t_L g1217 ( 
.A1(n_916),
.A2(n_613),
.B(n_621),
.C(n_622),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_916),
.A2(n_453),
.B(n_441),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_919),
.A2(n_461),
.B(n_453),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1029),
.A2(n_975),
.B(n_1006),
.C(n_923),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1032),
.A2(n_923),
.B(n_925),
.C(n_919),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1128),
.A2(n_950),
.B(n_929),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_SL g1223 ( 
.A1(n_1121),
.A2(n_274),
.B1(n_281),
.B2(n_276),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1056),
.A2(n_950),
.B(n_929),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1203),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1116),
.B(n_925),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1177),
.B(n_936),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1069),
.A2(n_938),
.B(n_936),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1055),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1080),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1116),
.B(n_938),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1052),
.B(n_939),
.Y(n_1232)
);

BUFx12f_ASAP7_75t_L g1233 ( 
.A(n_1071),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1130),
.B(n_946),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1047),
.A2(n_810),
.B1(n_327),
.B2(n_332),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1038),
.B(n_946),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1040),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1130),
.B(n_949),
.Y(n_1238)
);

AOI222xp33_ASAP7_75t_L g1239 ( 
.A1(n_1147),
.A2(n_289),
.B1(n_422),
.B2(n_425),
.C1(n_427),
.C2(n_430),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_SL g1240 ( 
.A(n_1163),
.B(n_810),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1082),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1065),
.B(n_1111),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1058),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1145),
.B(n_949),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1142),
.A2(n_621),
.B(n_613),
.C(n_622),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1203),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1203),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1105),
.B(n_954),
.Y(n_1248)
);

NAND3xp33_ASAP7_75t_L g1249 ( 
.A(n_1059),
.B(n_1034),
.C(n_1149),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1157),
.B(n_954),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1136),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1067),
.A2(n_613),
.B1(n_621),
.B2(n_1001),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1164),
.Y(n_1253)
);

NAND3xp33_ASAP7_75t_SL g1254 ( 
.A(n_1131),
.B(n_422),
.C(n_289),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1171),
.B(n_955),
.Y(n_1255)
);

INVx2_ASAP7_75t_SL g1256 ( 
.A(n_1101),
.Y(n_1256)
);

A2O1A1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_1178),
.A2(n_986),
.B(n_1009),
.C(n_1001),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1061),
.B(n_621),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1062),
.B(n_625),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1080),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1161),
.A2(n_955),
.B(n_1009),
.C(n_989),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1093),
.B(n_960),
.Y(n_1262)
);

NAND3xp33_ASAP7_75t_L g1263 ( 
.A(n_1209),
.B(n_341),
.C(n_334),
.Y(n_1263)
);

AOI21xp33_ASAP7_75t_L g1264 ( 
.A1(n_1086),
.A2(n_982),
.B(n_970),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1057),
.B(n_982),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1141),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1091),
.B(n_986),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_1103),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1057),
.B(n_1085),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1089),
.Y(n_1270)
);

NAND3xp33_ASAP7_75t_SL g1271 ( 
.A(n_1153),
.B(n_427),
.C(n_425),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1141),
.Y(n_1272)
);

NOR3xp33_ASAP7_75t_SL g1273 ( 
.A(n_1165),
.B(n_436),
.C(n_430),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1170),
.B(n_1108),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1046),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1091),
.B(n_989),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1113),
.B(n_618),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1129),
.A2(n_618),
.B(n_623),
.C(n_414),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1046),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1113),
.B(n_618),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1035),
.A2(n_432),
.B(n_457),
.C(n_409),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1139),
.A2(n_1160),
.B(n_1031),
.C(n_1051),
.Y(n_1282)
);

AND2x2_ASAP7_75t_SL g1283 ( 
.A(n_1098),
.B(n_413),
.Y(n_1283)
);

AO21x2_ASAP7_75t_L g1284 ( 
.A1(n_1074),
.A2(n_623),
.B(n_431),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1182),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1085),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1168),
.B(n_436),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1064),
.A2(n_442),
.B1(n_450),
.B2(n_465),
.Y(n_1288)
);

AO22x2_ASAP7_75t_L g1289 ( 
.A1(n_1202),
.A2(n_623),
.B1(n_424),
.B2(n_435),
.Y(n_1289)
);

A2O1A1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1195),
.A2(n_437),
.B(n_449),
.C(n_623),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1117),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1171),
.B(n_438),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1205),
.B(n_1024),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1124),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1156),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1169),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1098),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1185),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1036),
.A2(n_1112),
.A3(n_1166),
.B(n_1146),
.Y(n_1299)
);

AOI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1120),
.A2(n_1024),
.B(n_350),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1124),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_1214),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1078),
.A2(n_301),
.B(n_297),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1064),
.A2(n_438),
.B1(n_442),
.B2(n_443),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1107),
.B(n_443),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1205),
.B(n_611),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1167),
.B(n_611),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1126),
.B(n_611),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1125),
.Y(n_1309)
);

NOR3xp33_ASAP7_75t_SL g1310 ( 
.A(n_1087),
.B(n_446),
.C(n_444),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1188),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1125),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1192),
.Y(n_1313)
);

NOR2x1_ASAP7_75t_L g1314 ( 
.A(n_1107),
.B(n_269),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1126),
.B(n_611),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1199),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1132),
.A2(n_310),
.B(n_304),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1132),
.B(n_444),
.Y(n_1318)
);

NOR2xp67_ASAP7_75t_L g1319 ( 
.A(n_1049),
.B(n_611),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1210),
.A2(n_1201),
.B1(n_1140),
.B2(n_1155),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1148),
.A2(n_319),
.B(n_311),
.Y(n_1321)
);

O2A1O1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1190),
.A2(n_1072),
.B(n_1066),
.C(n_1087),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1127),
.B(n_446),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1066),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1141),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1154),
.B(n_450),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1159),
.B(n_1180),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1072),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1215),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1042),
.B(n_1211),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1154),
.B(n_611),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1150),
.A2(n_324),
.B(n_320),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1079),
.A2(n_330),
.B(n_325),
.Y(n_1333)
);

BUFx6f_ASAP7_75t_L g1334 ( 
.A(n_1159),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1033),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1094),
.A2(n_333),
.B(n_331),
.Y(n_1336)
);

AOI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1041),
.A2(n_350),
.B(n_611),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1143),
.A2(n_338),
.B(n_337),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1033),
.A2(n_452),
.B1(n_455),
.B2(n_460),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_1159),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1081),
.A2(n_345),
.B(n_343),
.Y(n_1341)
);

O2A1O1Ixp5_ASAP7_75t_SL g1342 ( 
.A1(n_1074),
.A2(n_350),
.B(n_465),
.C(n_452),
.Y(n_1342)
);

NOR3xp33_ASAP7_75t_SL g1343 ( 
.A(n_1092),
.B(n_460),
.C(n_455),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1155),
.A2(n_388),
.B1(n_347),
.B2(n_354),
.Y(n_1344)
);

OAI21xp33_ASAP7_75t_L g1345 ( 
.A1(n_1092),
.A2(n_419),
.B(n_355),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1050),
.A2(n_1054),
.B(n_1123),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1211),
.B(n_359),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1180),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1211),
.Y(n_1349)
);

A2O1A1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1181),
.A2(n_393),
.B(n_400),
.C(n_398),
.Y(n_1350)
);

NAND3xp33_ASAP7_75t_SL g1351 ( 
.A(n_1213),
.B(n_370),
.C(n_369),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1180),
.Y(n_1352)
);

BUFx6f_ASAP7_75t_L g1353 ( 
.A(n_1144),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1037),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1174),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1037),
.B(n_611),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1090),
.A2(n_394),
.B(n_348),
.Y(n_1357)
);

A2O1A1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1183),
.A2(n_1043),
.B(n_1194),
.C(n_1162),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1077),
.A2(n_406),
.B(n_372),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1197),
.B(n_461),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1039),
.A2(n_389),
.B1(n_377),
.B2(n_378),
.Y(n_1361)
);

BUFx4f_ASAP7_75t_L g1362 ( 
.A(n_1144),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1053),
.A2(n_350),
.B(n_269),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1039),
.B(n_384),
.Y(n_1364)
);

O2A1O1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1095),
.A2(n_395),
.B(n_416),
.C(n_417),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_R g1366 ( 
.A(n_1175),
.B(n_464),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1095),
.A2(n_418),
.B1(n_463),
.B2(n_462),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_1207),
.B(n_462),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1097),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1173),
.B(n_463),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1097),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1063),
.A2(n_3),
.B(n_4),
.C(n_6),
.Y(n_1372)
);

A2O1A1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1179),
.A2(n_464),
.B(n_421),
.C(n_420),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1207),
.B(n_350),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1073),
.A2(n_412),
.B(n_408),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1099),
.B(n_349),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1175),
.B(n_4),
.Y(n_1377)
);

O2A1O1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1075),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1099),
.B(n_351),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1102),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1102),
.Y(n_1381)
);

AOI21xp33_ASAP7_75t_L g1382 ( 
.A1(n_1137),
.A2(n_269),
.B(n_315),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1176),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1096),
.A2(n_407),
.B(n_404),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1044),
.B(n_350),
.Y(n_1385)
);

AND2x6_ASAP7_75t_L g1386 ( 
.A(n_1370),
.B(n_1075),
.Y(n_1386)
);

AO31x2_ASAP7_75t_L g1387 ( 
.A1(n_1220),
.A2(n_1076),
.A3(n_1118),
.B(n_1122),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1381),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1268),
.B(n_1048),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1234),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1227),
.A2(n_1133),
.B(n_1135),
.Y(n_1391)
);

CKINVDCx11_ASAP7_75t_R g1392 ( 
.A(n_1233),
.Y(n_1392)
);

AO21x1_ASAP7_75t_L g1393 ( 
.A1(n_1372),
.A2(n_1076),
.B(n_1212),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1227),
.A2(n_1346),
.B(n_1222),
.Y(n_1394)
);

O2A1O1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1282),
.A2(n_1219),
.B(n_1218),
.C(n_1198),
.Y(n_1395)
);

NOR2xp67_ASAP7_75t_L g1396 ( 
.A(n_1232),
.B(n_1184),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1241),
.Y(n_1397)
);

NAND2x1p5_ASAP7_75t_L g1398 ( 
.A(n_1362),
.B(n_1256),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1318),
.A2(n_1083),
.B(n_1204),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1362),
.Y(n_1400)
);

AO31x2_ASAP7_75t_L g1401 ( 
.A1(n_1358),
.A2(n_1196),
.A3(n_1200),
.B(n_1193),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1234),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1363),
.A2(n_1030),
.B(n_1186),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1224),
.A2(n_1070),
.B(n_1191),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1268),
.B(n_1172),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1337),
.A2(n_1187),
.B(n_1189),
.Y(n_1406)
);

NAND2x1p5_ASAP7_75t_L g1407 ( 
.A(n_1225),
.B(n_1176),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1322),
.A2(n_1138),
.B(n_1045),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_1340),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_SL g1410 ( 
.A1(n_1335),
.A2(n_1114),
.B(n_1110),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1368),
.A2(n_1217),
.B(n_1088),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1270),
.B(n_1274),
.Y(n_1412)
);

AOI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1385),
.A2(n_1115),
.B(n_1152),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1355),
.A2(n_1158),
.B(n_1119),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_SL g1415 ( 
.A(n_1283),
.B(n_1208),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1246),
.Y(n_1416)
);

AOI221x1_ASAP7_75t_L g1417 ( 
.A1(n_1249),
.A2(n_1216),
.B1(n_1206),
.B2(n_1084),
.C(n_1100),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1228),
.A2(n_1151),
.B(n_1060),
.Y(n_1418)
);

NOR2xp67_ASAP7_75t_SL g1419 ( 
.A(n_1251),
.B(n_1104),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1354),
.A2(n_1068),
.B(n_1109),
.Y(n_1420)
);

AO31x2_ASAP7_75t_L g1421 ( 
.A1(n_1385),
.A2(n_1106),
.A3(n_1134),
.B(n_350),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1270),
.B(n_9),
.Y(n_1422)
);

NAND3xp33_ASAP7_75t_L g1423 ( 
.A(n_1223),
.B(n_1273),
.C(n_1239),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1238),
.A2(n_315),
.B(n_397),
.Y(n_1424)
);

A2O1A1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1281),
.A2(n_403),
.B(n_396),
.C(n_382),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1376),
.A2(n_379),
.B(n_374),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1242),
.B(n_367),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1297),
.Y(n_1428)
);

AO21x1_ASAP7_75t_L g1429 ( 
.A1(n_1370),
.A2(n_315),
.B(n_15),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1238),
.A2(n_315),
.B(n_361),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1271),
.A2(n_365),
.B1(n_352),
.B2(n_23),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1286),
.B(n_13),
.Y(n_1432)
);

AO31x2_ASAP7_75t_L g1433 ( 
.A1(n_1257),
.A2(n_114),
.A3(n_223),
.B(n_220),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_SL g1434 ( 
.A(n_1246),
.Y(n_1434)
);

A2O1A1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1379),
.A2(n_1365),
.B(n_1345),
.C(n_1330),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1252),
.A2(n_112),
.B(n_215),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1246),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1300),
.A2(n_101),
.B(n_208),
.Y(n_1438)
);

INVxp67_ASAP7_75t_L g1439 ( 
.A(n_1236),
.Y(n_1439)
);

AO31x2_ASAP7_75t_L g1440 ( 
.A1(n_1221),
.A2(n_100),
.A3(n_207),
.B(n_205),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1252),
.A2(n_91),
.B(n_202),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1247),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1380),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1324),
.A2(n_90),
.B(n_201),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1254),
.B(n_13),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1326),
.B(n_16),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1374),
.A2(n_1342),
.B(n_1356),
.Y(n_1447)
);

AOI221xp5_ASAP7_75t_L g1448 ( 
.A1(n_1339),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.C(n_36),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1361),
.A2(n_36),
.B(n_37),
.Y(n_1449)
);

BUFx10_ASAP7_75t_L g1450 ( 
.A(n_1287),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1328),
.A2(n_1301),
.B(n_1294),
.Y(n_1451)
);

BUFx8_ASAP7_75t_L g1452 ( 
.A(n_1305),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1374),
.A2(n_129),
.B(n_196),
.Y(n_1453)
);

AO31x2_ASAP7_75t_L g1454 ( 
.A1(n_1290),
.A2(n_120),
.A3(n_188),
.B(n_187),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1356),
.A2(n_92),
.B(n_186),
.Y(n_1455)
);

INVx3_ASAP7_75t_SL g1456 ( 
.A(n_1247),
.Y(n_1456)
);

INVx4_ASAP7_75t_L g1457 ( 
.A(n_1247),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1289),
.A2(n_37),
.B1(n_42),
.B2(n_44),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1302),
.B(n_42),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1255),
.A2(n_130),
.B(n_182),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1366),
.B(n_44),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1269),
.B(n_1275),
.Y(n_1462)
);

AO31x2_ASAP7_75t_L g1463 ( 
.A1(n_1261),
.A2(n_88),
.A3(n_179),
.B(n_177),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1310),
.Y(n_1464)
);

AO21x2_ASAP7_75t_L g1465 ( 
.A1(n_1264),
.A2(n_87),
.B(n_176),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1255),
.A2(n_233),
.B(n_167),
.Y(n_1466)
);

OAI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1361),
.A2(n_47),
.B(n_49),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1327),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1266),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1309),
.A2(n_163),
.B(n_159),
.Y(n_1470)
);

AO31x2_ASAP7_75t_L g1471 ( 
.A1(n_1312),
.A2(n_157),
.A3(n_154),
.B(n_151),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1369),
.A2(n_148),
.B(n_144),
.Y(n_1472)
);

AO31x2_ASAP7_75t_L g1473 ( 
.A1(n_1331),
.A2(n_143),
.A3(n_142),
.B(n_141),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1331),
.A2(n_140),
.B(n_131),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1291),
.Y(n_1475)
);

INVxp67_ASAP7_75t_SL g1476 ( 
.A(n_1298),
.Y(n_1476)
);

INVxp67_ASAP7_75t_SL g1477 ( 
.A(n_1313),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1253),
.Y(n_1478)
);

AND2x6_ASAP7_75t_L g1479 ( 
.A(n_1353),
.B(n_47),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1371),
.A2(n_50),
.B(n_54),
.Y(n_1480)
);

AO31x2_ASAP7_75t_L g1481 ( 
.A1(n_1295),
.A2(n_50),
.A3(n_56),
.B(n_58),
.Y(n_1481)
);

O2A1O1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1339),
.A2(n_60),
.B(n_65),
.C(n_67),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1347),
.B(n_60),
.Y(n_1483)
);

BUFx2_ASAP7_75t_SL g1484 ( 
.A(n_1327),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1296),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1278),
.A2(n_65),
.B(n_68),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1239),
.B(n_68),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1266),
.Y(n_1488)
);

INVxp67_ASAP7_75t_SL g1489 ( 
.A(n_1262),
.Y(n_1489)
);

INVx2_ASAP7_75t_SL g1490 ( 
.A(n_1325),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1360),
.A2(n_70),
.B(n_71),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1266),
.Y(n_1492)
);

AO31x2_ASAP7_75t_L g1493 ( 
.A1(n_1311),
.A2(n_73),
.A3(n_76),
.B(n_79),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1343),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1359),
.A2(n_80),
.B(n_1375),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1292),
.B(n_1288),
.Y(n_1496)
);

O2A1O1Ixp33_ASAP7_75t_SL g1497 ( 
.A1(n_1350),
.A2(n_1351),
.B(n_1293),
.C(n_1373),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1308),
.A2(n_1263),
.B(n_1240),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1267),
.B(n_1276),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1285),
.Y(n_1500)
);

INVx5_ASAP7_75t_L g1501 ( 
.A(n_1272),
.Y(n_1501)
);

AOI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1240),
.A2(n_1230),
.B(n_1260),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1329),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1230),
.A2(n_1260),
.B(n_1248),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1306),
.A2(n_1317),
.B(n_1321),
.Y(n_1505)
);

AOI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1288),
.A2(n_1304),
.B1(n_1323),
.B2(n_1320),
.Y(n_1506)
);

BUFx10_ASAP7_75t_L g1507 ( 
.A(n_1272),
.Y(n_1507)
);

CKINVDCx8_ASAP7_75t_R g1508 ( 
.A(n_1272),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1367),
.A2(n_1364),
.B(n_1304),
.Y(n_1509)
);

AOI221x1_ASAP7_75t_L g1510 ( 
.A1(n_1289),
.A2(n_1382),
.B1(n_1264),
.B2(n_1377),
.C(n_1367),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1316),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1244),
.A2(n_1284),
.B1(n_1280),
.B2(n_1259),
.Y(n_1512)
);

AOI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1332),
.A2(n_1336),
.B(n_1338),
.Y(n_1513)
);

OAI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1235),
.A2(n_1277),
.B1(n_1243),
.B2(n_1237),
.Y(n_1514)
);

A2O1A1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1378),
.A2(n_1377),
.B(n_1245),
.C(n_1333),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1258),
.B(n_1250),
.Y(n_1516)
);

BUFx12f_ASAP7_75t_L g1517 ( 
.A(n_1334),
.Y(n_1517)
);

AO31x2_ASAP7_75t_L g1518 ( 
.A1(n_1349),
.A2(n_1284),
.A3(n_1384),
.B(n_1341),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1353),
.A2(n_1303),
.B(n_1357),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1267),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1276),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1314),
.A2(n_1226),
.B(n_1231),
.Y(n_1522)
);

BUFx2_ASAP7_75t_R g1523 ( 
.A(n_1265),
.Y(n_1523)
);

AO32x2_ASAP7_75t_L g1524 ( 
.A1(n_1299),
.A2(n_1382),
.A3(n_1383),
.B1(n_1319),
.B2(n_1348),
.Y(n_1524)
);

AO31x2_ASAP7_75t_L g1525 ( 
.A1(n_1299),
.A2(n_1352),
.A3(n_1383),
.B(n_1307),
.Y(n_1525)
);

AO31x2_ASAP7_75t_L g1526 ( 
.A1(n_1299),
.A2(n_1344),
.A3(n_1279),
.B(n_1315),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1334),
.B(n_1315),
.Y(n_1527)
);

NOR3xp33_ASAP7_75t_L g1528 ( 
.A(n_1334),
.B(n_973),
.C(n_951),
.Y(n_1528)
);

O2A1O1Ixp33_ASAP7_75t_SL g1529 ( 
.A1(n_1282),
.A2(n_874),
.B(n_862),
.C(n_873),
.Y(n_1529)
);

AO31x2_ASAP7_75t_L g1530 ( 
.A1(n_1220),
.A2(n_1036),
.A3(n_1358),
.B(n_1112),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1335),
.A2(n_1029),
.B1(n_1032),
.B2(n_973),
.Y(n_1531)
);

NOR3xp33_ASAP7_75t_L g1532 ( 
.A(n_1271),
.B(n_973),
.C(n_951),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1229),
.Y(n_1533)
);

A2O1A1Ixp33_ASAP7_75t_L g1534 ( 
.A1(n_1249),
.A2(n_1029),
.B(n_945),
.C(n_951),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1363),
.A2(n_1337),
.B(n_1346),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1363),
.A2(n_1337),
.B(n_1346),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1381),
.Y(n_1537)
);

INVx3_ASAP7_75t_SL g1538 ( 
.A(n_1241),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1268),
.B(n_876),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1268),
.B(n_1032),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1268),
.B(n_1032),
.Y(n_1541)
);

AO31x2_ASAP7_75t_L g1542 ( 
.A1(n_1220),
.A2(n_1036),
.A3(n_1358),
.B(n_1112),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1227),
.A2(n_733),
.B(n_874),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1274),
.B(n_808),
.Y(n_1544)
);

AOI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1227),
.A2(n_733),
.B(n_874),
.Y(n_1545)
);

OAI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1274),
.A2(n_1029),
.B1(n_1032),
.B2(n_973),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1227),
.A2(n_733),
.B(n_874),
.Y(n_1547)
);

AOI221x1_ASAP7_75t_L g1548 ( 
.A1(n_1249),
.A2(n_804),
.B1(n_759),
.B2(n_973),
.C(n_1289),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1227),
.A2(n_733),
.B(n_874),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1227),
.A2(n_733),
.B(n_874),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1381),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1340),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1237),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1227),
.A2(n_733),
.B(n_874),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1363),
.A2(n_1337),
.B(n_1346),
.Y(n_1555)
);

O2A1O1Ixp33_ASAP7_75t_L g1556 ( 
.A1(n_1282),
.A2(n_973),
.B(n_945),
.C(n_951),
.Y(n_1556)
);

O2A1O1Ixp33_ASAP7_75t_L g1557 ( 
.A1(n_1282),
.A2(n_973),
.B(n_945),
.C(n_951),
.Y(n_1557)
);

A2O1A1Ixp33_ASAP7_75t_L g1558 ( 
.A1(n_1249),
.A2(n_1029),
.B(n_945),
.C(n_951),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1381),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1274),
.A2(n_973),
.B1(n_998),
.B2(n_1029),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1381),
.Y(n_1561)
);

AOI221xp5_ASAP7_75t_SL g1562 ( 
.A1(n_1372),
.A2(n_973),
.B1(n_742),
.B2(n_913),
.C(n_951),
.Y(n_1562)
);

AOI221x1_ASAP7_75t_L g1563 ( 
.A1(n_1249),
.A2(n_804),
.B1(n_759),
.B2(n_973),
.C(n_1289),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1487),
.A2(n_1496),
.B1(n_1546),
.B2(n_1560),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1532),
.A2(n_1531),
.B1(n_1506),
.B2(n_1509),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1543),
.A2(n_1547),
.B(n_1545),
.Y(n_1566)
);

CKINVDCx14_ASAP7_75t_R g1567 ( 
.A(n_1392),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1538),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1416),
.Y(n_1569)
);

INVx6_ASAP7_75t_L g1570 ( 
.A(n_1501),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1397),
.Y(n_1571)
);

CKINVDCx16_ASAP7_75t_R g1572 ( 
.A(n_1434),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1409),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1478),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1552),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_1452),
.Y(n_1576)
);

AO22x1_ASAP7_75t_L g1577 ( 
.A1(n_1483),
.A2(n_1479),
.B1(n_1449),
.B2(n_1467),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_SL g1578 ( 
.A1(n_1423),
.A2(n_1446),
.B1(n_1489),
.B2(n_1479),
.Y(n_1578)
);

INVx4_ASAP7_75t_L g1579 ( 
.A(n_1517),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1478),
.Y(n_1580)
);

OAI21xp33_ASAP7_75t_SL g1581 ( 
.A1(n_1448),
.A2(n_1415),
.B(n_1486),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_SL g1582 ( 
.A1(n_1479),
.A2(n_1544),
.B1(n_1445),
.B2(n_1541),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1508),
.Y(n_1583)
);

OAI22xp33_ASAP7_75t_SL g1584 ( 
.A1(n_1412),
.A2(n_1461),
.B1(n_1459),
.B2(n_1422),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1452),
.Y(n_1585)
);

NAND2x1p5_ASAP7_75t_L g1586 ( 
.A(n_1501),
.B(n_1468),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1477),
.Y(n_1587)
);

INVx4_ASAP7_75t_L g1588 ( 
.A(n_1501),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_1428),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1458),
.A2(n_1528),
.B1(n_1429),
.B2(n_1514),
.Y(n_1590)
);

OAI21xp5_ASAP7_75t_SL g1591 ( 
.A1(n_1556),
.A2(n_1557),
.B(n_1534),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1558),
.A2(n_1431),
.B1(n_1540),
.B2(n_1435),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1479),
.A2(n_1512),
.B1(n_1561),
.B2(n_1388),
.Y(n_1593)
);

INVx8_ASAP7_75t_L g1594 ( 
.A(n_1434),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1456),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1388),
.A2(n_1537),
.B1(n_1561),
.B2(n_1551),
.Y(n_1596)
);

BUFx6f_ASAP7_75t_L g1597 ( 
.A(n_1416),
.Y(n_1597)
);

INVx4_ASAP7_75t_L g1598 ( 
.A(n_1400),
.Y(n_1598)
);

INVx6_ASAP7_75t_L g1599 ( 
.A(n_1507),
.Y(n_1599)
);

CKINVDCx11_ASAP7_75t_R g1600 ( 
.A(n_1450),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1537),
.A2(n_1559),
.B1(n_1551),
.B2(n_1516),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1559),
.A2(n_1539),
.B1(n_1443),
.B2(n_1439),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1464),
.Y(n_1603)
);

BUFx4_ASAP7_75t_R g1604 ( 
.A(n_1507),
.Y(n_1604)
);

AOI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1562),
.A2(n_1494),
.B1(n_1427),
.B2(n_1386),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1469),
.Y(n_1606)
);

BUFx12f_ASAP7_75t_L g1607 ( 
.A(n_1450),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1500),
.Y(n_1608)
);

CKINVDCx11_ASAP7_75t_R g1609 ( 
.A(n_1469),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1432),
.B(n_1490),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1500),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1443),
.A2(n_1386),
.B1(n_1389),
.B2(n_1503),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1468),
.B(n_1437),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1515),
.A2(n_1426),
.B1(n_1425),
.B2(n_1491),
.Y(n_1614)
);

INVx8_ASAP7_75t_L g1615 ( 
.A(n_1400),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1482),
.A2(n_1480),
.B1(n_1398),
.B2(n_1495),
.Y(n_1616)
);

INVx6_ASAP7_75t_L g1617 ( 
.A(n_1416),
.Y(n_1617)
);

CKINVDCx6p67_ASAP7_75t_R g1618 ( 
.A(n_1442),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1523),
.Y(n_1619)
);

INVx4_ASAP7_75t_L g1620 ( 
.A(n_1469),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1386),
.A2(n_1503),
.B1(n_1390),
.B2(n_1402),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1511),
.Y(n_1622)
);

AOI22x1_ASAP7_75t_SL g1623 ( 
.A1(n_1457),
.A2(n_1488),
.B1(n_1492),
.B2(n_1390),
.Y(n_1623)
);

BUFx4f_ASAP7_75t_SL g1624 ( 
.A(n_1457),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1451),
.B(n_1402),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1386),
.A2(n_1563),
.B1(n_1548),
.B2(n_1393),
.Y(n_1626)
);

CKINVDCx11_ASAP7_75t_R g1627 ( 
.A(n_1462),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1462),
.A2(n_1499),
.B1(n_1527),
.B2(n_1484),
.Y(n_1628)
);

BUFx6f_ASAP7_75t_L g1629 ( 
.A(n_1520),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1525),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1511),
.A2(n_1533),
.B1(n_1485),
.B2(n_1475),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1396),
.A2(n_1399),
.B1(n_1405),
.B2(n_1436),
.Y(n_1632)
);

CKINVDCx11_ASAP7_75t_R g1633 ( 
.A(n_1521),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1481),
.Y(n_1634)
);

INVx6_ASAP7_75t_L g1635 ( 
.A(n_1488),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1492),
.B(n_1510),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1465),
.A2(n_1410),
.B1(n_1411),
.B2(n_1441),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1502),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1525),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1465),
.A2(n_1444),
.B1(n_1470),
.B2(n_1419),
.Y(n_1640)
);

INVx4_ASAP7_75t_SL g1641 ( 
.A(n_1526),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_SL g1642 ( 
.A1(n_1481),
.A2(n_1493),
.B1(n_1408),
.B2(n_1472),
.Y(n_1642)
);

INVxp67_ASAP7_75t_SL g1643 ( 
.A(n_1414),
.Y(n_1643)
);

OAI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1417),
.A2(n_1498),
.B1(n_1549),
.B2(n_1554),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1493),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1493),
.B(n_1526),
.Y(n_1646)
);

BUFx12f_ASAP7_75t_L g1647 ( 
.A(n_1407),
.Y(n_1647)
);

OAI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1550),
.A2(n_1420),
.B1(n_1430),
.B2(n_1424),
.Y(n_1648)
);

OAI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1519),
.A2(n_1391),
.B1(n_1414),
.B2(n_1505),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1395),
.A2(n_1404),
.B1(n_1394),
.B2(n_1513),
.Y(n_1650)
);

OAI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1529),
.A2(n_1413),
.B1(n_1497),
.B2(n_1530),
.Y(n_1651)
);

BUFx10_ASAP7_75t_L g1652 ( 
.A(n_1504),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_SL g1653 ( 
.A1(n_1522),
.A2(n_1524),
.B(n_1518),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1524),
.Y(n_1654)
);

CKINVDCx6p67_ASAP7_75t_R g1655 ( 
.A(n_1473),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1524),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1447),
.A2(n_1460),
.B1(n_1466),
.B2(n_1453),
.Y(n_1657)
);

BUFx2_ASAP7_75t_SL g1658 ( 
.A(n_1473),
.Y(n_1658)
);

INVx6_ASAP7_75t_L g1659 ( 
.A(n_1518),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1530),
.B(n_1542),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_SL g1661 ( 
.A1(n_1471),
.A2(n_1473),
.B1(n_1454),
.B2(n_1440),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1471),
.Y(n_1662)
);

BUFx3_ASAP7_75t_L g1663 ( 
.A(n_1474),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1455),
.Y(n_1664)
);

BUFx12f_ASAP7_75t_L g1665 ( 
.A(n_1454),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1454),
.B(n_1440),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1440),
.B(n_1387),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1433),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1438),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1463),
.A2(n_1433),
.B1(n_1387),
.B2(n_1401),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1433),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1418),
.B(n_1403),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1463),
.Y(n_1673)
);

NAND2x1p5_ASAP7_75t_L g1674 ( 
.A(n_1406),
.B(n_1535),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1463),
.B(n_1387),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1401),
.A2(n_1421),
.B1(n_1536),
.B2(n_1555),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1421),
.A2(n_1487),
.B1(n_1017),
.B2(n_1018),
.Y(n_1677)
);

BUFx12f_ASAP7_75t_L g1678 ( 
.A(n_1401),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1487),
.B(n_1439),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1538),
.Y(n_1680)
);

BUFx12f_ASAP7_75t_L g1681 ( 
.A(n_1392),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1553),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1476),
.Y(n_1683)
);

CKINVDCx20_ASAP7_75t_R g1684 ( 
.A(n_1392),
.Y(n_1684)
);

BUFx3_ASAP7_75t_L g1685 ( 
.A(n_1538),
.Y(n_1685)
);

BUFx3_ASAP7_75t_L g1686 ( 
.A(n_1538),
.Y(n_1686)
);

BUFx12f_ASAP7_75t_L g1687 ( 
.A(n_1392),
.Y(n_1687)
);

NAND2x1p5_ASAP7_75t_L g1688 ( 
.A(n_1501),
.B(n_1468),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1553),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1487),
.A2(n_1017),
.B1(n_1018),
.B2(n_1011),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1553),
.Y(n_1691)
);

INVx4_ASAP7_75t_L g1692 ( 
.A(n_1538),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1553),
.Y(n_1693)
);

NAND2x1p5_ASAP7_75t_L g1694 ( 
.A(n_1501),
.B(n_1468),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1487),
.A2(n_1017),
.B1(n_1018),
.B2(n_1011),
.Y(n_1695)
);

BUFx12f_ASAP7_75t_L g1696 ( 
.A(n_1392),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1544),
.B2(n_1546),
.Y(n_1697)
);

BUFx4_ASAP7_75t_R g1698 ( 
.A(n_1428),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1487),
.B(n_1439),
.Y(n_1699)
);

BUFx4f_ASAP7_75t_L g1700 ( 
.A(n_1538),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1489),
.B(n_1412),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_1397),
.Y(n_1702)
);

BUFx6f_ASAP7_75t_L g1703 ( 
.A(n_1416),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_1392),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1553),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1544),
.B2(n_1546),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1553),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1487),
.A2(n_1017),
.B1(n_1018),
.B2(n_1011),
.Y(n_1708)
);

BUFx12f_ASAP7_75t_SL g1709 ( 
.A(n_1416),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_SL g1710 ( 
.A1(n_1544),
.A2(n_1423),
.B1(n_1283),
.B2(n_1560),
.Y(n_1710)
);

INVx4_ASAP7_75t_L g1711 ( 
.A(n_1538),
.Y(n_1711)
);

BUFx4f_ASAP7_75t_SL g1712 ( 
.A(n_1538),
.Y(n_1712)
);

BUFx10_ASAP7_75t_L g1713 ( 
.A(n_1544),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1544),
.B2(n_1546),
.Y(n_1714)
);

INVx4_ASAP7_75t_L g1715 ( 
.A(n_1538),
.Y(n_1715)
);

BUFx3_ASAP7_75t_L g1716 ( 
.A(n_1538),
.Y(n_1716)
);

BUFx8_ASAP7_75t_SL g1717 ( 
.A(n_1552),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_SL g1718 ( 
.A1(n_1487),
.A2(n_759),
.B1(n_1531),
.B2(n_804),
.Y(n_1718)
);

CKINVDCx11_ASAP7_75t_R g1719 ( 
.A(n_1392),
.Y(n_1719)
);

CKINVDCx11_ASAP7_75t_R g1720 ( 
.A(n_1392),
.Y(n_1720)
);

INVx6_ASAP7_75t_L g1721 ( 
.A(n_1501),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_SL g1722 ( 
.A1(n_1487),
.A2(n_759),
.B1(n_1531),
.B2(n_804),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1553),
.Y(n_1723)
);

INVx6_ASAP7_75t_L g1724 ( 
.A(n_1501),
.Y(n_1724)
);

INVx2_ASAP7_75t_SL g1725 ( 
.A(n_1397),
.Y(n_1725)
);

INVx6_ASAP7_75t_L g1726 ( 
.A(n_1501),
.Y(n_1726)
);

INVx3_ASAP7_75t_L g1727 ( 
.A(n_1508),
.Y(n_1727)
);

INVx6_ASAP7_75t_L g1728 ( 
.A(n_1501),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_1538),
.Y(n_1729)
);

BUFx2_ASAP7_75t_L g1730 ( 
.A(n_1476),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1487),
.A2(n_1017),
.B1(n_1018),
.B2(n_1011),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1489),
.B(n_1412),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1553),
.Y(n_1733)
);

BUFx10_ASAP7_75t_L g1734 ( 
.A(n_1544),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1489),
.B(n_1412),
.Y(n_1735)
);

CKINVDCx6p67_ASAP7_75t_R g1736 ( 
.A(n_1392),
.Y(n_1736)
);

INVx4_ASAP7_75t_SL g1737 ( 
.A(n_1479),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1553),
.Y(n_1738)
);

AOI21x1_ASAP7_75t_L g1739 ( 
.A1(n_1672),
.A2(n_1577),
.B(n_1650),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1574),
.B(n_1580),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1608),
.B(n_1611),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1634),
.Y(n_1742)
);

BUFx2_ASAP7_75t_L g1743 ( 
.A(n_1678),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1645),
.Y(n_1744)
);

BUFx8_ASAP7_75t_L g1745 ( 
.A(n_1681),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1625),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1622),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1587),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1663),
.Y(n_1749)
);

BUFx3_ASAP7_75t_L g1750 ( 
.A(n_1683),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1682),
.Y(n_1751)
);

BUFx3_ASAP7_75t_L g1752 ( 
.A(n_1730),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1689),
.Y(n_1753)
);

INVxp67_ASAP7_75t_L g1754 ( 
.A(n_1610),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1659),
.Y(n_1755)
);

BUFx3_ASAP7_75t_L g1756 ( 
.A(n_1638),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1652),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1738),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1691),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1693),
.Y(n_1760)
);

OR2x6_ASAP7_75t_L g1761 ( 
.A(n_1653),
.B(n_1665),
.Y(n_1761)
);

AO21x2_ASAP7_75t_L g1762 ( 
.A1(n_1651),
.A2(n_1675),
.B(n_1670),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1705),
.B(n_1707),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_1719),
.Y(n_1764)
);

INVx2_ASAP7_75t_SL g1765 ( 
.A(n_1594),
.Y(n_1765)
);

OA21x2_ASAP7_75t_L g1766 ( 
.A1(n_1566),
.A2(n_1660),
.B(n_1668),
.Y(n_1766)
);

BUFx3_ASAP7_75t_L g1767 ( 
.A(n_1570),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1723),
.Y(n_1768)
);

INVx3_ASAP7_75t_L g1769 ( 
.A(n_1669),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1733),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1630),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1701),
.Y(n_1772)
);

OAI21x1_ASAP7_75t_L g1773 ( 
.A1(n_1566),
.A2(n_1676),
.B(n_1674),
.Y(n_1773)
);

BUFx2_ASAP7_75t_L g1774 ( 
.A(n_1643),
.Y(n_1774)
);

AO21x2_ASAP7_75t_L g1775 ( 
.A1(n_1651),
.A2(n_1666),
.B(n_1649),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1679),
.B(n_1699),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1639),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1630),
.Y(n_1778)
);

OA21x2_ASAP7_75t_L g1779 ( 
.A1(n_1672),
.A2(n_1673),
.B(n_1637),
.Y(n_1779)
);

OAI21x1_ASAP7_75t_L g1780 ( 
.A1(n_1674),
.A2(n_1657),
.B(n_1640),
.Y(n_1780)
);

BUFx2_ASAP7_75t_L g1781 ( 
.A(n_1643),
.Y(n_1781)
);

BUFx3_ASAP7_75t_L g1782 ( 
.A(n_1570),
.Y(n_1782)
);

BUFx12f_ASAP7_75t_L g1783 ( 
.A(n_1719),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_SL g1784 ( 
.A1(n_1710),
.A2(n_1697),
.B1(n_1706),
.B2(n_1714),
.Y(n_1784)
);

NAND2x1_ASAP7_75t_L g1785 ( 
.A(n_1632),
.B(n_1669),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1646),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1654),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1656),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1591),
.A2(n_1565),
.B(n_1640),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1658),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1655),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1564),
.B(n_1565),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1667),
.Y(n_1793)
);

INVx1_ASAP7_75t_SL g1794 ( 
.A(n_1589),
.Y(n_1794)
);

HB1xp67_ASAP7_75t_L g1795 ( 
.A(n_1732),
.Y(n_1795)
);

OAI21x1_ASAP7_75t_L g1796 ( 
.A1(n_1657),
.A2(n_1637),
.B(n_1636),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1671),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1735),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1596),
.Y(n_1799)
);

OAI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1592),
.A2(n_1564),
.B(n_1614),
.Y(n_1800)
);

OR2x6_ASAP7_75t_L g1801 ( 
.A(n_1737),
.B(n_1594),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1596),
.Y(n_1802)
);

OAI21x1_ASAP7_75t_L g1803 ( 
.A1(n_1621),
.A2(n_1612),
.B(n_1616),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1662),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1648),
.A2(n_1649),
.B(n_1644),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1641),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1621),
.B(n_1612),
.Y(n_1807)
);

OAI21x1_ASAP7_75t_L g1808 ( 
.A1(n_1626),
.A2(n_1677),
.B(n_1593),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1602),
.B(n_1677),
.Y(n_1809)
);

BUFx12f_ASAP7_75t_L g1810 ( 
.A(n_1720),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1698),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1713),
.B(n_1734),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1582),
.B(n_1641),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1613),
.B(n_1601),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1698),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1718),
.A2(n_1722),
.B1(n_1708),
.B2(n_1731),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1601),
.B(n_1573),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1669),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1593),
.B(n_1590),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_SL g1820 ( 
.A1(n_1661),
.A2(n_1584),
.B1(n_1619),
.B2(n_1581),
.Y(n_1820)
);

OA21x2_ASAP7_75t_L g1821 ( 
.A1(n_1626),
.A2(n_1664),
.B(n_1590),
.Y(n_1821)
);

INVx2_ASAP7_75t_SL g1822 ( 
.A(n_1594),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1578),
.B(n_1575),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1644),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1737),
.B(n_1642),
.Y(n_1825)
);

AO21x2_ASAP7_75t_L g1826 ( 
.A1(n_1648),
.A2(n_1605),
.B(n_1628),
.Y(n_1826)
);

OAI21x1_ASAP7_75t_L g1827 ( 
.A1(n_1586),
.A2(n_1688),
.B(n_1694),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1629),
.Y(n_1828)
);

OAI21x1_ASAP7_75t_L g1829 ( 
.A1(n_1586),
.A2(n_1688),
.B(n_1694),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1642),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1569),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1631),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1631),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1737),
.Y(n_1834)
);

BUFx2_ASAP7_75t_L g1835 ( 
.A(n_1569),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1569),
.B(n_1597),
.Y(n_1836)
);

OAI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1690),
.A2(n_1708),
.B1(n_1695),
.B2(n_1700),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1623),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1597),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1713),
.B(n_1734),
.Y(n_1840)
);

AND2x4_ASAP7_75t_L g1841 ( 
.A(n_1597),
.B(n_1703),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1703),
.Y(n_1842)
);

INVx3_ASAP7_75t_L g1843 ( 
.A(n_1703),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1703),
.B(n_1598),
.Y(n_1844)
);

HB1xp67_ASAP7_75t_L g1845 ( 
.A(n_1606),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1606),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1635),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1635),
.Y(n_1848)
);

INVxp67_ASAP7_75t_L g1849 ( 
.A(n_1571),
.Y(n_1849)
);

AND2x4_ASAP7_75t_L g1850 ( 
.A(n_1620),
.B(n_1588),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1635),
.Y(n_1851)
);

INVx3_ASAP7_75t_L g1852 ( 
.A(n_1620),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1695),
.B(n_1627),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1583),
.B(n_1727),
.Y(n_1854)
);

O2A1O1Ixp33_ASAP7_75t_L g1855 ( 
.A1(n_1583),
.A2(n_1727),
.B(n_1702),
.C(n_1725),
.Y(n_1855)
);

OAI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1700),
.A2(n_1588),
.B(n_1598),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1617),
.Y(n_1857)
);

OAI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1680),
.A2(n_1729),
.B(n_1711),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1617),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1627),
.B(n_1617),
.Y(n_1860)
);

INVxp33_ASAP7_75t_L g1861 ( 
.A(n_1600),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1721),
.Y(n_1862)
);

NAND2x1p5_ASAP7_75t_L g1863 ( 
.A(n_1595),
.B(n_1579),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1721),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1724),
.Y(n_1865)
);

OAI21x1_ASAP7_75t_L g1866 ( 
.A1(n_1604),
.A2(n_1726),
.B(n_1724),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1726),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1728),
.Y(n_1868)
);

INVx2_ASAP7_75t_SL g1869 ( 
.A(n_1728),
.Y(n_1869)
);

INVx1_ASAP7_75t_SL g1870 ( 
.A(n_1600),
.Y(n_1870)
);

INVx2_ASAP7_75t_SL g1871 ( 
.A(n_1728),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1709),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1647),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1609),
.B(n_1618),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1599),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1572),
.B(n_1685),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1599),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1599),
.Y(n_1878)
);

INVx2_ASAP7_75t_SL g1879 ( 
.A(n_1568),
.Y(n_1879)
);

BUFx3_ASAP7_75t_L g1880 ( 
.A(n_1609),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1633),
.A2(n_1607),
.B1(n_1687),
.B2(n_1696),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1633),
.B(n_1716),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1615),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1615),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1751),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1819),
.A2(n_1567),
.B1(n_1736),
.B2(n_1720),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1750),
.B(n_1686),
.Y(n_1887)
);

AOI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1789),
.A2(n_1615),
.B(n_1579),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1776),
.B(n_1692),
.Y(n_1889)
);

O2A1O1Ixp33_ASAP7_75t_L g1890 ( 
.A1(n_1800),
.A2(n_1567),
.B(n_1576),
.C(n_1684),
.Y(n_1890)
);

NAND4xp25_ASAP7_75t_L g1891 ( 
.A(n_1784),
.B(n_1715),
.C(n_1692),
.D(n_1711),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1812),
.B(n_1712),
.Y(n_1892)
);

AO21x2_ASAP7_75t_L g1893 ( 
.A1(n_1791),
.A2(n_1717),
.B(n_1624),
.Y(n_1893)
);

OAI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1792),
.A2(n_1715),
.B(n_1585),
.Y(n_1894)
);

CKINVDCx11_ASAP7_75t_R g1895 ( 
.A(n_1783),
.Y(n_1895)
);

OAI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1792),
.A2(n_1603),
.B(n_1704),
.Y(n_1896)
);

AOI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1837),
.A2(n_1712),
.B1(n_1624),
.B2(n_1717),
.Y(n_1897)
);

AND2x4_ASAP7_75t_L g1898 ( 
.A(n_1750),
.B(n_1752),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1772),
.B(n_1795),
.Y(n_1899)
);

OA21x2_ASAP7_75t_L g1900 ( 
.A1(n_1796),
.A2(n_1805),
.B(n_1780),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1776),
.B(n_1752),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1753),
.Y(n_1902)
);

OAI22xp5_ASAP7_75t_SL g1903 ( 
.A1(n_1783),
.A2(n_1810),
.B1(n_1764),
.B2(n_1881),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1798),
.B(n_1748),
.Y(n_1904)
);

OR2x6_ASAP7_75t_L g1905 ( 
.A(n_1801),
.B(n_1866),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1811),
.B(n_1815),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1753),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1754),
.B(n_1756),
.Y(n_1908)
);

AOI211xp5_ASAP7_75t_L g1909 ( 
.A1(n_1824),
.A2(n_1823),
.B(n_1803),
.C(n_1807),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1758),
.Y(n_1910)
);

O2A1O1Ixp33_ASAP7_75t_L g1911 ( 
.A1(n_1824),
.A2(n_1855),
.B(n_1830),
.C(n_1840),
.Y(n_1911)
);

O2A1O1Ixp33_ASAP7_75t_L g1912 ( 
.A1(n_1830),
.A2(n_1854),
.B(n_1756),
.C(n_1826),
.Y(n_1912)
);

INVx2_ASAP7_75t_SL g1913 ( 
.A(n_1876),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1756),
.B(n_1860),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1743),
.B(n_1880),
.Y(n_1915)
);

AND2x4_ASAP7_75t_L g1916 ( 
.A(n_1743),
.B(n_1880),
.Y(n_1916)
);

O2A1O1Ixp33_ASAP7_75t_L g1917 ( 
.A1(n_1826),
.A2(n_1785),
.B(n_1807),
.C(n_1849),
.Y(n_1917)
);

O2A1O1Ixp33_ASAP7_75t_L g1918 ( 
.A1(n_1826),
.A2(n_1785),
.B(n_1858),
.C(n_1817),
.Y(n_1918)
);

AND2x4_ASAP7_75t_SL g1919 ( 
.A(n_1801),
.B(n_1874),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1860),
.B(n_1763),
.Y(n_1920)
);

OR2x6_ASAP7_75t_L g1921 ( 
.A(n_1801),
.B(n_1880),
.Y(n_1921)
);

NOR2x1_ASAP7_75t_SL g1922 ( 
.A(n_1801),
.B(n_1775),
.Y(n_1922)
);

NAND4xp25_ASAP7_75t_L g1923 ( 
.A(n_1820),
.B(n_1870),
.C(n_1856),
.D(n_1770),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1882),
.B(n_1740),
.Y(n_1924)
);

AND2x4_ASAP7_75t_L g1925 ( 
.A(n_1791),
.B(n_1825),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1838),
.B(n_1850),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1740),
.B(n_1741),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1882),
.B(n_1741),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1813),
.B(n_1767),
.Y(n_1929)
);

A2O1A1Ixp33_ASAP7_75t_L g1930 ( 
.A1(n_1803),
.A2(n_1808),
.B(n_1853),
.C(n_1809),
.Y(n_1930)
);

INVxp67_ASAP7_75t_L g1931 ( 
.A(n_1845),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1759),
.Y(n_1932)
);

AO32x2_ASAP7_75t_L g1933 ( 
.A1(n_1869),
.A2(n_1871),
.A3(n_1879),
.B1(n_1765),
.B2(n_1822),
.Y(n_1933)
);

AOI21xp5_ASAP7_75t_L g1934 ( 
.A1(n_1775),
.A2(n_1762),
.B(n_1779),
.Y(n_1934)
);

OA21x2_ASAP7_75t_L g1935 ( 
.A1(n_1796),
.A2(n_1780),
.B(n_1773),
.Y(n_1935)
);

AO32x2_ASAP7_75t_L g1936 ( 
.A1(n_1869),
.A2(n_1871),
.A3(n_1879),
.B1(n_1822),
.B2(n_1765),
.Y(n_1936)
);

INVxp67_ASAP7_75t_L g1937 ( 
.A(n_1831),
.Y(n_1937)
);

INVx1_ASAP7_75t_SL g1938 ( 
.A(n_1876),
.Y(n_1938)
);

HB1xp67_ASAP7_75t_L g1939 ( 
.A(n_1760),
.Y(n_1939)
);

OA21x2_ASAP7_75t_L g1940 ( 
.A1(n_1773),
.A2(n_1739),
.B(n_1808),
.Y(n_1940)
);

A2O1A1Ixp33_ASAP7_75t_L g1941 ( 
.A1(n_1853),
.A2(n_1809),
.B(n_1816),
.C(n_1838),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1760),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1782),
.B(n_1768),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1835),
.B(n_1874),
.Y(n_1944)
);

NOR2xp33_ASAP7_75t_SL g1945 ( 
.A(n_1810),
.B(n_1764),
.Y(n_1945)
);

OAI21xp5_ASAP7_75t_L g1946 ( 
.A1(n_1739),
.A2(n_1821),
.B(n_1846),
.Y(n_1946)
);

O2A1O1Ixp33_ASAP7_75t_SL g1947 ( 
.A1(n_1861),
.A2(n_1794),
.B(n_1844),
.C(n_1872),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1863),
.B(n_1872),
.Y(n_1948)
);

AO32x2_ASAP7_75t_L g1949 ( 
.A1(n_1786),
.A2(n_1814),
.A3(n_1821),
.B1(n_1799),
.B2(n_1802),
.Y(n_1949)
);

OAI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1821),
.A2(n_1846),
.B(n_1746),
.Y(n_1950)
);

OAI211xp5_ASAP7_75t_SL g1951 ( 
.A1(n_1883),
.A2(n_1878),
.B(n_1877),
.C(n_1875),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1839),
.B(n_1842),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1770),
.B(n_1747),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1842),
.B(n_1836),
.Y(n_1954)
);

NOR2xp33_ASAP7_75t_L g1955 ( 
.A(n_1863),
.B(n_1873),
.Y(n_1955)
);

AO32x2_ASAP7_75t_L g1956 ( 
.A1(n_1821),
.A2(n_1833),
.A3(n_1832),
.B1(n_1804),
.B2(n_1787),
.Y(n_1956)
);

OAI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1863),
.A2(n_1883),
.B1(n_1875),
.B2(n_1878),
.Y(n_1957)
);

O2A1O1Ixp33_ASAP7_75t_L g1958 ( 
.A1(n_1857),
.A2(n_1859),
.B(n_1847),
.C(n_1762),
.Y(n_1958)
);

OR2x6_ASAP7_75t_L g1959 ( 
.A(n_1834),
.B(n_1827),
.Y(n_1959)
);

AOI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1834),
.A2(n_1873),
.B1(n_1847),
.B2(n_1848),
.Y(n_1960)
);

AOI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1779),
.A2(n_1766),
.B(n_1781),
.Y(n_1961)
);

OAI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1746),
.A2(n_1827),
.B(n_1829),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1747),
.B(n_1848),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1836),
.B(n_1841),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1841),
.B(n_1851),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1857),
.B(n_1859),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1788),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1774),
.B(n_1781),
.Y(n_1968)
);

BUFx3_ASAP7_75t_L g1969 ( 
.A(n_1745),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1877),
.B(n_1868),
.Y(n_1970)
);

A2O1A1Ixp33_ASAP7_75t_L g1971 ( 
.A1(n_1829),
.A2(n_1793),
.B(n_1790),
.C(n_1806),
.Y(n_1971)
);

AOI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1862),
.A2(n_1864),
.B1(n_1868),
.B2(n_1867),
.Y(n_1972)
);

OAI22xp5_ASAP7_75t_SL g1973 ( 
.A1(n_1745),
.A2(n_1761),
.B1(n_1884),
.B2(n_1850),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1843),
.B(n_1828),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1901),
.B(n_1920),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1939),
.Y(n_1976)
);

CKINVDCx20_ASAP7_75t_R g1977 ( 
.A(n_1895),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1968),
.Y(n_1978)
);

HB1xp67_ASAP7_75t_L g1979 ( 
.A(n_1931),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1924),
.B(n_1749),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1928),
.B(n_1769),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1937),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1967),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1950),
.B(n_1927),
.Y(n_1984)
);

INVxp67_ASAP7_75t_SL g1985 ( 
.A(n_1961),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1885),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1902),
.Y(n_1987)
);

BUFx2_ASAP7_75t_L g1988 ( 
.A(n_1933),
.Y(n_1988)
);

AOI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1923),
.A2(n_1797),
.B1(n_1777),
.B2(n_1755),
.Y(n_1989)
);

BUFx2_ASAP7_75t_L g1990 ( 
.A(n_1933),
.Y(n_1990)
);

INVx2_ASAP7_75t_SL g1991 ( 
.A(n_1915),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1907),
.B(n_1778),
.Y(n_1992)
);

CKINVDCx6p67_ASAP7_75t_R g1993 ( 
.A(n_1969),
.Y(n_1993)
);

HB1xp67_ASAP7_75t_L g1994 ( 
.A(n_1904),
.Y(n_1994)
);

BUFx2_ASAP7_75t_L g1995 ( 
.A(n_1933),
.Y(n_1995)
);

BUFx2_ASAP7_75t_L g1996 ( 
.A(n_1936),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1910),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1898),
.B(n_1818),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1922),
.B(n_1757),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1932),
.Y(n_2000)
);

OR2x2_ASAP7_75t_L g2001 ( 
.A(n_1899),
.B(n_1778),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1942),
.B(n_1771),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1963),
.B(n_1912),
.Y(n_2003)
);

AND2x4_ASAP7_75t_L g2004 ( 
.A(n_1922),
.B(n_1757),
.Y(n_2004)
);

BUFx2_ASAP7_75t_L g2005 ( 
.A(n_1936),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1953),
.B(n_1771),
.Y(n_2006)
);

OAI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1941),
.A2(n_1884),
.B1(n_1852),
.B2(n_1850),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1935),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1918),
.B(n_1742),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1956),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1956),
.Y(n_2011)
);

BUFx2_ASAP7_75t_L g2012 ( 
.A(n_1936),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1956),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1949),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1949),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1949),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1966),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1900),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1970),
.Y(n_2019)
);

NAND3xp33_ASAP7_75t_L g2020 ( 
.A(n_1909),
.B(n_1790),
.C(n_1865),
.Y(n_2020)
);

BUFx6f_ASAP7_75t_L g2021 ( 
.A(n_1940),
.Y(n_2021)
);

INVxp67_ASAP7_75t_SL g2022 ( 
.A(n_1958),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1908),
.B(n_1818),
.Y(n_2023)
);

O2A1O1Ixp33_ASAP7_75t_L g2024 ( 
.A1(n_2022),
.A2(n_1917),
.B(n_1911),
.C(n_1930),
.Y(n_2024)
);

HB1xp67_ASAP7_75t_L g2025 ( 
.A(n_1978),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_2018),
.Y(n_2026)
);

AND2x4_ASAP7_75t_L g2027 ( 
.A(n_1999),
.B(n_1921),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1984),
.B(n_1938),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1992),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1988),
.B(n_1990),
.Y(n_2030)
);

INVx4_ASAP7_75t_L g2031 ( 
.A(n_1993),
.Y(n_2031)
);

HB1xp67_ASAP7_75t_L g2032 ( 
.A(n_1976),
.Y(n_2032)
);

AO21x2_ASAP7_75t_L g2033 ( 
.A1(n_1985),
.A2(n_1934),
.B(n_1946),
.Y(n_2033)
);

OA332x1_ASAP7_75t_L g2034 ( 
.A1(n_1979),
.A2(n_1945),
.A3(n_1903),
.B1(n_1957),
.B2(n_1886),
.B3(n_1890),
.C1(n_1896),
.C2(n_1889),
.Y(n_2034)
);

INVx1_ASAP7_75t_SL g2035 ( 
.A(n_1977),
.Y(n_2035)
);

OR2x6_ASAP7_75t_L g2036 ( 
.A(n_2020),
.B(n_1905),
.Y(n_2036)
);

OAI33xp33_ASAP7_75t_L g2037 ( 
.A1(n_2003),
.A2(n_1891),
.A3(n_1951),
.B1(n_1926),
.B2(n_1973),
.B3(n_1744),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1984),
.B(n_2017),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1992),
.Y(n_2039)
);

OAI31xp33_ASAP7_75t_L g2040 ( 
.A1(n_2020),
.A2(n_1971),
.A3(n_1888),
.B(n_1947),
.Y(n_2040)
);

OAI321xp33_ASAP7_75t_L g2041 ( 
.A1(n_2022),
.A2(n_1962),
.A3(n_1897),
.B1(n_1960),
.B2(n_1972),
.C(n_1959),
.Y(n_2041)
);

HB1xp67_ASAP7_75t_L g2042 ( 
.A(n_1976),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1988),
.B(n_1944),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2002),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1990),
.B(n_1914),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2002),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2017),
.B(n_1913),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1995),
.B(n_1906),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_L g2049 ( 
.A(n_1993),
.B(n_1892),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1983),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1983),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1986),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1995),
.B(n_1887),
.Y(n_2053)
);

AOI221xp5_ASAP7_75t_L g2054 ( 
.A1(n_2003),
.A2(n_1925),
.B1(n_1955),
.B2(n_1952),
.C(n_1894),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1986),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1996),
.B(n_1887),
.Y(n_2056)
);

INVxp67_ASAP7_75t_SL g2057 ( 
.A(n_2009),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1987),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1996),
.B(n_1964),
.Y(n_2059)
);

INVx2_ASAP7_75t_SL g2060 ( 
.A(n_1991),
.Y(n_2060)
);

OAI31xp33_ASAP7_75t_L g2061 ( 
.A1(n_2007),
.A2(n_1919),
.A3(n_1915),
.B(n_1916),
.Y(n_2061)
);

OR2x2_ASAP7_75t_L g2062 ( 
.A(n_2001),
.B(n_1954),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_2005),
.B(n_1916),
.Y(n_2063)
);

OR2x2_ASAP7_75t_L g2064 ( 
.A(n_2001),
.B(n_2005),
.Y(n_2064)
);

BUFx2_ASAP7_75t_L g2065 ( 
.A(n_2012),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2019),
.B(n_1994),
.Y(n_2066)
);

INVx1_ASAP7_75t_SL g2067 ( 
.A(n_1993),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2008),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1987),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_2012),
.B(n_1974),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1997),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_2021),
.Y(n_2072)
);

BUFx2_ASAP7_75t_L g2073 ( 
.A(n_1999),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_2008),
.Y(n_2074)
);

HB1xp67_ASAP7_75t_L g2075 ( 
.A(n_1982),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1975),
.B(n_1965),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1975),
.B(n_1929),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_2010),
.B(n_1940),
.Y(n_2078)
);

INVxp67_ASAP7_75t_L g2079 ( 
.A(n_2006),
.Y(n_2079)
);

OAI31xp33_ASAP7_75t_L g2080 ( 
.A1(n_2007),
.A2(n_1948),
.A3(n_1929),
.B(n_1943),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2000),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_2026),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2050),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_2064),
.B(n_2038),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_2026),
.Y(n_2085)
);

AND2x4_ASAP7_75t_L g2086 ( 
.A(n_2027),
.B(n_2073),
.Y(n_2086)
);

NAND3xp33_ASAP7_75t_SL g2087 ( 
.A(n_2040),
.B(n_2013),
.C(n_2011),
.Y(n_2087)
);

INVx4_ASAP7_75t_L g2088 ( 
.A(n_2031),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_2030),
.B(n_1991),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2057),
.B(n_2010),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2029),
.B(n_2011),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2030),
.B(n_1980),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2029),
.B(n_2011),
.Y(n_2093)
);

AND2x4_ASAP7_75t_L g2094 ( 
.A(n_2027),
.B(n_1999),
.Y(n_2094)
);

NAND3xp33_ASAP7_75t_L g2095 ( 
.A(n_2024),
.B(n_1985),
.C(n_2009),
.Y(n_2095)
);

OR2x2_ASAP7_75t_L g2096 ( 
.A(n_2064),
.B(n_2014),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_2065),
.B(n_2014),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2063),
.B(n_1980),
.Y(n_2098)
);

NOR2xp67_ASAP7_75t_L g2099 ( 
.A(n_2031),
.B(n_2041),
.Y(n_2099)
);

HB1xp67_ASAP7_75t_L g2100 ( 
.A(n_2075),
.Y(n_2100)
);

HB1xp67_ASAP7_75t_L g2101 ( 
.A(n_2025),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2039),
.B(n_2013),
.Y(n_2102)
);

INVxp67_ASAP7_75t_L g2103 ( 
.A(n_2037),
.Y(n_2103)
);

INVxp67_ASAP7_75t_SL g2104 ( 
.A(n_2026),
.Y(n_2104)
);

OR2x2_ASAP7_75t_L g2105 ( 
.A(n_2065),
.B(n_2066),
.Y(n_2105)
);

INVx1_ASAP7_75t_SL g2106 ( 
.A(n_2035),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2039),
.B(n_2013),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2053),
.B(n_1981),
.Y(n_2108)
);

HB1xp67_ASAP7_75t_L g2109 ( 
.A(n_2032),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2050),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2044),
.B(n_2015),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2053),
.B(n_2056),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2051),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2044),
.B(n_2046),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2056),
.B(n_1998),
.Y(n_2115)
);

INVx1_ASAP7_75t_SL g2116 ( 
.A(n_2067),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2073),
.B(n_2048),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2046),
.B(n_2015),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2051),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2048),
.B(n_1998),
.Y(n_2120)
);

INVx3_ASAP7_75t_L g2121 ( 
.A(n_2072),
.Y(n_2121)
);

NOR2xp33_ASAP7_75t_L g2122 ( 
.A(n_2049),
.B(n_1745),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2068),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2052),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2052),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2045),
.B(n_2059),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2043),
.B(n_2023),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_R g2128 ( 
.A(n_2034),
.B(n_1999),
.Y(n_2128)
);

AND2x4_ASAP7_75t_L g2129 ( 
.A(n_2027),
.B(n_2004),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_2079),
.B(n_2016),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2095),
.B(n_2028),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2126),
.B(n_2043),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2126),
.B(n_2077),
.Y(n_2133)
);

BUFx2_ASAP7_75t_L g2134 ( 
.A(n_2088),
.Y(n_2134)
);

OR2x2_ASAP7_75t_L g2135 ( 
.A(n_2084),
.B(n_2078),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_2082),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2083),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2095),
.B(n_2042),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2083),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2103),
.B(n_2081),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2110),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2110),
.Y(n_2142)
);

OR2x2_ASAP7_75t_L g2143 ( 
.A(n_2084),
.B(n_2078),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2113),
.Y(n_2144)
);

INVxp67_ASAP7_75t_L g2145 ( 
.A(n_2101),
.Y(n_2145)
);

HB1xp67_ASAP7_75t_L g2146 ( 
.A(n_2100),
.Y(n_2146)
);

OR2x2_ASAP7_75t_L g2147 ( 
.A(n_2090),
.B(n_2062),
.Y(n_2147)
);

OR2x2_ASAP7_75t_L g2148 ( 
.A(n_2090),
.B(n_2062),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2112),
.B(n_2077),
.Y(n_2149)
);

INVx1_ASAP7_75t_SL g2150 ( 
.A(n_2106),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2112),
.B(n_2031),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2113),
.Y(n_2152)
);

OR2x2_ASAP7_75t_L g2153 ( 
.A(n_2130),
.B(n_2055),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2086),
.B(n_2031),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2086),
.B(n_2076),
.Y(n_2155)
);

OAI21xp5_ASAP7_75t_L g2156 ( 
.A1(n_2087),
.A2(n_2099),
.B(n_2103),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2119),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2082),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2109),
.B(n_2116),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2119),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2086),
.B(n_2076),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2116),
.B(n_2055),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2086),
.B(n_2060),
.Y(n_2163)
);

NOR2xp67_ASAP7_75t_SL g2164 ( 
.A(n_2088),
.B(n_1745),
.Y(n_2164)
);

OR2x2_ASAP7_75t_L g2165 ( 
.A(n_2130),
.B(n_2058),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2087),
.B(n_2058),
.Y(n_2166)
);

AND2x4_ASAP7_75t_L g2167 ( 
.A(n_2094),
.B(n_2027),
.Y(n_2167)
);

NOR2x1_ASAP7_75t_L g2168 ( 
.A(n_2106),
.B(n_1893),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2124),
.Y(n_2169)
);

NOR2xp33_ASAP7_75t_L g2170 ( 
.A(n_2122),
.B(n_2060),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2117),
.B(n_2070),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2082),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2117),
.B(n_2094),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2124),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2105),
.B(n_2069),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2125),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2125),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2105),
.B(n_2069),
.Y(n_2178)
);

OR2x2_ASAP7_75t_L g2179 ( 
.A(n_2097),
.B(n_2081),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2114),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_L g2181 ( 
.A(n_2088),
.B(n_2047),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2114),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2152),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_2136),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2149),
.B(n_2094),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2152),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2149),
.B(n_2094),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2133),
.B(n_2129),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2133),
.B(n_2129),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2174),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2173),
.B(n_2129),
.Y(n_2191)
);

INVxp67_ASAP7_75t_L g2192 ( 
.A(n_2140),
.Y(n_2192)
);

AOI21xp5_ASAP7_75t_L g2193 ( 
.A1(n_2156),
.A2(n_2099),
.B(n_2040),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2174),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_2173),
.B(n_2129),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2155),
.B(n_2161),
.Y(n_2196)
);

NAND2x1p5_ASAP7_75t_L g2197 ( 
.A(n_2164),
.B(n_2088),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2137),
.Y(n_2198)
);

AOI22xp33_ASAP7_75t_L g2199 ( 
.A1(n_2166),
.A2(n_2036),
.B1(n_2033),
.B2(n_2016),
.Y(n_2199)
);

OR2x2_ASAP7_75t_L g2200 ( 
.A(n_2147),
.B(n_2097),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_2150),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2155),
.B(n_2089),
.Y(n_2202)
);

OAI22xp5_ASAP7_75t_L g2203 ( 
.A1(n_2131),
.A2(n_2036),
.B1(n_2128),
.B2(n_2089),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2136),
.Y(n_2204)
);

AOI22xp5_ASAP7_75t_L g2205 ( 
.A1(n_2168),
.A2(n_2033),
.B1(n_2036),
.B2(n_1989),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2146),
.B(n_2092),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2139),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2145),
.B(n_2092),
.Y(n_2208)
);

AND2x4_ASAP7_75t_L g2209 ( 
.A(n_2167),
.B(n_2121),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2141),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2142),
.Y(n_2211)
);

NAND4xp25_ASAP7_75t_L g2212 ( 
.A(n_2138),
.B(n_2128),
.C(n_2121),
.D(n_2061),
.Y(n_2212)
);

NOR2xp33_ASAP7_75t_L g2213 ( 
.A(n_2159),
.B(n_2115),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2144),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2158),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2161),
.B(n_2115),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2132),
.B(n_2120),
.Y(n_2217)
);

CKINVDCx16_ASAP7_75t_R g2218 ( 
.A(n_2154),
.Y(n_2218)
);

OR2x2_ASAP7_75t_L g2219 ( 
.A(n_2147),
.B(n_2096),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2162),
.B(n_2127),
.Y(n_2220)
);

AOI21xp5_ASAP7_75t_L g2221 ( 
.A1(n_2175),
.A2(n_2036),
.B(n_2033),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2132),
.B(n_2120),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2158),
.Y(n_2223)
);

NAND2xp33_ASAP7_75t_SL g2224 ( 
.A(n_2164),
.B(n_2127),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_2217),
.B(n_2154),
.Y(n_2225)
);

OAI21xp5_ASAP7_75t_L g2226 ( 
.A1(n_2193),
.A2(n_2181),
.B(n_2178),
.Y(n_2226)
);

OAI21xp33_ASAP7_75t_L g2227 ( 
.A1(n_2212),
.A2(n_2180),
.B(n_2182),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2183),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2183),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2186),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2217),
.B(n_2151),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2186),
.Y(n_2232)
);

NOR3xp33_ASAP7_75t_L g2233 ( 
.A(n_2192),
.B(n_2201),
.C(n_2203),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2190),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_2201),
.B(n_2170),
.Y(n_2235)
);

INVx1_ASAP7_75t_SL g2236 ( 
.A(n_2218),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2190),
.Y(n_2237)
);

NAND2x1p5_ASAP7_75t_L g2238 ( 
.A(n_2205),
.B(n_2134),
.Y(n_2238)
);

OAI22xp5_ASAP7_75t_L g2239 ( 
.A1(n_2218),
.A2(n_2167),
.B1(n_2036),
.B2(n_2171),
.Y(n_2239)
);

OAI32xp33_ASAP7_75t_L g2240 ( 
.A1(n_2212),
.A2(n_2143),
.A3(n_2135),
.B1(n_2148),
.B2(n_2182),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_2184),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2194),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2194),
.Y(n_2243)
);

OAI21xp5_ASAP7_75t_L g2244 ( 
.A1(n_2221),
.A2(n_2171),
.B(n_2121),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2213),
.B(n_2135),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2222),
.B(n_2143),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2222),
.B(n_2151),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2208),
.B(n_2148),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2198),
.Y(n_2249)
);

OAI221xp5_ASAP7_75t_L g2250 ( 
.A1(n_2199),
.A2(n_2104),
.B1(n_2096),
.B2(n_2165),
.C(n_2153),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2196),
.B(n_2206),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_2184),
.Y(n_2252)
);

INVx1_ASAP7_75t_SL g2253 ( 
.A(n_2224),
.Y(n_2253)
);

OAI21xp33_ASAP7_75t_L g2254 ( 
.A1(n_2220),
.A2(n_2163),
.B(n_2153),
.Y(n_2254)
);

AOI31xp33_ASAP7_75t_L g2255 ( 
.A1(n_2236),
.A2(n_2253),
.A3(n_2197),
.B(n_2235),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2225),
.B(n_2196),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2249),
.Y(n_2257)
);

OAI21xp5_ASAP7_75t_SL g2258 ( 
.A1(n_2226),
.A2(n_2197),
.B(n_2205),
.Y(n_2258)
);

AOI22xp5_ASAP7_75t_L g2259 ( 
.A1(n_2238),
.A2(n_2204),
.B1(n_2184),
.B2(n_2215),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_2225),
.B(n_2202),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2245),
.B(n_2235),
.Y(n_2261)
);

AOI32xp33_ASAP7_75t_L g2262 ( 
.A1(n_2250),
.A2(n_2200),
.A3(n_2219),
.B1(n_2207),
.B2(n_2198),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2249),
.Y(n_2263)
);

NOR3xp33_ASAP7_75t_L g2264 ( 
.A(n_2240),
.B(n_2210),
.C(n_2207),
.Y(n_2264)
);

INVx1_ASAP7_75t_SL g2265 ( 
.A(n_2231),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2228),
.Y(n_2266)
);

OR2x2_ASAP7_75t_L g2267 ( 
.A(n_2246),
.B(n_2200),
.Y(n_2267)
);

OR2x2_ASAP7_75t_L g2268 ( 
.A(n_2248),
.B(n_2219),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_2240),
.B(n_2251),
.Y(n_2269)
);

OAI211xp5_ASAP7_75t_SL g2270 ( 
.A1(n_2227),
.A2(n_2214),
.B(n_2211),
.C(n_2210),
.Y(n_2270)
);

AOI21xp33_ASAP7_75t_SL g2271 ( 
.A1(n_2238),
.A2(n_2197),
.B(n_2209),
.Y(n_2271)
);

AND2x4_ASAP7_75t_L g2272 ( 
.A(n_2231),
.B(n_2191),
.Y(n_2272)
);

INVx1_ASAP7_75t_SL g2273 ( 
.A(n_2247),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2229),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2238),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2241),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2230),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2276),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2276),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_SL g2280 ( 
.A(n_2264),
.B(n_2244),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_2272),
.Y(n_2281)
);

OAI22xp5_ASAP7_75t_L g2282 ( 
.A1(n_2269),
.A2(n_2167),
.B1(n_2239),
.B2(n_2195),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_SL g2283 ( 
.A(n_2264),
.B(n_2134),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2267),
.Y(n_2284)
);

INVx3_ASAP7_75t_L g2285 ( 
.A(n_2272),
.Y(n_2285)
);

OR2x2_ASAP7_75t_L g2286 ( 
.A(n_2265),
.B(n_2273),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2260),
.B(n_2247),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2256),
.Y(n_2288)
);

INVx1_ASAP7_75t_SL g2289 ( 
.A(n_2268),
.Y(n_2289)
);

OAI22xp33_ASAP7_75t_L g2290 ( 
.A1(n_2258),
.A2(n_2252),
.B1(n_2241),
.B2(n_2243),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2257),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2263),
.Y(n_2292)
);

AOI21xp33_ASAP7_75t_L g2293 ( 
.A1(n_2290),
.A2(n_2269),
.B(n_2275),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2286),
.Y(n_2294)
);

AOI221xp5_ASAP7_75t_L g2295 ( 
.A1(n_2280),
.A2(n_2262),
.B1(n_2275),
.B2(n_2270),
.C(n_2255),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_2285),
.B(n_2261),
.Y(n_2296)
);

OR2x6_ASAP7_75t_L g2297 ( 
.A(n_2278),
.B(n_2266),
.Y(n_2297)
);

OAI211xp5_ASAP7_75t_L g2298 ( 
.A1(n_2280),
.A2(n_2271),
.B(n_2270),
.C(n_2259),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2287),
.Y(n_2299)
);

NAND3xp33_ASAP7_75t_L g2300 ( 
.A(n_2283),
.B(n_2233),
.C(n_2274),
.Y(n_2300)
);

AOI221xp5_ASAP7_75t_L g2301 ( 
.A1(n_2290),
.A2(n_2277),
.B1(n_2232),
.B2(n_2242),
.C(n_2237),
.Y(n_2301)
);

AOI21xp5_ASAP7_75t_L g2302 ( 
.A1(n_2283),
.A2(n_2234),
.B(n_2252),
.Y(n_2302)
);

O2A1O1Ixp33_ASAP7_75t_L g2303 ( 
.A1(n_2289),
.A2(n_2211),
.B(n_2214),
.C(n_2254),
.Y(n_2303)
);

AOI211xp5_ASAP7_75t_L g2304 ( 
.A1(n_2282),
.A2(n_2209),
.B(n_2191),
.C(n_2195),
.Y(n_2304)
);

NOR3x1_ASAP7_75t_L g2305 ( 
.A(n_2284),
.B(n_2165),
.C(n_2160),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2296),
.B(n_2285),
.Y(n_2306)
);

AOI221xp5_ASAP7_75t_L g2307 ( 
.A1(n_2293),
.A2(n_2279),
.B1(n_2291),
.B2(n_2292),
.C(n_2288),
.Y(n_2307)
);

AOI211xp5_ASAP7_75t_L g2308 ( 
.A1(n_2298),
.A2(n_2281),
.B(n_2209),
.C(n_2187),
.Y(n_2308)
);

AOI21xp5_ASAP7_75t_L g2309 ( 
.A1(n_2295),
.A2(n_2302),
.B(n_2300),
.Y(n_2309)
);

AOI221xp5_ASAP7_75t_L g2310 ( 
.A1(n_2303),
.A2(n_2204),
.B1(n_2215),
.B2(n_2223),
.C(n_2172),
.Y(n_2310)
);

AOI21xp5_ASAP7_75t_L g2311 ( 
.A1(n_2301),
.A2(n_2209),
.B(n_2204),
.Y(n_2311)
);

AOI32xp33_ASAP7_75t_L g2312 ( 
.A1(n_2294),
.A2(n_2223),
.A3(n_2188),
.B1(n_2189),
.B2(n_2187),
.Y(n_2312)
);

AOI221xp5_ASAP7_75t_L g2313 ( 
.A1(n_2299),
.A2(n_2172),
.B1(n_2104),
.B2(n_2107),
.C(n_2102),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2297),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2305),
.B(n_2202),
.Y(n_2315)
);

OAI211xp5_ASAP7_75t_L g2316 ( 
.A1(n_2309),
.A2(n_2307),
.B(n_2306),
.C(n_2308),
.Y(n_2316)
);

AOI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_2315),
.A2(n_2297),
.B1(n_2304),
.B2(n_2189),
.Y(n_2317)
);

NOR2x1_ASAP7_75t_L g2318 ( 
.A(n_2314),
.B(n_2185),
.Y(n_2318)
);

CKINVDCx20_ASAP7_75t_R g2319 ( 
.A(n_2311),
.Y(n_2319)
);

AND5x1_ASAP7_75t_L g2320 ( 
.A(n_2312),
.B(n_2061),
.C(n_2054),
.D(n_2080),
.E(n_2185),
.Y(n_2320)
);

OAI211xp5_ASAP7_75t_L g2321 ( 
.A1(n_2310),
.A2(n_2188),
.B(n_2216),
.C(n_2163),
.Y(n_2321)
);

AOI21xp5_ASAP7_75t_L g2322 ( 
.A1(n_2313),
.A2(n_2216),
.B(n_2169),
.Y(n_2322)
);

AOI221xp5_ASAP7_75t_L g2323 ( 
.A1(n_2309),
.A2(n_2091),
.B1(n_2102),
.B2(n_2093),
.C(n_2107),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2306),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2318),
.Y(n_2325)
);

AOI22xp33_ASAP7_75t_L g2326 ( 
.A1(n_2319),
.A2(n_2021),
.B1(n_2072),
.B2(n_2085),
.Y(n_2326)
);

O2A1O1Ixp33_ASAP7_75t_L g2327 ( 
.A1(n_2316),
.A2(n_2179),
.B(n_2091),
.C(n_2093),
.Y(n_2327)
);

OAI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_2317),
.A2(n_2179),
.B1(n_2177),
.B2(n_2157),
.Y(n_2328)
);

NAND2x1p5_ASAP7_75t_L g2329 ( 
.A(n_2324),
.B(n_2320),
.Y(n_2329)
);

AND2x4_ASAP7_75t_L g2330 ( 
.A(n_2322),
.B(n_2176),
.Y(n_2330)
);

OR2x2_ASAP7_75t_L g2331 ( 
.A(n_2325),
.B(n_2321),
.Y(n_2331)
);

OR3x1_ASAP7_75t_L g2332 ( 
.A(n_2328),
.B(n_2323),
.C(n_2071),
.Y(n_2332)
);

AND2x4_ASAP7_75t_L g2333 ( 
.A(n_2330),
.B(n_2121),
.Y(n_2333)
);

NOR2x1_ASAP7_75t_L g2334 ( 
.A(n_2327),
.B(n_2111),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2332),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2335),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2336),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2336),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2337),
.Y(n_2339)
);

OAI22xp5_ASAP7_75t_SL g2340 ( 
.A1(n_2338),
.A2(n_2331),
.B1(n_2329),
.B2(n_2333),
.Y(n_2340)
);

AOI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_2339),
.A2(n_2334),
.B1(n_2326),
.B2(n_2111),
.Y(n_2341)
);

AOI22xp33_ASAP7_75t_SL g2342 ( 
.A1(n_2340),
.A2(n_2072),
.B1(n_2085),
.B2(n_2123),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_SL g2343 ( 
.A(n_2342),
.B(n_2072),
.Y(n_2343)
);

OAI21xp5_ASAP7_75t_L g2344 ( 
.A1(n_2343),
.A2(n_2341),
.B(n_2118),
.Y(n_2344)
);

XNOR2xp5_ASAP7_75t_L g2345 ( 
.A(n_2344),
.B(n_1921),
.Y(n_2345)
);

OAI221xp5_ASAP7_75t_R g2346 ( 
.A1(n_2345),
.A2(n_2072),
.B1(n_2118),
.B2(n_2108),
.C(n_2098),
.Y(n_2346)
);

AOI211xp5_ASAP7_75t_L g2347 ( 
.A1(n_2346),
.A2(n_2085),
.B(n_2080),
.C(n_2074),
.Y(n_2347)
);


endmodule