module real_jpeg_29375_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_0),
.B(n_107),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_3),
.A2(n_24),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_3),
.A2(n_22),
.B1(n_40),
.B2(n_43),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

AOI21xp33_ASAP7_75t_SL g19 ( 
.A1(n_4),
.A2(n_20),
.B(n_22),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_4),
.A2(n_17),
.B1(n_29),
.B2(n_30),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_4),
.A2(n_17),
.B1(n_24),
.B2(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_4),
.B(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_4),
.A2(n_17),
.B1(n_22),
.B2(n_43),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_4),
.A2(n_30),
.B(n_54),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_4),
.B(n_42),
.Y(n_100)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_8),
.A2(n_22),
.B1(n_43),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_8),
.A2(n_24),
.B1(n_41),
.B2(n_60),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_60),
.Y(n_79)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_9),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_88),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_87),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_61),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_14),
.B(n_61),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_36),
.C(n_49),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_15),
.B(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_16),
.B(n_27),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B(n_19),
.C(n_24),
.Y(n_16)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_17),
.A2(n_22),
.B(n_53),
.C(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_17),
.B(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_17),
.B(n_33),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_18),
.A2(n_20),
.B1(n_22),
.B2(n_43),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_18),
.A2(n_24),
.B(n_42),
.C(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_22),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_22),
.A2(n_43),
.B1(n_53),
.B2(n_54),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_24),
.B(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_24),
.A2(n_41),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_32),
.B(n_34),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_28),
.B(n_34),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_28),
.B(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_29),
.A2(n_30),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_29),
.B(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_32),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_32),
.B(n_34),
.Y(n_105)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_36),
.A2(n_37),
.B1(n_49),
.B2(n_50),
.Y(n_133)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_44),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_56),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_51),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_52),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_52),
.B(n_59),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_55),
.B(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_84),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_80),
.B2(n_81),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_77),
.B(n_112),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_106),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_130),
.B(n_134),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_108),
.B(n_129),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_91),
.B(n_97),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_104),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_102),
.C(n_104),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_118),
.B(n_128),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_116),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_110),
.B(n_116),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_123),
.B(n_127),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_120),
.B(n_122),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_131),
.B(n_132),
.Y(n_134)
);


endmodule