module fake_ibex_1786_n_1223 (n_151, n_147, n_85, n_167, n_128, n_208, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_201, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_215, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_214, n_79, n_81, n_35, n_159, n_202, n_158, n_211, n_132, n_174, n_210, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_207, n_54, n_19, n_1223);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_215;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_214;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_158;
input n_211;
input n_132;
input n_174;
input n_210;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_207;
input n_54;
input n_19;

output n_1223;

wire n_1084;
wire n_599;
wire n_822;
wire n_778;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1104;
wire n_1148;
wire n_992;
wire n_1011;
wire n_756;
wire n_529;
wire n_389;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_1090;
wire n_1110;
wire n_946;
wire n_1196;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_1182;
wire n_926;
wire n_1097;
wire n_1079;
wire n_1031;
wire n_1143;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_418;
wire n_256;
wire n_510;
wire n_845;
wire n_947;
wire n_981;
wire n_972;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_1080;
wire n_1162;
wire n_1199;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_1125;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_1152;
wire n_371;
wire n_1036;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_457;
wire n_412;
wire n_357;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1018;
wire n_1044;
wire n_1106;
wire n_1129;
wire n_449;
wire n_1131;
wire n_547;
wire n_1134;
wire n_727;
wire n_1138;
wire n_1077;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_1174;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1217;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_1147;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_1098;
wire n_377;
wire n_584;
wire n_1189;
wire n_647;
wire n_531;
wire n_1187;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_698;
wire n_901;
wire n_1096;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_1218;
wire n_1166;
wire n_1181;
wire n_1140;
wire n_327;
wire n_326;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_1144;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_1010;
wire n_1203;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_470;
wire n_276;
wire n_339;
wire n_770;
wire n_965;
wire n_348;
wire n_1109;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_1112;
wire n_1053;
wire n_1207;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_469;
wire n_323;
wire n_829;
wire n_1172;
wire n_1099;
wire n_598;
wire n_825;
wire n_740;
wire n_1169;
wire n_386;
wire n_549;
wire n_224;
wire n_1210;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_928;
wire n_655;
wire n_333;
wire n_898;
wire n_967;
wire n_1201;
wire n_400;
wire n_306;
wire n_550;
wire n_736;
wire n_1055;
wire n_673;
wire n_732;
wire n_832;
wire n_798;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_641;
wire n_557;
wire n_1103;
wire n_1161;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1177;
wire n_1068;
wire n_325;
wire n_301;
wire n_617;
wire n_496;
wire n_434;
wire n_1184;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_1195;
wire n_929;
wire n_604;
wire n_441;
wire n_315;
wire n_1024;
wire n_637;
wire n_1141;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_1075;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_1197;
wire n_574;
wire n_1168;
wire n_289;
wire n_716;
wire n_865;
wire n_1130;
wire n_1049;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_1179;
wire n_1192;
wire n_933;
wire n_1081;
wire n_1153;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_464;
wire n_669;
wire n_538;
wire n_838;
wire n_987;
wire n_1155;
wire n_750;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_1117;
wire n_1191;
wire n_1101;
wire n_518;
wire n_367;
wire n_221;
wire n_1052;
wire n_852;
wire n_789;
wire n_1133;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_1178;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_636;
wire n_594;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_1211;
wire n_570;
wire n_1116;
wire n_623;
wire n_585;
wire n_1030;
wire n_1094;
wire n_1020;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_1214;
wire n_420;
wire n_580;
wire n_483;
wire n_543;
wire n_487;
wire n_769;
wire n_1082;
wire n_222;
wire n_1137;
wire n_660;
wire n_1213;
wire n_524;
wire n_349;
wire n_857;
wire n_849;
wire n_765;
wire n_1070;
wire n_454;
wire n_1193;
wire n_1074;
wire n_777;
wire n_1200;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_1120;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_1180;
wire n_619;
wire n_1089;
wire n_536;
wire n_1124;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_1220;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_1064;
wire n_1071;
wire n_922;
wire n_1171;
wire n_438;
wire n_851;
wire n_1028;
wire n_1012;
wire n_993;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_1183;
wire n_253;
wire n_234;
wire n_1204;
wire n_300;
wire n_1151;
wire n_1135;
wire n_973;
wire n_1146;
wire n_358;
wire n_771;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_1038;
wire n_999;
wire n_1092;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_589;
wire n_648;
wire n_229;
wire n_472;
wire n_571;
wire n_783;
wire n_347;
wire n_1062;
wire n_847;
wire n_830;
wire n_1142;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_1215;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1173;
wire n_1069;
wire n_573;
wire n_1208;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_1007;
wire n_1126;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_837;
wire n_796;
wire n_797;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_699;
wire n_1063;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_1115;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1100;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_553;
wire n_554;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_1219;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_1170;
wire n_605;
wire n_539;
wire n_392;
wire n_354;
wire n_630;
wire n_567;
wire n_548;
wire n_516;
wire n_943;
wire n_1057;
wire n_1158;
wire n_763;
wire n_1086;
wire n_745;
wire n_329;
wire n_1149;
wire n_447;
wire n_1176;
wire n_940;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_788;
wire n_1202;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_1160;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_1216;
wire n_1222;
wire n_397;
wire n_283;
wire n_366;
wire n_803;
wire n_894;
wire n_1033;
wire n_1118;
wire n_692;
wire n_627;
wire n_990;
wire n_1198;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_1087;
wire n_757;
wire n_248;
wire n_702;
wire n_712;
wire n_451;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_1114;
wire n_409;
wire n_1093;
wire n_582;
wire n_978;
wire n_818;
wire n_1167;
wire n_653;
wire n_1205;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_1190;
wire n_517;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_1107;
wire n_223;
wire n_381;
wire n_1073;
wire n_1108;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_980;
wire n_681;
wire n_633;
wire n_1209;
wire n_1111;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_379;
wire n_320;
wire n_1128;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_440;
wire n_268;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_1145;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_1113;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_1164;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_1175;
wire n_485;
wire n_1139;
wire n_870;
wire n_1221;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_1212;
wire n_461;
wire n_575;
wire n_313;
wire n_1159;
wire n_1119;
wire n_903;
wire n_1154;
wire n_519;
wire n_345;
wire n_408;
wire n_1085;
wire n_361;
wire n_1095;
wire n_455;
wire n_1136;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_1091;
wire n_885;
wire n_513;
wire n_588;
wire n_877;
wire n_1121;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_1088;
wire n_896;
wire n_528;
wire n_1005;
wire n_1102;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_1150;
wire n_462;
wire n_1194;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_1165;
wire n_1185;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_1122;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_912;
wire n_874;
wire n_890;
wire n_921;
wire n_1105;
wire n_1058;
wire n_1163;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_1123;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_1000;
wire n_394;
wire n_984;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_231;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_1157;
wire n_751;
wire n_806;
wire n_1127;
wire n_932;
wire n_1186;
wire n_657;
wire n_764;
wire n_1156;
wire n_1206;
wire n_492;
wire n_649;
wire n_855;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

INVx1_ASAP7_75t_L g216 ( 
.A(n_61),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_115),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_80),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_12),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_36),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_124),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_117),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_102),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_38),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_63),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_75),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_96),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_71),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_127),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_89),
.Y(n_233)
);

NOR2xp67_ASAP7_75t_L g234 ( 
.A(n_100),
.B(n_155),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_193),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_46),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_74),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_153),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_26),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_60),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_162),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_16),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_99),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_116),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_55),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_187),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_104),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_56),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_171),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_134),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_90),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_76),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_18),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_137),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_94),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_93),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_205),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_113),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_11),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_58),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_95),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_182),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_146),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_161),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_87),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_107),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_135),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_210),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_72),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_65),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_27),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_154),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_106),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_152),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_142),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_40),
.Y(n_277)
);

INVxp33_ASAP7_75t_L g278 ( 
.A(n_145),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_42),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_8),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_16),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_81),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_194),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_3),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_36),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_212),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_44),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_130),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_82),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_120),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_163),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_37),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_52),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_207),
.Y(n_294)
);

BUFx2_ASAP7_75t_SL g295 ( 
.A(n_62),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_33),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_141),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_17),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_199),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_70),
.Y(n_300)
);

INVxp33_ASAP7_75t_L g301 ( 
.A(n_200),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_39),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_13),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_147),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_189),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_59),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_174),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_101),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_118),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_9),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_138),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_78),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_122),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_144),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_149),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_123),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_167),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_6),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_32),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_211),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_180),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_77),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_140),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_6),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_169),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_192),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_23),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_64),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_214),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_35),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_208),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_150),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_4),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_139),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_131),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_178),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_18),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_19),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_37),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_168),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_195),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_54),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_2),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_165),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_191),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_108),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_85),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_42),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_132),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_121),
.Y(n_350)
);

NOR2xp67_ASAP7_75t_L g351 ( 
.A(n_119),
.B(n_83),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_51),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_13),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_166),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_1),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_188),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_133),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_190),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_24),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_105),
.Y(n_360)
);

BUFx10_ASAP7_75t_L g361 ( 
.A(n_179),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_202),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_47),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_112),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_38),
.B(n_57),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_157),
.Y(n_366)
);

INVxp33_ASAP7_75t_L g367 ( 
.A(n_143),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_40),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_88),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_198),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_151),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_110),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_148),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_3),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_183),
.Y(n_375)
);

BUFx10_ASAP7_75t_L g376 ( 
.A(n_44),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_164),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_175),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_28),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_186),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_172),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_69),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_48),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_125),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_97),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_197),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_84),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_8),
.Y(n_388)
);

BUFx10_ASAP7_75t_L g389 ( 
.A(n_136),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_215),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_66),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_267),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_293),
.B(n_0),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_293),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_277),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_368),
.Y(n_396)
);

OAI21x1_ASAP7_75t_L g397 ( 
.A1(n_227),
.A2(n_111),
.B(n_213),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_272),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_227),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_262),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_278),
.B(n_0),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_300),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_235),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_272),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_314),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_296),
.Y(n_406)
);

BUFx12f_ASAP7_75t_L g407 ( 
.A(n_240),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_250),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_277),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_278),
.B(n_1),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_310),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_277),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_296),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_277),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_342),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_342),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_280),
.B(n_5),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_379),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_285),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_330),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_262),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_268),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_333),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_251),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_379),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_379),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_280),
.B(n_340),
.Y(n_428)
);

BUFx8_ASAP7_75t_SL g429 ( 
.A(n_285),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_370),
.B(n_10),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_379),
.Y(n_431)
);

INVx5_ASAP7_75t_L g432 ( 
.A(n_240),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_221),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_301),
.B(n_11),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_268),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_376),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_251),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_274),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_222),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_229),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_236),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_301),
.B(n_12),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_274),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_240),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_299),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_367),
.B(n_376),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_219),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_367),
.B(n_14),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_244),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_226),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_299),
.Y(n_452)
);

BUFx8_ASAP7_75t_SL g453 ( 
.A(n_324),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_317),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_275),
.B(n_15),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_229),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_375),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_375),
.Y(n_458)
);

BUFx12f_ASAP7_75t_L g459 ( 
.A(n_244),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_239),
.B(n_19),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_317),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_245),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_321),
.Y(n_463)
);

OAI22x1_ASAP7_75t_SL g464 ( 
.A1(n_324),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_244),
.B(n_20),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_321),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_307),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_343),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_378),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_378),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_307),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_286),
.B(n_24),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_383),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_284),
.B(n_25),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_242),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_307),
.B(n_25),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_302),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_361),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_216),
.Y(n_479)
);

OAI21x1_ASAP7_75t_L g480 ( 
.A1(n_218),
.A2(n_126),
.B(n_206),
.Y(n_480)
);

INVx5_ASAP7_75t_L g481 ( 
.A(n_361),
.Y(n_481)
);

BUFx12f_ASAP7_75t_L g482 ( 
.A(n_361),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_303),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_389),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_337),
.B(n_30),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_254),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_220),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_279),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_224),
.A2(n_128),
.B(n_204),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_352),
.B(n_353),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_355),
.B(n_31),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_230),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_389),
.B(n_32),
.Y(n_493)
);

INVx6_ASAP7_75t_L g494 ( 
.A(n_389),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_363),
.B(n_33),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_231),
.A2(n_129),
.B(n_196),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_304),
.B(n_34),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_374),
.B(n_34),
.Y(n_498)
);

INVx4_ASAP7_75t_L g499 ( 
.A(n_217),
.Y(n_499)
);

BUFx8_ASAP7_75t_L g500 ( 
.A(n_237),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_241),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_243),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_246),
.B(n_35),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_463),
.Y(n_504)
);

AO21x2_ASAP7_75t_L g505 ( 
.A1(n_397),
.A2(n_249),
.B(n_247),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_430),
.B(n_252),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_418),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_450),
.B(n_255),
.Y(n_508)
);

AND3x2_ASAP7_75t_L g509 ( 
.A(n_394),
.B(n_318),
.C(n_292),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_463),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_440),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_447),
.B(n_294),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_428),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_450),
.B(n_259),
.Y(n_514)
);

BUFx6f_ASAP7_75t_SL g515 ( 
.A(n_418),
.Y(n_515)
);

NOR2x1p5_ASAP7_75t_L g516 ( 
.A(n_407),
.B(n_281),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_433),
.Y(n_517)
);

NAND3xp33_ASAP7_75t_L g518 ( 
.A(n_410),
.B(n_327),
.C(n_298),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_418),
.Y(n_519)
);

BUFx6f_ASAP7_75t_SL g520 ( 
.A(n_445),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_433),
.Y(n_521)
);

BUFx6f_ASAP7_75t_SL g522 ( 
.A(n_445),
.Y(n_522)
);

AO21x2_ASAP7_75t_L g523 ( 
.A1(n_397),
.A2(n_264),
.B(n_263),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_441),
.Y(n_524)
);

OR2x6_ASAP7_75t_L g525 ( 
.A(n_407),
.B(n_295),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_474),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_484),
.B(n_382),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_474),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_463),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_485),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_466),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_425),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_485),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_467),
.B(n_269),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_466),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_498),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_432),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_466),
.Y(n_538)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_396),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_470),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_449),
.Y(n_541)
);

INVxp33_ASAP7_75t_L g542 ( 
.A(n_475),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_470),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_470),
.Y(n_544)
);

NOR2x1p5_ASAP7_75t_L g545 ( 
.A(n_459),
.B(n_338),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_479),
.B(n_276),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_SL g547 ( 
.A(n_393),
.B(n_253),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_441),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_406),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_432),
.B(n_339),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_414),
.Y(n_551)
);

BUFx10_ASAP7_75t_L g552 ( 
.A(n_438),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_416),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_494),
.Y(n_554)
);

INVx8_ASAP7_75t_L g555 ( 
.A(n_459),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_479),
.B(n_288),
.Y(n_556)
);

OAI22xp33_ASAP7_75t_L g557 ( 
.A1(n_411),
.A2(n_319),
.B1(n_287),
.B2(n_260),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_417),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_479),
.B(n_290),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_428),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_456),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_456),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_457),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_487),
.Y(n_564)
);

AO21x2_ASAP7_75t_L g565 ( 
.A1(n_480),
.A2(n_316),
.B(n_308),
.Y(n_565)
);

BUFx10_ASAP7_75t_L g566 ( 
.A(n_438),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_475),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_442),
.B(n_348),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_486),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_487),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_398),
.B(n_365),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_432),
.B(n_359),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_487),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_467),
.B(n_322),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_457),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_457),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_471),
.B(n_325),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_487),
.B(n_326),
.Y(n_578)
);

CKINVDCx6p67_ASAP7_75t_R g579 ( 
.A(n_482),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_486),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_398),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_457),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_412),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_492),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_471),
.B(n_329),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_478),
.B(n_334),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_395),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_395),
.Y(n_588)
);

BUFx10_ASAP7_75t_L g589 ( 
.A(n_494),
.Y(n_589)
);

BUFx16f_ASAP7_75t_R g590 ( 
.A(n_429),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_478),
.B(n_335),
.Y(n_591)
);

AO22x2_ASAP7_75t_L g592 ( 
.A1(n_451),
.A2(n_384),
.B1(n_381),
.B2(n_372),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_392),
.A2(n_253),
.B1(n_364),
.B2(n_258),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_L g594 ( 
.A(n_432),
.B(n_391),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_399),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_501),
.B(n_336),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_488),
.B(n_388),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_409),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_409),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_481),
.B(n_499),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_409),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_420),
.Y(n_602)
);

INVxp33_ASAP7_75t_SL g603 ( 
.A(n_403),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_488),
.B(n_223),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_494),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_481),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_409),
.Y(n_607)
);

AO21x2_ASAP7_75t_L g608 ( 
.A1(n_489),
.A2(n_350),
.B(n_349),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_502),
.B(n_354),
.Y(n_609)
);

AND2x2_ASAP7_75t_SL g610 ( 
.A(n_465),
.B(n_356),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_413),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_399),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_400),
.Y(n_613)
);

CKINVDCx11_ASAP7_75t_R g614 ( 
.A(n_473),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_400),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_422),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_412),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_402),
.A2(n_328),
.B1(n_258),
.B2(n_266),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_458),
.Y(n_619)
);

OAI21xp33_ASAP7_75t_SL g620 ( 
.A1(n_401),
.A2(n_360),
.B(n_357),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_423),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_436),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_436),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_421),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_502),
.B(n_362),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_413),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_439),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_408),
.Y(n_628)
);

BUFx16f_ASAP7_75t_R g629 ( 
.A(n_429),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_453),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_L g631 ( 
.A(n_481),
.B(n_390),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_415),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_415),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_421),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_415),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_408),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_405),
.A2(n_266),
.B1(n_283),
.B2(n_309),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_439),
.Y(n_638)
);

AND3x2_ASAP7_75t_L g639 ( 
.A(n_476),
.B(n_309),
.C(n_283),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_419),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_482),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_444),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_434),
.Y(n_643)
);

NOR2x1p5_ASAP7_75t_L g644 ( 
.A(n_434),
.B(n_437),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_437),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_419),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_499),
.B(n_225),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_446),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_581),
.B(n_404),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_555),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_583),
.B(n_448),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_617),
.B(n_462),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_539),
.B(n_493),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_513),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_624),
.B(n_634),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_541),
.B(n_435),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_560),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_624),
.B(n_490),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_512),
.B(n_443),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_619),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_634),
.B(n_500),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_515),
.A2(n_401),
.B1(n_503),
.B2(n_455),
.Y(n_662)
);

O2A1O1Ixp5_ASAP7_75t_L g663 ( 
.A1(n_506),
.A2(n_455),
.B(n_497),
.C(n_472),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_645),
.B(n_500),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_643),
.B(n_472),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_643),
.B(n_497),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_589),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_555),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_567),
.B(n_460),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_642),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_511),
.B(n_491),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_526),
.B(n_495),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_589),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_L g674 ( 
.A(n_555),
.B(n_528),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_549),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_551),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_553),
.Y(n_677)
);

OR2x6_ASAP7_75t_L g678 ( 
.A(n_525),
.B(n_468),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_569),
.B(n_228),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_580),
.B(n_232),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_558),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_530),
.B(n_452),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_580),
.B(n_233),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_527),
.B(n_238),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_554),
.B(n_257),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_595),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_508),
.B(n_248),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_568),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_604),
.B(n_256),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_612),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_613),
.Y(n_691)
);

NAND3xp33_ASAP7_75t_L g692 ( 
.A(n_518),
.B(n_424),
.C(n_477),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_548),
.Y(n_693)
);

BUFx6f_ASAP7_75t_SL g694 ( 
.A(n_641),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_615),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_616),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_533),
.B(n_454),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_621),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_622),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_514),
.B(n_261),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_536),
.B(n_454),
.Y(n_701)
);

INVx4_ASAP7_75t_L g702 ( 
.A(n_520),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_623),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_542),
.B(n_420),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_620),
.B(n_265),
.Y(n_705)
);

NOR2xp67_ASAP7_75t_L g706 ( 
.A(n_593),
.B(n_618),
.Y(n_706)
);

INVxp67_ASAP7_75t_SL g707 ( 
.A(n_542),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_507),
.B(n_461),
.Y(n_708)
);

AOI221xp5_ASAP7_75t_L g709 ( 
.A1(n_557),
.A2(n_483),
.B1(n_464),
.B2(n_461),
.C(n_469),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_597),
.B(n_473),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_519),
.B(n_469),
.Y(n_711)
);

OAI221xp5_ASAP7_75t_L g712 ( 
.A1(n_514),
.A2(n_306),
.B1(n_270),
.B2(n_271),
.C(n_273),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_537),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_534),
.B(n_282),
.Y(n_714)
);

NOR2x1p5_ASAP7_75t_L g715 ( 
.A(n_579),
.B(n_453),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_605),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_574),
.B(n_577),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_636),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_627),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_610),
.B(n_289),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_638),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_506),
.B(n_496),
.Y(n_722)
);

NAND3xp33_ASAP7_75t_L g723 ( 
.A(n_509),
.B(n_345),
.C(n_305),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_610),
.B(n_291),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_525),
.B(n_328),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_647),
.B(n_297),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_522),
.B(n_311),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_522),
.B(n_312),
.Y(n_728)
);

NOR3xp33_ASAP7_75t_L g729 ( 
.A(n_547),
.B(n_371),
.C(n_313),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_647),
.B(n_315),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_525),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_648),
.Y(n_732)
);

BUFx8_ASAP7_75t_L g733 ( 
.A(n_590),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_585),
.B(n_320),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_547),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_515),
.A2(n_347),
.B1(n_364),
.B2(n_331),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_586),
.B(n_323),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_637),
.A2(n_347),
.B1(n_332),
.B2(n_341),
.Y(n_738)
);

OAI221xp5_ASAP7_75t_L g739 ( 
.A1(n_586),
.A2(n_373),
.B1(n_344),
.B2(n_346),
.C(n_387),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_628),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_L g741 ( 
.A(n_509),
.B(n_377),
.C(n_358),
.Y(n_741)
);

OR2x6_ASAP7_75t_L g742 ( 
.A(n_516),
.B(n_234),
.Y(n_742)
);

INVx5_ASAP7_75t_L g743 ( 
.A(n_537),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_517),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_591),
.B(n_366),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_591),
.B(n_369),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_571),
.Y(n_747)
);

INVx8_ASAP7_75t_L g748 ( 
.A(n_532),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_552),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_550),
.B(n_572),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_592),
.A2(n_385),
.B1(n_380),
.B2(n_386),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_552),
.B(n_39),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_609),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_566),
.B(n_351),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_600),
.B(n_596),
.Y(n_755)
);

BUFx5_ASAP7_75t_L g756 ( 
.A(n_564),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_521),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_609),
.B(n_426),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_625),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_625),
.B(n_426),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_603),
.B(n_67),
.Y(n_761)
);

NAND2xp33_ASAP7_75t_L g762 ( 
.A(n_606),
.B(n_427),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_505),
.B(n_427),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_505),
.B(n_427),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_722),
.A2(n_523),
.B(n_565),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_653),
.B(n_639),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_671),
.B(n_740),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_722),
.A2(n_523),
.B(n_565),
.Y(n_768)
);

AOI21x1_ASAP7_75t_L g769 ( 
.A1(n_763),
.A2(n_556),
.B(n_546),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_656),
.B(n_644),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_749),
.B(n_545),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_656),
.B(n_524),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_743),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_672),
.A2(n_592),
.B1(n_578),
.B2(n_556),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_748),
.Y(n_775)
);

AO21x1_ASAP7_75t_L g776 ( 
.A1(n_763),
.A2(n_573),
.B(n_570),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_717),
.A2(n_608),
.B(n_559),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_707),
.B(n_614),
.Y(n_778)
);

BUFx4f_ASAP7_75t_L g779 ( 
.A(n_748),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_688),
.A2(n_706),
.B1(n_735),
.B2(n_669),
.Y(n_780)
);

NOR2xp67_ASAP7_75t_L g781 ( 
.A(n_702),
.B(n_630),
.Y(n_781)
);

A2O1A1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_663),
.A2(n_594),
.B(n_631),
.C(n_584),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_675),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_659),
.A2(n_540),
.B(n_504),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_755),
.A2(n_666),
.B(n_665),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_658),
.B(n_651),
.Y(n_786)
);

A2O1A1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_652),
.A2(n_576),
.B(n_575),
.C(n_563),
.Y(n_787)
);

AO21x1_ASAP7_75t_L g788 ( 
.A1(n_764),
.A2(n_562),
.B(n_561),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_750),
.A2(n_764),
.B(n_682),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_743),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_743),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_657),
.B(n_524),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_692),
.A2(n_602),
.B1(n_614),
.B2(n_582),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_676),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_677),
.B(n_41),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_681),
.B(n_43),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_708),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_729),
.A2(n_535),
.B1(n_510),
.B2(n_529),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_718),
.B(n_629),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_662),
.B(n_43),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_753),
.A2(n_529),
.B(n_531),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_708),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_711),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_654),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_697),
.A2(n_538),
.B(n_540),
.Y(n_805)
);

OAI21xp33_ASAP7_75t_L g806 ( 
.A1(n_679),
.A2(n_680),
.B(n_664),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_697),
.A2(n_701),
.B(n_711),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_720),
.B(n_45),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_704),
.B(n_45),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_701),
.A2(n_543),
.B(n_544),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_661),
.B(n_46),
.Y(n_811)
);

INVxp67_ASAP7_75t_SL g812 ( 
.A(n_650),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_725),
.B(n_47),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_668),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_686),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_736),
.A2(n_431),
.B1(n_646),
.B2(n_640),
.Y(n_816)
);

BUFx2_ASAP7_75t_SL g817 ( 
.A(n_694),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_746),
.B(n_48),
.Y(n_818)
);

O2A1O1Ixp5_ASAP7_75t_L g819 ( 
.A1(n_705),
.A2(n_754),
.B(n_730),
.C(n_726),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_690),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_684),
.A2(n_611),
.B(n_640),
.Y(n_821)
);

O2A1O1Ixp33_ASAP7_75t_SL g822 ( 
.A1(n_758),
.A2(n_760),
.B(n_700),
.C(n_714),
.Y(n_822)
);

NOR3xp33_ASAP7_75t_L g823 ( 
.A(n_709),
.B(n_632),
.C(n_588),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_L g824 ( 
.A1(n_759),
.A2(n_607),
.B(n_635),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_691),
.A2(n_607),
.B(n_633),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_724),
.B(n_49),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_695),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_689),
.B(n_50),
.Y(n_828)
);

CKINVDCx10_ASAP7_75t_R g829 ( 
.A(n_694),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_687),
.A2(n_601),
.B(n_587),
.Y(n_830)
);

CKINVDCx10_ASAP7_75t_R g831 ( 
.A(n_678),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_696),
.Y(n_832)
);

AO21x1_ASAP7_75t_L g833 ( 
.A1(n_751),
.A2(n_632),
.B(n_598),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_698),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_699),
.A2(n_599),
.B(n_588),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_751),
.A2(n_598),
.B(n_599),
.C(n_626),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_655),
.B(n_703),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_748),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_SL g839 ( 
.A1(n_725),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_731),
.B(n_53),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_683),
.B(n_53),
.Y(n_841)
);

NAND3xp33_ASAP7_75t_SL g842 ( 
.A(n_710),
.B(n_752),
.C(n_712),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_719),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_713),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_660),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_738),
.B(n_55),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_667),
.B(n_673),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_738),
.B(n_68),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_721),
.B(n_73),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_732),
.B(n_79),
.Y(n_850)
);

OR2x2_ASAP7_75t_SL g851 ( 
.A(n_733),
.B(n_86),
.Y(n_851)
);

BUFx12f_ASAP7_75t_L g852 ( 
.A(n_715),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_716),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_747),
.A2(n_91),
.B(n_92),
.C(n_98),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_678),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_670),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_649),
.B(n_103),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_734),
.A2(n_109),
.B(n_114),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_737),
.A2(n_745),
.B1(n_739),
.B2(n_761),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_674),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_693),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_727),
.B(n_728),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_822),
.A2(n_757),
.B(n_744),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_767),
.B(n_685),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_768),
.A2(n_741),
.B(n_723),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_777),
.A2(n_762),
.B(n_742),
.Y(n_866)
);

OAI21xp33_ASAP7_75t_L g867 ( 
.A1(n_786),
.A2(n_742),
.B(n_756),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_780),
.B(n_733),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_775),
.Y(n_869)
);

OAI22x1_ASAP7_75t_L g870 ( 
.A1(n_846),
.A2(n_848),
.B1(n_855),
.B2(n_813),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_802),
.B(n_803),
.Y(n_871)
);

OA22x2_ASAP7_75t_L g872 ( 
.A1(n_793),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_766),
.A2(n_160),
.B1(n_170),
.B2(n_173),
.Y(n_873)
);

AOI221xp5_ASAP7_75t_SL g874 ( 
.A1(n_836),
.A2(n_177),
.B1(n_181),
.B2(n_184),
.C(n_185),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_794),
.B(n_770),
.Y(n_875)
);

AND2x6_ASAP7_75t_L g876 ( 
.A(n_773),
.B(n_790),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_779),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_829),
.Y(n_878)
);

BUFx5_ASAP7_75t_L g879 ( 
.A(n_856),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_815),
.B(n_820),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_779),
.Y(n_881)
);

OAI21x1_ASAP7_75t_L g882 ( 
.A1(n_801),
.A2(n_824),
.B(n_825),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_774),
.A2(n_784),
.B(n_782),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_827),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_832),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_834),
.A2(n_843),
.B(n_837),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_805),
.A2(n_810),
.B(n_858),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_838),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_857),
.A2(n_862),
.B1(n_809),
.B2(n_859),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_795),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_842),
.B(n_828),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_831),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_796),
.A2(n_811),
.B1(n_818),
.B2(n_800),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_773),
.Y(n_894)
);

OAI21x1_ASAP7_75t_L g895 ( 
.A1(n_824),
.A2(n_825),
.B(n_835),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_841),
.A2(n_808),
.B(n_826),
.C(n_823),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_860),
.B(n_812),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_769),
.A2(n_787),
.B(n_835),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_849),
.A2(n_850),
.B(n_830),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_778),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_804),
.B(n_840),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_814),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_821),
.A2(n_772),
.B(n_792),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_853),
.B(n_839),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_771),
.B(n_790),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_791),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_852),
.Y(n_907)
);

OAI21x1_ASAP7_75t_L g908 ( 
.A1(n_798),
.A2(n_819),
.B(n_844),
.Y(n_908)
);

AO31x2_ASAP7_75t_L g909 ( 
.A1(n_816),
.A2(n_845),
.A3(n_861),
.B(n_851),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_847),
.A2(n_771),
.B(n_781),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_799),
.A2(n_845),
.B(n_861),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_845),
.B(n_817),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_767),
.B(n_725),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_783),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_779),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_806),
.A2(n_785),
.B(n_807),
.C(n_663),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_806),
.A2(n_785),
.B(n_807),
.C(n_663),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_767),
.B(n_541),
.Y(n_918)
);

BUFx2_ASAP7_75t_L g919 ( 
.A(n_779),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_775),
.B(n_749),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_767),
.B(n_541),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_806),
.A2(n_785),
.B(n_807),
.C(n_663),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_765),
.A2(n_768),
.B(n_789),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_806),
.A2(n_785),
.B(n_807),
.C(n_663),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_767),
.B(n_541),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_779),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_822),
.A2(n_785),
.B(n_777),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_767),
.B(n_653),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_767),
.B(n_653),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_822),
.A2(n_785),
.B(n_777),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_806),
.A2(n_785),
.B(n_807),
.C(n_663),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_767),
.B(n_541),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_767),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_783),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_767),
.B(n_541),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_822),
.A2(n_785),
.B(n_777),
.Y(n_936)
);

AO21x1_ASAP7_75t_L g937 ( 
.A1(n_765),
.A2(n_768),
.B(n_854),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_822),
.A2(n_785),
.B(n_777),
.Y(n_938)
);

NAND2x1p5_ASAP7_75t_L g939 ( 
.A(n_779),
.B(n_775),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_767),
.B(n_541),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_767),
.B(n_541),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_767),
.B(n_541),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_765),
.A2(n_768),
.B(n_789),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_838),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_797),
.A2(n_803),
.B1(n_802),
.B2(n_786),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_SL g946 ( 
.A1(n_846),
.A2(n_725),
.B1(n_420),
.B2(n_738),
.Y(n_946)
);

AO31x2_ASAP7_75t_L g947 ( 
.A1(n_788),
.A2(n_833),
.A3(n_776),
.B(n_768),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_767),
.B(n_541),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_829),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_767),
.B(n_541),
.Y(n_950)
);

AO31x2_ASAP7_75t_L g951 ( 
.A1(n_788),
.A2(n_833),
.A3(n_776),
.B(n_768),
.Y(n_951)
);

OAI21xp33_ASAP7_75t_SL g952 ( 
.A1(n_797),
.A2(n_803),
.B(n_802),
.Y(n_952)
);

AND3x4_ASAP7_75t_L g953 ( 
.A(n_781),
.B(n_629),
.C(n_590),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_767),
.B(n_541),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_767),
.B(n_653),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_767),
.B(n_541),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_767),
.B(n_653),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_822),
.A2(n_785),
.B(n_777),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_767),
.B(n_541),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_767),
.B(n_541),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_765),
.A2(n_768),
.B(n_789),
.Y(n_961)
);

OA21x2_ASAP7_75t_L g962 ( 
.A1(n_765),
.A2(n_768),
.B(n_764),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_829),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_806),
.A2(n_785),
.B(n_807),
.C(n_663),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_767),
.B(n_653),
.Y(n_965)
);

AO21x2_ASAP7_75t_L g966 ( 
.A1(n_765),
.A2(n_768),
.B(n_788),
.Y(n_966)
);

NOR2x1_ASAP7_75t_SL g967 ( 
.A(n_945),
.B(n_871),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_885),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_877),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_928),
.B(n_929),
.Y(n_970)
);

AOI21xp33_ASAP7_75t_L g971 ( 
.A1(n_889),
.A2(n_952),
.B(n_893),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_952),
.A2(n_930),
.B(n_927),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_869),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_881),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_915),
.B(n_919),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_939),
.Y(n_976)
);

AO31x2_ASAP7_75t_L g977 ( 
.A1(n_937),
.A2(n_958),
.A3(n_936),
.B(n_938),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_955),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_944),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_920),
.Y(n_980)
);

OA21x2_ASAP7_75t_L g981 ( 
.A1(n_923),
.A2(n_961),
.B(n_943),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_916),
.A2(n_922),
.B(n_917),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_926),
.B(n_920),
.Y(n_983)
);

NOR2x1_ASAP7_75t_R g984 ( 
.A(n_878),
.B(n_949),
.Y(n_984)
);

CKINVDCx16_ASAP7_75t_R g985 ( 
.A(n_907),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_888),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_905),
.B(n_886),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_957),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_963),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_965),
.Y(n_990)
);

BUFx8_ASAP7_75t_L g991 ( 
.A(n_900),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_914),
.Y(n_992)
);

BUFx4f_ASAP7_75t_L g993 ( 
.A(n_953),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_884),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_869),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_886),
.B(n_912),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_934),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_924),
.A2(n_931),
.B(n_964),
.Y(n_998)
);

OA21x2_ASAP7_75t_L g999 ( 
.A1(n_874),
.A2(n_883),
.B(n_887),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_913),
.B(n_933),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_876),
.Y(n_1001)
);

OA21x2_ASAP7_75t_L g1002 ( 
.A1(n_874),
.A2(n_883),
.B(n_887),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_912),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_946),
.A2(n_870),
.B1(n_891),
.B2(n_890),
.Y(n_1004)
);

OA21x2_ASAP7_75t_L g1005 ( 
.A1(n_898),
.A2(n_882),
.B(n_899),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_880),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_895),
.A2(n_896),
.B(n_898),
.Y(n_1007)
);

CKINVDCx20_ASAP7_75t_R g1008 ( 
.A(n_892),
.Y(n_1008)
);

BUFx8_ASAP7_75t_L g1009 ( 
.A(n_902),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_876),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_876),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_865),
.A2(n_893),
.B(n_908),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_906),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_SL g1014 ( 
.A1(n_911),
.A2(n_866),
.B(n_901),
.Y(n_1014)
);

AO21x2_ASAP7_75t_L g1015 ( 
.A1(n_966),
.A2(n_903),
.B(n_863),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_876),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_918),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_921),
.Y(n_1018)
);

OR2x6_ASAP7_75t_L g1019 ( 
.A(n_910),
.B(n_894),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_894),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_925),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_864),
.A2(n_904),
.B1(n_868),
.B2(n_875),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_932),
.Y(n_1023)
);

INVxp67_ASAP7_75t_SL g1024 ( 
.A(n_962),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_935),
.Y(n_1025)
);

INVxp67_ASAP7_75t_SL g1026 ( 
.A(n_879),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_940),
.B(n_960),
.Y(n_1027)
);

OR2x6_ASAP7_75t_L g1028 ( 
.A(n_910),
.B(n_959),
.Y(n_1028)
);

NAND2x1p5_ASAP7_75t_L g1029 ( 
.A(n_941),
.B(n_942),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_948),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_879),
.B(n_867),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_867),
.A2(n_897),
.B(n_872),
.Y(n_1032)
);

AND2x2_ASAP7_75t_SL g1033 ( 
.A(n_873),
.B(n_909),
.Y(n_1033)
);

NAND2x1p5_ASAP7_75t_L g1034 ( 
.A(n_950),
.B(n_954),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_879),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_956),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_947),
.A2(n_951),
.B(n_909),
.Y(n_1037)
);

BUFx10_ASAP7_75t_L g1038 ( 
.A(n_878),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_SL g1039 ( 
.A(n_952),
.B(n_945),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_928),
.B(n_767),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_928),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_945),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_928),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_928),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_928),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1024),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_1010),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_SL g1048 ( 
.A1(n_1039),
.A2(n_967),
.B1(n_1042),
.B2(n_991),
.Y(n_1048)
);

BUFx8_ASAP7_75t_L g1049 ( 
.A(n_979),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1024),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_973),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1026),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1006),
.B(n_968),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_1004),
.A2(n_1042),
.B1(n_971),
.B2(n_1028),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_994),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_989),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_981),
.Y(n_1057)
);

CKINVDCx11_ASAP7_75t_R g1058 ( 
.A(n_1038),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_989),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_997),
.Y(n_1060)
);

AO21x2_ASAP7_75t_L g1061 ( 
.A1(n_982),
.A2(n_998),
.B(n_972),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_1035),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1014),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1004),
.A2(n_971),
.B1(n_1036),
.B2(n_1022),
.Y(n_1064)
);

CKINVDCx9p33_ASAP7_75t_R g1065 ( 
.A(n_986),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_992),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_996),
.B(n_987),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_977),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_987),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_SL g1070 ( 
.A1(n_1039),
.A2(n_991),
.B1(n_1030),
.B2(n_996),
.Y(n_1070)
);

OAI222xp33_ASAP7_75t_L g1071 ( 
.A1(n_1028),
.A2(n_1022),
.B1(n_1034),
.B2(n_1029),
.C1(n_1030),
.C2(n_973),
.Y(n_1071)
);

OAI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_1029),
.A2(n_1034),
.B1(n_1028),
.B2(n_1036),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_974),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_978),
.B(n_988),
.Y(n_1074)
);

OA21x2_ASAP7_75t_L g1075 ( 
.A1(n_1012),
.A2(n_1037),
.B(n_1007),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_1000),
.A2(n_1045),
.B1(n_990),
.B2(n_1041),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1000),
.A2(n_1027),
.B1(n_1018),
.B2(n_1021),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_1043),
.A2(n_1044),
.B1(n_970),
.B2(n_1023),
.Y(n_1078)
);

BUFx4f_ASAP7_75t_L g1079 ( 
.A(n_1001),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1067),
.B(n_1002),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1061),
.B(n_1002),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_1062),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_1074),
.B(n_1040),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1046),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1057),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1064),
.B(n_1032),
.Y(n_1086)
);

INVx5_ASAP7_75t_L g1087 ( 
.A(n_1047),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1064),
.B(n_1055),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_1046),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_1065),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1055),
.B(n_1032),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_1062),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1050),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_1047),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1050),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1061),
.B(n_999),
.Y(n_1096)
);

OR2x2_ASAP7_75t_L g1097 ( 
.A(n_1069),
.B(n_1013),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1061),
.B(n_1005),
.Y(n_1098)
);

INVx5_ASAP7_75t_L g1099 ( 
.A(n_1047),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1077),
.A2(n_1070),
.B1(n_1048),
.B2(n_1054),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1063),
.B(n_1031),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1077),
.A2(n_1019),
.B1(n_1033),
.B2(n_1025),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1068),
.B(n_1015),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1067),
.B(n_1033),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_SL g1105 ( 
.A1(n_1056),
.A2(n_1008),
.B1(n_985),
.B2(n_974),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_1052),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1080),
.B(n_1075),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1080),
.B(n_1104),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1084),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1104),
.B(n_1075),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1088),
.B(n_1060),
.Y(n_1111)
);

INVxp67_ASAP7_75t_L g1112 ( 
.A(n_1083),
.Y(n_1112)
);

OR2x2_ASAP7_75t_L g1113 ( 
.A(n_1089),
.B(n_1092),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1088),
.B(n_1060),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1084),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1098),
.B(n_1075),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1093),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1098),
.B(n_1075),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1085),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_1092),
.Y(n_1120)
);

INVxp67_ASAP7_75t_L g1121 ( 
.A(n_1089),
.Y(n_1121)
);

INVxp67_ASAP7_75t_SL g1122 ( 
.A(n_1082),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_SL g1123 ( 
.A(n_1090),
.B(n_1071),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1095),
.B(n_1106),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_1105),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1101),
.B(n_1063),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1106),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1108),
.B(n_1081),
.Y(n_1128)
);

INVxp67_ASAP7_75t_L g1129 ( 
.A(n_1120),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1108),
.B(n_1081),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_1126),
.B(n_1103),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_1113),
.B(n_1091),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1119),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1110),
.B(n_1096),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_1113),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1109),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1125),
.B(n_1105),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1111),
.B(n_1051),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1110),
.B(n_1096),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1109),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_1124),
.B(n_1091),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1115),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1131),
.B(n_1126),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1134),
.B(n_1107),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1135),
.Y(n_1145)
);

OR2x2_ASAP7_75t_L g1146 ( 
.A(n_1128),
.B(n_1121),
.Y(n_1146)
);

NOR2x1_ASAP7_75t_L g1147 ( 
.A(n_1137),
.B(n_1090),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1133),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_1135),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1134),
.B(n_1139),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1136),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_1139),
.B(n_1116),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1136),
.Y(n_1153)
);

INVxp67_ASAP7_75t_L g1154 ( 
.A(n_1135),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1128),
.B(n_1130),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1130),
.B(n_1107),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1141),
.B(n_1138),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1150),
.B(n_1129),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1151),
.B(n_1141),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1153),
.B(n_1132),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1145),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1145),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1150),
.B(n_1132),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1143),
.B(n_1131),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1143),
.B(n_1131),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_1152),
.B(n_1116),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1147),
.A2(n_1100),
.B(n_1123),
.Y(n_1167)
);

AO221x1_ASAP7_75t_L g1168 ( 
.A1(n_1149),
.A2(n_1154),
.B1(n_1100),
.B2(n_1121),
.C(n_1102),
.Y(n_1168)
);

OAI221xp5_ASAP7_75t_L g1169 ( 
.A1(n_1157),
.A2(n_1123),
.B1(n_1112),
.B2(n_993),
.C(n_1114),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1143),
.B(n_1152),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1155),
.B(n_1118),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1167),
.A2(n_1146),
.B1(n_1144),
.B2(n_1156),
.Y(n_1172)
);

OAI21xp33_ASAP7_75t_L g1173 ( 
.A1(n_1167),
.A2(n_1131),
.B(n_1126),
.Y(n_1173)
);

NAND2x1p5_ASAP7_75t_L g1174 ( 
.A(n_1164),
.B(n_993),
.Y(n_1174)
);

XOR2x2_ASAP7_75t_L g1175 ( 
.A(n_1158),
.B(n_1058),
.Y(n_1175)
);

OAI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1166),
.A2(n_1094),
.B1(n_1087),
.B2(n_1099),
.Y(n_1176)
);

AO22x1_ASAP7_75t_L g1177 ( 
.A1(n_1164),
.A2(n_1049),
.B1(n_1059),
.B2(n_1122),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1169),
.A2(n_1073),
.B(n_1072),
.Y(n_1178)
);

AOI211xp5_ASAP7_75t_L g1179 ( 
.A1(n_1177),
.A2(n_1168),
.B(n_984),
.C(n_1102),
.Y(n_1179)
);

AOI22x1_ASAP7_75t_L g1180 ( 
.A1(n_1174),
.A2(n_1170),
.B1(n_1161),
.B2(n_1162),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1172),
.A2(n_1159),
.B1(n_1160),
.B2(n_1163),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1173),
.B(n_1159),
.Y(n_1182)
);

OAI211xp5_ASAP7_75t_L g1183 ( 
.A1(n_1178),
.A2(n_1008),
.B(n_1076),
.C(n_1078),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1176),
.A2(n_1160),
.B1(n_1165),
.B2(n_1171),
.Y(n_1184)
);

INVxp67_ASAP7_75t_L g1185 ( 
.A(n_1175),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1172),
.B(n_1140),
.Y(n_1186)
);

OAI21xp33_ASAP7_75t_L g1187 ( 
.A1(n_1182),
.A2(n_1114),
.B(n_1111),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1181),
.B(n_1140),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1186),
.B(n_1142),
.Y(n_1189)
);

OAI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_1179),
.A2(n_1086),
.B1(n_1124),
.B2(n_1142),
.C(n_1148),
.Y(n_1190)
);

NOR4xp25_ASAP7_75t_L g1191 ( 
.A(n_1185),
.B(n_1074),
.C(n_1066),
.D(n_995),
.Y(n_1191)
);

AOI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1183),
.A2(n_1049),
.B1(n_1126),
.B2(n_1086),
.Y(n_1192)
);

OAI322xp33_ASAP7_75t_L g1193 ( 
.A1(n_1184),
.A2(n_1127),
.A3(n_1148),
.B1(n_1097),
.B2(n_1051),
.C1(n_1115),
.C2(n_1117),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1180),
.A2(n_1094),
.B(n_1087),
.Y(n_1194)
);

NOR3xp33_ASAP7_75t_L g1195 ( 
.A(n_1190),
.B(n_984),
.C(n_969),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1189),
.Y(n_1196)
);

NAND3xp33_ASAP7_75t_L g1197 ( 
.A(n_1192),
.B(n_1049),
.C(n_1009),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_SL g1198 ( 
.A(n_1194),
.B(n_1038),
.Y(n_1198)
);

NOR3x1_ASAP7_75t_L g1199 ( 
.A(n_1188),
.B(n_1049),
.C(n_976),
.Y(n_1199)
);

NOR2x1_ASAP7_75t_L g1200 ( 
.A(n_1193),
.B(n_1016),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1187),
.B(n_1009),
.Y(n_1201)
);

NOR2xp67_ASAP7_75t_L g1202 ( 
.A(n_1196),
.B(n_1191),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1201),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1198),
.A2(n_1079),
.B(n_983),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1195),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1199),
.B(n_1118),
.Y(n_1206)
);

NAND4xp75_ASAP7_75t_L g1207 ( 
.A(n_1200),
.B(n_1003),
.C(n_1017),
.D(n_1053),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1197),
.B(n_983),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1202),
.B(n_1127),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1203),
.Y(n_1210)
);

NOR4xp25_ASAP7_75t_L g1211 ( 
.A(n_1205),
.B(n_1013),
.C(n_1066),
.D(n_1053),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1210),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1209),
.B(n_1208),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1212),
.B(n_1206),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1213),
.Y(n_1215)
);

XOR2xp5_ASAP7_75t_L g1216 ( 
.A(n_1215),
.B(n_1208),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1216),
.B(n_1214),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1216),
.A2(n_1214),
.B1(n_1213),
.B2(n_1204),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1218),
.A2(n_1207),
.B1(n_1211),
.B2(n_1079),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1219),
.A2(n_1217),
.B(n_975),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1220),
.Y(n_1221)
);

XOR2xp5_ASAP7_75t_L g1222 ( 
.A(n_1221),
.B(n_975),
.Y(n_1222)
);

AOI211xp5_ASAP7_75t_L g1223 ( 
.A1(n_1222),
.A2(n_980),
.B(n_1011),
.C(n_1020),
.Y(n_1223)
);


endmodule