module fake_jpeg_32016_n_548 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_548);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_548;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_52),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_59),
.B(n_65),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_11),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_66),
.Y(n_108)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_62),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_11),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_9),
.B(n_2),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_95),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_74),
.Y(n_160)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_79),
.Y(n_163)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_83),
.Y(n_165)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_85),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_86),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_9),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

HAxp5_ASAP7_75t_SL g100 ( 
.A(n_22),
.B(n_18),
.CON(n_100),
.SN(n_100)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_21),
.B1(n_46),
.B2(n_40),
.Y(n_124)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_25),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_48),
.B1(n_36),
.B2(n_34),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_109),
.A2(n_125),
.B1(n_130),
.B2(n_158),
.Y(n_184)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_95),
.B(n_21),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_118),
.B(n_124),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_89),
.A2(n_48),
.B1(n_36),
.B2(n_34),
.Y(n_125)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_48),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_129),
.B(n_132),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_36),
.B1(n_34),
.B2(n_26),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_54),
.A2(n_26),
.B1(n_22),
.B2(n_51),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_131),
.A2(n_140),
.B1(n_0),
.B2(n_3),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_53),
.B(n_26),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_102),
.A2(n_51),
.B1(n_46),
.B2(n_21),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_96),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_150),
.B(n_156),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_52),
.B(n_22),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_154),
.B(n_157),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_53),
.B(n_33),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_67),
.B(n_33),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_55),
.A2(n_51),
.B1(n_46),
.B2(n_40),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_82),
.A2(n_39),
.B1(n_37),
.B2(n_35),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_23),
.B1(n_37),
.B2(n_30),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_108),
.A2(n_74),
.B1(n_77),
.B2(n_57),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_169),
.Y(n_269)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

INVx3_ASAP7_75t_SL g247 ( 
.A(n_171),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_115),
.B(n_35),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_172),
.B(n_181),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_173),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_106),
.A2(n_71),
.B1(n_99),
.B2(n_93),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_174),
.A2(n_225),
.B1(n_229),
.B2(n_14),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

INVx11_ASAP7_75t_L g234 ( 
.A(n_176),
.Y(n_234)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_177),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_110),
.A2(n_86),
.B1(n_64),
.B2(n_35),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_178),
.A2(n_190),
.B1(n_193),
.B2(n_210),
.Y(n_244)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_179),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_114),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_180),
.B(n_187),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_124),
.B(n_20),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

A2O1A1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_124),
.A2(n_62),
.B(n_40),
.C(n_39),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_183),
.B(n_162),
.Y(n_231)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_185),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_108),
.A2(n_140),
.B1(n_130),
.B2(n_123),
.Y(n_186)
);

OR2x4_ASAP7_75t_L g276 ( 
.A(n_186),
.B(n_205),
.Y(n_276)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_116),
.A2(n_23),
.A3(n_30),
.B1(n_37),
.B2(n_39),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_188),
.A2(n_198),
.B1(n_206),
.B2(n_222),
.Y(n_251)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_189),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_110),
.A2(n_20),
.B1(n_30),
.B2(n_23),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_135),
.Y(n_191)
);

INVx11_ASAP7_75t_L g271 ( 
.A(n_191),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_165),
.A2(n_20),
.B1(n_70),
.B2(n_92),
.Y(n_193)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_145),
.Y(n_194)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_194),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_120),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_195),
.Y(n_272)
);

INVx11_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_196),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_125),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_197),
.B(n_203),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_109),
.A2(n_72),
.B1(n_63),
.B2(n_91),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_128),
.B(n_68),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_212),
.Y(n_236)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_138),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_200),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_201),
.Y(n_264)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_202),
.Y(n_266)
);

INVx4_ASAP7_75t_SL g203 ( 
.A(n_113),
.Y(n_203)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_111),
.Y(n_204)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_151),
.A2(n_33),
.B1(n_25),
.B2(n_42),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_158),
.A2(n_87),
.B1(n_79),
.B2(n_104),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_111),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_209),
.Y(n_253)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_133),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_166),
.Y(n_209)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_148),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_152),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_214),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_25),
.Y(n_212)
);

AOI21xp33_ASAP7_75t_L g213 ( 
.A1(n_127),
.A2(n_25),
.B(n_2),
.Y(n_213)
);

OR2x2_ASAP7_75t_SL g273 ( 
.A(n_213),
.B(n_0),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_160),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_113),
.A2(n_25),
.B(n_42),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_230),
.B(n_119),
.Y(n_233)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_161),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_217),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_135),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_218),
.A2(n_224),
.B1(n_148),
.B2(n_159),
.Y(n_246)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_107),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_219),
.B(n_220),
.Y(n_280)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_134),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_155),
.B(n_25),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_226),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_136),
.A2(n_97),
.B1(n_25),
.B2(n_42),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_137),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_160),
.B(n_12),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_136),
.A2(n_42),
.B1(n_3),
.B2(n_4),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_227),
.A2(n_141),
.B1(n_112),
.B2(n_153),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_163),
.A2(n_42),
.B1(n_3),
.B2(n_6),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_142),
.B1(n_141),
.B2(n_149),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_163),
.A2(n_42),
.B1(n_3),
.B2(n_6),
.Y(n_229)
);

NAND2x2_ASAP7_75t_SL g230 ( 
.A(n_151),
.B(n_0),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_231),
.A2(n_273),
.B(n_215),
.Y(n_295)
);

AND2x2_ASAP7_75t_SL g300 ( 
.A(n_233),
.B(n_189),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_246),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_216),
.B(n_133),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_250),
.B(n_219),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_181),
.B(n_159),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_255),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_170),
.B(n_226),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_230),
.A2(n_162),
.B1(n_120),
.B2(n_119),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_256),
.A2(n_259),
.B1(n_268),
.B2(n_279),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_212),
.B(n_147),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_258),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_175),
.B(n_142),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_230),
.A2(n_184),
.B1(n_203),
.B2(n_112),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_192),
.B(n_147),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_260),
.B(n_267),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_261),
.A2(n_278),
.B1(n_218),
.B2(n_191),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_262),
.A2(n_206),
.B1(n_198),
.B2(n_229),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_175),
.B(n_144),
.C(n_107),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_265),
.B(n_171),
.C(n_217),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_175),
.B(n_164),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_230),
.A2(n_144),
.B1(n_7),
.B2(n_8),
.Y(n_268)
);

O2A1O1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_183),
.A2(n_13),
.B(n_7),
.C(n_8),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_277),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_194),
.A2(n_14),
.B1(n_7),
.B2(n_9),
.Y(n_279)
);

AOI22x1_ASAP7_75t_L g281 ( 
.A1(n_186),
.A2(n_15),
.B1(n_12),
.B2(n_13),
.Y(n_281)
);

OA22x2_ASAP7_75t_L g302 ( 
.A1(n_281),
.A2(n_210),
.B1(n_204),
.B2(n_207),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_201),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_282),
.A2(n_208),
.B1(n_179),
.B2(n_176),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_199),
.B(n_0),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_283),
.B(n_17),
.Y(n_325)
);

OAI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_285),
.A2(n_296),
.B1(n_302),
.B2(n_288),
.Y(n_347)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_240),
.Y(n_286)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_286),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_232),
.B(n_255),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_287),
.B(n_235),
.C(n_272),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_251),
.A2(n_225),
.B1(n_169),
.B2(n_221),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_288),
.A2(n_298),
.B1(n_313),
.B2(n_316),
.Y(n_339)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_249),
.Y(n_289)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_289),
.Y(n_333)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_250),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_291),
.B(n_327),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_254),
.B(n_223),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_292),
.B(n_294),
.Y(n_345)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_249),
.Y(n_293)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_293),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_172),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_295),
.B(n_304),
.Y(n_356)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_266),
.Y(n_297)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_297),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_251),
.A2(n_187),
.B1(n_205),
.B2(n_185),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_266),
.Y(n_299)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_299),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_300),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_301),
.Y(n_370)
);

OAI21xp33_ASAP7_75t_SL g358 ( 
.A1(n_302),
.A2(n_241),
.B(n_264),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_305),
.A2(n_311),
.B1(n_257),
.B2(n_274),
.Y(n_338)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_280),
.Y(n_306)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_306),
.Y(n_350)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_240),
.Y(n_308)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_308),
.Y(n_335)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_245),
.Y(n_309)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_309),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_310),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_231),
.A2(n_224),
.B1(n_220),
.B2(n_177),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_312),
.B(n_317),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_239),
.A2(n_173),
.B1(n_182),
.B2(n_196),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_247),
.Y(n_314)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_314),
.Y(n_351)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_270),
.Y(n_315)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_315),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_L g316 ( 
.A1(n_269),
.A2(n_195),
.B1(n_0),
.B2(n_15),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_238),
.B(n_14),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_247),
.Y(n_318)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_318),
.Y(n_359)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_241),
.Y(n_319)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_319),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_264),
.Y(n_320)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_320),
.Y(n_366)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_247),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_321),
.B(n_323),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_252),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_322),
.A2(n_275),
.B1(n_274),
.B2(n_234),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_238),
.B(n_16),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_325),
.B(n_326),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_236),
.B(n_17),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_272),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_245),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_328),
.B(n_329),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_270),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_236),
.B(n_17),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_330),
.B(n_331),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_248),
.B(n_283),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_303),
.A2(n_277),
.B(n_267),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_332),
.A2(n_372),
.B(n_316),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_285),
.A2(n_276),
.B1(n_244),
.B2(n_269),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_337),
.A2(n_338),
.B1(n_344),
.B2(n_347),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_305),
.A2(n_276),
.B1(n_253),
.B2(n_242),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_300),
.A2(n_295),
.B(n_324),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_346),
.A2(n_348),
.B(n_365),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_296),
.A2(n_258),
.B(n_265),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_324),
.A2(n_248),
.B1(n_232),
.B2(n_273),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_349),
.A2(n_353),
.B1(n_354),
.B2(n_358),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_307),
.A2(n_278),
.B1(n_281),
.B2(n_261),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_307),
.A2(n_290),
.B1(n_284),
.B2(n_311),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_362),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_284),
.A2(n_281),
.B1(n_237),
.B2(n_275),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_306),
.B(n_237),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_367),
.B(n_319),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_304),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_300),
.A2(n_243),
.B(n_263),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_340),
.Y(n_373)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_373),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_350),
.B(n_287),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_374),
.B(n_389),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_376),
.A2(n_366),
.B(n_357),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_330),
.Y(n_377)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_377),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_367),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_379),
.B(n_407),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_341),
.B(n_326),
.Y(n_380)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_380),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_339),
.A2(n_370),
.B1(n_332),
.B2(n_365),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_381),
.A2(n_385),
.B1(n_393),
.B2(n_351),
.Y(n_416)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_340),
.Y(n_382)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_382),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_346),
.A2(n_302),
.B(n_297),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_383),
.A2(n_391),
.B(n_392),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_394),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_339),
.A2(n_302),
.B1(n_331),
.B2(n_299),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_386),
.A2(n_387),
.B(n_402),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_372),
.A2(n_348),
.B(n_370),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_343),
.Y(n_388)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_388),
.Y(n_438)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_368),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_341),
.B(n_367),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_390),
.Y(n_408)
);

A2O1A1Ixp33_ASAP7_75t_SL g391 ( 
.A1(n_337),
.A2(n_329),
.B(n_321),
.C(n_318),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_344),
.A2(n_314),
.B(n_320),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_353),
.A2(n_325),
.B1(n_329),
.B2(n_293),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_356),
.B(n_322),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_369),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_395),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_350),
.B(n_289),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_396),
.B(n_403),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_356),
.B(n_328),
.C(n_315),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_397),
.B(n_399),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_309),
.C(n_286),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_369),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_400),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_401),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_360),
.A2(n_343),
.B(n_354),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_333),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_363),
.A2(n_310),
.B1(n_243),
.B2(n_308),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_404),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_349),
.B(n_263),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_405),
.B(n_364),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_333),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_406),
.B(n_336),
.Y(n_421)
);

AO22x1_ASAP7_75t_L g407 ( 
.A1(n_362),
.A2(n_263),
.B1(n_235),
.B2(n_243),
.Y(n_407)
);

FAx1_ASAP7_75t_SL g413 ( 
.A(n_390),
.B(n_338),
.CI(n_345),
.CON(n_413),
.SN(n_413)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_413),
.B(n_423),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_416),
.A2(n_418),
.B1(n_430),
.B2(n_434),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_385),
.A2(n_351),
.B1(n_359),
.B2(n_336),
.Y(n_418)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_421),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_398),
.A2(n_355),
.B1(n_359),
.B2(n_342),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_377),
.B(n_352),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_427),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_398),
.A2(n_378),
.B1(n_375),
.B2(n_392),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_407),
.Y(n_460)
);

INVxp33_ASAP7_75t_L g427 ( 
.A(n_401),
.Y(n_427)
);

INVxp33_ASAP7_75t_L g428 ( 
.A(n_379),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_432),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_381),
.A2(n_342),
.B1(n_357),
.B2(n_363),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_431),
.A2(n_383),
.B(n_386),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_380),
.B(n_366),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_393),
.A2(n_364),
.B1(n_334),
.B2(n_335),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_435),
.B(n_399),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_429),
.B(n_384),
.C(n_397),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_452),
.C(n_458),
.Y(n_469)
);

AO21x2_ASAP7_75t_L g441 ( 
.A1(n_419),
.A2(n_415),
.B(n_437),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_441),
.A2(n_453),
.B(n_463),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_442),
.Y(n_472)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_415),
.Y(n_444)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_444),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g485 ( 
.A(n_445),
.B(n_434),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_415),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_447),
.B(n_449),
.Y(n_487)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_409),
.Y(n_448)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_448),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_426),
.Y(n_449)
);

INVxp33_ASAP7_75t_L g450 ( 
.A(n_412),
.Y(n_450)
);

INVxp33_ASAP7_75t_L g474 ( 
.A(n_450),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_429),
.B(n_376),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_451),
.B(n_454),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_422),
.B(n_394),
.C(n_405),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_436),
.A2(n_387),
.B(n_378),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_422),
.B(n_402),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_437),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_456),
.A2(n_465),
.B1(n_417),
.B2(n_438),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_395),
.C(n_400),
.Y(n_458)
);

OAI22xp33_ASAP7_75t_R g459 ( 
.A1(n_414),
.A2(n_407),
.B1(n_391),
.B2(n_375),
.Y(n_459)
);

AOI21xp33_ASAP7_75t_L g480 ( 
.A1(n_459),
.A2(n_461),
.B(n_423),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_460),
.B(n_464),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_410),
.B(n_406),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_408),
.B(n_403),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_462),
.B(n_418),
.Y(n_483)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_409),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_436),
.B(n_391),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_431),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_443),
.A2(n_433),
.B(n_425),
.Y(n_466)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_466),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_439),
.B(n_430),
.C(n_425),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_475),
.C(n_479),
.Y(n_490)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_471),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_445),
.B(n_416),
.C(n_417),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_454),
.B(n_451),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_450),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_458),
.B(n_419),
.C(n_413),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_480),
.A2(n_484),
.B1(n_472),
.B2(n_446),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_452),
.B(n_411),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_481),
.B(n_482),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_411),
.Y(n_482)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_483),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_413),
.C(n_408),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_484),
.B(n_457),
.C(n_440),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_485),
.B(n_486),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_442),
.B(n_410),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_487),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_492),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_483),
.A2(n_455),
.B1(n_444),
.B2(n_433),
.Y(n_493)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_493),
.Y(n_510)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_473),
.Y(n_494)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_494),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_468),
.B(n_446),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_501),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_499),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_SL g516 ( 
.A(n_498),
.B(n_502),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_467),
.A2(n_455),
.B1(n_440),
.B2(n_441),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_468),
.B(n_462),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_477),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_503),
.A2(n_441),
.B(n_448),
.Y(n_506)
);

XNOR2x1_ASAP7_75t_L g504 ( 
.A(n_479),
.B(n_460),
.Y(n_504)
);

OAI21xp33_ASAP7_75t_SL g512 ( 
.A1(n_504),
.A2(n_474),
.B(n_482),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_506),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_490),
.B(n_470),
.C(n_469),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_507),
.B(n_509),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_490),
.B(n_469),
.C(n_475),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_501),
.A2(n_472),
.B(n_441),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_511),
.A2(n_512),
.B(n_517),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_500),
.A2(n_476),
.B1(n_486),
.B2(n_441),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_514),
.B(n_518),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_495),
.A2(n_476),
.B(n_474),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_488),
.A2(n_463),
.B1(n_481),
.B2(n_391),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_509),
.A2(n_499),
.B(n_504),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_520),
.B(n_524),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_505),
.B(n_502),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_522),
.B(n_523),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_494),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_513),
.B(n_496),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_511),
.A2(n_489),
.B(n_493),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_526),
.B(n_513),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_510),
.A2(n_488),
.B1(n_491),
.B2(n_391),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_527),
.B(n_514),
.C(n_518),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_529),
.B(n_530),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_519),
.B(n_507),
.C(n_508),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_532),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_528),
.B(n_515),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_534),
.A2(n_521),
.B(n_524),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_537),
.A2(n_516),
.B(n_525),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_533),
.A2(n_527),
.B1(n_420),
.B2(n_438),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_538),
.B(n_525),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_539),
.A2(n_535),
.B(n_489),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_536),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_541),
.A2(n_542),
.B1(n_516),
.B2(n_420),
.Y(n_543)
);

OAI31xp33_ASAP7_75t_L g544 ( 
.A1(n_543),
.A2(n_491),
.A3(n_485),
.B(n_373),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_544),
.A2(n_388),
.B(n_382),
.Y(n_545)
);

OAI21xp33_ASAP7_75t_L g546 ( 
.A1(n_545),
.A2(n_334),
.B(n_335),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_546),
.B(n_243),
.C(n_234),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_547),
.A2(n_271),
.B(n_541),
.Y(n_548)
);


endmodule