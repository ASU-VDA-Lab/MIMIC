module fake_jpeg_31606_n_118 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_20),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx9p33_ASAP7_75t_R g54 ( 
.A(n_53),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_SL g72 ( 
.A(n_54),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_53),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_58),
.Y(n_68)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_4),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_61),
.B(n_5),
.C(n_6),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_26),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_52),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_61)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_67),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_41),
.B(n_14),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_50),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_57),
.Y(n_81)
);

INVxp33_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_74),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_30),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_80),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_79),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_68),
.A2(n_47),
.B1(n_44),
.B2(n_40),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_57),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_43),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_83),
.C(n_16),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_9),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_35),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_96),
.C(n_39),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_94),
.B1(n_99),
.B2(n_36),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_29),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_97),
.A2(n_37),
.B(n_38),
.Y(n_104)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_104),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_91),
.C(n_95),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_90),
.B1(n_95),
.B2(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

AO221x1_ASAP7_75t_L g113 ( 
.A1(n_111),
.A2(n_108),
.B1(n_107),
.B2(n_106),
.C(n_109),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_102),
.C(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_112),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_115),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_77),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_88),
.Y(n_118)
);


endmodule