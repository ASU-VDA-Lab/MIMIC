module fake_jpeg_22999_n_244 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_244);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_244;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_47),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_33),
.Y(n_77)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_56),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_26),
.B(n_24),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_54),
.B(n_69),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_25),
.B1(n_22),
.B2(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_46),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_22),
.B1(n_25),
.B2(n_34),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_5),
.B(n_9),
.C(n_11),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_72),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_0),
.Y(n_88)
);

AO22x1_ASAP7_75t_L g68 ( 
.A1(n_36),
.A2(n_26),
.B1(n_24),
.B2(n_18),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_68),
.A2(n_15),
.B(n_62),
.C(n_61),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_37),
.A2(n_22),
.B1(n_25),
.B2(n_17),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_41),
.A2(n_17),
.B1(n_31),
.B2(n_18),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_30),
.B(n_28),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_40),
.A2(n_35),
.B1(n_33),
.B2(n_19),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_30),
.B1(n_28),
.B2(n_20),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_79),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_9),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_46),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_83),
.A2(n_84),
.B1(n_104),
.B2(n_98),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_21),
.B1(n_16),
.B2(n_2),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_97),
.B1(n_78),
.B2(n_57),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_21),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_21),
.C(n_16),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_56),
.C(n_63),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_21),
.B1(n_16),
.B2(n_3),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_90),
.A2(n_94),
.B(n_104),
.C(n_91),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_21),
.B1(n_16),
.B2(n_4),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_81),
.B1(n_55),
.B2(n_64),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_1),
.B(n_2),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_106),
.B(n_102),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_9),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_80),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_53),
.A2(n_12),
.B(n_13),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_74),
.B(n_79),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_51),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_104)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_110),
.Y(n_112)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_51),
.B(n_67),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_101),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_113),
.B(n_137),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_115),
.B1(n_120),
.B2(n_121),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_116),
.B(n_117),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_57),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_56),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_118),
.B(n_119),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_82),
.A2(n_89),
.B1(n_100),
.B2(n_90),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_87),
.B(n_76),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_126),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_76),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_123),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_82),
.A2(n_52),
.B1(n_64),
.B2(n_84),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_85),
.B1(n_99),
.B2(n_121),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_92),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_52),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_129),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_83),
.C(n_97),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_135),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_136),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_88),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_108),
.B(n_99),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_93),
.B(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_109),
.Y(n_152)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_113),
.Y(n_159)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_119),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_155),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_152),
.A2(n_163),
.B(n_150),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_108),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_158),
.Y(n_165)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_156),
.A2(n_134),
.B1(n_132),
.B2(n_127),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_161),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_85),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_159),
.B(n_153),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_126),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_160),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_131),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_164),
.Y(n_168)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_166),
.B(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_183),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_129),
.B1(n_114),
.B2(n_139),
.Y(n_172)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_115),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_142),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_135),
.B1(n_133),
.B2(n_124),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_174),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_135),
.B(n_133),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_176),
.A2(n_177),
.B(n_182),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_178),
.B(n_179),
.Y(n_196)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_145),
.B(n_144),
.CI(n_156),
.CON(n_179),
.SN(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_161),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_181),
.Y(n_194)
);

OA21x2_ASAP7_75t_L g182 ( 
.A1(n_151),
.A2(n_164),
.B(n_155),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_140),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_SL g184 ( 
.A1(n_177),
.A2(n_142),
.B(n_145),
.Y(n_184)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_184),
.B(n_182),
.CI(n_174),
.CON(n_208),
.SN(n_208)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_189),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_158),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_198),
.C(n_153),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_171),
.B(n_147),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_195),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_148),
.Y(n_193)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_162),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_172),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_167),
.C(n_165),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_175),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_202),
.A2(n_205),
.B(n_206),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_191),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_204),
.A2(n_210),
.B1(n_190),
.B2(n_194),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_182),
.B(n_168),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_208),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_170),
.B1(n_166),
.B2(n_178),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_209),
.A2(n_199),
.B1(n_197),
.B2(n_179),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_186),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_189),
.C(n_185),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_149),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_188),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_217),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_221),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_215),
.A2(n_222),
.B(n_218),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_204),
.B(n_146),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_201),
.B(n_212),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_219),
.B(n_200),
.Y(n_228)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_199),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_179),
.B1(n_181),
.B2(n_141),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_227),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_201),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g233 ( 
.A(n_225),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_216),
.A2(n_206),
.B1(n_202),
.B2(n_208),
.Y(n_227)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_209),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_207),
.Y(n_238)
);

OAI221xp5_ASAP7_75t_L g231 ( 
.A1(n_228),
.A2(n_220),
.B1(n_200),
.B2(n_208),
.C(n_211),
.Y(n_231)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_231),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_229),
.Y(n_235)
);

OAI21x1_ASAP7_75t_L g239 ( 
.A1(n_235),
.A2(n_233),
.B(n_221),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_234),
.A2(n_226),
.B1(n_214),
.B2(n_216),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_239),
.A2(n_236),
.B(n_235),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_242),
.B(n_243),
.CI(n_240),
.CON(n_244),
.SN(n_244)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_141),
.Y(n_243)
);


endmodule