module fake_jpeg_22497_n_35 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_35);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_35;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

INVx4_ASAP7_75t_SL g15 ( 
.A(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_2),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_8),
.A2(n_10),
.B1(n_3),
.B2(n_13),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_16),
.A2(n_0),
.B(n_1),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_23),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_18),
.A2(n_1),
.B(n_5),
.C(n_6),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_11),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_19),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_17),
.Y(n_31)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_24),
.C(n_26),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_30),
.C(n_24),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_33),
.A2(n_18),
.B(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);


endmodule