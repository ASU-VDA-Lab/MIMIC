module fake_jpeg_27788_n_106 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_21),
.Y(n_35)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_0),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_26),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_10),
.B(n_1),
.Y(n_26)
);

CKINVDCx9p33_ASAP7_75t_R g27 ( 
.A(n_20),
.Y(n_27)
);

CKINVDCx12_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_14),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_15),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_24),
.A2(n_12),
.B1(n_13),
.B2(n_18),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_22),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_11),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_10),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_44),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_12),
.B1(n_18),
.B2(n_11),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_46),
.B1(n_50),
.B2(n_20),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_31),
.B(n_17),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_29),
.A2(n_17),
.B(n_13),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_23),
.C(n_19),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_52),
.B(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_60),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_51),
.B1(n_44),
.B2(n_49),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_57),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_51),
.A2(n_24),
.B1(n_28),
.B2(n_22),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

AND2x6_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_9),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_1),
.C(n_2),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_22),
.B1(n_23),
.B2(n_19),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_40),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_38),
.B1(n_41),
.B2(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_66),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_48),
.A2(n_23),
.B1(n_15),
.B2(n_16),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_71),
.Y(n_79)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_39),
.B(n_4),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_75),
.Y(n_84)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_77),
.A2(n_66),
.B1(n_60),
.B2(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_81),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_61),
.B1(n_63),
.B2(n_53),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_57),
.B1(n_53),
.B2(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_16),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_23),
.C(n_37),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_70),
.C(n_15),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_80),
.A2(n_76),
.B1(n_72),
.B2(n_67),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_89),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_77),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_91),
.C(n_85),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_79),
.B(n_78),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_91),
.C(n_87),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_95),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_81),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_21),
.C(n_4),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_93),
.B(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_97),
.B(n_98),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_21),
.C(n_4),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_5),
.C(n_6),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_2),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_2),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_104),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_101),
.Y(n_106)
);


endmodule