module fake_jpeg_23494_n_230 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_230);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_19),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_33),
.Y(n_41)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_36),
.B1(n_20),
.B2(n_25),
.Y(n_46)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_20),
.B1(n_16),
.B2(n_18),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_40),
.A2(n_43),
.B1(n_36),
.B2(n_29),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_27),
.A2(n_20),
.B1(n_25),
.B2(n_16),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_50),
.Y(n_66)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_26),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_53),
.Y(n_74)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_54),
.B(n_56),
.Y(n_81)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_63),
.Y(n_71)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_64),
.B1(n_45),
.B2(n_32),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_62),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_25),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

FAx1_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_51),
.CI(n_25),
.CON(n_65),
.SN(n_65)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_65),
.B(n_35),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_43),
.B1(n_32),
.B2(n_29),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_29),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_25),
.B(n_16),
.C(n_46),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_72),
.A2(n_79),
.B1(n_52),
.B2(n_60),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_50),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_78),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_80),
.B1(n_53),
.B2(n_36),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_50),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_36),
.B1(n_45),
.B2(n_35),
.Y(n_80)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_87),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_48),
.C(n_38),
.Y(n_109)
);

BUFx8_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_90),
.Y(n_91)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_65),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_0),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_56),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_54),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_67),
.B1(n_36),
.B2(n_65),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_102),
.B1(n_35),
.B2(n_55),
.Y(n_123)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_58),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_101),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_67),
.B1(n_60),
.B2(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_110),
.B(n_69),
.Y(n_125)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_77),
.Y(n_117)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_28),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_107),
.A2(n_86),
.B1(n_72),
.B2(n_71),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_121),
.B1(n_124),
.B2(n_125),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_81),
.C(n_87),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_115),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_87),
.C(n_33),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_122),
.B(n_17),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_72),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_120),
.B(n_126),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_105),
.A2(n_93),
.B1(n_96),
.B2(n_94),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_72),
.B(n_26),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_127),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_98),
.A2(n_44),
.B1(n_64),
.B2(n_83),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_103),
.A2(n_44),
.B1(n_17),
.B2(n_24),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_130),
.A2(n_17),
.B1(n_22),
.B2(n_24),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_132),
.A2(n_144),
.B1(n_15),
.B2(n_22),
.Y(n_160)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_116),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_134),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_102),
.B(n_92),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_138),
.B(n_140),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_121),
.Y(n_136)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_100),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_91),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_19),
.B1(n_21),
.B2(n_108),
.Y(n_158)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_92),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_91),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_150),
.B1(n_132),
.B2(n_135),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_104),
.B(n_101),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_146),
.A2(n_111),
.B1(n_114),
.B2(n_120),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_151),
.A2(n_161),
.B1(n_148),
.B2(n_147),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_127),
.C(n_126),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_154),
.C(n_164),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_99),
.C(n_33),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_108),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_162),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_142),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_159),
.B(n_160),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_69),
.B1(n_21),
.B2(n_23),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_141),
.B(n_28),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_28),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_28),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_37),
.C(n_61),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_168),
.B(n_151),
.Y(n_184)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_177),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_143),
.B1(n_148),
.B2(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_174),
.A2(n_180),
.B1(n_158),
.B2(n_161),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_133),
.B1(n_44),
.B2(n_37),
.Y(n_175)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_162),
.Y(n_186)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_61),
.C(n_31),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_179),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_31),
.C(n_30),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_15),
.B(n_27),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_173),
.A2(n_165),
.B(n_158),
.Y(n_185)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_186),
.B(n_192),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_191),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_164),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_155),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_178),
.C(n_171),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_196),
.C(n_197),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_172),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_172),
.C(n_176),
.Y(n_197)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_161),
.Y(n_207)
);

AOI21x1_ASAP7_75t_L g204 ( 
.A1(n_199),
.A2(n_193),
.B(n_183),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_207),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_201),
.A2(n_188),
.B(n_179),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_206),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_8),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_208),
.B(n_209),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_8),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_198),
.A2(n_8),
.B1(n_12),
.B2(n_4),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_211),
.A2(n_197),
.B1(n_196),
.B2(n_4),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_215),
.B(n_216),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_200),
.C(n_23),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_23),
.C(n_14),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_205),
.Y(n_220)
);

AOI31xp33_ASAP7_75t_L g219 ( 
.A1(n_213),
.A2(n_206),
.A3(n_216),
.B(n_214),
.Y(n_219)
);

OAI322xp33_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_218),
.A3(n_217),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_10),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_220),
.B(n_221),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_7),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_222),
.A2(n_10),
.B(n_11),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_6),
.C(n_7),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_0),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_226),
.C(n_223),
.Y(n_227)
);

AOI321xp33_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_1),
.C(n_0),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_11),
.B(n_12),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_0),
.C(n_1),
.Y(n_230)
);


endmodule