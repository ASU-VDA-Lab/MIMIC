module fake_jpeg_14322_n_510 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_510);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_510;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_15),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_57),
.B(n_83),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_59),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_6),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_62),
.B(n_64),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_21),
.B(n_6),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_65),
.Y(n_152)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

INVx5_ASAP7_75t_SL g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g137 ( 
.A(n_73),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_21),
.B(n_6),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_74),
.B(n_92),
.Y(n_147)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_76),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_82),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_20),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

BUFx4f_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx5_ASAP7_75t_SL g125 ( 
.A(n_88),
.Y(n_125)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_25),
.B(n_6),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_25),
.B(n_5),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_41),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_46),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g156 ( 
.A(n_98),
.B(n_99),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_56),
.B(n_29),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_103),
.B(n_104),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_29),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_54),
.A2(n_45),
.B1(n_46),
.B2(n_33),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_114),
.A2(n_148),
.B1(n_46),
.B2(n_42),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_63),
.A2(n_16),
.B1(n_45),
.B2(n_50),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_117),
.A2(n_28),
.B(n_32),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_58),
.A2(n_36),
.B1(n_45),
.B2(n_18),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_119),
.A2(n_36),
.B1(n_107),
.B2(n_27),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_73),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_126),
.B(n_140),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_65),
.B(n_35),
.C(n_40),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_41),
.C(n_47),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_100),
.C(n_127),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_66),
.A2(n_93),
.B1(n_97),
.B2(n_96),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_146),
.B1(n_85),
.B2(n_78),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_139),
.B(n_145),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_67),
.B(n_38),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_69),
.B(n_38),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_60),
.A2(n_45),
.B1(n_33),
.B2(n_24),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_77),
.A2(n_46),
.B1(n_33),
.B2(n_37),
.Y(n_148)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_158),
.A2(n_197),
.B1(n_200),
.B2(n_43),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_160),
.A2(n_153),
.B1(n_138),
.B2(n_115),
.Y(n_242)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_125),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_167),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_148),
.A2(n_80),
.B1(n_91),
.B2(n_95),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_163),
.A2(n_176),
.B1(n_179),
.B2(n_88),
.Y(n_236)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_118),
.Y(n_166)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_170),
.B(n_172),
.Y(n_233)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_173),
.Y(n_243)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_112),
.Y(n_174)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_114),
.A2(n_75),
.B1(n_70),
.B2(n_42),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_103),
.A2(n_42),
.B1(n_37),
.B2(n_88),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_180),
.A2(n_190),
.B1(n_199),
.B2(n_142),
.Y(n_241)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_101),
.Y(n_181)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

BUFx4f_ASAP7_75t_SL g219 ( 
.A(n_184),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_146),
.A2(n_37),
.B1(n_42),
.B2(n_81),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_185),
.A2(n_153),
.B1(n_116),
.B2(n_142),
.Y(n_238)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_123),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_188),
.Y(n_214)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_104),
.A2(n_40),
.B(n_35),
.C(n_49),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_26),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_101),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_191),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_131),
.B(n_26),
.C(n_49),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_192),
.B(n_141),
.C(n_86),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_147),
.A2(n_18),
.B1(n_99),
.B2(n_98),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_141),
.Y(n_234)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_143),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_196),
.Y(n_235)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_111),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_115),
.A2(n_47),
.B1(n_28),
.B2(n_32),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_L g200 ( 
.A1(n_119),
.A2(n_37),
.B1(n_18),
.B2(n_43),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_130),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_201),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_151),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_202),
.B(n_203),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_137),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_205),
.Y(n_230)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_113),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_198),
.B(n_156),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_193),
.C(n_179),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_213),
.B(n_175),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_34),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_215),
.B(n_225),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_220),
.A2(n_160),
.B1(n_163),
.B2(n_176),
.Y(n_249)
);

AO22x1_ASAP7_75t_L g221 ( 
.A1(n_170),
.A2(n_155),
.B1(n_124),
.B2(n_106),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_221),
.B(n_247),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_34),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_192),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_159),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_108),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_242),
.B1(n_158),
.B2(n_185),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_172),
.B(n_151),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_184),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_138),
.B1(n_173),
.B2(n_190),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_249),
.A2(n_260),
.B1(n_263),
.B2(n_266),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_200),
.B(n_165),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_235),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_251),
.B(n_255),
.Y(n_313)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_252),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_253),
.A2(n_258),
.B1(n_262),
.B2(n_264),
.Y(n_287)
);

XNOR2x1_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_269),
.Y(n_293)
);

BUFx24_ASAP7_75t_SL g255 ( 
.A(n_208),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_256),
.B(n_230),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_257),
.B(n_265),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_236),
.A2(n_102),
.B1(n_133),
.B2(n_205),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_261),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_237),
.A2(n_102),
.B1(n_133),
.B2(n_113),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_238),
.A2(n_202),
.B1(n_199),
.B2(n_164),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_213),
.A2(n_144),
.B1(n_124),
.B2(n_106),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_215),
.B(n_206),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_233),
.A2(n_144),
.B1(n_201),
.B2(n_181),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_225),
.B(n_184),
.Y(n_267)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_267),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_217),
.B(n_182),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_270),
.B(n_279),
.Y(n_306)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_209),
.Y(n_271)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_271),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_108),
.B1(n_105),
.B2(n_191),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_227),
.B1(n_246),
.B2(n_244),
.Y(n_290)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_212),
.Y(n_273)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_233),
.B(n_178),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_277),
.Y(n_291)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_281),
.C(n_285),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g276 ( 
.A(n_219),
.Y(n_276)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_233),
.B(n_177),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_207),
.Y(n_278)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_207),
.B(n_226),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_210),
.B(n_166),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_282),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_239),
.B(n_157),
.C(n_105),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_214),
.B(n_5),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_232),
.B(n_0),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_283),
.B(n_0),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_221),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_284),
.Y(n_317)
);

FAx1_ASAP7_75t_SL g285 ( 
.A(n_221),
.B(n_15),
.CI(n_5),
.CON(n_285),
.SN(n_285)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_284),
.A2(n_227),
.B1(n_245),
.B2(n_232),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_288),
.A2(n_250),
.B(n_274),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_290),
.A2(n_260),
.B1(n_263),
.B2(n_259),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_253),
.A2(n_258),
.B1(n_254),
.B2(n_262),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_294),
.A2(n_296),
.B1(n_222),
.B2(n_211),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_254),
.A2(n_240),
.B1(n_229),
.B2(n_239),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_297),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_270),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_305),
.Y(n_325)
);

OA22x2_ASAP7_75t_L g299 ( 
.A1(n_249),
.A2(n_240),
.B1(n_228),
.B2(n_223),
.Y(n_299)
);

OA22x2_ASAP7_75t_L g328 ( 
.A1(n_299),
.A2(n_321),
.B1(n_290),
.B2(n_287),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_300),
.B(n_279),
.Y(n_333)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_261),
.Y(n_301)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_301),
.Y(n_346)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_271),
.Y(n_304)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_304),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_283),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_280),
.B(n_219),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_307),
.B(n_318),
.Y(n_327)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_273),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_311),
.Y(n_331)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_252),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_321),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_248),
.A2(n_243),
.B1(n_216),
.B2(n_228),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_316),
.A2(n_260),
.B1(n_223),
.B2(n_218),
.Y(n_348)
);

XNOR2x1_ASAP7_75t_SL g318 ( 
.A(n_269),
.B(n_219),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_265),
.Y(n_326)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_248),
.C(n_277),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_322),
.B(n_324),
.C(n_332),
.Y(n_361)
);

INVxp33_ASAP7_75t_L g375 ( 
.A(n_323),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_275),
.C(n_256),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_330),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_328),
.B(n_339),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_329),
.A2(n_352),
.B1(n_319),
.B2(n_310),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_292),
.A2(n_275),
.B(n_257),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_272),
.C(n_281),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_347),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_300),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_336),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_268),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_300),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_337),
.B(n_338),
.Y(n_381)
);

NAND3xp33_ASAP7_75t_L g338 ( 
.A(n_309),
.B(n_267),
.C(n_268),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_291),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_317),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_340),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_303),
.B(n_282),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_341),
.B(n_343),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_285),
.Y(n_342)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_342),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_292),
.A2(n_317),
.B(n_288),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_291),
.B(n_281),
.C(n_251),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_344),
.B(n_355),
.C(n_332),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_318),
.A2(n_285),
.B(n_264),
.Y(n_347)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_348),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_313),
.B(n_285),
.Y(n_349)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_349),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_306),
.B(n_216),
.Y(n_350)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_350),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_289),
.A2(n_244),
.B1(n_222),
.B2(n_218),
.Y(n_351)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_351),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_306),
.B(n_276),
.Y(n_353)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_353),
.Y(n_384)
);

NAND2x1_ASAP7_75t_L g355 ( 
.A(n_299),
.B(n_276),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_324),
.B(n_302),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_358),
.B(n_364),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_359),
.A2(n_348),
.B1(n_328),
.B2(n_334),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_352),
.A2(n_294),
.B1(n_302),
.B2(n_287),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_362),
.A2(n_365),
.B1(n_377),
.B2(n_328),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_286),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_339),
.A2(n_329),
.B1(n_347),
.B2(n_337),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_367),
.B(n_336),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_344),
.B(n_296),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_369),
.B(n_370),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_286),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_327),
.B(n_308),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_371),
.B(n_379),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_325),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_374),
.B(n_378),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_342),
.A2(n_299),
.B1(n_304),
.B2(n_295),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_325),
.B(n_301),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_297),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_327),
.B(n_295),
.C(n_312),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_382),
.B(n_385),
.C(n_330),
.Y(n_388)
);

XNOR2x1_ASAP7_75t_SL g383 ( 
.A(n_335),
.B(n_299),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_383),
.B(n_355),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_353),
.B(n_311),
.C(n_315),
.Y(n_385)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_323),
.B(n_289),
.C(n_314),
.Y(n_387)
);

MAJx2_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_343),
.C(n_326),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_393),
.C(n_401),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_356),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_389),
.B(n_390),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_381),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_386),
.B(n_345),
.Y(n_391)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_391),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_360),
.A2(n_340),
.B1(n_328),
.B2(n_333),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_392),
.A2(n_395),
.B1(n_396),
.B2(n_413),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_375),
.A2(n_355),
.B(n_345),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_394),
.B(n_399),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_372),
.A2(n_363),
.B1(n_375),
.B2(n_368),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_372),
.A2(n_384),
.B1(n_369),
.B2(n_376),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_365),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_357),
.Y(n_400)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_400),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_361),
.B(n_367),
.C(n_364),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_402),
.B(n_410),
.C(n_414),
.Y(n_423)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_377),
.Y(n_404)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_404),
.Y(n_419)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_385),
.Y(n_405)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_405),
.Y(n_425)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_383),
.Y(n_406)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_406),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_408),
.A2(n_409),
.B1(n_411),
.B2(n_415),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_361),
.B(n_328),
.C(n_331),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_362),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_412),
.B(n_211),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_366),
.A2(n_354),
.B1(n_334),
.B2(n_346),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_382),
.B(n_331),
.C(n_346),
.Y(n_414)
);

INVx5_ASAP7_75t_L g415 ( 
.A(n_359),
.Y(n_415)
);

AO22x1_ASAP7_75t_L g424 ( 
.A1(n_404),
.A2(n_387),
.B1(n_380),
.B2(n_373),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_424),
.A2(n_8),
.B(n_12),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_401),
.B(n_358),
.C(n_379),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_428),
.C(n_429),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_402),
.B(n_370),
.C(n_371),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_388),
.B(n_414),
.C(n_398),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_398),
.B(n_354),
.C(n_349),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_430),
.B(n_432),
.C(n_437),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_391),
.B(n_341),
.Y(n_431)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_431),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_314),
.C(n_338),
.Y(n_432)
);

AND3x1_ASAP7_75t_L g434 ( 
.A(n_412),
.B(n_224),
.C(n_243),
.Y(n_434)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_434),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_407),
.B(n_224),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_435),
.B(n_436),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_397),
.B(n_0),
.C(n_1),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_422),
.A2(n_409),
.B1(n_415),
.B2(n_403),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_440),
.A2(n_433),
.B1(n_419),
.B2(n_432),
.Y(n_457)
);

FAx1_ASAP7_75t_L g441 ( 
.A(n_424),
.B(n_394),
.CI(n_393),
.CON(n_441),
.SN(n_441)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_441),
.B(n_447),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_421),
.B(n_396),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_442),
.B(n_452),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_426),
.A2(n_392),
.B1(n_395),
.B2(n_413),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_443),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_420),
.A2(n_397),
.B1(n_407),
.B2(n_9),
.Y(n_446)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_446),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_15),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_423),
.B(n_15),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_448),
.B(n_453),
.Y(n_456)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_431),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_454),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_418),
.B(n_14),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_451),
.B(n_455),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_425),
.B(n_14),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_423),
.B(n_14),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_429),
.B(n_0),
.C(n_1),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_457),
.A2(n_444),
.B1(n_446),
.B2(n_441),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_450),
.A2(n_417),
.B(n_427),
.Y(n_459)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_459),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_439),
.B(n_417),
.C(n_428),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_461),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_439),
.B(n_450),
.C(n_440),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_435),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_8),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_445),
.B(n_430),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_468),
.B(n_12),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_438),
.B(n_453),
.C(n_448),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_470),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_437),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_444),
.A2(n_434),
.B(n_436),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_471),
.A2(n_12),
.B(n_2),
.Y(n_482)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_472),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_461),
.B(n_451),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_473),
.B(n_465),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_447),
.Y(n_474)
);

OAI21x1_ASAP7_75t_SL g490 ( 
.A1(n_474),
.A2(n_483),
.B(n_464),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_463),
.A2(n_441),
.B1(n_455),
.B2(n_438),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_476),
.B(n_480),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_478),
.B(n_482),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_458),
.B(n_8),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_479),
.B(n_466),
.Y(n_486)
);

INVx3_ASAP7_75t_SL g481 ( 
.A(n_467),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_485),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_457),
.B(n_12),
.Y(n_483)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_464),
.Y(n_485)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_486),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_477),
.A2(n_460),
.B(n_463),
.Y(n_489)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_489),
.Y(n_500)
);

AO21x1_ASAP7_75t_L g496 ( 
.A1(n_490),
.A2(n_494),
.B(n_484),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_491),
.B(n_495),
.C(n_478),
.Y(n_498)
);

A2O1A1Ixp33_ASAP7_75t_SL g494 ( 
.A1(n_472),
.A2(n_471),
.B(n_469),
.C(n_456),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_456),
.Y(n_495)
);

AO21x1_ASAP7_75t_L g503 ( 
.A1(n_496),
.A2(n_497),
.B(n_488),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_493),
.Y(n_497)
);

INVxp33_ASAP7_75t_L g502 ( 
.A(n_498),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_493),
.A2(n_481),
.B1(n_474),
.B2(n_483),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_501),
.A2(n_492),
.B(n_494),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_503),
.B(n_499),
.C(n_487),
.Y(n_506)
);

AOI21xp33_ASAP7_75t_L g505 ( 
.A1(n_504),
.A2(n_500),
.B(n_496),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_505),
.A2(n_506),
.B(n_502),
.Y(n_507)
);

AOI21x1_ASAP7_75t_L g508 ( 
.A1(n_507),
.A2(n_482),
.B(n_3),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_1),
.C(n_3),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_509),
.A2(n_3),
.B(n_4),
.Y(n_510)
);


endmodule