module fake_jpeg_12410_n_417 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_417);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_417;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_40),
.B(n_43),
.Y(n_92)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_28),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_45),
.B(n_49),
.Y(n_90)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_14),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_47),
.B(n_61),
.Y(n_109)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_50),
.B(n_57),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_63),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_13),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_21),
.B(n_13),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_28),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_73),
.Y(n_101)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_25),
.B(n_0),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_51),
.Y(n_98)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_75),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_38),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_71),
.A2(n_19),
.B1(n_27),
.B2(n_26),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_77),
.B(n_36),
.C(n_27),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_34),
.B1(n_33),
.B2(n_31),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_79),
.A2(n_81),
.B1(n_87),
.B2(n_94),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_19),
.B1(n_27),
.B2(n_26),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_38),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_86),
.B(n_51),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_34),
.B1(n_33),
.B2(n_31),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_26),
.B1(n_19),
.B2(n_18),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_44),
.B(n_39),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_46),
.B(n_67),
.C(n_69),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_94),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_45),
.B(n_21),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_111),
.B(n_115),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_49),
.A2(n_35),
.B(n_32),
.Y(n_114)
);

OR2x2_ASAP7_75t_SL g156 ( 
.A(n_114),
.B(n_48),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_35),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_65),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_117),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_20),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_118),
.A2(n_122),
.B(n_150),
.Y(n_181)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g170 ( 
.A(n_121),
.Y(n_170)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_149),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_32),
.B1(n_20),
.B2(n_64),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_123),
.A2(n_129),
.B1(n_150),
.B2(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

INVxp67_ASAP7_75t_SL g163 ( 
.A(n_126),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_84),
.A2(n_42),
.B1(n_60),
.B2(n_52),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_50),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_137),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_108),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_132),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_135),
.Y(n_192)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g172 ( 
.A(n_136),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_81),
.B(n_40),
.Y(n_137)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_93),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_141),
.Y(n_180)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_140),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_97),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_43),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_90),
.B(n_66),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_88),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_77),
.A2(n_41),
.B1(n_53),
.B2(n_58),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_106),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_155),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_57),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_156),
.B(n_46),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_100),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_104),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_179),
.C(n_189),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_137),
.A2(n_78),
.B1(n_82),
.B2(n_62),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_161),
.A2(n_173),
.B1(n_175),
.B2(n_190),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_171),
.A2(n_126),
.B(n_144),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_78),
.B1(n_62),
.B2(n_56),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_130),
.A2(n_72),
.B1(n_56),
.B2(n_88),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_51),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_117),
.B(n_91),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_181),
.A2(n_184),
.B(n_150),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_122),
.B(n_127),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_125),
.B(n_134),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_195),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_119),
.B(n_91),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_119),
.A2(n_107),
.B1(n_18),
.B2(n_36),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_124),
.B(n_107),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_118),
.B1(n_140),
.B2(n_143),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_198),
.Y(n_246)
);

AND2x2_ASAP7_75t_SL g241 ( 
.A(n_199),
.B(n_166),
.Y(n_241)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_135),
.C(n_150),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_201),
.B(n_197),
.C(n_199),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_181),
.A2(n_151),
.B1(n_128),
.B2(n_148),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_202),
.A2(n_203),
.B1(n_209),
.B2(n_210),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_160),
.A2(n_121),
.B1(n_112),
.B2(n_147),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_204),
.B(n_186),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_195),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_205),
.B(n_207),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_154),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_206),
.B(n_208),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_180),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_120),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_160),
.A2(n_36),
.B1(n_18),
.B2(n_99),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_189),
.A2(n_112),
.B1(n_106),
.B2(n_99),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_187),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_212),
.B(n_216),
.Y(n_262)
);

OAI21xp33_ASAP7_75t_L g237 ( 
.A1(n_213),
.A2(n_221),
.B(n_226),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_182),
.A2(n_113),
.B1(n_85),
.B2(n_152),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_214),
.A2(n_223),
.B1(n_204),
.B2(n_210),
.Y(n_250)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_187),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_191),
.B(n_85),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_222),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_113),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_219),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_171),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_220),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_168),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_168),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_165),
.A2(n_158),
.B1(n_176),
.B2(n_179),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_175),
.A2(n_138),
.B1(n_136),
.B2(n_70),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_224),
.A2(n_163),
.B1(n_170),
.B2(n_166),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_158),
.A2(n_167),
.B1(n_165),
.B2(n_192),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_225),
.A2(n_174),
.B(n_193),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_194),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_194),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g267 ( 
.A1(n_227),
.A2(n_164),
.B(n_2),
.Y(n_267)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_172),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_231),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_159),
.B(n_153),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_232),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_162),
.B(n_169),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_235),
.Y(n_244)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_169),
.Y(n_234)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_174),
.B(n_153),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_233),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_238),
.B(n_239),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_206),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_263),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_214),
.A2(n_170),
.B1(n_185),
.B2(n_164),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_242),
.A2(n_224),
.B(n_216),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_250),
.A2(n_201),
.B1(n_220),
.B2(n_222),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_228),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_252),
.A2(n_202),
.B1(n_212),
.B2(n_221),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_185),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_257),
.C(n_197),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_235),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_265),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_219),
.Y(n_264)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_226),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_227),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_266),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_267),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_217),
.Y(n_269)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_203),
.B(n_193),
.Y(n_270)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_271),
.B(n_274),
.C(n_280),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_225),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_275),
.A2(n_286),
.B1(n_293),
.B2(n_270),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_277),
.A2(n_242),
.B(n_249),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_278),
.A2(n_236),
.B1(n_256),
.B2(n_238),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_239),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_279),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_251),
.C(n_261),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_282),
.Y(n_302)
);

XOR2x2_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_228),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_240),
.B(n_208),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_285),
.C(n_290),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_240),
.B(n_205),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_246),
.A2(n_218),
.B1(n_207),
.B2(n_211),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_243),
.B(n_209),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_262),
.Y(n_291)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_246),
.A2(n_218),
.B1(n_200),
.B2(n_215),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_243),
.B(n_230),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_298),
.Y(n_312)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_262),
.Y(n_295)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_245),
.Y(n_296)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_296),
.Y(n_319)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_245),
.Y(n_297)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_297),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_241),
.B(n_234),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_247),
.Y(n_299)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_299),
.Y(n_326)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_247),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_266),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_237),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_303),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_304),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_306),
.B(n_318),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_278),
.A2(n_236),
.B1(n_265),
.B2(n_256),
.Y(n_307)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_307),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_SL g308 ( 
.A1(n_277),
.A2(n_241),
.B(n_252),
.C(n_263),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_308),
.A2(n_316),
.B1(n_321),
.B2(n_322),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_310),
.A2(n_317),
.B1(n_292),
.B2(n_290),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_271),
.B(n_241),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_315),
.B(n_229),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_286),
.A2(n_293),
.B1(n_282),
.B2(n_273),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_287),
.A2(n_253),
.B1(n_258),
.B2(n_244),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_272),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g320 ( 
.A(n_272),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_320),
.B(n_1),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_279),
.A2(n_298),
.B1(n_289),
.B2(n_284),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_283),
.A2(n_270),
.B1(n_253),
.B2(n_244),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_276),
.A2(n_260),
.B1(n_248),
.B2(n_255),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_324),
.A2(n_70),
.B1(n_2),
.B2(n_3),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_260),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_248),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_305),
.B(n_259),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_328),
.B(n_331),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_294),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_285),
.Y(n_332)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_332),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_315),
.B(n_274),
.C(n_280),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_339),
.C(n_344),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_334),
.A2(n_346),
.B1(n_318),
.B2(n_320),
.Y(n_349)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_335),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_302),
.B(n_281),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_347),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_313),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_337),
.B(n_340),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_255),
.C(n_268),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_324),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_268),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_342),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_343),
.B(n_348),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_311),
.B(n_70),
.C(n_2),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_345),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_302),
.B(n_1),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_312),
.B(n_2),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_349),
.A2(n_338),
.B1(n_308),
.B2(n_327),
.Y(n_368)
);

AOI221xp5_ASAP7_75t_L g351 ( 
.A1(n_330),
.A2(n_322),
.B1(n_316),
.B2(n_321),
.C(n_310),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_351),
.B(n_3),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_303),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_359),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_339),
.B(n_312),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_5),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_329),
.B(n_326),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_330),
.B(n_323),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_361),
.B(n_5),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_338),
.A2(n_308),
.B1(n_301),
.B2(n_319),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_362),
.A2(n_301),
.B1(n_308),
.B2(n_346),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_327),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_365),
.A2(n_348),
.B(n_4),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_356),
.B(n_343),
.C(n_333),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_366),
.B(n_367),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_356),
.B(n_336),
.C(n_341),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_368),
.A2(n_376),
.B1(n_363),
.B2(n_352),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_327),
.C(n_344),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_373),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_371),
.A2(n_375),
.B1(n_7),
.B2(n_8),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_347),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_372),
.B(n_379),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_360),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_378),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_349),
.A2(n_358),
.B1(n_354),
.B2(n_365),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_377),
.B(n_7),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_364),
.B(n_5),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_373),
.B(n_350),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_380),
.B(n_382),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_367),
.C(n_370),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_362),
.C(n_352),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_383),
.A2(n_386),
.B(n_8),
.Y(n_396)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_385),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_355),
.C(n_359),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_369),
.B(n_355),
.Y(n_388)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_388),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_389),
.B(n_391),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_387),
.A2(n_377),
.B(n_9),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_394),
.B(n_399),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_396),
.B(n_384),
.C(n_386),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_382),
.B(n_8),
.C(n_9),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_397),
.B(n_11),
.Y(n_407)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_390),
.Y(n_398)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_398),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_383),
.A2(n_8),
.B(n_9),
.Y(n_399)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_401),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_395),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_404),
.B(n_405),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_400),
.A2(n_384),
.B(n_381),
.Y(n_405)
);

O2A1O1Ixp33_ASAP7_75t_SL g406 ( 
.A1(n_392),
.A2(n_9),
.B(n_11),
.C(n_12),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_406),
.B(n_407),
.Y(n_410)
);

NOR3xp33_ASAP7_75t_SL g409 ( 
.A(n_402),
.B(n_399),
.C(n_397),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_409),
.B(n_403),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_408),
.A2(n_403),
.B1(n_393),
.B2(n_12),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_412),
.A2(n_413),
.B(n_410),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_414),
.A2(n_411),
.B1(n_412),
.B2(n_393),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_415),
.B(n_11),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_416),
.B(n_12),
.Y(n_417)
);


endmodule