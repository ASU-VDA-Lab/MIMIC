module fake_jpeg_12619_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_6),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_1),
.B(n_30),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_13),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_54),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_18),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_48),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

OR2x2_ASAP7_75t_SL g66 ( 
.A(n_44),
.B(n_1),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_46),
.Y(n_70)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_17),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_40),
.B1(n_43),
.B2(n_50),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_73),
.B(n_64),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_78),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_40),
.B1(n_51),
.B2(n_43),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_58),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_52),
.B1(n_42),
.B2(n_41),
.Y(n_80)
);

AO22x1_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_81),
.B1(n_63),
.B2(n_64),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_62),
.A2(n_43),
.B1(n_22),
.B2(n_39),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_82),
.B(n_87),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_102)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_21),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_24),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_2),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_93),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_94),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_3),
.Y(n_93)
);

OR2x2_ASAP7_75t_SL g95 ( 
.A(n_69),
.B(n_3),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_25),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_27),
.C(n_37),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_68),
.B1(n_5),
.B2(n_7),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_12),
.B1(n_16),
.B2(n_29),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_110),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_105),
.B1(n_94),
.B2(n_97),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_4),
.B1(n_8),
.B2(n_10),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_11),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_11),
.Y(n_118)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_118),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_95),
.B(n_32),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_117),
.A2(n_109),
.B(n_100),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_34),
.C(n_14),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_105),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_121),
.B1(n_99),
.B2(n_109),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_125),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_103),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_106),
.A3(n_117),
.B1(n_126),
.B2(n_124),
.C1(n_120),
.C2(n_122),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_129),
.B(n_115),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_119),
.C(n_114),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_131),
.A2(n_108),
.B1(n_104),
.B2(n_101),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_104),
.Y(n_133)
);


endmodule