module fake_jpeg_26210_n_159 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_15),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_13),
.B(n_32),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_8),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_72),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_0),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_75),
.Y(n_79)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_63),
.Y(n_78)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_82),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_53),
.B1(n_47),
.B2(n_68),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_58),
.B1(n_54),
.B2(n_64),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_76),
.A2(n_53),
.B1(n_47),
.B2(n_69),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_91),
.B1(n_49),
.B2(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_61),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_51),
.B(n_60),
.C(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_90),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_61),
.B1(n_64),
.B2(n_59),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_59),
.B1(n_52),
.B2(n_62),
.Y(n_103)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_72),
.B(n_67),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_72),
.A2(n_52),
.B1(n_62),
.B2(n_48),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_62),
.B1(n_49),
.B2(n_2),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_94),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_114)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_0),
.Y(n_113)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_98),
.Y(n_110)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_66),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_106),
.B1(n_79),
.B2(n_1),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_104),
.A2(n_105),
.B1(n_81),
.B2(n_49),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_SL g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_79),
.Y(n_108)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_102),
.B1(n_93),
.B2(n_104),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_20),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_114),
.A2(n_105),
.B1(n_5),
.B2(n_6),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_121),
.B1(n_125),
.B2(n_107),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_24),
.B(n_45),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_92),
.B(n_99),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_126),
.B1(n_113),
.B2(n_14),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_110),
.A2(n_11),
.B(n_12),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_11),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_133),
.B1(n_135),
.B2(n_139),
.Y(n_143)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_128),
.B(n_129),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_116),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_132),
.Y(n_145)
);

NAND2xp33_ASAP7_75t_SL g134 ( 
.A(n_124),
.B(n_107),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_136),
.Y(n_146)
);

OAI22x1_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_115),
.B1(n_116),
.B2(n_13),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_17),
.C(n_18),
.Y(n_136)
);

NOR2x1_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_19),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_129),
.Y(n_142)
);

BUFx12_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_142),
.C(n_147),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_146),
.B(n_138),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_146),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_150),
.A2(n_144),
.B(n_130),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_148),
.C(n_142),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_141),
.B(n_145),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_25),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_27),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_143),
.C(n_140),
.Y(n_157)
);

AOI31xp33_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_37),
.A3(n_40),
.B(n_41),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_42),
.Y(n_159)
);


endmodule