module fake_jpeg_12346_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_12),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_23),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_1),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_33),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_35),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_78),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_2),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_3),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_2),
.Y(n_78)
);

BUFx8_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_3),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_74),
.Y(n_86)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_50),
.B1(n_64),
.B2(n_58),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_64),
.B1(n_60),
.B2(n_56),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_89),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_80),
.A2(n_63),
.B1(n_70),
.B2(n_73),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_28),
.B1(n_47),
.B2(n_46),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_94),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_83),
.Y(n_89)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_62),
.C(n_65),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_51),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_78),
.Y(n_94)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_69),
.B1(n_55),
.B2(n_54),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_95),
.B(n_70),
.Y(n_104)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NAND3xp33_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_72),
.C(n_67),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_98),
.A2(n_106),
.B(n_100),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_111),
.Y(n_121)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

NOR2xp67_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_52),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_13),
.B1(n_15),
.B2(n_17),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_87),
.B(n_56),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_9),
.C(n_10),
.Y(n_126)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_60),
.A3(n_57),
.B1(n_6),
.B2(n_7),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_21),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_4),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_113),
.B(n_5),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_127),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_120),
.Y(n_145)
);

CKINVDCx12_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_119),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_104),
.A2(n_5),
.B(n_7),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_44),
.C(n_48),
.Y(n_143)
);

NOR2x1_ASAP7_75t_R g124 ( 
.A(n_106),
.B(n_8),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_124),
.B(n_118),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_126),
.A2(n_42),
.B(n_43),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_11),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_129),
.A2(n_19),
.B1(n_32),
.B2(n_34),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_110),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_36),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_114),
.B1(n_20),
.B2(n_31),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_135),
.B(n_136),
.Y(n_153)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_138),
.B(n_143),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_139),
.A2(n_125),
.B(n_131),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_38),
.C(n_40),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_141),
.C(n_144),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_144),
.C(n_140),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_146),
.C(n_134),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_116),
.B(n_118),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_148),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_158),
.A2(n_157),
.B(n_156),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_159),
.B(n_151),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_153),
.B(n_149),
.Y(n_163)
);

FAx1_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_145),
.CI(n_121),
.CON(n_164),
.SN(n_164)
);


endmodule