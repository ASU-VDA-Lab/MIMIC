module real_aes_2613_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_288;
wire n_147;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g245 ( .A(n_0), .B(n_160), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_1), .B(n_802), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_2), .B(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g151 ( .A(n_3), .Y(n_151) );
NAND2xp33_ASAP7_75t_SL g230 ( .A(n_4), .B(n_150), .Y(n_230) );
INVx1_ASAP7_75t_L g221 ( .A(n_5), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_6), .B(n_164), .Y(n_489) );
INVx1_ASAP7_75t_L g532 ( .A(n_7), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g802 ( .A(n_8), .Y(n_802) );
AND2x2_ASAP7_75t_L g138 ( .A(n_9), .B(n_139), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_10), .Y(n_546) );
INVx2_ASAP7_75t_L g140 ( .A(n_11), .Y(n_140) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_12), .Y(n_116) );
AND3x1_ASAP7_75t_L g799 ( .A(n_12), .B(n_35), .C(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g497 ( .A(n_13), .Y(n_497) );
AOI221x1_ASAP7_75t_L g224 ( .A1(n_14), .A2(n_153), .B1(n_225), .B2(n_227), .C(n_229), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_15), .B(n_144), .Y(n_211) );
INVx1_ASAP7_75t_L g120 ( .A(n_16), .Y(n_120) );
NOR2xp33_ASAP7_75t_SL g797 ( .A(n_16), .B(n_121), .Y(n_797) );
INVx1_ASAP7_75t_L g495 ( .A(n_17), .Y(n_495) );
INVx1_ASAP7_75t_SL g482 ( .A(n_18), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_19), .B(n_145), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_20), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_21), .A2(n_153), .B(n_158), .Y(n_152) );
AOI221xp5_ASAP7_75t_SL g235 ( .A1(n_22), .A2(n_40), .B1(n_144), .B2(n_153), .C(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_23), .B(n_160), .Y(n_159) );
AOI33xp33_ASAP7_75t_L g512 ( .A1(n_24), .A2(n_52), .A3(n_197), .B1(n_204), .B2(n_513), .B3(n_514), .Y(n_512) );
AOI22x1_ASAP7_75t_R g124 ( .A1(n_25), .A2(n_37), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_25), .Y(n_126) );
INVx1_ASAP7_75t_L g540 ( .A(n_26), .Y(n_540) );
OR2x2_ASAP7_75t_L g141 ( .A(n_27), .B(n_89), .Y(n_141) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_27), .A2(n_89), .B(n_140), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_28), .B(n_162), .Y(n_215) );
INVxp67_ASAP7_75t_L g223 ( .A(n_29), .Y(n_223) );
AND2x2_ASAP7_75t_L g184 ( .A(n_30), .B(n_174), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_31), .B(n_195), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_32), .A2(n_153), .B(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_33), .B(n_162), .Y(n_237) );
AND2x2_ASAP7_75t_L g150 ( .A(n_34), .B(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g154 ( .A(n_34), .B(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g203 ( .A(n_34), .Y(n_203) );
OR2x6_ASAP7_75t_L g118 ( .A(n_35), .B(n_119), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_36), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_37), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_38), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_39), .B(n_195), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_41), .A2(n_164), .B1(n_228), .B2(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_42), .B(n_464), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_43), .A2(n_81), .B1(n_153), .B2(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_44), .B(n_145), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_45), .B(n_160), .Y(n_182) );
XOR2xp5_ASAP7_75t_L g446 ( .A(n_46), .B(n_447), .Y(n_446) );
AOI22x1_ASAP7_75t_SL g784 ( .A1(n_46), .A2(n_67), .B1(n_785), .B2(n_786), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_46), .Y(n_785) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_47), .B(n_191), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_48), .B(n_145), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_49), .Y(n_459) );
AND2x2_ASAP7_75t_L g248 ( .A(n_50), .B(n_174), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_51), .B(n_174), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_53), .B(n_145), .Y(n_524) );
INVx1_ASAP7_75t_L g147 ( .A(n_54), .Y(n_147) );
INVx1_ASAP7_75t_L g157 ( .A(n_54), .Y(n_157) );
AND2x2_ASAP7_75t_L g525 ( .A(n_55), .B(n_174), .Y(n_525) );
AOI221xp5_ASAP7_75t_L g530 ( .A1(n_56), .A2(n_74), .B1(n_195), .B2(n_201), .C(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_57), .B(n_195), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_58), .B(n_144), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_59), .B(n_228), .Y(n_548) );
AOI21xp5_ASAP7_75t_SL g469 ( .A1(n_60), .A2(n_201), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g175 ( .A(n_61), .B(n_174), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_62), .B(n_162), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_63), .B(n_160), .Y(n_171) );
AND2x2_ASAP7_75t_SL g216 ( .A(n_64), .B(n_139), .Y(n_216) );
INVx1_ASAP7_75t_L g492 ( .A(n_65), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_66), .A2(n_153), .B(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_67), .Y(n_786) );
INVx1_ASAP7_75t_L g523 ( .A(n_68), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_69), .B(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_SL g206 ( .A(n_70), .B(n_191), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_71), .A2(n_201), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g149 ( .A(n_72), .Y(n_149) );
INVx1_ASAP7_75t_L g155 ( .A(n_72), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_73), .B(n_195), .Y(n_515) );
AND2x2_ASAP7_75t_L g484 ( .A(n_75), .B(n_227), .Y(n_484) );
INVx1_ASAP7_75t_L g493 ( .A(n_76), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_77), .A2(n_201), .B(n_481), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_78), .A2(n_190), .B(n_201), .C(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_79), .B(n_144), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_80), .A2(n_84), .B1(n_144), .B2(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g121 ( .A(n_82), .Y(n_121) );
AND2x2_ASAP7_75t_SL g467 ( .A(n_83), .B(n_227), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_85), .A2(n_201), .B1(n_510), .B2(n_511), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_86), .B(n_160), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_87), .B(n_160), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_88), .A2(n_153), .B(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g471 ( .A(n_90), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_91), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_92), .B(n_162), .Y(n_170) );
AND2x2_ASAP7_75t_L g516 ( .A(n_93), .B(n_227), .Y(n_516) );
OAI22xp33_ASAP7_75t_SL g782 ( .A1(n_94), .A2(n_783), .B1(n_784), .B2(n_787), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_94), .Y(n_787) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_95), .A2(n_538), .B(n_539), .C(n_541), .Y(n_537) );
INVxp67_ASAP7_75t_L g226 ( .A(n_96), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_97), .B(n_144), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_98), .B(n_162), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_99), .A2(n_153), .B(n_213), .Y(n_212) );
BUFx2_ASAP7_75t_L g108 ( .A(n_100), .Y(n_108) );
BUFx2_ASAP7_75t_SL g778 ( .A(n_100), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_101), .B(n_145), .Y(n_472) );
AOI21xp33_ASAP7_75t_SL g102 ( .A1(n_103), .A2(n_792), .B(n_803), .Y(n_102) );
OA21x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_123), .B(n_776), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_105), .B(n_109), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_110), .A2(n_780), .B(n_789), .Y(n_779) );
NOR2xp33_ASAP7_75t_SL g110 ( .A(n_111), .B(n_122), .Y(n_110) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g791 ( .A(n_115), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
OR2x6_ASAP7_75t_SL g444 ( .A(n_116), .B(n_117), .Y(n_444) );
AND2x6_ASAP7_75t_SL g767 ( .A(n_116), .B(n_118), .Y(n_767) );
OR2x2_ASAP7_75t_L g775 ( .A(n_116), .B(n_118), .Y(n_775) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_127), .B(n_768), .Y(n_123) );
AOI21xp33_ASAP7_75t_L g768 ( .A1(n_124), .A2(n_769), .B(n_771), .Y(n_768) );
INVx1_ASAP7_75t_SL g127 ( .A(n_128), .Y(n_127) );
OAI22x1_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_442), .B1(n_445), .B2(n_766), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g770 ( .A(n_130), .Y(n_770) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_364), .Y(n_130) );
NOR3xp33_ASAP7_75t_SL g131 ( .A(n_132), .B(n_288), .C(n_338), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_268), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_207), .B(n_249), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_185), .Y(n_135) );
INVx1_ASAP7_75t_SL g374 ( .A(n_136), .Y(n_374) );
AOI32xp33_ASAP7_75t_L g405 ( .A1(n_136), .A2(n_387), .A3(n_406), .B1(n_407), .B2(n_408), .Y(n_405) );
AND2x2_ASAP7_75t_L g407 ( .A(n_136), .B(n_264), .Y(n_407) );
AND2x4_ASAP7_75t_SL g136 ( .A(n_137), .B(n_165), .Y(n_136) );
HB1xp67_ASAP7_75t_L g186 ( .A(n_137), .Y(n_186) );
INVx5_ASAP7_75t_L g267 ( .A(n_137), .Y(n_267) );
OR2x2_ASAP7_75t_L g274 ( .A(n_137), .B(n_266), .Y(n_274) );
INVx2_ASAP7_75t_L g279 ( .A(n_137), .Y(n_279) );
AND2x2_ASAP7_75t_L g291 ( .A(n_137), .B(n_166), .Y(n_291) );
AND2x2_ASAP7_75t_L g296 ( .A(n_137), .B(n_176), .Y(n_296) );
OR2x2_ASAP7_75t_L g303 ( .A(n_137), .B(n_188), .Y(n_303) );
AND2x4_ASAP7_75t_L g312 ( .A(n_137), .B(n_177), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_SL g354 ( .A1(n_137), .A2(n_270), .B(n_305), .C(n_343), .Y(n_354) );
OR2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_142), .Y(n_137) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_139), .Y(n_174) );
AND2x2_ASAP7_75t_SL g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x4_ASAP7_75t_L g164 ( .A(n_140), .B(n_141), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_152), .B(n_164), .Y(n_142) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_150), .Y(n_144) );
INVx1_ASAP7_75t_L g231 ( .A(n_145), .Y(n_231) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
AND2x6_ASAP7_75t_L g160 ( .A(n_146), .B(n_155), .Y(n_160) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x4_ASAP7_75t_L g162 ( .A(n_148), .B(n_157), .Y(n_162) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx5_ASAP7_75t_L g163 ( .A(n_150), .Y(n_163) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_150), .Y(n_541) );
AND2x2_ASAP7_75t_L g156 ( .A(n_151), .B(n_157), .Y(n_156) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_151), .Y(n_198) );
AND2x6_ASAP7_75t_L g153 ( .A(n_154), .B(n_156), .Y(n_153) );
BUFx3_ASAP7_75t_L g199 ( .A(n_154), .Y(n_199) );
INVx2_ASAP7_75t_L g205 ( .A(n_155), .Y(n_205) );
AND2x4_ASAP7_75t_L g201 ( .A(n_156), .B(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g197 ( .A(n_157), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_161), .B(n_163), .Y(n_158) );
INVxp67_ASAP7_75t_L g496 ( .A(n_160), .Y(n_496) );
INVxp67_ASAP7_75t_L g498 ( .A(n_162), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_163), .A2(n_170), .B(n_171), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_163), .A2(n_181), .B(n_182), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_163), .A2(n_214), .B(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_163), .A2(n_237), .B(n_238), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_163), .A2(n_245), .B(n_246), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_163), .A2(n_462), .B(n_463), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_163), .A2(n_465), .B(n_471), .C(n_472), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_SL g481 ( .A1(n_163), .A2(n_465), .B(n_482), .C(n_483), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_163), .B(n_164), .Y(n_499) );
INVx1_ASAP7_75t_L g510 ( .A(n_163), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_163), .A2(n_465), .B(n_523), .C(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_SL g531 ( .A1(n_163), .A2(n_465), .B(n_532), .C(n_533), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_164), .B(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_164), .B(n_223), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_164), .B(n_226), .Y(n_225) );
NOR3xp33_ASAP7_75t_L g229 ( .A(n_164), .B(n_230), .C(n_231), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_164), .A2(n_469), .B(n_473), .Y(n_468) );
INVx3_ASAP7_75t_SL g304 ( .A(n_165), .Y(n_304) );
AND2x2_ASAP7_75t_L g350 ( .A(n_165), .B(n_267), .Y(n_350) );
AND2x4_ASAP7_75t_L g165 ( .A(n_166), .B(n_176), .Y(n_165) );
AND2x2_ASAP7_75t_L g187 ( .A(n_166), .B(n_188), .Y(n_187) );
OR2x2_ASAP7_75t_L g281 ( .A(n_166), .B(n_177), .Y(n_281) );
AND2x2_ASAP7_75t_L g285 ( .A(n_166), .B(n_264), .Y(n_285) );
INVx1_ASAP7_75t_L g311 ( .A(n_166), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_166), .B(n_177), .Y(n_333) );
INVx2_ASAP7_75t_L g337 ( .A(n_166), .Y(n_337) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_166), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_166), .B(n_267), .Y(n_414) );
AO21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_173), .B(n_175), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_172), .Y(n_167) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_173), .A2(n_178), .B(n_184), .Y(n_177) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_173), .A2(n_178), .B(n_184), .Y(n_266) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_173), .A2(n_478), .B(n_484), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_174), .Y(n_173) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_174), .A2(n_235), .B(n_239), .Y(n_234) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g348 ( .A(n_177), .B(n_188), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_183), .Y(n_178) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
INVx1_ASAP7_75t_L g358 ( .A(n_186), .Y(n_358) );
NAND2xp33_ASAP7_75t_SL g383 ( .A(n_186), .B(n_275), .Y(n_383) );
AND2x2_ASAP7_75t_L g425 ( .A(n_187), .B(n_267), .Y(n_425) );
AND2x2_ASAP7_75t_L g336 ( .A(n_188), .B(n_337), .Y(n_336) );
BUFx2_ASAP7_75t_L g399 ( .A(n_188), .Y(n_399) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_189), .Y(n_264) );
AOI21x1_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_193), .B(n_206), .Y(n_189) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_190), .A2(n_508), .B(n_516), .Y(n_507) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_190), .A2(n_508), .B(n_516), .Y(n_556) );
INVx2_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_191), .A2(n_211), .B(n_212), .Y(n_210) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_191), .A2(n_530), .B(n_534), .Y(n_529) );
BUFx4f_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx3_ASAP7_75t_L g228 ( .A(n_192), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_200), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_195), .A2(n_201), .B1(n_220), .B2(n_222), .Y(n_219) );
INVx1_ASAP7_75t_L g549 ( .A(n_195), .Y(n_549) );
AND2x4_ASAP7_75t_L g195 ( .A(n_196), .B(n_199), .Y(n_195) );
INVx1_ASAP7_75t_L g457 ( .A(n_196), .Y(n_457) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
OR2x6_ASAP7_75t_L g465 ( .A(n_197), .B(n_205), .Y(n_465) );
INVxp33_ASAP7_75t_L g513 ( .A(n_197), .Y(n_513) );
INVx1_ASAP7_75t_L g458 ( .A(n_199), .Y(n_458) );
INVxp67_ASAP7_75t_L g547 ( .A(n_201), .Y(n_547) );
NOR2x1p5_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
INVx1_ASAP7_75t_L g514 ( .A(n_204), .Y(n_514) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_207), .A2(n_290), .B1(n_392), .B2(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_232), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_208), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_208), .B(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_217), .Y(n_208) );
INVx2_ASAP7_75t_L g255 ( .A(n_209), .Y(n_255) );
OR2x2_ASAP7_75t_L g259 ( .A(n_209), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_209), .B(n_272), .Y(n_277) );
AND2x4_ASAP7_75t_SL g287 ( .A(n_209), .B(n_218), .Y(n_287) );
OR2x2_ASAP7_75t_L g294 ( .A(n_209), .B(n_234), .Y(n_294) );
OR2x2_ASAP7_75t_L g306 ( .A(n_209), .B(n_218), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_209), .B(n_234), .Y(n_320) );
INVx1_ASAP7_75t_L g325 ( .A(n_209), .Y(n_325) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_209), .Y(n_343) );
AND2x2_ASAP7_75t_L g406 ( .A(n_209), .B(n_326), .Y(n_406) );
INVx2_ASAP7_75t_L g410 ( .A(n_209), .Y(n_410) );
OR2x2_ASAP7_75t_L g417 ( .A(n_209), .B(n_307), .Y(n_417) );
OR2x2_ASAP7_75t_L g439 ( .A(n_209), .B(n_440), .Y(n_439) );
OR2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_216), .Y(n_209) );
AND2x2_ASAP7_75t_L g256 ( .A(n_217), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_217), .B(n_240), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_217), .B(n_316), .Y(n_378) );
INVx3_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g275 ( .A(n_218), .Y(n_275) );
AND2x4_ASAP7_75t_L g326 ( .A(n_218), .B(n_327), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_218), .B(n_271), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_218), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_218), .B(n_260), .Y(n_419) );
AND2x4_ASAP7_75t_L g218 ( .A(n_219), .B(n_224), .Y(n_218) );
INVx3_ASAP7_75t_L g518 ( .A(n_227), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_227), .A2(n_518), .B1(n_537), .B2(n_542), .Y(n_536) );
INVx4_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AOI21x1_ASAP7_75t_L g241 ( .A1(n_228), .A2(n_242), .B(n_248), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_228), .B(n_545), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_231), .A2(n_465), .B1(n_492), .B2(n_493), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_231), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g286 ( .A(n_232), .B(n_287), .Y(n_286) );
AO221x1_ASAP7_75t_L g360 ( .A1(n_232), .A2(n_275), .B1(n_306), .B2(n_361), .C(n_362), .Y(n_360) );
OAI322xp33_ASAP7_75t_L g412 ( .A1(n_232), .A2(n_332), .A3(n_413), .B1(n_415), .B2(n_416), .C1(n_417), .C2(n_418), .Y(n_412) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_240), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
BUFx3_ASAP7_75t_L g254 ( .A(n_234), .Y(n_254) );
INVx2_ASAP7_75t_L g260 ( .A(n_234), .Y(n_260) );
AND2x2_ASAP7_75t_L g272 ( .A(n_234), .B(n_240), .Y(n_272) );
INVx1_ASAP7_75t_L g317 ( .A(n_234), .Y(n_317) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_234), .Y(n_373) );
INVx1_ASAP7_75t_L g257 ( .A(n_240), .Y(n_257) );
OR2x2_ASAP7_75t_L g307 ( .A(n_240), .B(n_260), .Y(n_307) );
INVx2_ASAP7_75t_L g327 ( .A(n_240), .Y(n_327) );
INVx1_ASAP7_75t_L g380 ( .A(n_240), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_240), .B(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_247), .Y(n_242) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OAI21xp33_ASAP7_75t_SL g250 ( .A1(n_251), .A2(n_258), .B(n_261), .Y(n_250) );
AOI221xp5_ASAP7_75t_L g289 ( .A1(n_251), .A2(n_290), .B1(n_292), .B2(n_296), .C(n_297), .Y(n_289) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_256), .Y(n_252) );
NOR2x1p5_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g376 ( .A(n_255), .Y(n_376) );
INVx1_ASAP7_75t_SL g295 ( .A(n_256), .Y(n_295) );
OAI21xp5_ASAP7_75t_L g400 ( .A1(n_256), .A2(n_401), .B(n_403), .Y(n_400) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_257), .Y(n_300) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_260), .Y(n_363) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
OAI211xp5_ASAP7_75t_L g338 ( .A1(n_263), .A2(n_339), .B(n_344), .C(n_355), .Y(n_338) );
OR2x2_ASAP7_75t_L g428 ( .A(n_263), .B(n_333), .Y(n_428) );
AND2x2_ASAP7_75t_L g430 ( .A(n_263), .B(n_296), .Y(n_430) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g270 ( .A(n_264), .B(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g332 ( .A(n_264), .B(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g370 ( .A(n_264), .B(n_337), .Y(n_370) );
OA33x2_ASAP7_75t_L g377 ( .A1(n_264), .A2(n_294), .A3(n_378), .B1(n_379), .B2(n_381), .B3(n_383), .Y(n_377) );
OR2x2_ASAP7_75t_L g388 ( .A(n_264), .B(n_373), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_264), .B(n_312), .Y(n_402) );
AND2x4_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
AND2x2_ASAP7_75t_L g290 ( .A(n_266), .B(n_291), .Y(n_290) );
AOI22xp33_ASAP7_75t_SL g339 ( .A1(n_266), .A2(n_296), .B1(n_340), .B2(n_341), .Y(n_339) );
NAND3xp33_ASAP7_75t_L g379 ( .A(n_267), .B(n_347), .C(n_380), .Y(n_379) );
AOI322xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_273), .A3(n_275), .B1(n_276), .B2(n_278), .C1(n_282), .C2(n_286), .Y(n_268) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g375 ( .A(n_271), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g330 ( .A1(n_272), .A2(n_287), .B(n_331), .C(n_334), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_273), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
NAND4xp25_ASAP7_75t_SL g394 ( .A(n_274), .B(n_303), .C(n_395), .D(n_397), .Y(n_394) );
INVx1_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx2_ASAP7_75t_L g284 ( .A(n_279), .Y(n_284) );
OR2x2_ASAP7_75t_L g329 ( .A(n_279), .B(n_281), .Y(n_329) );
AND2x2_ASAP7_75t_L g398 ( .A(n_280), .B(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x2_ASAP7_75t_L g403 ( .A(n_284), .B(n_398), .Y(n_403) );
BUFx2_ASAP7_75t_L g396 ( .A(n_285), .Y(n_396) );
INVx1_ASAP7_75t_SL g426 ( .A(n_286), .Y(n_426) );
AND2x4_ASAP7_75t_L g362 ( .A(n_287), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g415 ( .A(n_287), .Y(n_415) );
NAND3xp33_ASAP7_75t_L g288 ( .A(n_289), .B(n_308), .C(n_330), .Y(n_288) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
INVx1_ASAP7_75t_SL g352 ( .A(n_294), .Y(n_352) );
OAI211xp5_ASAP7_75t_L g420 ( .A1(n_294), .A2(n_421), .B(n_422), .C(n_431), .Y(n_420) );
OR2x2_ASAP7_75t_L g342 ( .A(n_295), .B(n_343), .Y(n_342) );
OAI22xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_301), .B1(n_304), .B2(n_305), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_299), .B(n_382), .Y(n_381) );
INVxp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_302), .B(n_359), .Y(n_441) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g416 ( .A(n_303), .B(n_304), .Y(n_416) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g361 ( .A(n_307), .Y(n_361) );
AOI222xp33_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_313), .B1(n_318), .B2(n_322), .C1(n_323), .C2(n_328), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_311), .Y(n_322) );
AND2x2_ASAP7_75t_L g369 ( .A(n_312), .B(n_370), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_312), .A2(n_385), .B1(n_390), .B2(n_394), .Y(n_384) );
INVx2_ASAP7_75t_SL g437 ( .A(n_312), .Y(n_437) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVxp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g393 ( .A(n_317), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_317), .B(n_380), .Y(n_440) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g353 ( .A(n_321), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_323), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g391 ( .A(n_325), .Y(n_391) );
AND2x2_ASAP7_75t_SL g392 ( .A(n_326), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g434 ( .A(n_326), .B(n_363), .Y(n_434) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g359 ( .A(n_333), .Y(n_359) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g438 ( .A(n_336), .Y(n_438) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_337), .Y(n_382) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
O2A1O1Ixp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_349), .B(n_351), .C(n_354), .Y(n_344) );
AND2x2_ASAP7_75t_SL g345 ( .A(n_346), .B(n_348), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g389 ( .A(n_351), .Y(n_389) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_360), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_SL g357 ( .A(n_358), .B(n_359), .Y(n_357) );
NOR3xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_404), .C(n_420), .Y(n_364) );
NAND3xp33_ASAP7_75t_L g365 ( .A(n_366), .B(n_384), .C(n_400), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_371), .B1(n_374), .B2(n_375), .C(n_377), .Y(n_367) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_386), .B(n_389), .Y(n_385) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g413 ( .A(n_399), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g421 ( .A(n_403), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_411), .Y(n_404) );
INVx2_ASAP7_75t_L g427 ( .A(n_406), .Y(n_427) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g418 ( .A(n_409), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B1(n_427), .B2(n_428), .C(n_429), .Y(n_423) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_435), .B1(n_439), .B2(n_441), .Y(n_432) );
INVx1_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
CKINVDCx11_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_444), .A2(n_446), .B1(n_766), .B2(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AO22x1_ASAP7_75t_L g780 ( .A1(n_447), .A2(n_781), .B1(n_782), .B2(n_788), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_447), .Y(n_781) );
NAND4xp75_ASAP7_75t_L g447 ( .A(n_448), .B(n_617), .C(n_683), .D(n_746), .Y(n_447) );
NOR2x1_ASAP7_75t_L g448 ( .A(n_449), .B(n_580), .Y(n_448) );
OR3x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_550), .C(n_577), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_485), .B(n_505), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_474), .Y(n_452) );
AND2x2_ASAP7_75t_L g680 ( .A(n_453), .B(n_650), .Y(n_680) );
INVx1_ASAP7_75t_L g753 ( .A(n_453), .Y(n_753) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_466), .Y(n_453) );
INVx2_ASAP7_75t_L g504 ( .A(n_454), .Y(n_504) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_454), .Y(n_568) );
AND2x2_ASAP7_75t_L g572 ( .A(n_454), .B(n_488), .Y(n_572) );
AND2x4_ASAP7_75t_L g588 ( .A(n_454), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g592 ( .A(n_454), .Y(n_592) );
AND2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_460), .Y(n_454) );
NOR3xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .C(n_459), .Y(n_456) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVxp67_ASAP7_75t_L g538 ( .A(n_465), .Y(n_538) );
AND2x2_ASAP7_75t_L g486 ( .A(n_466), .B(n_487), .Y(n_486) );
INVx4_ASAP7_75t_L g569 ( .A(n_466), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_466), .B(n_559), .Y(n_573) );
INVx2_ASAP7_75t_L g587 ( .A(n_466), .Y(n_587) );
AND2x4_ASAP7_75t_L g591 ( .A(n_466), .B(n_592), .Y(n_591) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_466), .Y(n_626) );
OR2x2_ASAP7_75t_L g632 ( .A(n_466), .B(n_477), .Y(n_632) );
NOR2x1_ASAP7_75t_SL g661 ( .A(n_466), .B(n_488), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g763 ( .A(n_466), .B(n_735), .Y(n_763) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
AND2x2_ASAP7_75t_L g660 ( .A(n_474), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2x1_ASAP7_75t_L g694 ( .A(n_475), .B(n_487), .Y(n_694) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g501 ( .A(n_477), .Y(n_501) );
INVx2_ASAP7_75t_L g560 ( .A(n_477), .Y(n_560) );
AND2x2_ASAP7_75t_L g583 ( .A(n_477), .B(n_488), .Y(n_583) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_477), .Y(n_610) );
INVx1_ASAP7_75t_L g651 ( .A(n_477), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_500), .Y(n_485) );
AND2x2_ASAP7_75t_L g663 ( .A(n_486), .B(n_558), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_487), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g730 ( .A(n_487), .Y(n_730) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g589 ( .A(n_488), .Y(n_589) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_494), .B(n_499), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B1(n_497), .B2(n_498), .Y(n_494) );
OAI211xp5_ASAP7_75t_SL g666 ( .A1(n_500), .A2(n_667), .B(n_671), .C(n_677), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_501), .B(n_502), .Y(n_500) );
AND2x2_ASAP7_75t_SL g582 ( .A(n_502), .B(n_583), .Y(n_582) );
INVx2_ASAP7_75t_SL g713 ( .A(n_502), .Y(n_713) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g635 ( .A(n_504), .B(n_589), .Y(n_635) );
OR2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_526), .Y(n_505) );
AOI32xp33_ASAP7_75t_L g671 ( .A1(n_506), .A2(n_655), .A3(n_672), .B1(n_673), .B2(n_675), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_517), .Y(n_506) );
INVx2_ASAP7_75t_L g597 ( .A(n_507), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_507), .B(n_529), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_509), .B(n_515), .Y(n_508) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx3_ASAP7_75t_L g609 ( .A(n_517), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_517), .B(n_535), .Y(n_640) );
AND2x2_ASAP7_75t_L g645 ( .A(n_517), .B(n_646), .Y(n_645) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_517), .Y(n_727) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_525), .Y(n_517) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_518), .A2(n_519), .B(n_525), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
OR2x2_ASAP7_75t_L g628 ( .A(n_526), .B(n_629), .Y(n_628) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g579 ( .A(n_527), .B(n_553), .Y(n_579) );
AND2x2_ASAP7_75t_L g728 ( .A(n_527), .B(n_726), .Y(n_728) );
AND2x4_ASAP7_75t_L g527 ( .A(n_528), .B(n_535), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g565 ( .A(n_529), .Y(n_565) );
AND2x4_ASAP7_75t_L g604 ( .A(n_529), .B(n_605), .Y(n_604) );
INVxp67_ASAP7_75t_L g638 ( .A(n_529), .Y(n_638) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_529), .Y(n_646) );
AND2x2_ASAP7_75t_L g655 ( .A(n_529), .B(n_535), .Y(n_655) );
INVx1_ASAP7_75t_L g739 ( .A(n_529), .Y(n_739) );
INVx2_ASAP7_75t_L g576 ( .A(n_535), .Y(n_576) );
INVx1_ASAP7_75t_L g603 ( .A(n_535), .Y(n_603) );
INVx1_ASAP7_75t_L g670 ( .A(n_535), .Y(n_670) );
OR2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_543), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_547), .B1(n_548), .B2(n_549), .Y(n_543) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OAI32xp33_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_561), .A3(n_566), .B1(n_570), .B2(n_574), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_552), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_557), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_553), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g654 ( .A(n_553), .B(n_655), .Y(n_654) );
INVxp67_ASAP7_75t_L g679 ( .A(n_553), .Y(n_679) );
AND2x2_ASAP7_75t_L g760 ( .A(n_553), .B(n_602), .Y(n_760) );
AND2x4_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g575 ( .A(n_555), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g674 ( .A(n_555), .B(n_597), .Y(n_674) );
NOR2xp67_ASAP7_75t_L g696 ( .A(n_555), .B(n_576), .Y(n_696) );
NOR2x1_ASAP7_75t_L g738 ( .A(n_555), .B(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g605 ( .A(n_556), .Y(n_605) );
INVx1_ASAP7_75t_L g629 ( .A(n_556), .Y(n_629) );
AND2x2_ASAP7_75t_L g644 ( .A(n_556), .B(n_576), .Y(n_644) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g672 ( .A(n_558), .B(n_661), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_558), .B(n_591), .Y(n_742) );
INVx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_559), .Y(n_711) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_560), .Y(n_693) );
INVxp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g594 ( .A(n_563), .B(n_595), .Y(n_594) );
NOR2xp67_ASAP7_75t_L g678 ( .A(n_563), .B(n_679), .Y(n_678) );
NOR2xp67_ASAP7_75t_SL g765 ( .A(n_563), .B(n_703), .Y(n_765) );
INVx3_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g622 ( .A(n_565), .B(n_576), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_566), .B(n_632), .Y(n_690) );
INVx2_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_SL g656 ( .A(n_567), .B(n_583), .Y(n_656) );
AND2x4_ASAP7_75t_SL g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NOR2x1_ASAP7_75t_L g615 ( .A(n_569), .B(n_616), .Y(n_615) );
AND2x4_ASAP7_75t_L g721 ( .A(n_569), .B(n_592), .Y(n_721) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_569), .Y(n_750) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_570), .B(n_742), .Y(n_741) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
OR2x2_ASAP7_75t_L g692 ( .A(n_571), .B(n_693), .Y(n_692) );
NOR2x1_ASAP7_75t_L g757 ( .A(n_571), .B(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g681 ( .A(n_572), .B(n_626), .Y(n_681) );
INVxp33_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2x1p5_ASAP7_75t_L g595 ( .A(n_575), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g755 ( .A(n_575), .B(n_637), .Y(n_755) );
INVx2_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_598), .Y(n_580) );
OAI21xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_584), .B(n_593), .Y(n_581) );
AND2x2_ASAP7_75t_L g716 ( .A(n_583), .B(n_591), .Y(n_716) );
NAND2xp33_ASAP7_75t_R g584 ( .A(n_585), .B(n_590), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g758 ( .A(n_587), .Y(n_758) );
INVx4_ASAP7_75t_L g616 ( .A(n_588), .Y(n_616) );
INVx1_ASAP7_75t_L g735 ( .A(n_589), .Y(n_735) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g729 ( .A(n_591), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_SL g733 ( .A(n_591), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_594), .A2(n_659), .B1(n_763), .B2(n_764), .Y(n_762) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x4_ASAP7_75t_L g623 ( .A(n_597), .B(n_609), .Y(n_623) );
AND2x2_ASAP7_75t_L g637 ( .A(n_597), .B(n_638), .Y(n_637) );
A2O1A1Ixp33_ASAP7_75t_SL g598 ( .A1(n_599), .A2(n_606), .B(n_611), .C(n_614), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx3_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g685 ( .A(n_601), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx1_ASAP7_75t_L g613 ( .A(n_602), .Y(n_613) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g673 ( .A(n_603), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g682 ( .A(n_603), .B(n_604), .Y(n_682) );
INVx1_ASAP7_75t_L g714 ( .A(n_603), .Y(n_714) );
AND2x4_ASAP7_75t_L g695 ( .A(n_604), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g717 ( .A(n_604), .B(n_608), .Y(n_717) );
AND2x2_ASAP7_75t_L g725 ( .A(n_604), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx1_ASAP7_75t_L g700 ( .A(n_608), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_608), .B(n_622), .Y(n_702) );
AND2x2_ASAP7_75t_L g705 ( .A(n_608), .B(n_655), .Y(n_705) );
INVx3_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_609), .B(n_670), .Y(n_719) );
AND2x2_ASAP7_75t_L g647 ( .A(n_610), .B(n_635), .Y(n_647) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g743 ( .A(n_613), .B(n_623), .Y(n_743) );
BUFx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_615), .B(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g627 ( .A(n_616), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_616), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_657), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_641), .Y(n_618) );
OAI222xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_624), .B1(n_628), .B2(n_630), .C1(n_633), .C2(n_636), .Y(n_619) );
INVx1_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_SL g634 ( .A(n_626), .B(n_635), .Y(n_634) );
OR2x6_ASAP7_75t_L g706 ( .A(n_626), .B(n_676), .Y(n_706) );
NAND5xp2_ASAP7_75t_L g709 ( .A(n_626), .B(n_629), .C(n_645), .D(n_710), .E(n_712), .Y(n_709) );
NAND2x1_ASAP7_75t_L g745 ( .A(n_627), .B(n_631), .Y(n_745) );
INVx2_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
NOR2x1_ASAP7_75t_L g675 ( .A(n_632), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_634), .A2(n_725), .B1(n_728), .B2(n_729), .Y(n_724) );
INVx2_ASAP7_75t_L g676 ( .A(n_635), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_635), .B(n_651), .Y(n_688) );
INVx3_ASAP7_75t_L g723 ( .A(n_636), .Y(n_723) );
NAND2x1p5_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
AND2x2_ASAP7_75t_L g668 ( .A(n_637), .B(n_669), .Y(n_668) );
BUFx2_ASAP7_75t_L g701 ( .A(n_637), .Y(n_701) );
INVx2_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g664 ( .A(n_640), .B(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_642), .B(n_653), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_647), .B(n_648), .Y(n_642) );
AND2x4_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
INVx1_ASAP7_75t_L g652 ( .A(n_644), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_647), .A2(n_654), .B1(n_655), .B2(n_656), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_652), .Y(n_648) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x4_ASAP7_75t_SL g734 ( .A(n_651), .B(n_735), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_658), .B(n_666), .Y(n_657) );
AOI21xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_662), .B(n_664), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
BUFx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g703 ( .A(n_674), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .B1(n_681), .B2(n_682), .Y(n_677) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_707), .Y(n_683) );
NOR3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_689), .C(n_697), .Y(n_684) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
BUFx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OA21x2_ASAP7_75t_SL g689 ( .A1(n_690), .A2(n_691), .B(n_695), .Y(n_689) );
NAND2xp33_ASAP7_75t_SL g691 ( .A(n_692), .B(n_694), .Y(n_691) );
AOI21xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_704), .B(n_706), .Y(n_697) );
OAI211xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_701), .B(n_702), .C(n_703), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_701), .A2(n_741), .B1(n_743), .B2(n_744), .Y(n_740) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_731), .Y(n_707) );
NAND4xp25_ASAP7_75t_L g708 ( .A(n_709), .B(n_715), .C(n_722), .D(n_724), .Y(n_708) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g720 ( .A(n_711), .B(n_721), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx1_ASAP7_75t_L g751 ( .A(n_714), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_718), .B2(n_720), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_720), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI21xp5_ASAP7_75t_SL g731 ( .A1(n_732), .A2(n_736), .B(n_740), .Y(n_731) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
INVxp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g746 ( .A(n_747), .B(n_761), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_751), .B(n_752), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B1(n_756), .B2(n_759), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
CKINVDCx11_ASAP7_75t_R g766 ( .A(n_767), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
INVx1_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_779), .Y(n_776) );
CKINVDCx5p33_ASAP7_75t_R g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g788 ( .A(n_782), .Y(n_788) );
CKINVDCx16_ASAP7_75t_R g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_SL g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_SL g792 ( .A(n_793), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_SL g794 ( .A(n_795), .Y(n_794) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_795), .Y(n_806) );
OR2x2_ASAP7_75t_L g795 ( .A(n_796), .B(n_798), .Y(n_795) );
CKINVDCx16_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
endmodule