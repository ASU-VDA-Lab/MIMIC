module real_aes_5941_n_10 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
output n_10;
wire n_17;
wire n_13;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_20;
wire n_18;
CKINVDCx5p33_ASAP7_75t_R g20 ( .A(n_0), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_1), .Y(n_19) );
NOR2xp33_ASAP7_75t_R g13 ( .A(n_2), .B(n_14), .Y(n_13) );
NAND2xp33_ASAP7_75t_R g12 ( .A(n_3), .B(n_13), .Y(n_12) );
NAND2xp33_ASAP7_75t_R g10 ( .A(n_4), .B(n_11), .Y(n_10) );
NAND3xp33_ASAP7_75t_SL g14 ( .A(n_5), .B(n_15), .C(n_16), .Y(n_14) );
NOR2xp33_ASAP7_75t_R g18 ( .A(n_6), .B(n_7), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_8), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_9), .Y(n_16) );
NOR4xp25_ASAP7_75t_SL g11 ( .A(n_12), .B(n_17), .C(n_19), .D(n_20), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_18), .Y(n_17) );
endmodule