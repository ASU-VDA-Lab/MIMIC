module fake_netlist_6_2834_n_781 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_781);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_781;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_208;
wire n_462;
wire n_607;
wire n_726;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_6),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_72),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_16),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_89),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_119),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_57),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_120),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_161),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_46),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_98),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_87),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_60),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_127),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_146),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_14),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_76),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_30),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_0),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_82),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_15),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_13),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_84),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_18),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_40),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_49),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_90),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_48),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_50),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_132),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_10),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_35),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_22),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_152),
.Y(n_201)
);

NOR2xp67_ASAP7_75t_L g202 ( 
.A(n_75),
.B(n_140),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_21),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_66),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_37),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_114),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_25),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_53),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_52),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_97),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_43),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_150),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_108),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_113),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_99),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_62),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_0),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_47),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_41),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_221),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_221),
.Y(n_225)
);

OAI21x1_ASAP7_75t_L g226 ( 
.A1(n_182),
.A2(n_81),
.B(n_157),
.Y(n_226)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_221),
.Y(n_227)
);

OA21x2_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_1),
.B(n_2),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

AND2x4_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_1),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_165),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_179),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_221),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_191),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_193),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_173),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

OAI22x1_ASAP7_75t_L g244 ( 
.A1(n_190),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_162),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_199),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_205),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

AND2x4_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_5),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_184),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_252)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_215),
.Y(n_255)
);

OA21x2_ASAP7_75t_L g256 ( 
.A1(n_202),
.A2(n_7),
.B(n_8),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_163),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_200),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_164),
.Y(n_259)
);

BUFx8_ASAP7_75t_SL g260 ( 
.A(n_203),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_166),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_167),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_168),
.Y(n_263)
);

BUFx8_ASAP7_75t_SL g264 ( 
.A(n_170),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_171),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_172),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_224),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_R g269 ( 
.A(n_259),
.B(n_174),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_260),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_259),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_260),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_264),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_264),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_261),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_222),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_261),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_258),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_242),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_176),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_229),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_262),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_257),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_266),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_229),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_224),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_224),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_263),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_265),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_222),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_227),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_253),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_253),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_227),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_253),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_232),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_232),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_254),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_238),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_240),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_233),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_227),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_233),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_248),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_248),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_233),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_234),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_246),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_234),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_234),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_L g312 ( 
.A(n_230),
.B(n_177),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_235),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_235),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_246),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_235),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_237),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_237),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_L g319 ( 
.A1(n_280),
.A2(n_231),
.B(n_251),
.C(n_225),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_251),
.Y(n_320)
);

BUFx6f_ASAP7_75t_SL g321 ( 
.A(n_271),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_301),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_281),
.Y(n_324)
);

OR2x6_ASAP7_75t_L g325 ( 
.A(n_276),
.B(n_244),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_294),
.B(n_231),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_297),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_283),
.B(n_237),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_298),
.B(n_230),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_296),
.B(n_178),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_300),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_288),
.B(n_241),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_307),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_289),
.B(n_241),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_303),
.B(n_241),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_282),
.B(n_313),
.Y(n_337)
);

NAND3xp33_ASAP7_75t_L g338 ( 
.A(n_305),
.B(n_252),
.C(n_255),
.Y(n_338)
);

NAND2xp33_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_180),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_290),
.B(n_247),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_281),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_299),
.B(n_183),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_285),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_285),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_276),
.B(n_247),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_317),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_285),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_318),
.B(n_247),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_302),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_312),
.B(n_236),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_304),
.B(n_249),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_268),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_286),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_287),
.Y(n_354)
);

BUFx8_ASAP7_75t_L g355 ( 
.A(n_273),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_302),
.Y(n_356)
);

OR2x6_ASAP7_75t_L g357 ( 
.A(n_278),
.B(n_236),
.Y(n_357)
);

AND2x6_ASAP7_75t_SL g358 ( 
.A(n_309),
.B(n_252),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_275),
.Y(n_359)
);

AO21x1_ASAP7_75t_L g360 ( 
.A1(n_308),
.A2(n_226),
.B(n_225),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_269),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_311),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_316),
.B(n_249),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_314),
.B(n_249),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_L g365 ( 
.A(n_269),
.B(n_186),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_277),
.B(n_250),
.Y(n_366)
);

NAND2xp33_ASAP7_75t_L g367 ( 
.A(n_292),
.B(n_187),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_314),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_302),
.B(n_250),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_284),
.B(n_188),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_293),
.B(n_250),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_279),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_295),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_274),
.B(n_194),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_315),
.B(n_255),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_270),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_272),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_297),
.B(n_195),
.Y(n_378)
);

BUFx5_ASAP7_75t_L g379 ( 
.A(n_267),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_281),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_281),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_281),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_291),
.B(n_255),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_301),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_384),
.Y(n_385)
);

NAND2x1p5_ASAP7_75t_L g386 ( 
.A(n_327),
.B(n_228),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_323),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_368),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_352),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_366),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_328),
.B(n_256),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_333),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_384),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_336),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_335),
.B(n_256),
.Y(n_395)
);

NAND3xp33_ASAP7_75t_SL g396 ( 
.A(n_338),
.B(n_214),
.C(n_201),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_349),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_319),
.B(n_228),
.Y(n_398)
);

AND3x2_ASAP7_75t_SL g399 ( 
.A(n_358),
.B(n_9),
.C(n_10),
.Y(n_399)
);

NOR3xp33_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_213),
.C(n_204),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_322),
.B(n_9),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_362),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_337),
.B(n_196),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_353),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_339),
.A2(n_220),
.B1(n_211),
.B2(n_212),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_383),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_350),
.B(n_326),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_351),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_320),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_361),
.B(n_207),
.Y(n_410)
);

OAI22xp33_ASAP7_75t_L g411 ( 
.A1(n_325),
.A2(n_217),
.B1(n_245),
.B2(n_239),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_364),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_R g413 ( 
.A(n_365),
.B(n_12),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_324),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_340),
.B(n_223),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_330),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_357),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_345),
.B(n_243),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g419 ( 
.A(n_371),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_369),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_348),
.B(n_17),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_347),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_363),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_332),
.B(n_19),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_349),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_334),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_378),
.B(n_11),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_379),
.B(n_20),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_379),
.B(n_23),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_379),
.B(n_24),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_347),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_347),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_329),
.Y(n_433)
);

INVxp33_ASAP7_75t_SL g434 ( 
.A(n_374),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_346),
.B(n_357),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_349),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_370),
.B(n_331),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_381),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_343),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_356),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_381),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_354),
.B(n_26),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_344),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_380),
.Y(n_444)
);

OR2x2_ASAP7_75t_L g445 ( 
.A(n_325),
.B(n_11),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_321),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_382),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_321),
.Y(n_448)
);

OR2x6_ASAP7_75t_L g449 ( 
.A(n_372),
.B(n_359),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_379),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_341),
.Y(n_451)
);

OAI21xp33_ASAP7_75t_L g452 ( 
.A1(n_427),
.A2(n_342),
.B(n_367),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_446),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_397),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_385),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_391),
.A2(n_360),
.B(n_373),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_385),
.Y(n_457)
);

O2A1O1Ixp33_ASAP7_75t_L g458 ( 
.A1(n_409),
.A2(n_377),
.B(n_376),
.C(n_379),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_407),
.B(n_356),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_387),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_393),
.A2(n_356),
.B1(n_355),
.B2(n_29),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_395),
.A2(n_27),
.B(n_28),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_390),
.B(n_31),
.Y(n_463)
);

OA22x2_ASAP7_75t_L g464 ( 
.A1(n_416),
.A2(n_355),
.B1(n_33),
.B2(n_34),
.Y(n_464)
);

O2A1O1Ixp33_ASAP7_75t_SL g465 ( 
.A1(n_398),
.A2(n_32),
.B(n_36),
.C(n_38),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_392),
.B(n_39),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_403),
.B(n_42),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_450),
.A2(n_44),
.B(n_45),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_419),
.B(n_51),
.Y(n_469)
);

AOI21x1_ASAP7_75t_L g470 ( 
.A1(n_415),
.A2(n_54),
.B(n_55),
.Y(n_470)
);

NAND2x1p5_ASAP7_75t_L g471 ( 
.A(n_426),
.B(n_56),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_434),
.B(n_58),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_402),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_435),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_437),
.B(n_59),
.Y(n_475)
);

O2A1O1Ixp33_ASAP7_75t_L g476 ( 
.A1(n_396),
.A2(n_61),
.B(n_63),
.C(n_64),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_389),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_386),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_449),
.Y(n_479)
);

NAND3xp33_ASAP7_75t_SL g480 ( 
.A(n_417),
.B(n_69),
.C(n_70),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_449),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_424),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_412),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_423),
.B(n_77),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_404),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_420),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_486)
);

CKINVDCx14_ASAP7_75t_R g487 ( 
.A(n_445),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_401),
.B(n_83),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_397),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_442),
.B(n_85),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_442),
.B(n_424),
.Y(n_491)
);

OAI21x1_ASAP7_75t_SL g492 ( 
.A1(n_421),
.A2(n_428),
.B(n_429),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_397),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_394),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_425),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_408),
.B(n_86),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_425),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_411),
.B(n_88),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_414),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_406),
.B(n_91),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_450),
.A2(n_92),
.B(n_93),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_400),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_418),
.A2(n_100),
.B(n_101),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_410),
.B(n_102),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_425),
.B(n_103),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_451),
.B(n_388),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_422),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_498),
.A2(n_413),
.B1(n_447),
.B2(n_444),
.Y(n_508)
);

CKINVDCx6p67_ASAP7_75t_R g509 ( 
.A(n_453),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_448),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_456),
.A2(n_430),
.B(n_414),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_482),
.B(n_443),
.Y(n_512)
);

INVx4_ASAP7_75t_SL g513 ( 
.A(n_474),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_454),
.Y(n_514)
);

INVx8_ASAP7_75t_L g515 ( 
.A(n_454),
.Y(n_515)
);

BUFx12f_ASAP7_75t_L g516 ( 
.A(n_479),
.Y(n_516)
);

AOI22x1_ASAP7_75t_L g517 ( 
.A1(n_492),
.A2(n_433),
.B1(n_439),
.B2(n_441),
.Y(n_517)
);

BUFx12f_ASAP7_75t_L g518 ( 
.A(n_481),
.Y(n_518)
);

BUFx2_ASAP7_75t_SL g519 ( 
.A(n_454),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_497),
.B(n_440),
.Y(n_520)
);

NAND2x1p5_ASAP7_75t_L g521 ( 
.A(n_497),
.B(n_440),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_489),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g523 ( 
.A1(n_496),
.A2(n_439),
.B(n_438),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_489),
.Y(n_524)
);

NAND2x1p5_ASAP7_75t_L g525 ( 
.A(n_489),
.B(n_440),
.Y(n_525)
);

BUFx5_ASAP7_75t_L g526 ( 
.A(n_455),
.Y(n_526)
);

AO21x2_ASAP7_75t_L g527 ( 
.A1(n_467),
.A2(n_432),
.B(n_431),
.Y(n_527)
);

BUFx2_ASAP7_75t_SL g528 ( 
.A(n_493),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_457),
.Y(n_529)
);

AO21x2_ASAP7_75t_L g530 ( 
.A1(n_500),
.A2(n_405),
.B(n_436),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_487),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_SL g532 ( 
.A1(n_464),
.A2(n_399),
.B1(n_436),
.B2(n_107),
.Y(n_532)
);

NAND2x1p5_ASAP7_75t_L g533 ( 
.A(n_493),
.B(n_436),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_484),
.A2(n_104),
.B(n_105),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_493),
.Y(n_535)
);

NAND2x1p5_ASAP7_75t_L g536 ( 
.A(n_495),
.B(n_491),
.Y(n_536)
);

OAI21x1_ASAP7_75t_SL g537 ( 
.A1(n_458),
.A2(n_109),
.B(n_110),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_473),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_463),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_462),
.A2(n_112),
.B(n_115),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_495),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_460),
.B(n_116),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_466),
.A2(n_118),
.B(n_121),
.Y(n_543)
);

INVx3_ASAP7_75t_SL g544 ( 
.A(n_488),
.Y(n_544)
);

AO21x2_ASAP7_75t_L g545 ( 
.A1(n_459),
.A2(n_122),
.B(n_124),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_506),
.B(n_125),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_495),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_477),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_485),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_499),
.Y(n_550)
);

AO21x2_ASAP7_75t_L g551 ( 
.A1(n_452),
.A2(n_126),
.B(n_128),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_539),
.B(n_490),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_529),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_543),
.A2(n_469),
.B(n_504),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_526),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_515),
.Y(n_556)
);

AO21x1_ASAP7_75t_L g557 ( 
.A1(n_543),
.A2(n_475),
.B(n_476),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_538),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_541),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_526),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_526),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_539),
.B(n_506),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_526),
.Y(n_563)
);

OAI22xp33_ASAP7_75t_L g564 ( 
.A1(n_544),
.A2(n_472),
.B1(n_507),
.B2(n_471),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g565 ( 
.A1(n_523),
.A2(n_470),
.B(n_501),
.Y(n_565)
);

CKINVDCx11_ASAP7_75t_R g566 ( 
.A(n_509),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_550),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_549),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_532),
.A2(n_461),
.B1(n_480),
.B2(n_502),
.Y(n_569)
);

BUFx12f_ASAP7_75t_L g570 ( 
.A(n_516),
.Y(n_570)
);

OAI21x1_ASAP7_75t_L g571 ( 
.A1(n_511),
.A2(n_468),
.B(n_503),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_513),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_548),
.Y(n_573)
);

OA21x2_ASAP7_75t_L g574 ( 
.A1(n_517),
.A2(n_483),
.B(n_505),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_515),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_540),
.A2(n_478),
.B(n_486),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_541),
.Y(n_577)
);

AO21x1_ASAP7_75t_SL g578 ( 
.A1(n_508),
.A2(n_514),
.B(n_537),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_532),
.A2(n_465),
.B1(n_130),
.B2(n_131),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_550),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_546),
.A2(n_129),
.B1(n_133),
.B2(n_134),
.Y(n_581)
);

OAI21x1_ASAP7_75t_L g582 ( 
.A1(n_534),
.A2(n_135),
.B(n_136),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_514),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_515),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_527),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_546),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_527),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_510),
.B(n_137),
.Y(n_588)
);

BUFx10_ASAP7_75t_L g589 ( 
.A(n_542),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_542),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_525),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_575),
.Y(n_592)
);

O2A1O1Ixp33_ASAP7_75t_SL g593 ( 
.A1(n_554),
.A2(n_547),
.B(n_535),
.C(n_536),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_575),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_R g595 ( 
.A(n_566),
.B(n_518),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_562),
.B(n_568),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_572),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_SL g598 ( 
.A1(n_552),
.A2(n_551),
.B1(n_531),
.B2(n_512),
.Y(n_598)
);

BUFx4f_ASAP7_75t_SL g599 ( 
.A(n_570),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_553),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_586),
.B(n_513),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_R g602 ( 
.A(n_566),
.B(n_524),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_575),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_552),
.B(n_512),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_575),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_559),
.B(n_536),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_584),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_R g608 ( 
.A(n_588),
.B(n_535),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_583),
.B(n_547),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_559),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_573),
.B(n_522),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_558),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_R g613 ( 
.A(n_584),
.B(n_508),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_590),
.B(n_528),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_569),
.A2(n_520),
.B(n_521),
.Y(n_615)
);

CKINVDCx16_ASAP7_75t_R g616 ( 
.A(n_570),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_584),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_564),
.B(n_519),
.Y(n_618)
);

AND2x4_ASAP7_75t_SL g619 ( 
.A(n_589),
.B(n_521),
.Y(n_619)
);

NOR3xp33_ASAP7_75t_SL g620 ( 
.A(n_591),
.B(n_545),
.C(n_551),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_577),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_584),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_580),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_556),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_579),
.A2(n_530),
.B1(n_545),
.B2(n_520),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_556),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_589),
.B(n_581),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_R g628 ( 
.A(n_574),
.B(n_138),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_580),
.B(n_530),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_567),
.B(n_533),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_555),
.B(n_533),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_576),
.A2(n_525),
.B(n_142),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_555),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_567),
.B(n_139),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_589),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_567),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_578),
.B(n_560),
.Y(n_637)
);

AO31x2_ASAP7_75t_L g638 ( 
.A1(n_557),
.A2(n_143),
.A3(n_144),
.B(n_145),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_600),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_637),
.B(n_561),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_609),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_596),
.B(n_557),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_604),
.B(n_563),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_633),
.Y(n_644)
);

CKINVDCx6p67_ASAP7_75t_R g645 ( 
.A(n_616),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_612),
.Y(n_646)
);

BUFx2_ASAP7_75t_SL g647 ( 
.A(n_592),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_629),
.B(n_587),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_602),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_629),
.B(n_587),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_594),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_621),
.B(n_585),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_605),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_607),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_610),
.B(n_574),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_623),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_618),
.B(n_574),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_606),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_606),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_611),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_617),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_636),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_631),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_598),
.B(n_582),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_593),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_622),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_638),
.B(n_582),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_638),
.B(n_565),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_624),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_631),
.Y(n_670)
);

NOR2x1_ASAP7_75t_L g671 ( 
.A(n_635),
.B(n_571),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_627),
.B(n_614),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_630),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_626),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_638),
.B(n_565),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_634),
.Y(n_676)
);

NOR2xp67_ASAP7_75t_L g677 ( 
.A(n_603),
.B(n_147),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_642),
.B(n_615),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_639),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_646),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_658),
.Y(n_681)
);

NAND3xp33_ASAP7_75t_L g682 ( 
.A(n_657),
.B(n_608),
.C(n_628),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_672),
.B(n_597),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_673),
.B(n_632),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_641),
.B(n_601),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_656),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_659),
.Y(n_687)
);

OAI22xp33_ASAP7_75t_L g688 ( 
.A1(n_645),
.A2(n_615),
.B1(n_599),
.B2(n_603),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_662),
.B(n_625),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_640),
.B(n_601),
.Y(n_690)
);

AOI21xp33_ASAP7_75t_L g691 ( 
.A1(n_657),
.A2(n_571),
.B(n_620),
.Y(n_691)
);

NOR2xp67_ASAP7_75t_L g692 ( 
.A(n_660),
.B(n_149),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_663),
.B(n_619),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_656),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_652),
.B(n_613),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_652),
.B(n_595),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_644),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_644),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_645),
.A2(n_151),
.B1(n_153),
.B2(n_155),
.Y(n_699)
);

AND2x4_ASAP7_75t_SL g700 ( 
.A(n_640),
.B(n_670),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_648),
.B(n_156),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_640),
.B(n_158),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_681),
.B(n_655),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_683),
.B(n_696),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_684),
.B(n_664),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_679),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_680),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_697),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_696),
.B(n_648),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_695),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_678),
.B(n_650),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_698),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_678),
.B(n_695),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_686),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_693),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_685),
.B(n_650),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_693),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_710),
.B(n_700),
.Y(n_718)
);

INVxp67_ASAP7_75t_SL g719 ( 
.A(n_703),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_710),
.B(n_687),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_713),
.B(n_689),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_711),
.B(n_694),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_706),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_707),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_705),
.B(n_700),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_705),
.A2(n_688),
.B1(n_682),
.B2(n_699),
.Y(n_726)
);

XOR2x2_ASAP7_75t_L g727 ( 
.A(n_726),
.B(n_704),
.Y(n_727)
);

OAI22xp33_ASAP7_75t_SL g728 ( 
.A1(n_721),
.A2(n_717),
.B1(n_703),
.B2(n_715),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_L g729 ( 
.A(n_720),
.B(n_699),
.Y(n_729)
);

INVxp33_ASAP7_75t_L g730 ( 
.A(n_718),
.Y(n_730)
);

A2O1A1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_719),
.A2(n_692),
.B(n_691),
.C(n_666),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_720),
.B(n_709),
.Y(n_732)
);

NAND3xp33_ASAP7_75t_L g733 ( 
.A(n_729),
.B(n_691),
.C(n_724),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_732),
.B(n_722),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_730),
.B(n_725),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_727),
.Y(n_736)
);

NOR3xp33_ASAP7_75t_L g737 ( 
.A(n_731),
.B(n_688),
.C(n_701),
.Y(n_737)
);

NOR2xp67_ASAP7_75t_L g738 ( 
.A(n_736),
.B(n_723),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_735),
.B(n_649),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_734),
.Y(n_740)
);

AOI211xp5_ASAP7_75t_L g741 ( 
.A1(n_733),
.A2(n_728),
.B(n_664),
.C(n_661),
.Y(n_741)
);

OAI21xp5_ASAP7_75t_SL g742 ( 
.A1(n_737),
.A2(n_702),
.B(n_690),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_740),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_738),
.B(n_716),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_743),
.B(n_739),
.Y(n_745)
);

OAI221xp5_ASAP7_75t_L g746 ( 
.A1(n_744),
.A2(n_741),
.B1(n_742),
.B2(n_669),
.C(n_674),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_743),
.B(n_669),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_747),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_745),
.B(n_674),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_746),
.B(n_666),
.Y(n_750)
);

NOR2x1_ASAP7_75t_L g751 ( 
.A(n_747),
.B(n_661),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_745),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_748),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_752),
.A2(n_701),
.B1(n_667),
.B2(n_653),
.Y(n_754)
);

NAND4xp75_ASAP7_75t_L g755 ( 
.A(n_751),
.B(n_677),
.C(n_671),
.D(n_665),
.Y(n_755)
);

OAI21x1_ASAP7_75t_SL g756 ( 
.A1(n_749),
.A2(n_715),
.B(n_712),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_750),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_752),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_758),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_753),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_757),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_755),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_756),
.Y(n_763)
);

AOI22x1_ASAP7_75t_L g764 ( 
.A1(n_759),
.A2(n_754),
.B1(n_647),
.B2(n_651),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_760),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_763),
.B(n_754),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_763),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_761),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_765),
.B(n_762),
.Y(n_769)
);

AO22x2_ASAP7_75t_L g770 ( 
.A1(n_767),
.A2(n_763),
.B1(n_653),
.B2(n_708),
.Y(n_770)
);

OAI31xp33_ASAP7_75t_L g771 ( 
.A1(n_766),
.A2(n_667),
.A3(n_675),
.B(n_668),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_769),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_770),
.B(n_768),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_771),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_769),
.B(n_764),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_SL g776 ( 
.A1(n_770),
.A2(n_654),
.B1(n_651),
.B2(n_676),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_772),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_777),
.B(n_773),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_778),
.A2(n_774),
.B1(n_775),
.B2(n_776),
.Y(n_779)
);

AOI221xp5_ASAP7_75t_L g780 ( 
.A1(n_779),
.A2(n_654),
.B1(n_651),
.B2(n_714),
.C(n_643),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_780),
.A2(n_654),
.B1(n_651),
.B2(n_714),
.Y(n_781)
);


endmodule