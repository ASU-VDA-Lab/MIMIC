module fake_jpeg_29969_n_112 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_51),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_2),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_47),
.B1(n_45),
.B2(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_1),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_47),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_59),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_58),
.A2(n_61),
.B(n_63),
.C(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_55),
.B(n_41),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_5),
.Y(n_83)
);

NOR2x1_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_41),
.Y(n_61)
);

NAND4xp25_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_4),
.C(n_5),
.D(n_7),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_48),
.B(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_68),
.Y(n_77)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_45),
.B1(n_44),
.B2(n_43),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_39),
.B1(n_43),
.B2(n_6),
.Y(n_71)
);

INVx2_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

NOR3xp33_ASAP7_75t_SL g87 ( 
.A(n_73),
.B(n_8),
.C(n_9),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_39),
.B1(n_20),
.B2(n_21),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_10),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_4),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_19),
.B1(n_33),
.B2(n_32),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_35),
.B1(n_16),
.B2(n_17),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_84),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_90),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_22),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_89),
.C(n_92),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_23),
.C(n_29),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_12),
.C(n_13),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_96),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_78),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_82),
.B(n_14),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_81),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_99),
.C(n_94),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_81),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_24),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_SL g107 ( 
.A(n_104),
.B(n_105),
.C(n_106),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_85),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_105),
.C(n_101),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_91),
.C(n_103),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_102),
.B(n_95),
.C(n_30),
.D(n_25),
.Y(n_112)
);


endmodule