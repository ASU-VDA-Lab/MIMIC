module fake_jpeg_13902_n_557 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_557);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_557;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_12),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_60),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_22),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_61),
.B(n_63),
.Y(n_128)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_22),
.B(n_1),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_64),
.B(n_68),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_1),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_65),
.B(n_77),
.Y(n_150)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_66),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_67),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_19),
.B(n_1),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_23),
.B(n_1),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_70),
.B(n_96),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_75),
.Y(n_193)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_76),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_24),
.B(n_2),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_40),
.Y(n_79)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_79),
.Y(n_166)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_82),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_83),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_84),
.Y(n_164)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_86),
.Y(n_198)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_89),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_18),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_93),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_3),
.Y(n_96)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_97),
.Y(n_194)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_98),
.Y(n_169)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

BUFx10_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g171 ( 
.A(n_101),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_32),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_106),
.Y(n_136)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_37),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_37),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_110),
.Y(n_139)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_27),
.Y(n_108)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_31),
.Y(n_109)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_37),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_20),
.B(n_3),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_5),
.Y(n_149)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_31),
.Y(n_112)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_20),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_116),
.Y(n_140)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_26),
.Y(n_115)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_26),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_27),
.Y(n_117)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_117),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_24),
.B(n_4),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_118),
.B(n_41),
.Y(n_167)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_119),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_124),
.Y(n_143)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_122),
.Y(n_196)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_27),
.Y(n_123)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_35),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_36),
.B(n_44),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_130),
.B(n_150),
.C(n_128),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_76),
.A2(n_58),
.B1(n_59),
.B2(n_55),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_137),
.A2(n_148),
.B1(n_176),
.B2(n_180),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_71),
.A2(n_43),
.B1(n_54),
.B2(n_49),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_149),
.B(n_201),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_62),
.B(n_66),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_151),
.B(n_152),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_59),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_96),
.B(n_56),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_154),
.A2(n_101),
.B(n_82),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_39),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_158),
.B(n_181),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_80),
.B(n_39),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_165),
.B(n_190),
.Y(n_249)
);

NAND3xp33_ASAP7_75t_L g256 ( 
.A(n_167),
.B(n_175),
.C(n_8),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_98),
.A2(n_41),
.B1(n_55),
.B2(n_34),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_168),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_120),
.A2(n_85),
.B1(n_87),
.B2(n_67),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_174),
.A2(n_84),
.B1(n_89),
.B2(n_91),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_115),
.B(n_34),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_71),
.A2(n_27),
.B1(n_54),
.B2(n_43),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_121),
.A2(n_43),
.B1(n_54),
.B2(n_49),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_73),
.B(n_33),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_81),
.B(n_33),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_182),
.B(n_189),
.Y(n_261)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_90),
.B(n_54),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_171),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_92),
.B(n_29),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_95),
.B(n_29),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_121),
.A2(n_49),
.B1(n_43),
.B2(n_35),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_191),
.A2(n_192),
.B1(n_204),
.B2(n_82),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_104),
.A2(n_49),
.B1(n_36),
.B2(n_44),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_78),
.B(n_53),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_119),
.B(n_53),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_6),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_60),
.A2(n_83),
.B1(n_69),
.B2(n_74),
.Y(n_204)
);

BUFx2_ASAP7_75t_SL g205 ( 
.A(n_172),
.Y(n_205)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_205),
.Y(n_309)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_206),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_141),
.A2(n_114),
.B1(n_79),
.B2(n_90),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_207),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_155),
.A2(n_38),
.B1(n_101),
.B2(n_122),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_208),
.A2(n_241),
.B1(n_248),
.B2(n_262),
.Y(n_292)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_209),
.Y(n_319)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_210),
.Y(n_316)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_211),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_126),
.Y(n_212)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_212),
.Y(n_321)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_126),
.Y(n_213)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_213),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_214),
.B(n_240),
.Y(n_324)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_215),
.Y(n_325)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_216),
.Y(n_282)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_217),
.Y(n_286)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_218),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_219),
.A2(n_220),
.B1(n_270),
.B2(n_131),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_134),
.A2(n_123),
.B1(n_99),
.B2(n_108),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_221),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_154),
.A2(n_101),
.B(n_105),
.C(n_103),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_223),
.B(n_266),
.Y(n_274)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_224),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_225),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_125),
.Y(n_226)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_226),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_162),
.A2(n_51),
.B1(n_50),
.B2(n_38),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_227),
.A2(n_250),
.B1(n_183),
.B2(n_156),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_173),
.B(n_82),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_229),
.B(n_231),
.Y(n_306)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_140),
.Y(n_230)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_230),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_232),
.A2(n_242),
.B1(n_264),
.B2(n_131),
.Y(n_294)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_136),
.Y(n_233)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_233),
.Y(n_313)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_138),
.Y(n_235)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_235),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_129),
.Y(n_236)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_236),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_133),
.B(n_117),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_237),
.B(n_239),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_184),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_243),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_143),
.B(n_94),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_184),
.B(n_88),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_135),
.A2(n_100),
.B1(n_97),
.B2(n_50),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_174),
.A2(n_93),
.B1(n_86),
.B2(n_75),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_127),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_144),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_244),
.B(n_245),
.Y(n_290)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_171),
.Y(n_245)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_145),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_247),
.B(n_252),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_135),
.A2(n_51),
.B1(n_57),
.B2(n_72),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_196),
.A2(n_6),
.B(n_7),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_251),
.A2(n_159),
.B(n_178),
.Y(n_301)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_163),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_253),
.B(n_255),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_147),
.B(n_6),
.Y(n_254)
);

NOR2x1p5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_269),
.Y(n_275)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_166),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_256),
.B(n_257),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_157),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_191),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_258),
.B(n_259),
.Y(n_312)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_127),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_148),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_260),
.Y(n_287)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_163),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_129),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_263),
.A2(n_267),
.B1(n_272),
.B2(n_273),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_192),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_166),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_265),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_202),
.B(n_9),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_142),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_142),
.B(n_11),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_271),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_161),
.B(n_11),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_176),
.A2(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_L g271 ( 
.A1(n_180),
.A2(n_12),
.B(n_187),
.C(n_198),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_188),
.Y(n_272)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_156),
.Y(n_273)
);

OA21x2_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_183),
.B(n_178),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_277),
.A2(n_304),
.B1(n_307),
.B2(n_318),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_160),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_281),
.B(n_283),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_254),
.B(n_179),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_179),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_284),
.B(n_285),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_177),
.Y(n_285)
);

AO22x2_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_132),
.B1(n_200),
.B2(n_164),
.Y(n_288)
);

AO21x2_ASAP7_75t_L g332 ( 
.A1(n_288),
.A2(n_320),
.B(n_223),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_294),
.A2(n_296),
.B1(n_300),
.B2(n_272),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_299),
.A2(n_273),
.B1(n_193),
.B2(n_198),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_219),
.A2(n_177),
.B1(n_132),
.B2(n_199),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_301),
.A2(n_238),
.B(n_240),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_260),
.A2(n_186),
.B1(n_164),
.B2(n_199),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_229),
.A2(n_200),
.B1(n_186),
.B2(n_146),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_269),
.B(n_195),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_315),
.B(n_323),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_250),
.A2(n_195),
.B1(n_159),
.B2(n_146),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_220),
.A2(n_194),
.B1(n_188),
.B2(n_193),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_222),
.B(n_12),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_231),
.B(n_194),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_326),
.B(n_245),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_296),
.A2(n_294),
.B1(n_276),
.B2(n_274),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_328),
.A2(n_337),
.B1(n_350),
.B2(n_367),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_317),
.Y(n_330)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_321),
.Y(n_331)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_331),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_332),
.A2(n_349),
.B1(n_358),
.B2(n_364),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_310),
.B(n_234),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g370 ( 
.A(n_333),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_289),
.B(n_246),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_334),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_336),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_276),
.A2(n_228),
.B1(n_261),
.B2(n_270),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_297),
.B(n_226),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_338),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_225),
.C(n_240),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_341),
.B(n_279),
.C(n_275),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_327),
.Y(n_342)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_342),
.Y(n_369)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_321),
.Y(n_343)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_343),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_290),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_344),
.B(n_346),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_306),
.B(n_225),
.Y(n_345)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_345),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_281),
.B(n_255),
.Y(n_346)
);

INVx8_ASAP7_75t_L g347 ( 
.A(n_317),
.Y(n_347)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_347),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_301),
.A2(n_251),
.B(n_212),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_348),
.A2(n_352),
.B(n_359),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_287),
.A2(n_235),
.B1(n_244),
.B2(n_247),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_274),
.A2(n_263),
.B1(n_236),
.B2(n_211),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_291),
.Y(n_351)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_351),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_313),
.B(n_265),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_353),
.B(n_356),
.Y(n_380)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_291),
.Y(n_354)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_354),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_295),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_355),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_293),
.B(n_216),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_280),
.Y(n_357)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_357),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_278),
.A2(n_221),
.B1(n_218),
.B2(n_217),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_323),
.B(n_209),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_298),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_360),
.A2(n_361),
.B1(n_309),
.B2(n_319),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_314),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_275),
.B(n_212),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_362),
.B(n_366),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_308),
.B(n_213),
.Y(n_363)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_363),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_277),
.A2(n_210),
.B1(n_224),
.B2(n_215),
.Y(n_364)
);

AND2x2_ASAP7_75t_SL g365 ( 
.A(n_324),
.B(n_283),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_365),
.B(n_277),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_275),
.B(n_243),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_368),
.A2(n_332),
.B1(n_340),
.B2(n_364),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_324),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_371),
.B(n_378),
.C(n_379),
.Y(n_427)
);

OAI32xp33_ASAP7_75t_L g372 ( 
.A1(n_329),
.A2(n_312),
.A3(n_284),
.B1(n_315),
.B2(n_285),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_372),
.B(n_329),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_374),
.A2(n_376),
.B1(n_403),
.B2(n_362),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_332),
.A2(n_300),
.B1(n_292),
.B2(n_303),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_353),
.B(n_365),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_383),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_384),
.B(n_385),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_365),
.B(n_304),
.Y(n_385)
);

AOI322xp5_ASAP7_75t_L g386 ( 
.A1(n_337),
.A2(n_328),
.A3(n_345),
.B1(n_367),
.B2(n_363),
.C1(n_350),
.C2(n_333),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_386),
.B(n_355),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_365),
.B(n_303),
.C(n_314),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_388),
.B(n_389),
.C(n_331),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_336),
.B(n_282),
.C(n_286),
.Y(n_389)
);

OAI22x1_ASAP7_75t_L g399 ( 
.A1(n_340),
.A2(n_288),
.B1(n_311),
.B2(n_325),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_399),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_332),
.A2(n_288),
.B1(n_322),
.B2(n_316),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_373),
.Y(n_404)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_404),
.Y(n_453)
);

FAx1_ASAP7_75t_L g405 ( 
.A(n_384),
.B(n_348),
.CI(n_332),
.CON(n_405),
.SN(n_405)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_405),
.A2(n_395),
.B(n_381),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_390),
.A2(n_332),
.B1(n_392),
.B2(n_374),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_406),
.A2(n_413),
.B1(n_401),
.B2(n_399),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_407),
.B(n_409),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_385),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_408),
.B(n_421),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_382),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_398),
.Y(n_410)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_410),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_412),
.A2(n_349),
.B1(n_396),
.B2(n_387),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_390),
.A2(n_335),
.B1(n_346),
.B2(n_368),
.Y(n_413)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_398),
.Y(n_415)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_415),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_371),
.B(n_339),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_416),
.B(n_432),
.C(n_433),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_400),
.B(n_344),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_417),
.B(n_419),
.Y(n_442)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_377),
.Y(n_418)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_418),
.Y(n_447)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_394),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_366),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_420),
.A2(n_423),
.B1(n_429),
.B2(n_430),
.Y(n_445)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_369),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_422),
.B(n_380),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_403),
.A2(n_335),
.B1(n_360),
.B2(n_288),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_382),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_424),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_375),
.B(n_356),
.Y(n_425)
);

XNOR2x2_ASAP7_75t_SL g450 ( 
.A(n_425),
.B(n_426),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_375),
.B(n_339),
.Y(n_426)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_369),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_370),
.A2(n_359),
.B1(n_352),
.B2(n_343),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_388),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_431),
.A2(n_395),
.B1(n_389),
.B2(n_376),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_379),
.B(n_358),
.Y(n_432)
);

OA22x2_ASAP7_75t_L g434 ( 
.A1(n_412),
.A2(n_423),
.B1(n_405),
.B2(n_428),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_434),
.B(n_459),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_427),
.B(n_378),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_435),
.B(n_437),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_427),
.B(n_380),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_439),
.A2(n_456),
.B(n_414),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_440),
.B(n_458),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_441),
.B(n_411),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_443),
.A2(n_448),
.B1(n_452),
.B2(n_440),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_406),
.A2(n_381),
.B1(n_397),
.B2(n_372),
.Y(n_448)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_449),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_396),
.C(n_351),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_454),
.C(n_460),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_428),
.A2(n_387),
.B1(n_391),
.B2(n_393),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_433),
.B(n_393),
.C(n_361),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_414),
.A2(n_253),
.B(n_262),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_416),
.B(n_327),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_407),
.A2(n_391),
.B1(n_347),
.B2(n_330),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_286),
.C(n_282),
.Y(n_460)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_447),
.Y(n_463)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_463),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_464),
.B(n_465),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_441),
.B(n_411),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_SL g467 ( 
.A(n_439),
.B(n_405),
.C(n_420),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_467),
.A2(n_479),
.B(n_482),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_446),
.B(n_426),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_468),
.B(n_473),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_435),
.B(n_408),
.C(n_425),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_436),
.C(n_460),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_445),
.B(n_413),
.Y(n_470)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_470),
.Y(n_488)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_438),
.Y(n_471)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_471),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_442),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_447),
.Y(n_474)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_474),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_457),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_475),
.B(n_477),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_454),
.B(n_404),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_458),
.Y(n_493)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_453),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_480),
.A2(n_449),
.B1(n_434),
.B2(n_455),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_437),
.B(n_305),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_481),
.B(n_450),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_448),
.A2(n_410),
.B(n_415),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_459),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_483),
.B(n_443),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_486),
.B(n_494),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_483),
.Y(n_487)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_487),
.Y(n_510)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_490),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_462),
.B(n_436),
.C(n_451),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_491),
.B(n_502),
.C(n_466),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_493),
.B(n_481),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_462),
.B(n_455),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_495),
.A2(n_487),
.B1(n_502),
.B2(n_499),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_469),
.B(n_450),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_497),
.B(n_501),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_467),
.A2(n_444),
.B(n_452),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_500),
.A2(n_461),
.B(n_456),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_466),
.B(n_434),
.C(n_438),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_479),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_503),
.A2(n_515),
.B1(n_512),
.B2(n_510),
.Y(n_522)
);

AND2x4_ASAP7_75t_SL g504 ( 
.A(n_484),
.B(n_472),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_504),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_496),
.A2(n_470),
.B1(n_495),
.B2(n_490),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_507),
.B(n_508),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_500),
.A2(n_461),
.B1(n_472),
.B2(n_482),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_509),
.B(n_516),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_511),
.B(n_513),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_489),
.B(n_498),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_512),
.B(n_514),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_475),
.Y(n_513)
);

NAND3xp33_ASAP7_75t_SL g514 ( 
.A(n_489),
.B(n_484),
.C(n_434),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_517),
.A2(n_478),
.B1(n_471),
.B2(n_485),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_504),
.B(n_517),
.Y(n_519)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_519),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_521),
.B(n_526),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_522),
.B(n_525),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_504),
.B(n_497),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_503),
.A2(n_477),
.B1(n_463),
.B2(n_474),
.Y(n_526)
);

AOI221xp5_ASAP7_75t_L g527 ( 
.A1(n_516),
.A2(n_478),
.B1(n_501),
.B2(n_465),
.C(n_464),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_527),
.A2(n_508),
.B1(n_492),
.B2(n_506),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_505),
.B(n_491),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_511),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_530),
.B(n_534),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_524),
.B(n_505),
.Y(n_533)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_533),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_518),
.B(n_486),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_535),
.A2(n_519),
.B1(n_520),
.B2(n_527),
.Y(n_543)
);

OAI221xp5_ASAP7_75t_L g536 ( 
.A1(n_525),
.A2(n_506),
.B1(n_492),
.B2(n_347),
.C(n_330),
.Y(n_536)
);

OA21x2_ASAP7_75t_SL g541 ( 
.A1(n_536),
.A2(n_528),
.B(n_520),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_523),
.B(n_357),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_538),
.A2(n_319),
.B(n_302),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_528),
.A2(n_357),
.B(n_354),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_539),
.A2(n_325),
.B(n_305),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_541),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_531),
.A2(n_537),
.B(n_532),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_542),
.B(n_543),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_545),
.B(n_546),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_540),
.B(n_531),
.Y(n_548)
);

OAI321xp33_ASAP7_75t_L g552 ( 
.A1(n_548),
.A2(n_153),
.A3(n_163),
.B1(n_302),
.B2(n_544),
.C(n_549),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_544),
.A2(n_539),
.B1(n_316),
.B2(n_280),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_551),
.B(n_153),
.C(n_550),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_552),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_554),
.B(n_553),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_555),
.B(n_547),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_556),
.B(n_153),
.Y(n_557)
);


endmodule