module real_aes_4140_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_1289, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_1287, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_1288, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_1289;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_1287;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_1288;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_592;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_400;
wire n_1160;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_417;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_552;
wire n_590;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_859;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1161;
wire n_686;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_837;
wire n_829;
wire n_1030;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_580;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1162;
wire n_762;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_414;
wire n_776;
wire n_1138;
wire n_890;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_577;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_937;
wire n_773;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_816;
wire n_625;
wire n_953;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_609;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1054;
wire n_1050;
wire n_426;
wire n_1134;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1060;
wire n_1154;
wire n_632;
wire n_714;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1033;
wire n_1028;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1240;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_974;
wire n_857;
wire n_376;
wire n_491;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1198;
wire n_993;
wire n_819;
wire n_737;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_449;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1273;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_698;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_483;
wire n_394;
wire n_1280;
wire n_729;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_603;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_855;
wire n_429;
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_0), .A2(n_231), .B1(n_574), .B2(n_669), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_1), .A2(n_327), .B1(n_524), .B2(n_534), .Y(n_697) );
INVx1_ASAP7_75t_L g558 ( .A(n_2), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_3), .A2(n_272), .B1(n_497), .B2(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g1270 ( .A(n_4), .Y(n_1270) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_5), .A2(n_253), .B1(n_514), .B2(n_534), .Y(n_822) );
INVx1_ASAP7_75t_L g894 ( .A(n_6), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_7), .A2(n_183), .B1(n_436), .B2(n_653), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_8), .A2(n_311), .B1(n_459), .B2(n_572), .Y(n_797) );
AOI22xp33_ASAP7_75t_SL g508 ( .A1(n_9), .A2(n_296), .B1(n_509), .B2(n_511), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g1275 ( .A1(n_10), .A2(n_144), .B1(n_736), .B2(n_850), .Y(n_1275) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_11), .A2(n_212), .B1(n_497), .B2(n_968), .Y(n_967) );
AOI221xp5_ASAP7_75t_L g1267 ( .A1(n_12), .A2(n_285), .B1(n_594), .B2(n_1268), .C(n_1269), .Y(n_1267) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_13), .A2(n_83), .B1(n_486), .B2(n_665), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_14), .A2(n_234), .B1(n_515), .B2(n_690), .Y(n_877) );
INVx1_ASAP7_75t_L g562 ( .A(n_15), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_16), .A2(n_302), .B1(n_484), .B2(n_486), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_17), .A2(n_19), .B1(n_484), .B2(n_669), .Y(n_923) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_18), .A2(n_80), .B1(n_614), .B2(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_20), .B(n_394), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_21), .A2(n_137), .B1(n_496), .B2(n_690), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g1246 ( .A1(n_22), .A2(n_176), .B1(n_757), .B2(n_1247), .Y(n_1246) );
AOI21xp33_ASAP7_75t_L g931 ( .A1(n_23), .A2(n_436), .B(n_932), .Y(n_931) );
AOI22xp5_ASAP7_75t_L g808 ( .A1(n_24), .A2(n_239), .B1(n_497), .B2(n_579), .Y(n_808) );
INVx1_ASAP7_75t_L g814 ( .A(n_25), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g1251 ( .A1(n_26), .A2(n_300), .B1(n_479), .B2(n_481), .Y(n_1251) );
INVx1_ASAP7_75t_L g555 ( .A(n_27), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g1243 ( .A1(n_28), .A2(n_291), .B1(n_594), .B2(n_841), .C(n_1244), .Y(n_1243) );
AOI221x1_ASAP7_75t_L g499 ( .A1(n_29), .A2(n_96), .B1(n_500), .B2(n_501), .C(n_502), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_30), .A2(n_355), .B1(n_624), .B2(n_625), .Y(n_638) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_31), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_32), .A2(n_38), .B1(n_574), .B2(n_669), .Y(n_798) );
INVx1_ASAP7_75t_L g654 ( .A(n_33), .Y(n_654) );
INVx1_ASAP7_75t_L g958 ( .A(n_34), .Y(n_958) );
AOI22xp5_ASAP7_75t_L g1012 ( .A1(n_34), .A2(n_267), .B1(n_1013), .B2(n_1015), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_35), .A2(n_372), .B1(n_445), .B2(n_454), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_36), .A2(n_276), .B1(n_614), .B2(n_906), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_37), .A2(n_94), .B1(n_770), .B2(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g869 ( .A(n_39), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g1030 ( .A1(n_39), .A2(n_193), .B1(n_1013), .B2(n_1015), .Y(n_1030) );
AOI21xp33_ASAP7_75t_L g977 ( .A1(n_40), .A2(n_701), .B(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g704 ( .A(n_41), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_42), .A2(n_148), .B1(n_740), .B2(n_810), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_43), .A2(n_354), .B1(n_1017), .B2(n_1023), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_44), .A2(n_246), .B1(n_852), .B2(n_930), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_45), .A2(n_203), .B1(n_1000), .B2(n_1004), .Y(n_999) );
INVxp33_ASAP7_75t_SL g1057 ( .A(n_46), .Y(n_1057) );
AOI22xp33_ASAP7_75t_SL g758 ( .A1(n_47), .A2(n_299), .B1(n_438), .B2(n_759), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_48), .A2(n_116), .B1(n_692), .B2(n_693), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_49), .A2(n_62), .B1(n_1007), .B2(n_1010), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_50), .B(n_651), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_51), .A2(n_312), .B1(n_459), .B2(n_475), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g1252 ( .A1(n_52), .A2(n_361), .B1(n_466), .B2(n_497), .Y(n_1252) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_53), .A2(n_304), .B1(n_609), .B2(n_757), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_54), .A2(n_229), .B1(n_497), .B2(n_625), .Y(n_921) );
AOI22xp5_ASAP7_75t_L g969 ( .A1(n_55), .A2(n_60), .B1(n_574), .B2(n_970), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_56), .A2(n_135), .B1(n_692), .B2(n_693), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_57), .A2(n_342), .B1(n_769), .B2(n_770), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_58), .A2(n_243), .B1(n_459), .B2(n_475), .Y(n_924) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_59), .A2(n_358), .B1(n_566), .B2(n_567), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_61), .A2(n_343), .B1(n_527), .B2(n_566), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_63), .A2(n_112), .B1(n_624), .B2(n_625), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_64), .B(n_610), .Y(n_649) );
AOI21xp33_ASAP7_75t_L g760 ( .A1(n_65), .A2(n_761), .B(n_762), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_66), .A2(n_368), .B1(n_479), .B2(n_481), .Y(n_667) );
OA22x2_ASAP7_75t_L g399 ( .A1(n_67), .A2(n_157), .B1(n_394), .B2(n_398), .Y(n_399) );
INVx1_ASAP7_75t_L g434 ( .A(n_67), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_68), .A2(n_141), .B1(n_692), .B2(n_693), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g1016 ( .A1(n_69), .A2(n_288), .B1(n_1017), .B2(n_1018), .Y(n_1016) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_70), .A2(n_322), .B1(n_515), .B2(n_519), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g1250 ( .A1(n_71), .A2(n_106), .B1(n_475), .B2(n_943), .Y(n_1250) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_72), .A2(n_115), .B1(n_560), .B2(n_852), .Y(n_975) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_73), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g1253 ( .A1(n_74), .A2(n_190), .B1(n_669), .B2(n_773), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_75), .A2(n_147), .B1(n_454), .B2(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_76), .A2(n_363), .B1(n_496), .B2(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g1135 ( .A(n_77), .Y(n_1135) );
AOI22xp5_ASAP7_75t_L g972 ( .A1(n_78), .A2(n_222), .B1(n_459), .B2(n_572), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_79), .B(n_557), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_81), .A2(n_316), .B1(n_459), .B2(n_466), .Y(n_458) );
INVx1_ASAP7_75t_L g397 ( .A(n_82), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_82), .B(n_175), .Y(n_428) );
OAI21xp33_ASAP7_75t_L g442 ( .A1(n_82), .A2(n_157), .B(n_443), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_84), .A2(n_337), .B1(n_479), .B2(n_481), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_85), .A2(n_263), .B1(n_479), .B2(n_481), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_86), .A2(n_219), .B1(n_481), .B2(n_740), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_87), .A2(n_235), .B1(n_609), .B2(n_610), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_88), .A2(n_177), .B1(n_594), .B2(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g897 ( .A(n_89), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_90), .A2(n_224), .B1(n_621), .B2(n_622), .Y(n_637) );
AOI21xp33_ASAP7_75t_L g676 ( .A1(n_91), .A2(n_594), .B(n_677), .Y(n_676) );
XOR2x2_ASAP7_75t_L g881 ( .A(n_92), .B(n_882), .Y(n_881) );
INVxp33_ASAP7_75t_L g1049 ( .A(n_92), .Y(n_1049) );
AND2x4_ASAP7_75t_L g1003 ( .A(n_93), .B(n_270), .Y(n_1003) );
INVx1_ASAP7_75t_L g1009 ( .A(n_93), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_95), .A2(n_228), .B1(n_616), .B2(n_858), .Y(n_857) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_97), .A2(n_294), .B1(n_479), .B2(n_481), .Y(n_799) );
INVx1_ASAP7_75t_L g592 ( .A(n_98), .Y(n_592) );
INVx1_ASAP7_75t_L g900 ( .A(n_99), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_100), .A2(n_357), .B1(n_479), .B2(n_614), .Y(n_613) );
AO22x1_ASAP7_75t_L g664 ( .A1(n_101), .A2(n_319), .B1(n_486), .B2(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_102), .A2(n_174), .B1(n_610), .B2(n_733), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_103), .A2(n_125), .B1(n_509), .B2(n_511), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_104), .A2(n_146), .B1(n_454), .B2(n_674), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_105), .A2(n_323), .B1(n_674), .B2(n_953), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_107), .B(n_388), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_108), .A2(n_226), .B1(n_454), .B2(n_560), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g1274 ( .A1(n_109), .A2(n_119), .B1(n_757), .B2(n_890), .Y(n_1274) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_110), .A2(n_142), .B1(n_574), .B2(n_575), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_111), .A2(n_201), .B1(n_624), .B2(n_625), .Y(n_941) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_113), .A2(n_332), .B1(n_665), .B2(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g1002 ( .A(n_114), .Y(n_1002) );
AND2x4_ASAP7_75t_L g1005 ( .A(n_114), .B(n_989), .Y(n_1005) );
INVx1_ASAP7_75t_SL g1014 ( .A(n_114), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1264 ( .A1(n_117), .A2(n_353), .B1(n_943), .B2(n_1265), .Y(n_1264) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_118), .B(n_388), .Y(n_679) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_120), .A2(n_124), .B1(n_621), .B2(n_622), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g1034 ( .A1(n_121), .A2(n_238), .B1(n_1017), .B2(n_1018), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_122), .B(n_699), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_123), .A2(n_197), .B1(n_575), .B2(n_864), .Y(n_863) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_126), .A2(n_413), .B(n_419), .Y(n_412) );
AOI33xp33_ASAP7_75t_R g742 ( .A1(n_127), .A2(n_251), .A3(n_391), .B1(n_441), .B2(n_743), .B3(n_1289), .Y(n_742) );
INVx1_ASAP7_75t_L g917 ( .A(n_128), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_129), .A2(n_273), .B1(n_1000), .B2(n_1004), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_130), .A2(n_328), .B1(n_514), .B2(n_515), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_131), .A2(n_265), .B1(n_514), .B2(n_518), .Y(n_694) );
AO22x1_ASAP7_75t_L g1277 ( .A1(n_132), .A2(n_321), .B1(n_616), .B2(n_624), .Y(n_1277) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_133), .A2(n_163), .B1(n_860), .B2(n_861), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_134), .A2(n_240), .B1(n_754), .B2(n_755), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_136), .A2(n_227), .B1(n_616), .B2(n_782), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_138), .A2(n_161), .B1(n_572), .B2(n_719), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_139), .A2(n_262), .B1(n_518), .B2(n_690), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_140), .A2(n_188), .B1(n_651), .B2(n_653), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g812 ( .A1(n_143), .A2(n_307), .B1(n_531), .B2(n_701), .C(n_813), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_145), .A2(n_290), .B1(n_551), .B2(n_713), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_149), .B(n_388), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_150), .A2(n_277), .B1(n_621), .B2(n_943), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_151), .A2(n_371), .B1(n_1007), .B2(n_1010), .Y(n_1037) );
AOI22xp5_ASAP7_75t_L g971 ( .A1(n_152), .A2(n_310), .B1(n_479), .B2(n_481), .Y(n_971) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_153), .A2(n_169), .B1(n_486), .B2(n_625), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_154), .A2(n_336), .B1(n_564), .B2(n_794), .Y(n_793) );
CKINVDCx6p67_ASAP7_75t_R g588 ( .A(n_155), .Y(n_588) );
INVx1_ASAP7_75t_L g411 ( .A(n_156), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_156), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_156), .B(n_216), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_157), .B(n_284), .Y(n_427) );
XNOR2x1_ASAP7_75t_L g686 ( .A(n_158), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g964 ( .A(n_159), .Y(n_964) );
AOI22xp5_ASAP7_75t_L g1033 ( .A1(n_159), .A2(n_168), .B1(n_1013), .B2(n_1015), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_160), .A2(n_181), .B1(n_852), .B2(n_853), .Y(n_851) );
INVx1_ASAP7_75t_L g948 ( .A(n_162), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_164), .A2(n_172), .B1(n_572), .B2(n_719), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_165), .B(n_701), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_166), .A2(n_180), .B1(n_496), .B2(n_519), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_167), .A2(n_257), .B1(n_616), .B2(n_624), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_170), .A2(n_280), .B1(n_484), .B2(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g892 ( .A(n_171), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_173), .A2(n_186), .B1(n_825), .B2(n_890), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_175), .B(n_404), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_178), .A2(n_204), .B1(n_622), .B2(n_625), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_179), .A2(n_345), .B1(n_616), .B2(n_618), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_182), .A2(n_370), .B1(n_777), .B2(n_778), .Y(n_776) );
INVx1_ASAP7_75t_L g951 ( .A(n_184), .Y(n_951) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_185), .A2(n_309), .B1(n_616), .B2(n_618), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_187), .Y(n_529) );
INVx1_ASAP7_75t_L g979 ( .A(n_189), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_191), .B(n_736), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_192), .A2(n_362), .B1(n_496), .B2(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_194), .A2(n_338), .B1(n_454), .B2(n_609), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_195), .A2(n_374), .B1(n_454), .B2(n_674), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_196), .A2(n_260), .B1(n_1023), .B2(n_1054), .Y(n_1137) );
AOI22xp33_ASAP7_75t_SL g1031 ( .A1(n_198), .A2(n_271), .B1(n_1017), .B2(n_1018), .Y(n_1031) );
INVx1_ASAP7_75t_L g549 ( .A(n_199), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_200), .A2(n_236), .B1(n_518), .B2(n_719), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_202), .A2(n_365), .B1(n_701), .B2(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g957 ( .A(n_205), .Y(n_957) );
INVx1_ASAP7_75t_L g710 ( .A(n_206), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_207), .A2(n_320), .B1(n_575), .B2(n_621), .Y(n_1278) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_208), .A2(n_249), .B1(n_780), .B2(n_781), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_209), .A2(n_281), .B1(n_518), .B2(n_519), .Y(n_517) );
XOR2x2_ASAP7_75t_L g726 ( .A(n_210), .B(n_727), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_211), .A2(n_301), .B1(n_860), .B2(n_906), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_213), .A2(n_279), .B1(n_496), .B2(n_531), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_214), .B(n_765), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_215), .A2(n_356), .B1(n_692), .B2(n_693), .Y(n_880) );
INVx1_ASAP7_75t_L g395 ( .A(n_216), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g1024 ( .A1(n_217), .A2(n_221), .B1(n_1013), .B2(n_1015), .Y(n_1024) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_218), .A2(n_335), .B1(n_445), .B2(n_454), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_220), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_223), .A2(n_352), .B1(n_514), .B2(n_518), .Y(n_878) );
INVx1_ASAP7_75t_L g803 ( .A(n_225), .Y(n_803) );
XNOR2x1_ASAP7_75t_L g750 ( .A(n_230), .B(n_751), .Y(n_750) );
XNOR2x2_ASAP7_75t_SL g831 ( .A(n_230), .B(n_751), .Y(n_831) );
INVx1_ASAP7_75t_L g648 ( .A(n_232), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g1260 ( .A1(n_233), .A2(n_1261), .B1(n_1279), .B2(n_1280), .Y(n_1260) );
CKINVDCx5p33_ASAP7_75t_R g1280 ( .A(n_233), .Y(n_1280) );
AOI22xp33_ASAP7_75t_SL g469 ( .A1(n_237), .A2(n_293), .B1(n_470), .B2(n_475), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g838 ( .A1(n_241), .A2(n_839), .B(n_842), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_242), .A2(n_339), .B1(n_848), .B2(n_849), .Y(n_847) );
INVx1_ASAP7_75t_L g1136 ( .A(n_244), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_245), .A2(n_360), .B1(n_527), .B2(n_701), .Y(n_700) );
OAI21x1_ASAP7_75t_L g659 ( .A1(n_247), .A2(n_660), .B(n_680), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_247), .B(n_663), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_248), .A2(n_340), .B1(n_531), .B2(n_699), .C(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_250), .A2(n_259), .B1(n_712), .B2(n_713), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_252), .A2(n_292), .B1(n_713), .B2(n_736), .Y(n_1248) );
INVx1_ASAP7_75t_L g843 ( .A(n_254), .Y(n_843) );
INVx1_ASAP7_75t_L g604 ( .A(n_255), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_256), .B(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g933 ( .A(n_258), .Y(n_933) );
INVx1_ASAP7_75t_L g763 ( .A(n_261), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_264), .A2(n_298), .B1(n_459), .B2(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g885 ( .A(n_266), .Y(n_885) );
INVx1_ASAP7_75t_L g384 ( .A(n_268), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_268), .B(n_477), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_269), .A2(n_645), .B(n_647), .Y(n_644) );
HB1xp67_ASAP7_75t_L g991 ( .A(n_270), .Y(n_991) );
AND2x4_ASAP7_75t_L g1008 ( .A(n_270), .B(n_1009), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_274), .A2(n_283), .B1(n_515), .B2(n_519), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_275), .Y(n_525) );
XNOR2x1_ASAP7_75t_L g705 ( .A(n_278), .B(n_706), .Y(n_705) );
AOI211x1_ASAP7_75t_L g944 ( .A1(n_282), .A2(n_945), .B(n_947), .C(n_954), .Y(n_944) );
INVx1_ASAP7_75t_L g409 ( .A(n_284), .Y(n_409) );
INVxp67_ASAP7_75t_L g453 ( .A(n_284), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_286), .A2(n_364), .B1(n_772), .B2(n_774), .Y(n_771) );
INVx1_ASAP7_75t_L g678 ( .A(n_287), .Y(n_678) );
INVx1_ASAP7_75t_L g595 ( .A(n_289), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g1263 ( .A1(n_295), .A2(n_331), .B1(n_614), .B2(n_906), .Y(n_1263) );
INVx2_ASAP7_75t_L g989 ( .A(n_297), .Y(n_989) );
INVx1_ASAP7_75t_L g1051 ( .A(n_303), .Y(n_1051) );
INVx1_ASAP7_75t_SL g498 ( .A(n_305), .Y(n_498) );
NOR3xp33_ASAP7_75t_L g539 ( .A(n_305), .B(n_540), .C(n_541), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_306), .A2(n_347), .B1(n_436), .B2(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g552 ( .A(n_308), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_313), .A2(n_314), .B1(n_527), .B2(n_534), .Y(n_873) );
AOI21xp33_ASAP7_75t_L g702 ( .A1(n_315), .A2(n_531), .B(n_703), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_317), .A2(n_333), .B1(n_551), .B2(n_560), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_318), .A2(n_329), .B1(n_531), .B2(n_566), .Y(n_872) );
INVx1_ASAP7_75t_L g420 ( .A(n_324), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_325), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g600 ( .A(n_326), .Y(n_600) );
XOR2xp5_ASAP7_75t_L g818 ( .A(n_330), .B(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g1055 ( .A(n_334), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_341), .A2(n_346), .B1(n_557), .B2(n_560), .Y(n_672) );
INVx1_ASAP7_75t_L g800 ( .A(n_344), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_348), .A2(n_369), .B1(n_610), .B2(n_699), .Y(n_874) );
AO22x2_ASAP7_75t_L g543 ( .A1(n_349), .A2(n_544), .B1(n_545), .B2(n_546), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_349), .Y(n_544) );
AND2x2_ASAP7_75t_L g502 ( .A(n_350), .B(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_351), .A2(n_366), .B1(n_618), .B2(n_903), .Y(n_902) );
CKINVDCx5p33_ASAP7_75t_R g1240 ( .A(n_354), .Y(n_1240) );
AOI22xp33_ASAP7_75t_L g1258 ( .A1(n_354), .A2(n_1259), .B1(n_1281), .B2(n_1283), .Y(n_1258) );
INVx1_ASAP7_75t_L g956 ( .A(n_359), .Y(n_956) );
INVx1_ASAP7_75t_L g606 ( .A(n_367), .Y(n_606) );
XOR2x2_ASAP7_75t_L g835 ( .A(n_371), .B(n_836), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g1245 ( .A(n_373), .Y(n_1245) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_984), .B(n_992), .Y(n_375) );
XNOR2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_745), .Y(n_376) );
XNOR2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_628), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AO22x2_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B1(n_583), .B2(n_627), .Y(n_379) );
INVx2_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
AO22x2_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_542), .B1(n_580), .B2(n_581), .Y(n_381) );
INVx1_ASAP7_75t_L g580 ( .A(n_382), .Y(n_580) );
XNOR2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_492), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B(n_489), .Y(n_383) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_456), .Y(n_385) );
NAND3xp33_ASAP7_75t_L g489 ( .A(n_386), .B(n_490), .C(n_491), .Y(n_489) );
AND4x1_ASAP7_75t_L g386 ( .A(n_387), .B(n_412), .C(n_435), .D(n_444), .Y(n_386) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_388), .Y(n_761) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g501 ( .A(n_389), .Y(n_501) );
INVx2_ASAP7_75t_L g712 ( .A(n_389), .Y(n_712) );
INVx2_ASAP7_75t_L g841 ( .A(n_389), .Y(n_841) );
INVx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx3_ASAP7_75t_L g564 ( .A(n_390), .Y(n_564) );
INVx2_ASAP7_75t_L g734 ( .A(n_390), .Y(n_734) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_400), .Y(n_390) );
AND2x2_ASAP7_75t_L g455 ( .A(n_391), .B(n_418), .Y(n_455) );
AND2x2_ASAP7_75t_L g485 ( .A(n_391), .B(n_473), .Y(n_485) );
AND2x4_ASAP7_75t_L g487 ( .A(n_391), .B(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g496 ( .A(n_391), .B(n_473), .Y(n_496) );
AND2x4_ASAP7_75t_L g534 ( .A(n_391), .B(n_418), .Y(n_534) );
AND2x2_ASAP7_75t_L g617 ( .A(n_391), .B(n_473), .Y(n_617) );
AND2x4_ASAP7_75t_L g690 ( .A(n_391), .B(n_463), .Y(n_690) );
AND2x2_ASAP7_75t_L g701 ( .A(n_391), .B(n_400), .Y(n_701) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_399), .Y(n_391) );
INVx1_ASAP7_75t_L g417 ( .A(n_392), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_396), .Y(n_392) );
NAND2xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx2_ASAP7_75t_L g398 ( .A(n_394), .Y(n_398) );
INVx3_ASAP7_75t_L g404 ( .A(n_394), .Y(n_404) );
NAND2xp33_ASAP7_75t_L g410 ( .A(n_394), .B(n_411), .Y(n_410) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_394), .Y(n_425) );
INVx1_ASAP7_75t_L g443 ( .A(n_394), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_395), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
OAI21xp5_ASAP7_75t_L g452 ( .A1(n_397), .A2(n_443), .B(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g416 ( .A(n_399), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g451 ( .A(n_399), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g462 ( .A(n_399), .Y(n_462) );
AND2x4_ASAP7_75t_L g437 ( .A(n_400), .B(n_416), .Y(n_437) );
AND2x4_ASAP7_75t_L g440 ( .A(n_400), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g480 ( .A(n_400), .B(n_461), .Y(n_480) );
AND2x4_ASAP7_75t_L g527 ( .A(n_400), .B(n_441), .Y(n_527) );
AND2x4_ASAP7_75t_L g693 ( .A(n_400), .B(n_461), .Y(n_693) );
AND2x2_ASAP7_75t_L g699 ( .A(n_400), .B(n_416), .Y(n_699) );
AND2x4_ASAP7_75t_L g400 ( .A(n_401), .B(n_406), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g418 ( .A(n_402), .B(n_406), .Y(n_418) );
AND2x2_ASAP7_75t_L g448 ( .A(n_402), .B(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g464 ( .A(n_402), .B(n_465), .Y(n_464) );
AND2x4_ASAP7_75t_L g473 ( .A(n_402), .B(n_474), .Y(n_473) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_405), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_404), .B(n_409), .Y(n_408) );
INVxp67_ASAP7_75t_L g431 ( .A(n_404), .Y(n_431) );
NAND3xp33_ASAP7_75t_L g429 ( .A(n_405), .B(n_430), .C(n_432), .Y(n_429) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g465 ( .A(n_407), .Y(n_465) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g899 ( .A(n_414), .Y(n_899) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx3_ASAP7_75t_L g551 ( .A(n_415), .Y(n_551) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_415), .Y(n_594) );
BUFx3_ASAP7_75t_L g852 ( .A(n_415), .Y(n_852) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
AND2x4_ASAP7_75t_L g531 ( .A(n_416), .B(n_418), .Y(n_531) );
AND2x4_ASAP7_75t_L g461 ( .A(n_417), .B(n_462), .Y(n_461) );
AND2x4_ASAP7_75t_L g482 ( .A(n_418), .B(n_461), .Y(n_482) );
AND2x4_ASAP7_75t_L g692 ( .A(n_418), .B(n_461), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_421), .B(n_678), .Y(n_677) );
NOR2xp67_ASAP7_75t_SL g709 ( .A(n_421), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g794 ( .A(n_421), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_421), .B(n_814), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g978 ( .A(n_421), .B(n_979), .Y(n_978) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_422), .Y(n_568) );
INVx2_ASAP7_75t_L g610 ( .A(n_422), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_422), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_SL g825 ( .A(n_422), .Y(n_825) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx3_ASAP7_75t_L g505 ( .A(n_423), .Y(n_505) );
AO21x2_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B(n_429), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_425), .B(n_450), .Y(n_449) );
HB1xp67_ASAP7_75t_L g990 ( .A(n_426), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_431), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g441 ( .A(n_432), .B(n_442), .Y(n_441) );
BUFx3_ASAP7_75t_L g759 ( .A(n_436), .Y(n_759) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx8_ASAP7_75t_SL g500 ( .A(n_437), .Y(n_500) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_437), .Y(n_557) );
INVx2_ASAP7_75t_L g603 ( .A(n_437), .Y(n_603) );
INVx2_ASAP7_75t_L g652 ( .A(n_437), .Y(n_652) );
BUFx3_ASAP7_75t_L g736 ( .A(n_437), .Y(n_736) );
INVx1_ASAP7_75t_L g955 ( .A(n_438), .Y(n_955) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_439), .A2(n_600), .B1(n_601), .B2(n_604), .Y(n_599) );
INVx3_ASAP7_75t_L g653 ( .A(n_439), .Y(n_653) );
INVx2_ASAP7_75t_L g713 ( .A(n_439), .Y(n_713) );
INVx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_440), .Y(n_560) );
BUFx6f_ASAP7_75t_L g850 ( .A(n_440), .Y(n_850) );
AND2x4_ASAP7_75t_L g468 ( .A(n_441), .B(n_463), .Y(n_468) );
AND2x4_ASAP7_75t_L g472 ( .A(n_441), .B(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g515 ( .A(n_441), .B(n_463), .Y(n_515) );
AND2x4_ASAP7_75t_L g519 ( .A(n_441), .B(n_473), .Y(n_519) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g647 ( .A1(n_446), .A2(n_648), .B(n_649), .Y(n_647) );
OAI21xp5_ASAP7_75t_L g762 ( .A1(n_446), .A2(n_763), .B(n_764), .Y(n_762) );
INVx2_ASAP7_75t_L g890 ( .A(n_446), .Y(n_890) );
INVx4_ASAP7_75t_L g930 ( .A(n_446), .Y(n_930) );
INVx2_ASAP7_75t_L g1247 ( .A(n_446), .Y(n_1247) );
INVx5_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx2_ASAP7_75t_L g609 ( .A(n_447), .Y(n_609) );
BUFx4f_ASAP7_75t_L g674 ( .A(n_447), .Y(n_674) );
BUFx2_ASAP7_75t_L g731 ( .A(n_447), .Y(n_731) );
AND2x4_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .Y(n_447) );
AND2x4_ASAP7_75t_L g524 ( .A(n_448), .B(n_451), .Y(n_524) );
AND2x2_ASAP7_75t_L g566 ( .A(n_448), .B(n_451), .Y(n_566) );
INVx3_ASAP7_75t_L g553 ( .A(n_454), .Y(n_553) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g598 ( .A(n_455), .Y(n_598) );
BUFx3_ASAP7_75t_L g757 ( .A(n_455), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_477), .Y(n_456) );
INVxp67_ASAP7_75t_SL g491 ( .A(n_457), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_469), .Y(n_457) );
BUFx3_ASAP7_75t_L g856 ( .A(n_459), .Y(n_856) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_460), .Y(n_622) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_460), .Y(n_719) );
BUFx6f_ASAP7_75t_L g943 ( .A(n_460), .Y(n_943) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_463), .Y(n_460) );
AND2x4_ASAP7_75t_L g476 ( .A(n_461), .B(n_473), .Y(n_476) );
AND2x4_ASAP7_75t_L g514 ( .A(n_461), .B(n_488), .Y(n_514) );
AND2x4_ASAP7_75t_L g518 ( .A(n_461), .B(n_473), .Y(n_518) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g488 ( .A(n_464), .Y(n_488) );
INVx1_ASAP7_75t_L g474 ( .A(n_465), .Y(n_474) );
BUFx2_ASAP7_75t_L g770 ( .A(n_466), .Y(n_770) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx3_ASAP7_75t_L g579 ( .A(n_467), .Y(n_579) );
INVx5_ASAP7_75t_L g665 ( .A(n_467), .Y(n_665) );
INVx2_ASAP7_75t_L g968 ( .A(n_467), .Y(n_968) );
INVx1_ASAP7_75t_L g1265 ( .A(n_467), .Y(n_1265) );
INVx6_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx12f_ASAP7_75t_L g625 ( .A(n_468), .Y(n_625) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx4_ASAP7_75t_L g575 ( .A(n_471), .Y(n_575) );
INVx4_ASAP7_75t_L g618 ( .A(n_471), .Y(n_618) );
INVx4_ASAP7_75t_L g669 ( .A(n_471), .Y(n_669) );
INVx1_ASAP7_75t_L g782 ( .A(n_471), .Y(n_782) );
INVx2_ASAP7_75t_SL g970 ( .A(n_471), .Y(n_970) );
INVx8_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_473), .Y(n_743) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx12f_ASAP7_75t_L g572 ( .A(n_476), .Y(n_572) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_476), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_483), .Y(n_477) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g512 ( .A(n_480), .Y(n_512) );
BUFx3_ASAP7_75t_L g740 ( .A(n_480), .Y(n_740) );
BUFx5_ASAP7_75t_L g906 ( .A(n_480), .Y(n_906) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_481), .Y(n_777) );
BUFx12f_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g510 ( .A(n_482), .Y(n_510) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_482), .Y(n_614) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx4f_ASAP7_75t_L g574 ( .A(n_485), .Y(n_574) );
BUFx3_ASAP7_75t_L g858 ( .A(n_486), .Y(n_858) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_487), .Y(n_497) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_487), .Y(n_624) );
BUFx12f_ASAP7_75t_L g775 ( .A(n_487), .Y(n_775) );
INVx1_ASAP7_75t_L g586 ( .A(n_492), .Y(n_586) );
NAND2x1_ASAP7_75t_L g492 ( .A(n_493), .B(n_535), .Y(n_492) );
NOR3xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_506), .C(n_516), .Y(n_493) );
OAI22xp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_498), .B1(n_499), .B2(n_1287), .Y(n_494) );
INVx1_ASAP7_75t_L g540 ( .A(n_495), .Y(n_540) );
NOR2xp67_ASAP7_75t_L g506 ( .A(n_498), .B(n_507), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_498), .A2(n_517), .B1(n_520), .B2(n_1288), .Y(n_516) );
INVx1_ASAP7_75t_L g537 ( .A(n_499), .Y(n_537) );
INVx1_ASAP7_75t_L g607 ( .A(n_501), .Y(n_607) );
INVx1_ASAP7_75t_L g646 ( .A(n_501), .Y(n_646) );
INVx4_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx4_ASAP7_75t_L g766 ( .A(n_505), .Y(n_766) );
NAND3xp33_ASAP7_75t_L g535 ( .A(n_507), .B(n_536), .C(n_539), .Y(n_535) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_513), .Y(n_507) );
BUFx4f_ASAP7_75t_L g860 ( .A(n_509), .Y(n_860) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g810 ( .A(n_510), .Y(n_810) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_511), .Y(n_636) );
INVx1_ASAP7_75t_L g862 ( .A(n_511), .Y(n_862) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g541 ( .A(n_517), .Y(n_541) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_519), .Y(n_717) );
INVx1_ASAP7_75t_L g538 ( .A(n_520), .Y(n_538) );
NOR2x1_ASAP7_75t_L g520 ( .A(n_521), .B(n_528), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B1(n_525), .B2(n_526), .Y(n_521) );
INVx4_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B1(n_532), .B2(n_533), .Y(n_528) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g582 ( .A(n_543), .Y(n_582) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_569), .Y(n_546) );
NOR3xp33_ASAP7_75t_SL g547 ( .A(n_548), .B(n_554), .C(n_561), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .B1(n_552), .B2(n_553), .Y(n_548) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx2_ASAP7_75t_L g754 ( .A(n_551), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_556), .B1(n_558), .B2(n_559), .Y(n_554) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OAI21xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B(n_565), .Y(n_561) );
INVx2_ASAP7_75t_L g1268 ( .A(n_563), .Y(n_1268) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g1244 ( .A(n_568), .B(n_1245), .Y(n_1244) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_576), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
BUFx6f_ASAP7_75t_L g780 ( .A(n_572), .Y(n_780) );
INVx1_ASAP7_75t_L g865 ( .A(n_572), .Y(n_865) );
BUFx12f_ASAP7_75t_L g903 ( .A(n_572), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_584), .Y(n_627) );
OAI22xp5_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_586), .B1(n_587), .B2(n_626), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVxp67_ASAP7_75t_SL g626 ( .A(n_587), .Y(n_626) );
XNOR2x1_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
NAND2x1_ASAP7_75t_L g589 ( .A(n_590), .B(n_611), .Y(n_589) );
NOR3xp33_ASAP7_75t_SL g590 ( .A(n_591), .B(n_599), .C(n_605), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B1(n_595), .B2(n_596), .Y(n_591) );
INVx4_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_598), .Y(n_643) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
OAI21xp5_ASAP7_75t_SL g950 ( .A1(n_603), .A2(n_951), .B(n_952), .Y(n_950) );
OAI21xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_607), .B(n_608), .Y(n_605) );
NOR2x1_ASAP7_75t_L g611 ( .A(n_612), .B(n_619), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
BUFx8_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
BUFx6f_ASAP7_75t_L g773 ( .A(n_617), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_623), .Y(n_619) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_622), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B1(n_655), .B2(n_744), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
XOR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_654), .Y(n_632) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_634), .B(n_640), .Y(n_633) );
NAND4xp25_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .C(n_638), .D(n_639), .Y(n_634) );
NAND3xp33_ASAP7_75t_L g640 ( .A(n_641), .B(n_644), .C(n_650), .Y(n_640) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx3_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g848 ( .A(n_652), .Y(n_848) );
INVx1_ASAP7_75t_L g744 ( .A(n_655), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_657), .B1(n_723), .B2(n_724), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OA22x2_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_684), .B1(n_685), .B2(n_722), .Y(n_657) );
INVx2_ASAP7_75t_L g722 ( .A(n_658), .Y(n_722) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_670), .Y(n_660) );
NOR3xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .C(n_666), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NOR3xp33_ASAP7_75t_L g682 ( .A(n_664), .B(n_675), .C(n_683), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_666), .B(n_671), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_675), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx2_ASAP7_75t_SL g844 ( .A(n_674), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_679), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
XNOR2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_705), .Y(n_685) );
OR2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_696), .Y(n_687) );
NAND4xp25_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .C(n_694), .D(n_695), .Y(n_688) );
NAND4xp25_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .C(n_700), .D(n_702), .Y(n_696) );
NOR2x1_ASAP7_75t_L g706 ( .A(n_707), .B(n_715), .Y(n_706) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_711), .C(n_714), .Y(n_707) );
NAND4xp25_ASAP7_75t_L g715 ( .A(n_716), .B(n_718), .C(n_720), .D(n_721), .Y(n_715) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_728), .B(n_737), .Y(n_727) );
NAND4xp25_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .C(n_732), .D(n_735), .Y(n_728) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx6f_ASAP7_75t_L g888 ( .A(n_734), .Y(n_888) );
INVx2_ASAP7_75t_L g893 ( .A(n_736), .Y(n_893) );
NAND4xp25_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .C(n_741), .D(n_742), .Y(n_737) );
BUFx2_ASAP7_75t_L g778 ( .A(n_740), .Y(n_778) );
XNOR2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_911), .Y(n_745) );
OAI21xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_832), .B(n_909), .Y(n_746) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_748), .B(n_910), .Y(n_909) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_783), .B1(n_784), .B2(n_831), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
OR2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_767), .Y(n_751) );
NAND3xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_758), .C(n_760), .Y(n_752) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OAI22xp33_ASAP7_75t_L g896 ( .A1(n_756), .A2(n_897), .B1(n_898), .B2(n_900), .Y(n_896) );
OAI22xp5_ASAP7_75t_L g954 ( .A1(n_756), .A2(n_955), .B1(n_956), .B2(n_957), .Y(n_954) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
BUFx2_ASAP7_75t_L g853 ( .A(n_757), .Y(n_853) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g846 ( .A(n_766), .Y(n_846) );
NOR2xp33_ASAP7_75t_L g932 ( .A(n_766), .B(n_933), .Y(n_932) );
INVx4_ASAP7_75t_L g953 ( .A(n_766), .Y(n_953) );
NOR2xp33_ASAP7_75t_L g1269 ( .A(n_766), .B(n_1270), .Y(n_1269) );
NAND4xp25_ASAP7_75t_L g767 ( .A(n_768), .B(n_771), .C(n_776), .D(n_779), .Y(n_767) );
BUFx3_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
BUFx3_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
BUFx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
XNOR2x1_ASAP7_75t_L g784 ( .A(n_785), .B(n_801), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
XOR2x2_ASAP7_75t_L g787 ( .A(n_788), .B(n_800), .Y(n_787) );
NOR2x1_ASAP7_75t_L g788 ( .A(n_789), .B(n_795), .Y(n_788) );
NAND4xp25_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .C(n_792), .D(n_793), .Y(n_789) );
NAND4xp25_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .C(n_798), .D(n_799), .Y(n_795) );
XNOR2x1_ASAP7_75t_L g801 ( .A(n_802), .B(n_817), .Y(n_801) );
XNOR2x1_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
NOR2x1_ASAP7_75t_L g804 ( .A(n_805), .B(n_811), .Y(n_804) );
NAND4xp25_ASAP7_75t_SL g805 ( .A(n_806), .B(n_807), .C(n_808), .D(n_809), .Y(n_805) );
NAND3xp33_ASAP7_75t_L g811 ( .A(n_812), .B(n_815), .C(n_816), .Y(n_811) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
OR2x2_ASAP7_75t_L g819 ( .A(n_820), .B(n_826), .Y(n_819) );
NAND4xp25_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .C(n_823), .D(n_824), .Y(n_820) );
NAND4xp25_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .C(n_829), .D(n_830), .Y(n_826) );
INVx2_ASAP7_75t_SL g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g910 ( .A(n_833), .Y(n_910) );
AO22x2_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_835), .B1(n_866), .B2(n_908), .Y(n_833) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
NOR2x1_ASAP7_75t_L g836 ( .A(n_837), .B(n_854), .Y(n_836) );
NAND3xp33_ASAP7_75t_L g837 ( .A(n_838), .B(n_847), .C(n_851), .Y(n_837) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OAI21xp5_ASAP7_75t_L g947 ( .A1(n_840), .A2(n_948), .B(n_949), .Y(n_947) );
INVx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
OAI21xp33_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_844), .B(n_845), .Y(n_842) );
BUFx3_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx4_ASAP7_75t_L g895 ( .A(n_850), .Y(n_895) );
INVx2_ASAP7_75t_L g946 ( .A(n_852), .Y(n_946) );
NAND4xp25_ASAP7_75t_L g854 ( .A(n_855), .B(n_857), .C(n_859), .D(n_863), .Y(n_854) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx2_ASAP7_75t_L g908 ( .A(n_866), .Y(n_908) );
XNOR2x1_ASAP7_75t_L g866 ( .A(n_867), .B(n_881), .Y(n_866) );
AOI22x1_ASAP7_75t_L g960 ( .A1(n_867), .A2(n_961), .B1(n_980), .B2(n_981), .Y(n_960) );
INVx2_ASAP7_75t_L g981 ( .A(n_867), .Y(n_981) );
INVx3_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
XNOR2x1_ASAP7_75t_L g868 ( .A(n_869), .B(n_870), .Y(n_868) );
OR2x2_ASAP7_75t_L g870 ( .A(n_871), .B(n_876), .Y(n_870) );
NAND4xp25_ASAP7_75t_L g871 ( .A(n_872), .B(n_873), .C(n_874), .D(n_875), .Y(n_871) );
NAND4xp25_ASAP7_75t_L g876 ( .A(n_877), .B(n_878), .C(n_879), .D(n_880), .Y(n_876) );
NAND2x1_ASAP7_75t_L g882 ( .A(n_883), .B(n_901), .Y(n_882) );
NOR3xp33_ASAP7_75t_L g883 ( .A(n_884), .B(n_891), .C(n_896), .Y(n_883) );
OAI21xp5_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_886), .B(n_889), .Y(n_884) );
INVx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_892), .A2(n_893), .B1(n_894), .B2(n_895), .Y(n_891) );
INVx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
AND4x1_ASAP7_75t_L g901 ( .A(n_902), .B(n_904), .C(n_905), .D(n_907), .Y(n_901) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
AOI22xp5_ASAP7_75t_L g912 ( .A1(n_913), .A2(n_914), .B1(n_934), .B2(n_983), .Y(n_912) );
INVx2_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
BUFx3_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
XNOR2xp5_ASAP7_75t_L g916 ( .A(n_917), .B(n_918), .Y(n_916) );
NOR4xp75_ASAP7_75t_L g918 ( .A(n_919), .B(n_922), .C(n_925), .D(n_928), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_920), .B(n_921), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_923), .B(n_924), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_926), .B(n_927), .Y(n_925) );
NAND2xp5_ASAP7_75t_SL g928 ( .A(n_929), .B(n_931), .Y(n_928) );
INVx2_ASAP7_75t_SL g983 ( .A(n_934), .Y(n_983) );
OA22x2_ASAP7_75t_L g934 ( .A1(n_935), .A2(n_959), .B1(n_960), .B2(n_982), .Y(n_934) );
HB1xp67_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
INVx1_ASAP7_75t_L g982 ( .A(n_936), .Y(n_982) );
XNOR2x1_ASAP7_75t_L g936 ( .A(n_937), .B(n_958), .Y(n_936) );
NAND2x1_ASAP7_75t_L g937 ( .A(n_938), .B(n_944), .Y(n_937) );
AND4x1_ASAP7_75t_L g938 ( .A(n_939), .B(n_940), .C(n_941), .D(n_942), .Y(n_938) );
INVx2_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVxp67_ASAP7_75t_SL g961 ( .A(n_962), .Y(n_961) );
BUFx2_ASAP7_75t_L g980 ( .A(n_962), .Y(n_980) );
XNOR2x1_ASAP7_75t_L g962 ( .A(n_963), .B(n_965), .Y(n_962) );
CKINVDCx5p33_ASAP7_75t_R g963 ( .A(n_964), .Y(n_963) );
NOR2x1_ASAP7_75t_L g965 ( .A(n_966), .B(n_973), .Y(n_965) );
NAND4xp25_ASAP7_75t_L g966 ( .A(n_967), .B(n_969), .C(n_971), .D(n_972), .Y(n_966) );
NAND4xp25_ASAP7_75t_L g973 ( .A(n_974), .B(n_975), .C(n_976), .D(n_977), .Y(n_973) );
INVx2_ASAP7_75t_R g984 ( .A(n_985), .Y(n_984) );
BUFx4_ASAP7_75t_SL g985 ( .A(n_986), .Y(n_985) );
NAND3xp33_ASAP7_75t_L g986 ( .A(n_987), .B(n_990), .C(n_991), .Y(n_986) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_987), .B(n_1256), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_987), .B(n_1257), .Y(n_1282) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
OA21x2_ASAP7_75t_L g1284 ( .A1(n_988), .A2(n_1014), .B(n_1285), .Y(n_1284) );
HB1xp67_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_989), .B(n_1002), .Y(n_1001) );
AND3x4_ASAP7_75t_L g1013 ( .A(n_989), .B(n_1008), .C(n_1014), .Y(n_1013) );
NOR2xp33_ASAP7_75t_L g1256 ( .A(n_990), .B(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g1257 ( .A(n_991), .Y(n_1257) );
OAI221xp5_ASAP7_75t_L g992 ( .A1(n_993), .A2(n_1234), .B1(n_1236), .B2(n_1254), .C(n_1258), .Y(n_992) );
AOI211xp5_ASAP7_75t_L g993 ( .A1(n_994), .A2(n_1133), .B(n_1138), .C(n_1206), .Y(n_993) );
NAND4xp25_ASAP7_75t_L g994 ( .A(n_995), .B(n_1078), .C(n_1101), .D(n_1122), .Y(n_994) );
AOI211xp5_ASAP7_75t_L g995 ( .A1(n_996), .A2(n_1019), .B(n_1039), .C(n_1065), .Y(n_995) );
AOI21xp33_ASAP7_75t_L g1175 ( .A1(n_996), .A2(n_1176), .B(n_1177), .Y(n_1175) );
INVx1_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
NOR2xp33_ASAP7_75t_L g1097 ( .A(n_997), .B(n_1077), .Y(n_1097) );
OR2x2_ASAP7_75t_L g997 ( .A(n_998), .B(n_1011), .Y(n_997) );
INVx1_ASAP7_75t_L g1060 ( .A(n_998), .Y(n_1060) );
INVx1_ASAP7_75t_L g1068 ( .A(n_998), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_999), .B(n_1006), .Y(n_998) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1003), .Y(n_1000) );
AND2x4_ASAP7_75t_L g1007 ( .A(n_1001), .B(n_1008), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_1001), .B(n_1003), .Y(n_1017) );
AND2x4_ASAP7_75t_L g1054 ( .A(n_1001), .B(n_1003), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_1003), .B(n_1005), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_1003), .B(n_1005), .Y(n_1018) );
AND2x4_ASAP7_75t_L g1023 ( .A(n_1003), .B(n_1005), .Y(n_1023) );
CKINVDCx5p33_ASAP7_75t_R g1285 ( .A(n_1003), .Y(n_1285) );
AND2x4_ASAP7_75t_L g1010 ( .A(n_1005), .B(n_1008), .Y(n_1010) );
AND2x4_ASAP7_75t_L g1015 ( .A(n_1005), .B(n_1008), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_1005), .B(n_1008), .Y(n_1050) );
INVx3_ASAP7_75t_L g1048 ( .A(n_1007), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_1011), .B(n_1059), .Y(n_1058) );
OR2x2_ASAP7_75t_L g1061 ( .A(n_1011), .B(n_1046), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1011), .B(n_1077), .Y(n_1076) );
INVx2_ASAP7_75t_L g1093 ( .A(n_1011), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1011), .B(n_1060), .Y(n_1100) );
OR2x2_ASAP7_75t_L g1105 ( .A(n_1011), .B(n_1077), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1011), .B(n_1046), .Y(n_1118) );
OR2x2_ASAP7_75t_L g1131 ( .A(n_1011), .B(n_1060), .Y(n_1131) );
HB1xp67_ASAP7_75t_L g1153 ( .A(n_1011), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1016), .Y(n_1011) );
NOR2x1_ASAP7_75t_R g1019 ( .A(n_1020), .B(n_1025), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_1020), .B(n_1029), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_1020), .B(n_1064), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1020), .B(n_1071), .Y(n_1095) );
NOR2xp33_ASAP7_75t_L g1110 ( .A(n_1020), .B(n_1111), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1020), .B(n_1032), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1020), .B(n_1109), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1020), .B(n_1028), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1020), .B(n_1176), .Y(n_1211) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_SL g1074 ( .A(n_1021), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1021), .B(n_1109), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_1021), .B(n_1144), .Y(n_1143) );
OR2x2_ASAP7_75t_L g1158 ( .A(n_1021), .B(n_1083), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_1021), .B(n_1029), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1021), .B(n_1176), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1024), .Y(n_1021) );
INVx2_ASAP7_75t_L g1056 ( .A(n_1023), .Y(n_1056) );
BUFx2_ASAP7_75t_L g1235 ( .A(n_1023), .Y(n_1235) );
NAND2xp5_ASAP7_75t_SL g1025 ( .A(n_1026), .B(n_1035), .Y(n_1025) );
INVx3_ASAP7_75t_SL g1026 ( .A(n_1027), .Y(n_1026) );
NOR2x1_ASAP7_75t_L g1176 ( .A(n_1027), .B(n_1035), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1032), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_1028), .B(n_1032), .Y(n_1071) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_1029), .B(n_1032), .Y(n_1064) );
OR2x2_ASAP7_75t_L g1083 ( .A(n_1029), .B(n_1032), .Y(n_1083) );
AOI221xp5_ASAP7_75t_L g1196 ( .A1(n_1029), .A2(n_1044), .B1(n_1126), .B2(n_1197), .C(n_1199), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1031), .Y(n_1029) );
O2A1O1Ixp33_ASAP7_75t_L g1065 ( .A1(n_1032), .A2(n_1066), .B(n_1069), .C(n_1075), .Y(n_1065) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1032), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1032), .B(n_1073), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1034), .Y(n_1032) );
NAND2xp5_ASAP7_75t_SL g1040 ( .A(n_1035), .B(n_1041), .Y(n_1040) );
NOR2xp33_ASAP7_75t_L g1067 ( .A(n_1035), .B(n_1068), .Y(n_1067) );
INVx2_ASAP7_75t_L g1080 ( .A(n_1035), .Y(n_1080) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1035), .Y(n_1114) );
INVx2_ASAP7_75t_L g1117 ( .A(n_1035), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1035), .B(n_1071), .Y(n_1144) );
BUFx6f_ASAP7_75t_L g1156 ( .A(n_1035), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_1035), .B(n_1180), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1035), .B(n_1045), .Y(n_1191) );
INVx4_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
OR2x2_ASAP7_75t_L g1072 ( .A(n_1036), .B(n_1073), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1036), .B(n_1077), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1036), .B(n_1046), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1038), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_1040), .A2(n_1043), .B1(n_1061), .B2(n_1062), .Y(n_1039) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1058), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_1044), .B(n_1089), .Y(n_1088) );
INVx2_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1045), .B(n_1103), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1045), .B(n_1079), .Y(n_1219) );
INVx1_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
INVx2_ASAP7_75t_L g1077 ( .A(n_1046), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1046), .B(n_1100), .Y(n_1099) );
OR2x2_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1052), .Y(n_1046) );
OAI22xp5_ASAP7_75t_L g1047 ( .A1(n_1048), .A2(n_1049), .B1(n_1050), .B2(n_1051), .Y(n_1047) );
OAI221xp5_ASAP7_75t_L g1134 ( .A1(n_1048), .A2(n_1050), .B1(n_1135), .B2(n_1136), .C(n_1137), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_1053), .A2(n_1055), .B1(n_1056), .B2(n_1057), .Y(n_1052) );
INVx3_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
AOI221xp5_ASAP7_75t_L g1161 ( .A1(n_1058), .A2(n_1162), .B1(n_1164), .B2(n_1167), .C(n_1174), .Y(n_1161) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1059), .Y(n_1089) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
NOR2xp33_ASAP7_75t_L g1113 ( .A(n_1061), .B(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1061), .Y(n_1166) );
NOR2xp33_ASAP7_75t_L g1182 ( .A(n_1061), .B(n_1068), .Y(n_1182) );
OAI22xp5_ASAP7_75t_L g1224 ( .A1(n_1061), .A2(n_1225), .B1(n_1226), .B2(n_1228), .Y(n_1224) );
OAI221xp5_ASAP7_75t_L g1174 ( .A1(n_1062), .A2(n_1133), .B1(n_1175), .B2(n_1181), .C(n_1183), .Y(n_1174) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1063), .B(n_1076), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_1064), .B(n_1086), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1064), .B(n_1099), .Y(n_1098) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1064), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1064), .B(n_1073), .Y(n_1121) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
INVx2_ASAP7_75t_L g1103 ( .A(n_1068), .Y(n_1103) );
BUFx3_ASAP7_75t_L g1165 ( .A(n_1068), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1068), .B(n_1077), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1072), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1071), .B(n_1073), .Y(n_1126) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1072), .Y(n_1086) );
AND2x4_ASAP7_75t_L g1081 ( .A(n_1073), .B(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
INVx2_ASAP7_75t_L g1124 ( .A(n_1077), .Y(n_1124) );
AOI21xp33_ASAP7_75t_SL g1210 ( .A1(n_1077), .A2(n_1211), .B(n_1212), .Y(n_1210) );
O2A1O1Ixp33_ASAP7_75t_L g1078 ( .A1(n_1079), .A2(n_1084), .B(n_1087), .C(n_1090), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1081), .Y(n_1079) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1080), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_1080), .B(n_1108), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1080), .B(n_1095), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1080), .B(n_1173), .Y(n_1172) );
NOR2xp33_ASAP7_75t_L g1232 ( .A(n_1080), .B(n_1083), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_1081), .B(n_1092), .Y(n_1091) );
INVx2_ASAP7_75t_SL g1170 ( .A(n_1081), .Y(n_1170) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1083), .B(n_1112), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_1084), .A2(n_1100), .B1(n_1187), .B2(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
NOR2xp33_ASAP7_75t_L g1202 ( .A(n_1089), .B(n_1150), .Y(n_1202) );
OAI221xp5_ASAP7_75t_L g1090 ( .A1(n_1091), .A2(n_1093), .B1(n_1094), .B2(n_1096), .C(n_1098), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1092), .B(n_1121), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1093), .B(n_1198), .Y(n_1197) );
CKINVDCx14_ASAP7_75t_R g1223 ( .A(n_1093), .Y(n_1223) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_1093), .B(n_1227), .Y(n_1226) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1099), .Y(n_1233) );
AOI211xp5_ASAP7_75t_L g1122 ( .A1(n_1100), .A2(n_1123), .B(n_1127), .C(n_1130), .Y(n_1122) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1100), .Y(n_1178) );
AOI221xp5_ASAP7_75t_L g1101 ( .A1(n_1102), .A2(n_1106), .B1(n_1110), .B2(n_1113), .C(n_1115), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1104), .Y(n_1102) );
NOR2xp33_ASAP7_75t_L g1192 ( .A(n_1103), .B(n_1133), .Y(n_1192) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1103), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1103), .B(n_1134), .Y(n_1213) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
NOR2xp33_ASAP7_75t_L g1217 ( .A(n_1105), .B(n_1114), .Y(n_1217) );
INVxp67_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1109), .B(n_1156), .Y(n_1163) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1113), .Y(n_1203) );
AOI21xp5_ASAP7_75t_L g1115 ( .A1(n_1116), .A2(n_1119), .B(n_1120), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1117), .B(n_1118), .Y(n_1116) );
NAND2xp67_ASAP7_75t_L g1125 ( .A(n_1117), .B(n_1126), .Y(n_1125) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1118), .Y(n_1157) );
AOI221xp5_ASAP7_75t_SL g1193 ( .A1(n_1118), .A2(n_1142), .B1(n_1172), .B2(n_1194), .C(n_1195), .Y(n_1193) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1119), .Y(n_1205) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
NOR2xp33_ASAP7_75t_L g1225 ( .A(n_1121), .B(n_1173), .Y(n_1225) );
NOR2xp67_ASAP7_75t_SL g1123 ( .A(n_1124), .B(n_1125), .Y(n_1123) );
INVx2_ASAP7_75t_L g1128 ( .A(n_1124), .Y(n_1128) );
NOR2xp33_ASAP7_75t_L g1169 ( .A(n_1124), .B(n_1170), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_1124), .B(n_1172), .Y(n_1171) );
AOI221xp5_ASAP7_75t_L g1214 ( .A1(n_1124), .A2(n_1190), .B1(n_1215), .B2(n_1217), .C(n_1218), .Y(n_1214) );
NOR2xp33_ASAP7_75t_L g1221 ( .A(n_1125), .B(n_1128), .Y(n_1221) );
NOR2xp33_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1129), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1128), .B(n_1209), .Y(n_1208) );
AOI21xp33_ASAP7_75t_L g1230 ( .A1(n_1129), .A2(n_1231), .B(n_1233), .Y(n_1230) );
NOR2xp33_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1132), .Y(n_1130) );
OAI211xp5_ASAP7_75t_L g1162 ( .A1(n_1133), .A2(n_1143), .B(n_1158), .C(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1133), .Y(n_1227) );
INVx2_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
HB1xp67_ASAP7_75t_L g1140 ( .A(n_1134), .Y(n_1140) );
OAI211xp5_ASAP7_75t_L g1138 ( .A1(n_1139), .A2(n_1141), .B(n_1161), .C(n_1193), .Y(n_1138) );
INVx2_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
O2A1O1Ixp33_ASAP7_75t_L g1141 ( .A1(n_1142), .A2(n_1145), .B(n_1151), .C(n_1154), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
NAND3xp33_ASAP7_75t_L g1167 ( .A(n_1143), .B(n_1168), .C(n_1171), .Y(n_1167) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1144), .Y(n_1216) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1146 ( .A(n_1147), .B(n_1149), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
NOR2xp33_ASAP7_75t_L g1184 ( .A(n_1148), .B(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
A2O1A1Ixp33_ASAP7_75t_L g1154 ( .A1(n_1155), .A2(n_1157), .B(n_1158), .C(n_1159), .Y(n_1154) );
AOI221xp5_ASAP7_75t_L g1220 ( .A1(n_1155), .A2(n_1221), .B1(n_1222), .B2(n_1224), .C(n_1230), .Y(n_1220) );
INVx2_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1158), .Y(n_1173) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1158), .B(n_1216), .Y(n_1215) );
CKINVDCx5p33_ASAP7_75t_R g1159 ( .A(n_1160), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1165), .B(n_1166), .Y(n_1164) );
OAI321xp33_ASAP7_75t_L g1206 ( .A1(n_1166), .A2(n_1207), .A3(n_1210), .B1(n_1213), .B2(n_1214), .C(n_1220), .Y(n_1206) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
NOR2xp33_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1179), .Y(n_1177) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
OAI21xp33_ASAP7_75t_L g1183 ( .A1(n_1184), .A2(n_1187), .B(n_1192), .Y(n_1183) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1191), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1192), .Y(n_1200) );
OAI221xp5_ASAP7_75t_L g1195 ( .A1(n_1196), .A2(n_1200), .B1(n_1201), .B2(n_1203), .C(n_1204), .Y(n_1195) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1199), .Y(n_1209) );
INVxp67_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
INVxp67_ASAP7_75t_SL g1207 ( .A(n_1208), .Y(n_1207) );
INVxp67_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
CKINVDCx14_ASAP7_75t_R g1222 ( .A(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
CKINVDCx5p33_ASAP7_75t_R g1234 ( .A(n_1235), .Y(n_1234) );
INVx2_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
INVxp67_ASAP7_75t_SL g1238 ( .A(n_1239), .Y(n_1238) );
XNOR2x1_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1241), .Y(n_1239) );
OR2x2_ASAP7_75t_L g1241 ( .A(n_1242), .B(n_1249), .Y(n_1241) );
NAND3xp33_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1246), .C(n_1248), .Y(n_1242) );
NAND4xp25_ASAP7_75t_SL g1249 ( .A(n_1250), .B(n_1251), .C(n_1252), .D(n_1253), .Y(n_1249) );
CKINVDCx16_ASAP7_75t_R g1254 ( .A(n_1255), .Y(n_1254) );
INVxp67_ASAP7_75t_SL g1259 ( .A(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1261), .Y(n_1279) );
NAND5xp2_ASAP7_75t_L g1261 ( .A(n_1262), .B(n_1266), .C(n_1271), .D(n_1276), .E(n_1278), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1263), .B(n_1264), .Y(n_1262) );
BUFx2_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVxp67_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1274), .B(n_1275), .Y(n_1273) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
BUFx2_ASAP7_75t_SL g1281 ( .A(n_1282), .Y(n_1281) );
HB1xp67_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
endmodule