module fake_netlist_6_4702_n_1761 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1761);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1761;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g160 ( 
.A(n_51),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_35),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_145),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_125),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_10),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_71),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_48),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_63),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_5),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_91),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_117),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_4),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_57),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_53),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_74),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_12),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_77),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_33),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_121),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_76),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_114),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_6),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_60),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_98),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_40),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_42),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_156),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_102),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_81),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_148),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_110),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_42),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_35),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_43),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_23),
.Y(n_196)
);

BUFx2_ASAP7_75t_SL g197 ( 
.A(n_29),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_92),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_15),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_64),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_47),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_39),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_79),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_52),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_84),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_9),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_105),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_13),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_29),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_65),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_82),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_39),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_101),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_36),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_158),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_15),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_67),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_157),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_24),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_68),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_85),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_143),
.Y(n_223)
);

BUFx2_ASAP7_75t_SL g224 ( 
.A(n_62),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_48),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_80),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_142),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_153),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_134),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_89),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_108),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_11),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_9),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_70),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_123),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_45),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_27),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_118),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_58),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_72),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_126),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_4),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_124),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_104),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_37),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_66),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_24),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_23),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_109),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_144),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_13),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_100),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_130),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_40),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_22),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_20),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_150),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_1),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_131),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_127),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_113),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_46),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_26),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_107),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_17),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_21),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_88),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_16),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_8),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_7),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_36),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_45),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_38),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_5),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_22),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_20),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_159),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_49),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_152),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_8),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_59),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_54),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_46),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_47),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_3),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_116),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_50),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_141),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_99),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_93),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_1),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_96),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_17),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_6),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_133),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_34),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_73),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_69),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_137),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_86),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_61),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_78),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_83),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_147),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_132),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_41),
.Y(n_306)
);

BUFx5_ASAP7_75t_L g307 ( 
.A(n_14),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_18),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_115),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_37),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_154),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_129),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_14),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_2),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_38),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_30),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_49),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_188),
.B(n_0),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_305),
.Y(n_319)
);

INVxp33_ASAP7_75t_SL g320 ( 
.A(n_161),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_284),
.Y(n_321)
);

BUFx10_ASAP7_75t_L g322 ( 
.A(n_169),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_192),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_309),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_307),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_171),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_198),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_185),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_0),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_204),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_307),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_205),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_307),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_307),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_211),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_307),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_271),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_307),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_175),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_282),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_214),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_187),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_178),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_216),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_218),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_178),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_227),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_229),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_228),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_178),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_174),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_230),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_309),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_178),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_241),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_250),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_279),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_178),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_199),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_199),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_R g362 ( 
.A(n_163),
.B(n_170),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_229),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_197),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_243),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_268),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_244),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_246),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_290),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_160),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_169),
.B(n_2),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_194),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_189),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_249),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_268),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_312),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_291),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_291),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_252),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_196),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_202),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_165),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_161),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_234),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_281),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_253),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_209),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_257),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_259),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_215),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_181),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_217),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_232),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_329),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_340),
.Y(n_395)
);

OAI21x1_ASAP7_75t_L g396 ( 
.A1(n_330),
.A2(n_222),
.B(n_175),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_340),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_344),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_323),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_352),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_338),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_344),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_340),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_347),
.Y(n_404)
);

NAND2xp33_ASAP7_75t_R g405 ( 
.A(n_320),
.B(n_163),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_357),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_328),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_340),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_340),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_R g410 ( 
.A(n_362),
.B(n_203),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_331),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_347),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_351),
.Y(n_413)
);

NAND2xp33_ASAP7_75t_R g414 ( 
.A(n_333),
.B(n_170),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_336),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_340),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_342),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_354),
.B(n_233),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_324),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_345),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_351),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_324),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_358),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_346),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_R g425 ( 
.A(n_391),
.B(n_264),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_355),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_359),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_348),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_359),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_326),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_326),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_332),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_350),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_353),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_332),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_334),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_334),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_335),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_335),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_337),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_369),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_376),
.Y(n_443)
);

NAND2x1_ASAP7_75t_L g444 ( 
.A(n_371),
.B(n_183),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_383),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_356),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_337),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_339),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_339),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_349),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_384),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_385),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_365),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_367),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_343),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_368),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_349),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_374),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_325),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_349),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_325),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_363),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_380),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_380),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_379),
.Y(n_465)
);

NAND2xp33_ASAP7_75t_SL g466 ( 
.A(n_410),
.B(n_237),
.Y(n_466)
);

AND3x2_ASAP7_75t_L g467 ( 
.A(n_394),
.B(n_318),
.C(n_201),
.Y(n_467)
);

OR2x6_ASAP7_75t_L g468 ( 
.A(n_461),
.B(n_224),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_432),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_408),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_461),
.A2(n_341),
.B1(n_319),
.B2(n_343),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_459),
.B(n_386),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_459),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_418),
.A2(n_382),
.B1(n_373),
.B2(n_370),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_450),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_455),
.Y(n_476)
);

INVx6_ASAP7_75t_L g477 ( 
.A(n_437),
.Y(n_477)
);

BUFx8_ASAP7_75t_SL g478 ( 
.A(n_451),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_388),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_418),
.A2(n_433),
.B1(n_436),
.B2(n_432),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_399),
.B(n_389),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_402),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_433),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_463),
.B(n_325),
.Y(n_484)
);

INVx4_ASAP7_75t_SL g485 ( 
.A(n_437),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_394),
.B(n_321),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_402),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_436),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_438),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_438),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_439),
.B(n_370),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_460),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_463),
.B(n_370),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_464),
.B(n_360),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_439),
.B(n_322),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_464),
.B(n_360),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_407),
.A2(n_364),
.B1(n_266),
.B2(n_269),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_462),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_401),
.B(n_327),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_450),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_440),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_450),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_440),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_411),
.B(n_322),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_431),
.B(n_322),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_401),
.B(n_372),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_449),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_431),
.B(n_322),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_449),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_450),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_431),
.B(n_183),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_408),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_L g513 ( 
.A(n_437),
.B(n_229),
.Y(n_513)
);

OR2x6_ASAP7_75t_L g514 ( 
.A(n_444),
.B(n_381),
.Y(n_514)
);

INVx5_ASAP7_75t_L g515 ( 
.A(n_437),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_462),
.Y(n_516)
);

NAND3xp33_ASAP7_75t_L g517 ( 
.A(n_414),
.B(n_195),
.C(n_193),
.Y(n_517)
);

AND2x6_ASAP7_75t_L g518 ( 
.A(n_431),
.B(n_222),
.Y(n_518)
);

OAI21xp33_ASAP7_75t_SL g519 ( 
.A1(n_396),
.A2(n_286),
.B(n_200),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_398),
.B(n_361),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_396),
.B(n_387),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_448),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_425),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_448),
.B(n_200),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_462),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_448),
.B(n_286),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_415),
.B(n_162),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_448),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_419),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_417),
.B(n_308),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_405),
.A2(n_301),
.B1(n_191),
.B2(n_190),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_420),
.B(n_219),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_419),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_445),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_422),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_422),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_424),
.B(n_172),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_429),
.B(n_172),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_444),
.A2(n_287),
.B1(n_255),
.B2(n_256),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_450),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_SL g542 ( 
.A1(n_434),
.A2(n_186),
.B1(n_285),
.B2(n_316),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_437),
.Y(n_543)
);

BUFx4f_ASAP7_75t_L g544 ( 
.A(n_437),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_422),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_441),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_447),
.B(n_267),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_441),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_447),
.Y(n_549)
);

AND2x2_ASAP7_75t_SL g550 ( 
.A(n_451),
.B(n_167),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_398),
.Y(n_551)
);

BUFx4f_ASAP7_75t_L g552 ( 
.A(n_447),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_404),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_447),
.B(n_450),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_404),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_447),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_447),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_412),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_412),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_413),
.Y(n_560)
);

OR2x6_ASAP7_75t_L g561 ( 
.A(n_413),
.B(n_254),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_421),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_421),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_426),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_426),
.B(n_361),
.Y(n_565)
);

BUFx8_ASAP7_75t_SL g566 ( 
.A(n_400),
.Y(n_566)
);

NAND2x1p5_ASAP7_75t_L g567 ( 
.A(n_457),
.B(n_173),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_427),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_427),
.Y(n_569)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_457),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_428),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_465),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_428),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_408),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_430),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_435),
.B(n_177),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_446),
.B(n_453),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_406),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_430),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_457),
.A2(n_294),
.B1(n_270),
.B2(n_274),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_454),
.B(n_177),
.Y(n_581)
);

INVxp67_ASAP7_75t_SL g582 ( 
.A(n_457),
.Y(n_582)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_457),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_395),
.B(n_366),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_452),
.Y(n_585)
);

BUFx4f_ASAP7_75t_L g586 ( 
.A(n_457),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_L g587 ( 
.A(n_408),
.B(n_229),
.Y(n_587)
);

INVx4_ASAP7_75t_SL g588 ( 
.A(n_408),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_395),
.B(n_277),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_395),
.Y(n_590)
);

INVx6_ASAP7_75t_L g591 ( 
.A(n_408),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_397),
.A2(n_275),
.B1(n_296),
.B2(n_293),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_397),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_456),
.B(n_179),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_397),
.B(n_207),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_403),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_403),
.B(n_366),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_458),
.B(n_179),
.Y(n_598)
);

AND2x2_ASAP7_75t_SL g599 ( 
.A(n_403),
.B(n_210),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_409),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_409),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_423),
.A2(n_220),
.B1(n_317),
.B2(n_236),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_442),
.B(n_182),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_409),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_409),
.A2(n_283),
.B1(n_265),
.B2(n_310),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_409),
.B(n_212),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_409),
.Y(n_607)
);

INVx5_ASAP7_75t_L g608 ( 
.A(n_416),
.Y(n_608)
);

AND2x2_ASAP7_75t_SL g609 ( 
.A(n_416),
.B(n_221),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_416),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_416),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_416),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_416),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_489),
.B(n_223),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_499),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_609),
.B(n_229),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_489),
.B(n_226),
.Y(n_617)
);

AND2x6_ASAP7_75t_SL g618 ( 
.A(n_527),
.B(n_387),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_492),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_490),
.B(n_231),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_499),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_533),
.B(n_314),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_561),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_490),
.B(n_235),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_483),
.B(n_488),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_483),
.B(n_238),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_494),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_609),
.A2(n_180),
.B1(n_184),
.B2(n_190),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_517),
.B(n_180),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_473),
.Y(n_630)
);

NOR2xp67_ASAP7_75t_L g631 ( 
.A(n_523),
.B(n_184),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_494),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_506),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_488),
.B(n_240),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_521),
.A2(n_229),
.B1(n_260),
.B2(n_261),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_561),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_469),
.B(n_288),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_521),
.B(n_229),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_532),
.B(n_191),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_506),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_570),
.A2(n_363),
.B(n_303),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_480),
.B(n_300),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_560),
.B(n_239),
.Y(n_643)
);

AOI22x1_ASAP7_75t_L g644 ( 
.A1(n_521),
.A2(n_363),
.B1(n_239),
.B2(n_297),
.Y(n_644)
);

INVx8_ASAP7_75t_L g645 ( 
.A(n_468),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_496),
.Y(n_646)
);

NOR2xp67_ASAP7_75t_L g647 ( 
.A(n_523),
.B(n_289),
.Y(n_647)
);

AOI221xp5_ASAP7_75t_L g648 ( 
.A1(n_542),
.A2(n_164),
.B1(n_166),
.B2(n_168),
.C(n_176),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_473),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_498),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_L g651 ( 
.A(n_518),
.B(n_229),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_496),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_560),
.B(n_289),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_484),
.B(n_390),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_498),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_584),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_538),
.B(n_292),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_562),
.B(n_579),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_599),
.A2(n_280),
.B1(n_166),
.B2(n_168),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_539),
.B(n_576),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_562),
.B(n_292),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_599),
.A2(n_280),
.B1(n_176),
.B2(n_186),
.Y(n_662)
);

BUFx6f_ASAP7_75t_SL g663 ( 
.A(n_572),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_505),
.B(n_295),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_579),
.B(n_295),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_484),
.B(n_390),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_508),
.B(n_297),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_495),
.B(n_522),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_486),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_558),
.B(n_298),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_561),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_476),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_584),
.Y(n_673)
);

A2O1A1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_519),
.A2(n_392),
.B(n_393),
.C(n_164),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_528),
.B(n_298),
.Y(n_675)
);

A2O1A1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_559),
.A2(n_392),
.B(n_393),
.C(n_299),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_561),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_566),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_516),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_597),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_564),
.B(n_299),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_491),
.B(n_301),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_514),
.A2(n_550),
.B1(n_466),
.B2(n_468),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_597),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_568),
.B(n_302),
.Y(n_685)
);

A2O1A1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_569),
.A2(n_302),
.B(n_304),
.C(n_311),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_573),
.B(n_304),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_SL g688 ( 
.A(n_572),
.B(n_443),
.Y(n_688)
);

NAND3xp33_ASAP7_75t_L g689 ( 
.A(n_474),
.B(n_272),
.C(n_208),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_518),
.A2(n_285),
.B1(n_306),
.B2(n_313),
.Y(n_690)
);

OAI221xp5_ASAP7_75t_L g691 ( 
.A1(n_592),
.A2(n_263),
.B1(n_213),
.B2(n_225),
.C(n_242),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_468),
.A2(n_311),
.B1(n_206),
.B2(n_273),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_571),
.B(n_278),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_571),
.B(n_276),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_581),
.B(n_245),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_493),
.B(n_551),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_514),
.A2(n_247),
.B1(n_248),
.B2(n_251),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_493),
.B(n_258),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_516),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_486),
.B(n_315),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_520),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_594),
.B(n_262),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_566),
.Y(n_703)
);

INVx5_ASAP7_75t_L g704 ( 
.A(n_518),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_525),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_472),
.B(n_306),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_582),
.A2(n_378),
.B(n_377),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_551),
.B(n_316),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_520),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_604),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_479),
.B(n_313),
.Y(n_711)
);

OR2x6_ASAP7_75t_L g712 ( 
.A(n_585),
.B(n_378),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_583),
.A2(n_377),
.B(n_375),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_553),
.B(n_375),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_565),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_525),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_598),
.B(n_315),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_553),
.B(n_55),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_536),
.Y(n_719)
);

BUFx5_ASAP7_75t_L g720 ( 
.A(n_518),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_536),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_555),
.B(n_151),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_555),
.B(n_149),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_563),
.B(n_146),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_471),
.B(n_497),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_546),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_565),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_563),
.B(n_140),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_547),
.A2(n_139),
.B(n_138),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_575),
.B(n_136),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_575),
.B(n_128),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_507),
.B(n_120),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_509),
.B(n_119),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_501),
.Y(n_734)
);

AND2x6_ASAP7_75t_L g735 ( 
.A(n_600),
.B(n_112),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_535),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_468),
.A2(n_111),
.B1(n_106),
.B2(n_103),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_476),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_501),
.B(n_97),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_503),
.B(n_95),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_585),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_481),
.B(n_3),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_602),
.B(n_7),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_503),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_510),
.B(n_549),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_518),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_596),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_546),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_554),
.B(n_94),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_514),
.A2(n_90),
.B1(n_87),
.B2(n_75),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_511),
.A2(n_16),
.B(n_18),
.C(n_19),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_514),
.A2(n_56),
.B1(n_21),
.B2(n_25),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_596),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_482),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_510),
.B(n_19),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_467),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_510),
.B(n_50),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_548),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_482),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_550),
.B(n_524),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_578),
.Y(n_761)
);

BUFx12f_ASAP7_75t_L g762 ( 
.A(n_478),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_556),
.B(n_25),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_L g764 ( 
.A(n_577),
.B(n_26),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_540),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_526),
.B(n_28),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_504),
.B(n_31),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_557),
.B(n_31),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_466),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_603),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_589),
.B(n_32),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_518),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_530),
.B(n_32),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_548),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_580),
.B(n_33),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_543),
.B(n_34),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_487),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_531),
.B(n_41),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_543),
.B(n_43),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_531),
.B(n_534),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_777),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_746),
.A2(n_605),
.B1(n_595),
.B2(n_606),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_660),
.B(n_534),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_746),
.A2(n_552),
.B1(n_544),
.B2(n_545),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_710),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_635),
.A2(n_725),
.B1(n_622),
.B2(n_742),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_719),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_734),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_627),
.B(n_613),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_721),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_696),
.A2(n_544),
.B(n_552),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_660),
.B(n_537),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_760),
.A2(n_477),
.B1(n_529),
.B2(n_607),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_622),
.B(n_610),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_657),
.B(n_610),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_668),
.A2(n_552),
.B(n_544),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_744),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_657),
.B(n_600),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_695),
.B(n_702),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_742),
.B(n_586),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_656),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_625),
.B(n_590),
.Y(n_802)
);

NOR2x1p5_ASAP7_75t_SL g803 ( 
.A(n_720),
.B(n_601),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_741),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_725),
.A2(n_593),
.B(n_590),
.C(n_601),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_695),
.B(n_613),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_726),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_638),
.A2(n_586),
.B(n_611),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_630),
.Y(n_809)
);

O2A1O1Ixp5_ASAP7_75t_L g810 ( 
.A1(n_760),
.A2(n_586),
.B(n_502),
.C(n_475),
.Y(n_810)
);

NOR3xp33_ASAP7_75t_L g811 ( 
.A(n_702),
.B(n_513),
.C(n_587),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_633),
.B(n_478),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_668),
.A2(n_502),
.B(n_475),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_683),
.B(n_485),
.Y(n_814)
);

O2A1O1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_778),
.A2(n_513),
.B(n_587),
.C(n_487),
.Y(n_815)
);

CKINVDCx11_ASAP7_75t_R g816 ( 
.A(n_762),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_748),
.Y(n_817)
);

NOR2x1_ASAP7_75t_R g818 ( 
.A(n_703),
.B(n_477),
.Y(n_818)
);

NOR2xp67_ASAP7_75t_R g819 ( 
.A(n_772),
.B(n_477),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_673),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_706),
.A2(n_477),
.B1(n_475),
.B2(n_541),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_635),
.A2(n_567),
.B1(n_591),
.B2(n_604),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_658),
.A2(n_541),
.B(n_502),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_640),
.B(n_567),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_639),
.A2(n_612),
.B(n_470),
.C(n_512),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_639),
.A2(n_612),
.B(n_470),
.C(n_512),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_745),
.A2(n_541),
.B(n_500),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_717),
.A2(n_470),
.B(n_574),
.C(n_512),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_710),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_669),
.B(n_500),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_706),
.B(n_485),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_R g832 ( 
.A(n_738),
.B(n_591),
.Y(n_832)
);

NAND3xp33_ASAP7_75t_L g833 ( 
.A(n_717),
.B(n_500),
.C(n_470),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_615),
.B(n_567),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_767),
.A2(n_591),
.B1(n_470),
.B2(n_512),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_638),
.A2(n_515),
.B(n_608),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_621),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_704),
.A2(n_574),
.B(n_512),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_674),
.A2(n_616),
.B(n_780),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_704),
.A2(n_574),
.B(n_515),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_711),
.B(n_574),
.Y(n_841)
);

AOI21x1_ASAP7_75t_L g842 ( 
.A1(n_616),
.A2(n_753),
.B(n_747),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_758),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_674),
.A2(n_515),
.B(n_608),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_774),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_711),
.B(n_574),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_654),
.B(n_485),
.Y(n_847)
);

O2A1O1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_778),
.A2(n_44),
.B(n_485),
.C(n_588),
.Y(n_848)
);

OAI21x1_ASAP7_75t_L g849 ( 
.A1(n_619),
.A2(n_588),
.B(n_591),
.Y(n_849)
);

AOI21xp33_ASAP7_75t_L g850 ( 
.A1(n_767),
.A2(n_44),
.B(n_515),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_704),
.A2(n_515),
.B(n_608),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_743),
.A2(n_588),
.B1(n_608),
.B2(n_690),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_680),
.B(n_588),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_704),
.A2(n_608),
.B(n_649),
.Y(n_854)
);

INVxp67_ASAP7_75t_SL g855 ( 
.A(n_649),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_684),
.A2(n_667),
.B(n_651),
.Y(n_856)
);

AO21x1_ASAP7_75t_L g857 ( 
.A1(n_771),
.A2(n_749),
.B(n_755),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_643),
.A2(n_661),
.B(n_665),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_630),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_736),
.Y(n_860)
);

INVx6_ASAP7_75t_L g861 ( 
.A(n_741),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_653),
.A2(n_723),
.B(n_722),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_642),
.A2(n_646),
.B(n_652),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_663),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_632),
.A2(n_709),
.B(n_701),
.Y(n_865)
);

AO21x1_ASAP7_75t_L g866 ( 
.A1(n_749),
.A2(n_757),
.B(n_776),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_712),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_724),
.A2(n_731),
.B(n_728),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_768),
.A2(n_766),
.B(n_765),
.C(n_751),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_730),
.A2(n_698),
.B(n_617),
.Y(n_870)
);

NAND3xp33_ASAP7_75t_L g871 ( 
.A(n_648),
.B(n_629),
.C(n_773),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_614),
.A2(n_620),
.B(n_624),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_739),
.A2(n_710),
.B(n_732),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_666),
.B(n_715),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_650),
.Y(n_875)
);

AO21x1_ASAP7_75t_L g876 ( 
.A1(n_779),
.A2(n_629),
.B(n_773),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_770),
.B(n_769),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_727),
.B(n_754),
.Y(n_878)
);

AO21x1_ASAP7_75t_L g879 ( 
.A1(n_740),
.A2(n_768),
.B(n_718),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_710),
.A2(n_759),
.B(n_655),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_700),
.Y(n_881)
);

BUFx12f_ASAP7_75t_L g882 ( 
.A(n_761),
.Y(n_882)
);

AND2x6_ASAP7_75t_L g883 ( 
.A(n_772),
.B(n_775),
.Y(n_883)
);

AOI21x1_ASAP7_75t_L g884 ( 
.A1(n_626),
.A2(n_634),
.B(n_637),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_630),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_630),
.B(n_636),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_679),
.A2(n_716),
.B(n_705),
.Y(n_887)
);

OAI21xp33_ASAP7_75t_L g888 ( 
.A1(n_659),
.A2(n_662),
.B(n_689),
.Y(n_888)
);

O2A1O1Ixp33_ASAP7_75t_SL g889 ( 
.A1(n_740),
.A2(n_718),
.B(n_733),
.C(n_686),
.Y(n_889)
);

AOI21x1_ASAP7_75t_L g890 ( 
.A1(n_699),
.A2(n_641),
.B(n_664),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_712),
.B(n_647),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_623),
.B(n_671),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_714),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_697),
.B(n_688),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_733),
.A2(n_664),
.B(n_694),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_735),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_628),
.A2(n_764),
.B(n_693),
.C(n_690),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_670),
.A2(n_685),
.B(n_687),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_735),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_682),
.B(n_681),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_675),
.A2(n_682),
.B(n_763),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_675),
.A2(n_729),
.B(n_707),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_631),
.B(n_623),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_708),
.B(n_676),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_672),
.B(n_712),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_713),
.A2(n_708),
.B(n_636),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_671),
.B(n_677),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_766),
.B(n_720),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_618),
.B(n_663),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_677),
.A2(n_737),
.B(n_645),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_756),
.B(n_692),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_645),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_678),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_659),
.B(n_662),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_645),
.A2(n_720),
.B(n_750),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_735),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_678),
.B(n_735),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_L g918 ( 
.A1(n_644),
.A2(n_752),
.B(n_691),
.Y(n_918)
);

BUFx8_ASAP7_75t_L g919 ( 
.A(n_735),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_720),
.B(n_660),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_720),
.Y(n_921)
);

AOI21x1_ASAP7_75t_L g922 ( 
.A1(n_720),
.A2(n_638),
.B(n_668),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_760),
.A2(n_622),
.B1(n_660),
.B2(n_695),
.Y(n_923)
);

NAND2x2_ASAP7_75t_L g924 ( 
.A(n_678),
.B(n_756),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_734),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_660),
.B(n_622),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_777),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_660),
.B(n_622),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_696),
.A2(n_552),
.B(n_544),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_710),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_622),
.A2(n_660),
.B(n_725),
.C(n_702),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_696),
.A2(n_552),
.B(n_544),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_696),
.A2(n_552),
.B(n_544),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_660),
.B(n_622),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_622),
.A2(n_660),
.B(n_725),
.C(n_702),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_660),
.B(n_572),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_710),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_622),
.A2(n_660),
.B(n_725),
.C(n_702),
.Y(n_938)
);

AO21x1_ASAP7_75t_L g939 ( 
.A1(n_616),
.A2(n_742),
.B(n_760),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_734),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_638),
.A2(n_674),
.B(n_519),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_710),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_660),
.B(n_622),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_696),
.A2(n_552),
.B(n_544),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_696),
.A2(n_552),
.B(n_544),
.Y(n_945)
);

AO21x1_ASAP7_75t_L g946 ( 
.A1(n_616),
.A2(n_742),
.B(n_760),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_696),
.A2(n_552),
.B(n_544),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_746),
.A2(n_635),
.B1(n_725),
.B2(n_622),
.Y(n_948)
);

OAI21xp33_ASAP7_75t_L g949 ( 
.A1(n_622),
.A2(n_662),
.B(n_659),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_696),
.A2(n_552),
.B(n_544),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_696),
.A2(n_552),
.B(n_544),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_760),
.A2(n_622),
.B1(n_660),
.B2(n_695),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_696),
.A2(n_552),
.B(n_544),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_746),
.A2(n_635),
.B1(n_725),
.B2(n_622),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_660),
.B(n_622),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_660),
.B(n_622),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_622),
.B(n_633),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_696),
.A2(n_552),
.B(n_544),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_696),
.A2(n_552),
.B(n_544),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_777),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_622),
.B(n_633),
.Y(n_961)
);

OA22x2_ASAP7_75t_L g962 ( 
.A1(n_683),
.A2(n_633),
.B1(n_640),
.B2(n_669),
.Y(n_962)
);

BUFx5_ASAP7_75t_L g963 ( 
.A(n_735),
.Y(n_963)
);

AOI21xp33_ASAP7_75t_L g964 ( 
.A1(n_622),
.A2(n_742),
.B(n_725),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_738),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_760),
.A2(n_622),
.B1(n_660),
.B2(n_695),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_696),
.B(n_660),
.Y(n_967)
);

OAI21x1_ASAP7_75t_L g968 ( 
.A1(n_849),
.A2(n_873),
.B(n_922),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_926),
.B(n_955),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_931),
.A2(n_938),
.B(n_935),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_928),
.B(n_934),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_813),
.A2(n_827),
.B(n_823),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_809),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_872),
.A2(n_870),
.B(n_862),
.Y(n_974)
);

AOI21xp33_ASAP7_75t_L g975 ( 
.A1(n_799),
.A2(n_956),
.B(n_943),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_920),
.A2(n_858),
.B(n_868),
.Y(n_976)
);

AOI221xp5_ASAP7_75t_SL g977 ( 
.A1(n_948),
.A2(n_954),
.B1(n_786),
.B2(n_949),
.C(n_888),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_890),
.A2(n_842),
.B(n_902),
.Y(n_978)
);

AO31x2_ASAP7_75t_L g979 ( 
.A1(n_939),
.A2(n_946),
.A3(n_876),
.B(n_866),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_788),
.Y(n_980)
);

AOI211x1_ASAP7_75t_L g981 ( 
.A1(n_964),
.A2(n_914),
.B(n_786),
.C(n_954),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_967),
.B(n_923),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_952),
.B(n_966),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_964),
.A2(n_948),
.B(n_871),
.C(n_869),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_967),
.B(n_792),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_936),
.B(n_957),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_806),
.A2(n_846),
.B(n_841),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_881),
.B(n_961),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_856),
.A2(n_908),
.B(n_791),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_783),
.B(n_874),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_794),
.B(n_893),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_897),
.A2(n_894),
.B(n_898),
.C(n_863),
.Y(n_992)
);

AND3x4_ASAP7_75t_L g993 ( 
.A(n_892),
.B(n_913),
.C(n_917),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_797),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_941),
.A2(n_839),
.B(n_805),
.Y(n_995)
);

BUFx2_ASAP7_75t_R g996 ( 
.A(n_965),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_900),
.B(n_865),
.Y(n_997)
);

AO31x2_ASAP7_75t_L g998 ( 
.A1(n_828),
.A2(n_857),
.A3(n_826),
.B(n_825),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_905),
.B(n_804),
.Y(n_999)
);

NOR2xp67_ASAP7_75t_L g1000 ( 
.A(n_859),
.B(n_895),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_865),
.B(n_863),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_908),
.A2(n_933),
.B(n_932),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_929),
.A2(n_951),
.B(n_944),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_795),
.A2(n_915),
.B1(n_798),
.B2(n_855),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_911),
.B(n_860),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_839),
.A2(n_941),
.B(n_811),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_809),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_801),
.B(n_820),
.Y(n_1008)
);

INVxp67_ASAP7_75t_L g1009 ( 
.A(n_877),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_891),
.B(n_824),
.Y(n_1010)
);

AO31x2_ASAP7_75t_L g1011 ( 
.A1(n_879),
.A2(n_784),
.A3(n_782),
.B(n_901),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_945),
.A2(n_950),
.B(n_947),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_787),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_L g1014 ( 
.A(n_918),
.B(n_850),
.C(n_904),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_832),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_810),
.A2(n_796),
.B(n_880),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_953),
.A2(n_958),
.B(n_959),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_808),
.A2(n_838),
.B(n_887),
.Y(n_1018)
);

AOI21x1_ASAP7_75t_SL g1019 ( 
.A1(n_847),
.A2(n_853),
.B(n_878),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_809),
.Y(n_1020)
);

O2A1O1Ixp5_ASAP7_75t_L g1021 ( 
.A1(n_800),
.A2(n_918),
.B(n_831),
.C(n_814),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_861),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_790),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_808),
.A2(n_840),
.B(n_836),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_782),
.A2(n_784),
.B(n_815),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_837),
.B(n_892),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_836),
.A2(n_854),
.B(n_844),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_861),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_878),
.B(n_925),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_844),
.A2(n_884),
.B(n_899),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_883),
.A2(n_962),
.B1(n_940),
.B2(n_850),
.Y(n_1031)
);

AO31x2_ASAP7_75t_L g1032 ( 
.A1(n_835),
.A2(n_822),
.A3(n_852),
.B(n_906),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_802),
.A2(n_848),
.B(n_822),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_807),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_883),
.B(n_830),
.Y(n_1035)
);

BUFx4f_ASAP7_75t_L g1036 ( 
.A(n_882),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_802),
.A2(n_962),
.B(n_852),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_883),
.B(n_789),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_921),
.A2(n_889),
.B(n_835),
.Y(n_1039)
);

AO31x2_ASAP7_75t_L g1040 ( 
.A1(n_853),
.A2(n_910),
.A3(n_845),
.B(n_843),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_899),
.A2(n_851),
.B(n_793),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_817),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_886),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_833),
.A2(n_819),
.B(n_821),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_886),
.B(n_867),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_896),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_819),
.A2(n_930),
.B(n_785),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_917),
.B(n_912),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_834),
.A2(n_789),
.B(n_960),
.C(n_781),
.Y(n_1049)
);

INVx8_ASAP7_75t_L g1050 ( 
.A(n_883),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_SL g1051 ( 
.A1(n_859),
.A2(n_927),
.B(n_875),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_885),
.B(n_785),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_829),
.A2(n_942),
.B(n_937),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_829),
.A2(n_942),
.B(n_937),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_907),
.B(n_812),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_803),
.A2(n_903),
.B(n_909),
.C(n_896),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_885),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_930),
.A2(n_963),
.B(n_864),
.Y(n_1058)
);

INVx5_ASAP7_75t_L g1059 ( 
.A(n_896),
.Y(n_1059)
);

AOI21x1_ASAP7_75t_SL g1060 ( 
.A1(n_963),
.A2(n_919),
.B(n_916),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_963),
.A2(n_919),
.B(n_916),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_963),
.B(n_916),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_816),
.B(n_924),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_818),
.B(n_926),
.Y(n_1064)
);

BUFx12f_ASAP7_75t_L g1065 ( 
.A(n_816),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_872),
.A2(n_552),
.B(n_544),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_926),
.B(n_955),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_849),
.A2(n_873),
.B(n_922),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_872),
.A2(n_552),
.B(n_544),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_926),
.B(n_955),
.Y(n_1070)
);

O2A1O1Ixp5_ASAP7_75t_L g1071 ( 
.A1(n_799),
.A2(n_964),
.B(n_931),
.C(n_938),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_849),
.A2(n_873),
.B(n_922),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_926),
.B(n_955),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_804),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_SL g1075 ( 
.A1(n_879),
.A2(n_915),
.B(n_910),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_931),
.A2(n_938),
.B(n_935),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_849),
.A2(n_873),
.B(n_922),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_849),
.A2(n_873),
.B(n_922),
.Y(n_1078)
);

AO31x2_ASAP7_75t_L g1079 ( 
.A1(n_939),
.A2(n_946),
.A3(n_876),
.B(n_866),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_849),
.A2(n_873),
.B(n_922),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_804),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_787),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_872),
.A2(n_552),
.B(n_544),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_872),
.A2(n_552),
.B(n_544),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_872),
.A2(n_552),
.B(n_544),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_931),
.A2(n_938),
.B(n_935),
.C(n_926),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_804),
.Y(n_1087)
);

AO31x2_ASAP7_75t_L g1088 ( 
.A1(n_939),
.A2(n_946),
.A3(n_876),
.B(n_866),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_809),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_886),
.B(n_912),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_957),
.B(n_961),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_849),
.A2(n_873),
.B(n_922),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_926),
.B(n_955),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_931),
.A2(n_935),
.B1(n_938),
.B2(n_926),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_931),
.A2(n_938),
.B(n_935),
.C(n_926),
.Y(n_1095)
);

AOI21x1_ASAP7_75t_L g1096 ( 
.A1(n_831),
.A2(n_846),
.B(n_841),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_926),
.B(n_955),
.Y(n_1097)
);

AOI21xp33_ASAP7_75t_L g1098 ( 
.A1(n_926),
.A2(n_955),
.B(n_799),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_788),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_849),
.A2(n_873),
.B(n_922),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_809),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_787),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_788),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_886),
.B(n_912),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_931),
.A2(n_938),
.B(n_935),
.C(n_926),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_787),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_872),
.A2(n_552),
.B(n_544),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_861),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_809),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_788),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_849),
.A2(n_873),
.B(n_922),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_788),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_926),
.B(n_955),
.Y(n_1113)
);

AOI21x1_ASAP7_75t_L g1114 ( 
.A1(n_831),
.A2(n_846),
.B(n_841),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_872),
.A2(n_552),
.B(n_544),
.Y(n_1115)
);

INVxp67_ASAP7_75t_SL g1116 ( 
.A(n_809),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_788),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_926),
.B(n_955),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_980),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_973),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_1074),
.Y(n_1121)
);

AOI21xp33_ASAP7_75t_SL g1122 ( 
.A1(n_1113),
.A2(n_1067),
.B(n_969),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_1074),
.Y(n_1123)
);

NOR2xp67_ASAP7_75t_L g1124 ( 
.A(n_1015),
.B(n_1064),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1070),
.B(n_1073),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_994),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_1065),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1071),
.A2(n_1095),
.B(n_1086),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1093),
.B(n_1097),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_SL g1130 ( 
.A(n_1022),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1118),
.B(n_971),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_1090),
.B(n_1104),
.Y(n_1132)
);

BUFx4f_ASAP7_75t_L g1133 ( 
.A(n_993),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_985),
.B(n_982),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_974),
.A2(n_976),
.B(n_987),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1090),
.B(n_1104),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_992),
.A2(n_1069),
.B(n_1066),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1083),
.A2(n_1084),
.B(n_1085),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_1028),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1099),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_1010),
.B(n_1045),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1081),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1098),
.A2(n_1105),
.B(n_1094),
.C(n_975),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_1081),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_973),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1107),
.A2(n_1115),
.B(n_983),
.Y(n_1146)
);

AO21x1_ASAP7_75t_L g1147 ( 
.A1(n_970),
.A2(n_1076),
.B(n_1025),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_970),
.A2(n_1076),
.B(n_984),
.C(n_1025),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1004),
.A2(n_1006),
.B(n_1039),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1091),
.A2(n_986),
.B1(n_1014),
.B2(n_1055),
.Y(n_1150)
);

OA21x2_ASAP7_75t_L g1151 ( 
.A1(n_995),
.A2(n_1030),
.B(n_978),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1103),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1009),
.B(n_988),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_1108),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1087),
.B(n_999),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_1036),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_SL g1157 ( 
.A1(n_1037),
.A2(n_995),
.B(n_1033),
.C(n_1012),
.Y(n_1157)
);

INVx1_ASAP7_75t_SL g1158 ( 
.A(n_1087),
.Y(n_1158)
);

BUFx10_ASAP7_75t_L g1159 ( 
.A(n_1043),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_1026),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_990),
.B(n_991),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1005),
.B(n_1043),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1043),
.B(n_1013),
.Y(n_1163)
);

INVx1_ASAP7_75t_SL g1164 ( 
.A(n_996),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1110),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1112),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1117),
.Y(n_1167)
);

BUFx4_ASAP7_75t_SL g1168 ( 
.A(n_1048),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1029),
.B(n_997),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_1008),
.B(n_1023),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1048),
.B(n_1061),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_973),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1014),
.A2(n_977),
.B(n_1021),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_SL g1174 ( 
.A1(n_1037),
.A2(n_1033),
.B(n_1003),
.C(n_1017),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_977),
.A2(n_1031),
.B(n_1001),
.C(n_1049),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1034),
.B(n_1082),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_968),
.A2(n_1078),
.B(n_1068),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1042),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1007),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1102),
.B(n_1106),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_1050),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_981),
.A2(n_1031),
.B1(n_1050),
.B2(n_1038),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_1007),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1057),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1050),
.A2(n_1075),
.B1(n_1048),
.B2(n_1058),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_1036),
.Y(n_1186)
);

BUFx12f_ASAP7_75t_L g1187 ( 
.A(n_1063),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_1007),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1056),
.A2(n_1035),
.B(n_1058),
.C(n_1061),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_989),
.A2(n_1000),
.B(n_1002),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_981),
.B(n_1011),
.Y(n_1191)
);

INVxp33_ASAP7_75t_L g1192 ( 
.A(n_1046),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1011),
.B(n_1079),
.Y(n_1193)
);

AND2x4_ASAP7_75t_SL g1194 ( 
.A(n_1046),
.B(n_1020),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_1020),
.B(n_1089),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_R g1196 ( 
.A(n_1059),
.B(n_1101),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1044),
.A2(n_1051),
.B(n_1062),
.C(n_1052),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1059),
.Y(n_1198)
);

AOI21xp33_ASAP7_75t_L g1199 ( 
.A1(n_1018),
.A2(n_1016),
.B(n_1027),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1024),
.A2(n_1041),
.B(n_1114),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1059),
.B(n_1089),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1101),
.B(n_1109),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1116),
.B(n_1096),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1040),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1040),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_979),
.B(n_1079),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1000),
.A2(n_1054),
.B1(n_1053),
.B2(n_1047),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_972),
.A2(n_1072),
.B(n_1100),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1040),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_979),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1077),
.A2(n_1111),
.B(n_1092),
.C(n_1080),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1011),
.B(n_979),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1060),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1079),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1088),
.B(n_1032),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1019),
.B(n_1088),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1032),
.A2(n_1113),
.B1(n_954),
.B2(n_948),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1088),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1032),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_998),
.Y(n_1220)
);

NAND2x1p5_ASAP7_75t_L g1221 ( 
.A(n_998),
.B(n_1059),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_998),
.A2(n_974),
.B(n_976),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1050),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_969),
.B(n_1067),
.Y(n_1224)
);

OR2x6_ASAP7_75t_L g1225 ( 
.A(n_1050),
.B(n_861),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1113),
.B(n_969),
.Y(n_1226)
);

OAI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_969),
.A2(n_928),
.B1(n_943),
.B2(n_934),
.Y(n_1227)
);

OR2x6_ASAP7_75t_L g1228 ( 
.A(n_1050),
.B(n_861),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_974),
.A2(n_976),
.B(n_799),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1113),
.A2(n_955),
.B(n_926),
.C(n_935),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1113),
.A2(n_954),
.B1(n_948),
.B2(n_969),
.Y(n_1231)
);

INVx1_ASAP7_75t_SL g1232 ( 
.A(n_1074),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1090),
.B(n_1104),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1113),
.B(n_926),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1113),
.B(n_969),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_973),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1090),
.B(n_1104),
.Y(n_1237)
);

AOI221x1_ASAP7_75t_L g1238 ( 
.A1(n_1094),
.A2(n_964),
.B1(n_938),
.B2(n_935),
.C(n_931),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1065),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1113),
.B(n_969),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1074),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_980),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_1074),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1113),
.B(n_969),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_980),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1113),
.B(n_969),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1113),
.A2(n_954),
.B1(n_948),
.B2(n_969),
.Y(n_1247)
);

NAND2x1p5_ASAP7_75t_L g1248 ( 
.A(n_1059),
.B(n_859),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_980),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_1015),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1090),
.B(n_1104),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1113),
.B(n_969),
.Y(n_1252)
);

INVx2_ASAP7_75t_SL g1253 ( 
.A(n_1022),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1113),
.B(n_1091),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1022),
.Y(n_1255)
);

OR2x6_ASAP7_75t_L g1256 ( 
.A(n_1050),
.B(n_861),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_980),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_1015),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1113),
.B(n_969),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_974),
.A2(n_976),
.B(n_799),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1119),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1234),
.A2(n_1247),
.B1(n_1231),
.B2(n_1217),
.Y(n_1262)
);

INVx6_ASAP7_75t_L g1263 ( 
.A(n_1225),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1225),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1231),
.A2(n_1247),
.B1(n_1147),
.B2(n_1217),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1121),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1126),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1225),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1228),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1227),
.A2(n_1246),
.B1(n_1259),
.B2(n_1235),
.Y(n_1270)
);

BUFx12f_ASAP7_75t_L g1271 ( 
.A(n_1127),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1181),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1226),
.A2(n_1244),
.B1(n_1259),
.B2(n_1252),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1242),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_SL g1275 ( 
.A1(n_1226),
.A2(n_1252),
.B1(n_1246),
.B2(n_1244),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1249),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1230),
.A2(n_1235),
.B1(n_1240),
.B2(n_1224),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1240),
.A2(n_1128),
.B1(n_1133),
.B2(n_1125),
.Y(n_1278)
);

INVx6_ASAP7_75t_L g1279 ( 
.A(n_1228),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1140),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1169),
.B(n_1134),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1128),
.A2(n_1133),
.B1(n_1129),
.B2(n_1125),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_SL g1283 ( 
.A1(n_1189),
.A2(n_1143),
.B(n_1197),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1123),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1155),
.Y(n_1285)
);

AO21x1_ASAP7_75t_L g1286 ( 
.A1(n_1149),
.A2(n_1216),
.B(n_1173),
.Y(n_1286)
);

AO21x1_ASAP7_75t_SL g1287 ( 
.A1(n_1193),
.A2(n_1212),
.B(n_1191),
.Y(n_1287)
);

AO21x2_ASAP7_75t_L g1288 ( 
.A1(n_1138),
.A2(n_1137),
.B(n_1208),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_SL g1289 ( 
.A1(n_1210),
.A2(n_1173),
.B(n_1185),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1152),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1129),
.A2(n_1131),
.B1(n_1161),
.B2(n_1150),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1165),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1166),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1171),
.B(n_1181),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1167),
.Y(n_1295)
);

BUFx12f_ASAP7_75t_L g1296 ( 
.A(n_1239),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1177),
.A2(n_1200),
.B(n_1190),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1254),
.A2(n_1141),
.B1(n_1131),
.B2(n_1134),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1142),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1144),
.Y(n_1300)
);

AO21x2_ASAP7_75t_L g1301 ( 
.A1(n_1135),
.A2(n_1260),
.B(n_1229),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1156),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1245),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1161),
.B(n_1148),
.Y(n_1304)
);

OAI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1238),
.A2(n_1122),
.B1(n_1164),
.B2(n_1232),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1141),
.A2(n_1182),
.B1(n_1220),
.B2(n_1160),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1257),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1206),
.B(n_1171),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1191),
.B(n_1215),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_1198),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1228),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1158),
.A2(n_1232),
.B1(n_1243),
.B2(n_1256),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1178),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_R g1314 ( 
.A(n_1250),
.B(n_1258),
.Y(n_1314)
);

INVx5_ASAP7_75t_L g1315 ( 
.A(n_1223),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_1164),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1170),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1158),
.A2(n_1243),
.B1(n_1256),
.B2(n_1241),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1256),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1184),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1182),
.A2(n_1153),
.B1(n_1162),
.B2(n_1237),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1163),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1218),
.A2(n_1175),
.B1(n_1237),
.B2(n_1132),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1176),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1180),
.Y(n_1325)
);

BUFx10_ASAP7_75t_L g1326 ( 
.A(n_1130),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1172),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1195),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1203),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1193),
.B(n_1212),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1202),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1202),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1219),
.B(n_1214),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1198),
.Y(n_1334)
);

INVxp33_ASAP7_75t_L g1335 ( 
.A(n_1132),
.Y(n_1335)
);

BUFx12f_ASAP7_75t_L g1336 ( 
.A(n_1187),
.Y(n_1336)
);

NAND2x1p5_ASAP7_75t_L g1337 ( 
.A(n_1219),
.B(n_1151),
.Y(n_1337)
);

AO21x1_ASAP7_75t_SL g1338 ( 
.A1(n_1204),
.A2(n_1200),
.B(n_1207),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1222),
.A2(n_1146),
.B(n_1199),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1157),
.A2(n_1174),
.B(n_1199),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1221),
.B(n_1251),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1186),
.Y(n_1342)
);

BUFx12f_ASAP7_75t_L g1343 ( 
.A(n_1159),
.Y(n_1343)
);

OA21x2_ASAP7_75t_L g1344 ( 
.A1(n_1211),
.A2(n_1209),
.B(n_1205),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1151),
.Y(n_1345)
);

INVx11_ASAP7_75t_L g1346 ( 
.A(n_1168),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1136),
.B(n_1233),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1248),
.Y(n_1348)
);

NAND2x1p5_ASAP7_75t_L g1349 ( 
.A(n_1213),
.B(n_1198),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1136),
.B(n_1251),
.Y(n_1350)
);

BUFx12f_ASAP7_75t_L g1351 ( 
.A(n_1154),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1201),
.Y(n_1352)
);

NAND2x1p5_ASAP7_75t_L g1353 ( 
.A(n_1201),
.B(n_1233),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1124),
.A2(n_1130),
.B1(n_1179),
.B2(n_1192),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1196),
.A2(n_1194),
.B(n_1188),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1120),
.Y(n_1356)
);

NAND2xp33_ASAP7_75t_SL g1357 ( 
.A(n_1120),
.B(n_1145),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1120),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1139),
.A2(n_1255),
.B1(n_1183),
.B2(n_1236),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1253),
.A2(n_1145),
.B1(n_1183),
.B2(n_1236),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1145),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1183),
.B(n_1236),
.Y(n_1362)
);

AOI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1208),
.A2(n_1149),
.B(n_987),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1156),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1234),
.A2(n_926),
.B1(n_955),
.B2(n_1113),
.Y(n_1365)
);

INVx4_ASAP7_75t_L g1366 ( 
.A(n_1198),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1119),
.Y(n_1367)
);

BUFx12f_ASAP7_75t_L g1368 ( 
.A(n_1127),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1234),
.A2(n_926),
.B1(n_955),
.B2(n_949),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1119),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1181),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1177),
.A2(n_1208),
.B(n_1016),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1234),
.A2(n_926),
.B1(n_955),
.B2(n_1113),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1121),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1234),
.A2(n_926),
.B1(n_955),
.B2(n_1113),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1234),
.A2(n_926),
.B1(n_955),
.B2(n_1113),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1229),
.A2(n_1260),
.B(n_974),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1234),
.A2(n_926),
.B1(n_955),
.B2(n_1113),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1119),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_1155),
.Y(n_1380)
);

BUFx2_ASAP7_75t_SL g1381 ( 
.A(n_1130),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1119),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1308),
.B(n_1281),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1369),
.A2(n_1373),
.B(n_1365),
.Y(n_1384)
);

AO21x2_ASAP7_75t_L g1385 ( 
.A1(n_1377),
.A2(n_1340),
.B(n_1283),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1308),
.B(n_1281),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1375),
.B(n_1378),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1304),
.B(n_1262),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1345),
.Y(n_1389)
);

CKINVDCx6p67_ASAP7_75t_R g1390 ( 
.A(n_1336),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1309),
.B(n_1330),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1345),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1338),
.Y(n_1393)
);

AO21x2_ASAP7_75t_L g1394 ( 
.A1(n_1363),
.A2(n_1289),
.B(n_1286),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1333),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1304),
.B(n_1291),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1333),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1265),
.B(n_1309),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1287),
.B(n_1329),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1337),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_1374),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1270),
.B(n_1273),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1287),
.B(n_1330),
.Y(n_1403)
);

INVx4_ASAP7_75t_L g1404 ( 
.A(n_1315),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1337),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1372),
.A2(n_1297),
.B(n_1337),
.Y(n_1406)
);

OAI21xp33_ASAP7_75t_L g1407 ( 
.A1(n_1376),
.A2(n_1275),
.B(n_1277),
.Y(n_1407)
);

OR2x6_ASAP7_75t_L g1408 ( 
.A(n_1297),
.B(n_1286),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1344),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1344),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1288),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1374),
.Y(n_1412)
);

INVxp67_ASAP7_75t_SL g1413 ( 
.A(n_1292),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1282),
.B(n_1278),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1317),
.B(n_1298),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1314),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1372),
.A2(n_1306),
.B(n_1321),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1305),
.B(n_1328),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1266),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1301),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1280),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1290),
.B(n_1293),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1339),
.A2(n_1355),
.B(n_1323),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1284),
.Y(n_1424)
);

AO21x2_ASAP7_75t_L g1425 ( 
.A1(n_1320),
.A2(n_1307),
.B(n_1303),
.Y(n_1425)
);

AO21x2_ASAP7_75t_L g1426 ( 
.A1(n_1295),
.A2(n_1313),
.B(n_1382),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1341),
.B(n_1274),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1299),
.Y(n_1428)
);

AO21x2_ASAP7_75t_L g1429 ( 
.A1(n_1261),
.A2(n_1370),
.B(n_1379),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1300),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1355),
.A2(n_1272),
.B(n_1371),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1276),
.B(n_1322),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1267),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1367),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1324),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1325),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1341),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1294),
.B(n_1338),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1285),
.B(n_1380),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1335),
.B(n_1350),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_1327),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_1364),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1318),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1272),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1371),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1348),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1347),
.B(n_1332),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1347),
.B(n_1331),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1403),
.B(n_1389),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_L g1450 ( 
.A(n_1387),
.B(n_1312),
.C(n_1354),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1403),
.B(n_1361),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1384),
.A2(n_1335),
.B(n_1360),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1389),
.B(n_1361),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1391),
.B(n_1352),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1391),
.B(n_1396),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1409),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1408),
.B(n_1358),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1410),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1392),
.B(n_1352),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1409),
.Y(n_1460)
);

OAI221xp5_ASAP7_75t_L g1461 ( 
.A1(n_1407),
.A2(n_1384),
.B1(n_1414),
.B2(n_1402),
.C(n_1396),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1394),
.B(n_1353),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1431),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1394),
.B(n_1353),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1408),
.B(n_1362),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1408),
.B(n_1349),
.Y(n_1466)
);

NOR2x1_ASAP7_75t_L g1467 ( 
.A(n_1429),
.B(n_1385),
.Y(n_1467)
);

INVx5_ASAP7_75t_L g1468 ( 
.A(n_1408),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1400),
.B(n_1319),
.Y(n_1469)
);

AOI211xp5_ASAP7_75t_L g1470 ( 
.A1(n_1407),
.A2(n_1350),
.B(n_1264),
.C(n_1268),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1437),
.B(n_1385),
.Y(n_1471)
);

INVxp67_ASAP7_75t_SL g1472 ( 
.A(n_1413),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1408),
.B(n_1311),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1385),
.B(n_1356),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1408),
.B(n_1311),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1423),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1425),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1405),
.B(n_1399),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1414),
.A2(n_1263),
.B1(n_1279),
.B2(n_1316),
.Y(n_1479)
);

BUFx2_ASAP7_75t_L g1480 ( 
.A(n_1423),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1398),
.B(n_1310),
.Y(n_1481)
);

NAND3xp33_ASAP7_75t_L g1482 ( 
.A(n_1461),
.B(n_1443),
.C(n_1418),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1461),
.A2(n_1402),
.B1(n_1388),
.B2(n_1443),
.Y(n_1483)
);

NAND3xp33_ASAP7_75t_L g1484 ( 
.A(n_1450),
.B(n_1418),
.C(n_1415),
.Y(n_1484)
);

OAI221xp5_ASAP7_75t_SL g1485 ( 
.A1(n_1450),
.A2(n_1388),
.B1(n_1415),
.B2(n_1398),
.C(n_1359),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1449),
.B(n_1395),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1452),
.A2(n_1470),
.B(n_1479),
.Y(n_1487)
);

AOI221x1_ASAP7_75t_SL g1488 ( 
.A1(n_1470),
.A2(n_1436),
.B1(n_1435),
.B2(n_1422),
.C(n_1421),
.Y(n_1488)
);

OAI221xp5_ASAP7_75t_L g1489 ( 
.A1(n_1479),
.A2(n_1452),
.B1(n_1440),
.B2(n_1430),
.C(n_1401),
.Y(n_1489)
);

OAI221xp5_ASAP7_75t_L g1490 ( 
.A1(n_1473),
.A2(n_1430),
.B1(n_1401),
.B2(n_1419),
.C(n_1424),
.Y(n_1490)
);

NAND3xp33_ASAP7_75t_L g1491 ( 
.A(n_1467),
.B(n_1399),
.C(n_1428),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1481),
.A2(n_1263),
.B1(n_1279),
.B2(n_1393),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1455),
.B(n_1393),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1449),
.B(n_1478),
.Y(n_1494)
);

OAI221xp5_ASAP7_75t_SL g1495 ( 
.A1(n_1473),
.A2(n_1390),
.B1(n_1439),
.B2(n_1424),
.C(n_1419),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_SL g1496 ( 
.A1(n_1473),
.A2(n_1438),
.B(n_1393),
.Y(n_1496)
);

OAI221xp5_ASAP7_75t_L g1497 ( 
.A1(n_1475),
.A2(n_1412),
.B1(n_1441),
.B2(n_1316),
.C(n_1269),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1454),
.A2(n_1279),
.B1(n_1393),
.B2(n_1390),
.Y(n_1498)
);

NAND3xp33_ASAP7_75t_L g1499 ( 
.A(n_1467),
.B(n_1432),
.C(n_1446),
.Y(n_1499)
);

AOI221xp5_ASAP7_75t_L g1500 ( 
.A1(n_1454),
.A2(n_1441),
.B1(n_1383),
.B2(n_1386),
.C(n_1435),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1469),
.A2(n_1439),
.B1(n_1417),
.B2(n_1447),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_L g1502 ( 
.A(n_1457),
.B(n_1432),
.C(n_1446),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1465),
.B(n_1397),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1451),
.B(n_1386),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1475),
.A2(n_1393),
.B1(n_1390),
.B2(n_1442),
.Y(n_1505)
);

AOI221xp5_ASAP7_75t_L g1506 ( 
.A1(n_1471),
.A2(n_1436),
.B1(n_1422),
.B2(n_1434),
.C(n_1433),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1478),
.B(n_1397),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1469),
.B(n_1427),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1469),
.B(n_1426),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1478),
.B(n_1405),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1469),
.B(n_1426),
.Y(n_1511)
);

NOR3xp33_ASAP7_75t_L g1512 ( 
.A(n_1457),
.B(n_1357),
.C(n_1366),
.Y(n_1512)
);

OA211x2_ASAP7_75t_L g1513 ( 
.A1(n_1468),
.A2(n_1404),
.B(n_1423),
.C(n_1431),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1453),
.B(n_1426),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1453),
.B(n_1425),
.Y(n_1515)
);

NOR3xp33_ASAP7_75t_L g1516 ( 
.A(n_1457),
.B(n_1366),
.C(n_1420),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1453),
.B(n_1425),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1476),
.A2(n_1406),
.B(n_1411),
.Y(n_1518)
);

NAND3xp33_ASAP7_75t_L g1519 ( 
.A(n_1474),
.B(n_1445),
.C(n_1444),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1459),
.B(n_1425),
.Y(n_1520)
);

NAND3xp33_ASAP7_75t_L g1521 ( 
.A(n_1474),
.B(n_1445),
.C(n_1444),
.Y(n_1521)
);

OAI221xp5_ASAP7_75t_SL g1522 ( 
.A1(n_1466),
.A2(n_1448),
.B1(n_1433),
.B2(n_1434),
.C(n_1421),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1515),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1494),
.B(n_1468),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1509),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1511),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1494),
.B(n_1468),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1501),
.B(n_1510),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1487),
.B(n_1468),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1503),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1517),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1501),
.B(n_1468),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1520),
.B(n_1456),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1514),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1506),
.B(n_1456),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1516),
.B(n_1468),
.Y(n_1536)
);

A2O1A1Ixp33_ASAP7_75t_L g1537 ( 
.A1(n_1488),
.A2(n_1468),
.B(n_1472),
.C(n_1464),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1519),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1502),
.B(n_1460),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1521),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1486),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1499),
.B(n_1460),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1512),
.B(n_1468),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1518),
.B(n_1471),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1486),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1518),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1513),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1507),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1508),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1504),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1493),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1491),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1496),
.B(n_1476),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1522),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1492),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1505),
.B(n_1480),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1538),
.B(n_1500),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1538),
.B(n_1477),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1524),
.B(n_1527),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1541),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1538),
.B(n_1477),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1541),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1541),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1546),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1546),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1545),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1540),
.B(n_1490),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1524),
.B(n_1480),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1545),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1545),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1546),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1524),
.B(n_1480),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1524),
.B(n_1463),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1548),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1540),
.B(n_1458),
.Y(n_1575)
);

INVxp67_ASAP7_75t_SL g1576 ( 
.A(n_1542),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1539),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1546),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1540),
.B(n_1533),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1555),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1527),
.B(n_1462),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1544),
.Y(n_1582)
);

NOR3xp33_ASAP7_75t_L g1583 ( 
.A(n_1529),
.B(n_1484),
.C(n_1482),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1544),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1533),
.B(n_1465),
.Y(n_1585)
);

INVxp67_ASAP7_75t_L g1586 ( 
.A(n_1554),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1560),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1560),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1562),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1580),
.B(n_1528),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1580),
.B(n_1528),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1567),
.B(n_1530),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1567),
.B(n_1530),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1579),
.B(n_1549),
.Y(n_1594)
);

OAI221xp5_ASAP7_75t_L g1595 ( 
.A1(n_1583),
.A2(n_1483),
.B1(n_1485),
.B2(n_1529),
.C(n_1554),
.Y(n_1595)
);

NAND2xp33_ASAP7_75t_R g1596 ( 
.A(n_1557),
.B(n_1416),
.Y(n_1596)
);

A2O1A1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1583),
.A2(n_1554),
.B(n_1537),
.C(n_1552),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1562),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1559),
.B(n_1543),
.Y(n_1599)
);

NOR2xp67_ASAP7_75t_L g1600 ( 
.A(n_1586),
.B(n_1551),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1563),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1579),
.B(n_1549),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1563),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1559),
.B(n_1543),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1566),
.Y(n_1605)
);

INVx5_ASAP7_75t_L g1606 ( 
.A(n_1564),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1557),
.B(n_1552),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1566),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1569),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_SL g1610 ( 
.A(n_1586),
.B(n_1495),
.Y(n_1610)
);

AND3x2_ASAP7_75t_L g1611 ( 
.A(n_1576),
.B(n_1552),
.C(n_1547),
.Y(n_1611)
);

OAI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1576),
.A2(n_1537),
.B(n_1552),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1577),
.B(n_1523),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1559),
.B(n_1528),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1581),
.B(n_1550),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1577),
.B(n_1523),
.Y(n_1616)
);

NOR2xp67_ASAP7_75t_L g1617 ( 
.A(n_1575),
.B(n_1551),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1558),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1569),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1581),
.B(n_1550),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1570),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1570),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1575),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1558),
.B(n_1523),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1585),
.B(n_1555),
.Y(n_1625)
);

NOR2x1_ASAP7_75t_L g1626 ( 
.A(n_1561),
.B(n_1547),
.Y(n_1626)
);

INVxp67_ASAP7_75t_L g1627 ( 
.A(n_1561),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1585),
.B(n_1549),
.Y(n_1628)
);

CKINVDCx16_ASAP7_75t_R g1629 ( 
.A(n_1581),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1629),
.B(n_1568),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1590),
.B(n_1568),
.Y(n_1631)
);

NAND3xp33_ASAP7_75t_L g1632 ( 
.A(n_1607),
.B(n_1483),
.C(n_1547),
.Y(n_1632)
);

BUFx4f_ASAP7_75t_SL g1633 ( 
.A(n_1592),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1591),
.B(n_1568),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1607),
.B(n_1610),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1599),
.B(n_1543),
.Y(n_1636)
);

INVx1_ASAP7_75t_SL g1637 ( 
.A(n_1593),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1587),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1588),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1589),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1601),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1611),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1614),
.B(n_1572),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1623),
.B(n_1594),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1625),
.B(n_1550),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1599),
.B(n_1572),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1603),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1604),
.B(n_1543),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1602),
.B(n_1574),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1625),
.B(n_1531),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1597),
.B(n_1617),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1606),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1595),
.A2(n_1612),
.B1(n_1604),
.B2(n_1543),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1613),
.B(n_1574),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1595),
.B(n_1531),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1600),
.B(n_1606),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1611),
.B(n_1531),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1605),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_1596),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1618),
.B(n_1534),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1608),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1618),
.B(n_1534),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1615),
.B(n_1572),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1606),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1609),
.Y(n_1665)
);

INVx3_ASAP7_75t_L g1666 ( 
.A(n_1656),
.Y(n_1666)
);

AO22x1_ASAP7_75t_L g1667 ( 
.A1(n_1642),
.A2(n_1626),
.B1(n_1606),
.B2(n_1547),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1664),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1637),
.B(n_1620),
.Y(n_1669)
);

AOI21xp33_ASAP7_75t_SL g1670 ( 
.A1(n_1651),
.A2(n_1302),
.B(n_1497),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1630),
.B(n_1573),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1638),
.Y(n_1672)
);

OAI22xp33_ASAP7_75t_SL g1673 ( 
.A1(n_1635),
.A2(n_1627),
.B1(n_1613),
.B2(n_1616),
.Y(n_1673)
);

AND4x1_ASAP7_75t_L g1674 ( 
.A(n_1635),
.B(n_1653),
.C(n_1632),
.D(n_1655),
.Y(n_1674)
);

OAI322xp33_ASAP7_75t_L g1675 ( 
.A1(n_1657),
.A2(n_1627),
.A3(n_1535),
.B1(n_1616),
.B2(n_1624),
.C1(n_1622),
.C2(n_1619),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1633),
.B(n_1534),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1639),
.B(n_1624),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_SL g1678 ( 
.A(n_1659),
.B(n_1543),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1640),
.B(n_1598),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_1656),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1650),
.A2(n_1656),
.B(n_1660),
.Y(n_1681)
);

AOI222xp33_ASAP7_75t_L g1682 ( 
.A1(n_1641),
.A2(n_1535),
.B1(n_1489),
.B2(n_1532),
.C1(n_1556),
.C2(n_1542),
.Y(n_1682)
);

XNOR2xp5_ASAP7_75t_L g1683 ( 
.A(n_1630),
.B(n_1302),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1631),
.B(n_1526),
.Y(n_1684)
);

NAND4xp25_ASAP7_75t_SL g1685 ( 
.A(n_1646),
.B(n_1532),
.C(n_1553),
.D(n_1556),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_SL g1686 ( 
.A1(n_1636),
.A2(n_1648),
.B1(n_1532),
.B2(n_1631),
.Y(n_1686)
);

XNOR2x1_ASAP7_75t_L g1687 ( 
.A(n_1636),
.B(n_1381),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1645),
.B(n_1628),
.Y(n_1688)
);

AOI21xp33_ASAP7_75t_L g1689 ( 
.A1(n_1652),
.A2(n_1621),
.B(n_1539),
.Y(n_1689)
);

OAI21xp5_ASAP7_75t_SL g1690 ( 
.A1(n_1636),
.A2(n_1556),
.B(n_1536),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1666),
.B(n_1646),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1674),
.B(n_1271),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1666),
.B(n_1634),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1680),
.B(n_1669),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1679),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1680),
.B(n_1634),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1688),
.B(n_1644),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1679),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1672),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1668),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1681),
.B(n_1647),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1677),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1671),
.B(n_1648),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1667),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1677),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1686),
.B(n_1648),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1683),
.B(n_1658),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1676),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1682),
.A2(n_1536),
.B1(n_1661),
.B2(n_1665),
.Y(n_1709)
);

NAND4xp25_ASAP7_75t_L g1710 ( 
.A(n_1692),
.B(n_1678),
.C(n_1682),
.D(n_1689),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1697),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1694),
.B(n_1673),
.Y(n_1712)
);

NOR3xp33_ASAP7_75t_L g1713 ( 
.A(n_1692),
.B(n_1675),
.C(n_1670),
.Y(n_1713)
);

O2A1O1Ixp33_ASAP7_75t_L g1714 ( 
.A1(n_1701),
.A2(n_1689),
.B(n_1652),
.C(n_1664),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1694),
.B(n_1687),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1704),
.A2(n_1685),
.B(n_1662),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1706),
.A2(n_1684),
.B1(n_1644),
.B2(n_1643),
.Y(n_1717)
);

OAI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1709),
.A2(n_1690),
.B1(n_1664),
.B2(n_1584),
.Y(n_1718)
);

NAND4xp25_ASAP7_75t_L g1719 ( 
.A(n_1707),
.B(n_1643),
.C(n_1654),
.D(n_1663),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1691),
.A2(n_1536),
.B1(n_1556),
.B2(n_1553),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1712),
.A2(n_1704),
.B1(n_1693),
.B2(n_1708),
.Y(n_1721)
);

NAND4xp75_ASAP7_75t_L g1722 ( 
.A(n_1711),
.B(n_1700),
.C(n_1706),
.D(n_1696),
.Y(n_1722)
);

NOR3xp33_ASAP7_75t_L g1723 ( 
.A(n_1714),
.B(n_1698),
.C(n_1695),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1719),
.B(n_1697),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1715),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_SL g1726 ( 
.A(n_1713),
.B(n_1696),
.C(n_1691),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1720),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1717),
.Y(n_1728)
);

BUFx2_ASAP7_75t_L g1729 ( 
.A(n_1710),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1718),
.B(n_1703),
.Y(n_1730)
);

NOR3xp33_ASAP7_75t_L g1731 ( 
.A(n_1729),
.B(n_1721),
.C(n_1725),
.Y(n_1731)
);

NAND3xp33_ASAP7_75t_L g1732 ( 
.A(n_1723),
.B(n_1716),
.C(n_1699),
.Y(n_1732)
);

INVx3_ASAP7_75t_L g1733 ( 
.A(n_1722),
.Y(n_1733)
);

NAND3xp33_ASAP7_75t_L g1734 ( 
.A(n_1721),
.B(n_1705),
.C(n_1702),
.Y(n_1734)
);

NOR2xp67_ASAP7_75t_SL g1735 ( 
.A(n_1724),
.B(n_1271),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1733),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1731),
.A2(n_1726),
.B1(n_1730),
.B2(n_1728),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1732),
.A2(n_1727),
.B1(n_1703),
.B2(n_1663),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1734),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1735),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1731),
.A2(n_1342),
.B1(n_1364),
.B2(n_1553),
.Y(n_1741)
);

NOR3x2_ASAP7_75t_L g1742 ( 
.A(n_1737),
.B(n_1368),
.C(n_1296),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1738),
.B(n_1649),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1736),
.Y(n_1744)
);

OAI31xp33_ASAP7_75t_L g1745 ( 
.A1(n_1739),
.A2(n_1654),
.A3(n_1649),
.B(n_1334),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1741),
.B(n_1525),
.Y(n_1746)
);

NOR2x1_ASAP7_75t_L g1747 ( 
.A(n_1744),
.B(n_1740),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1743),
.B(n_1296),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1746),
.Y(n_1749)
);

AOI22x1_ASAP7_75t_L g1750 ( 
.A1(n_1748),
.A2(n_1368),
.B1(n_1742),
.B2(n_1336),
.Y(n_1750)
);

OAI211xp5_ASAP7_75t_SL g1751 ( 
.A1(n_1750),
.A2(n_1747),
.B(n_1749),
.C(n_1745),
.Y(n_1751)
);

AOI221x1_ASAP7_75t_L g1752 ( 
.A1(n_1751),
.A2(n_1564),
.B1(n_1565),
.B2(n_1578),
.C(n_1571),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1751),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1753),
.Y(n_1754)
);

AOI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1752),
.A2(n_1564),
.B1(n_1565),
.B2(n_1571),
.C(n_1578),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1754),
.A2(n_1326),
.B(n_1565),
.Y(n_1756)
);

AOI221x1_ASAP7_75t_L g1757 ( 
.A1(n_1755),
.A2(n_1571),
.B1(n_1578),
.B2(n_1326),
.C(n_1582),
.Y(n_1757)
);

OAI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1756),
.A2(n_1326),
.B(n_1346),
.Y(n_1758)
);

AOI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1758),
.A2(n_1757),
.B1(n_1351),
.B2(n_1343),
.Y(n_1759)
);

OAI221xp5_ASAP7_75t_R g1760 ( 
.A1(n_1759),
.A2(n_1346),
.B1(n_1351),
.B2(n_1343),
.C(n_1582),
.Y(n_1760)
);

AOI211xp5_ASAP7_75t_L g1761 ( 
.A1(n_1760),
.A2(n_1334),
.B(n_1310),
.C(n_1498),
.Y(n_1761)
);


endmodule