module fake_jpeg_24561_n_177 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_13),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_44),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_42),
.Y(n_51)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_19),
.B1(n_46),
.B2(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_46),
.Y(n_57)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_17),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_17),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_40),
.B(n_26),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_63),
.B(n_20),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_24),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_24),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_15),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_69),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_27),
.B1(n_18),
.B2(n_32),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_80),
.B1(n_83),
.B2(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_82),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_41),
.B1(n_45),
.B2(n_31),
.Y(n_80)
);

MAJx2_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_44),
.C(n_43),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_6),
.B(n_58),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_31),
.B1(n_25),
.B2(n_23),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_23),
.B1(n_15),
.B2(n_25),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_SL g87 ( 
.A(n_53),
.B(n_43),
.C(n_3),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_87),
.B(n_49),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_62),
.A2(n_1),
.B(n_4),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_88),
.Y(n_96)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_89),
.B(n_92),
.Y(n_112)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_98),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_56),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_58),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_105),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_5),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_103),
.C(n_75),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_6),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_58),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_106),
.B(n_114),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_105),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_78),
.A2(n_50),
.B1(n_55),
.B2(n_66),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_92),
.B1(n_93),
.B2(n_52),
.Y(n_128)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_91),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_55),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_60),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_112),
.Y(n_116)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_121),
.Y(n_135)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_120),
.B(n_122),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_95),
.C(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_89),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_111),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_88),
.B1(n_78),
.B2(n_75),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_60),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_127),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_128),
.A2(n_96),
.B(n_106),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_86),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_97),
.C(n_100),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_116),
.B1(n_102),
.B2(n_117),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_140),
.C(n_131),
.Y(n_145)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_137),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_103),
.C(n_102),
.Y(n_137)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_103),
.B(n_111),
.C(n_104),
.D(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_114),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_142),
.A2(n_144),
.B1(n_130),
.B2(n_94),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_152),
.Y(n_160)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_129),
.B(n_130),
.C(n_118),
.D(n_119),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_129),
.B(n_128),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_153),
.B(n_144),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_139),
.B1(n_135),
.B2(n_138),
.Y(n_157)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_65),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_90),
.C(n_94),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_156),
.Y(n_165)
);

BUFx24_ASAP7_75t_SL g156 ( 
.A(n_154),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_161),
.Y(n_163)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_166),
.Y(n_168)
);

FAx1_ASAP7_75t_SL g164 ( 
.A(n_160),
.B(n_145),
.CI(n_147),
.CON(n_164),
.SN(n_164)
);

OAI21x1_ASAP7_75t_SL g167 ( 
.A1(n_164),
.A2(n_143),
.B(n_158),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_149),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_167),
.A2(n_169),
.B(n_170),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_152),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_140),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_168),
.A2(n_163),
.B1(n_164),
.B2(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_164),
.A3(n_148),
.B1(n_93),
.B2(n_10),
.C1(n_11),
.C2(n_7),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_8),
.Y(n_174)
);

A2O1A1O1Ixp25_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_173),
.B(n_171),
.C(n_12),
.D(n_14),
.Y(n_176)
);

AOI221xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_175),
.B1(n_9),
.B2(n_14),
.C(n_8),
.Y(n_177)
);


endmodule