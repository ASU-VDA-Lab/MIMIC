module fake_jpeg_3599_n_615 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_615);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_615;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_4),
.B(n_3),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_18),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_59),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_60),
.Y(n_143)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_62),
.Y(n_151)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g187 ( 
.A(n_65),
.Y(n_187)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_67),
.Y(n_189)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_69),
.Y(n_217)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g175 ( 
.A(n_70),
.Y(n_175)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

BUFx12f_ASAP7_75t_SL g73 ( 
.A(n_39),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_73),
.B(n_80),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_74),
.Y(n_167)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_77),
.Y(n_176)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_36),
.B(n_11),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_37),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_82),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_83),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_84),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_36),
.B(n_11),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_91),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_47),
.Y(n_87)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_88),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_19),
.B(n_11),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g170 ( 
.A(n_92),
.Y(n_170)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_93),
.Y(n_199)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_94),
.Y(n_180)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_19),
.B(n_12),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_109),
.Y(n_149)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_97),
.Y(n_181)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx5_ASAP7_75t_SL g210 ( 
.A(n_98),
.Y(n_210)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_100),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_101),
.Y(n_204)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_102),
.Y(n_203)
);

INVx4_ASAP7_75t_SL g103 ( 
.A(n_53),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_103),
.Y(n_169)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_104),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_105),
.Y(n_211)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_41),
.Y(n_107)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_23),
.B(n_12),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_121),
.Y(n_147)
);

BUFx4f_ASAP7_75t_SL g109 ( 
.A(n_53),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_110),
.Y(n_205)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

INVx3_ASAP7_75t_SL g112 ( 
.A(n_22),
.Y(n_112)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_23),
.B(n_10),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_128),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_22),
.Y(n_118)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_29),
.Y(n_120)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_38),
.B(n_13),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_122),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_123),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_126),
.Y(n_208)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_56),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_54),
.B1(n_28),
.B2(n_32),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g244 ( 
.A1(n_131),
.A2(n_146),
.B1(n_156),
.B2(n_173),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_80),
.A2(n_54),
.B1(n_56),
.B2(n_38),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_137),
.A2(n_210),
.B1(n_170),
.B2(n_204),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_58),
.A2(n_54),
.B1(n_28),
.B2(n_24),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_139),
.A2(n_196),
.B1(n_116),
.B2(n_107),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_91),
.A2(n_42),
.B1(n_40),
.B2(n_48),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_145),
.A2(n_183),
.B1(n_193),
.B2(n_198),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_65),
.A2(n_60),
.B1(n_87),
.B2(n_81),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_65),
.A2(n_24),
.B1(n_32),
.B2(n_50),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_108),
.B(n_55),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_159),
.B(n_171),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_121),
.B(n_55),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_81),
.A2(n_57),
.B1(n_50),
.B2(n_49),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_109),
.B(n_49),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_174),
.B(n_188),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_67),
.A2(n_57),
.B1(n_48),
.B2(n_42),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_59),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_186),
.B(n_197),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_110),
.B(n_40),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_69),
.A2(n_30),
.B1(n_14),
.B2(n_3),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_72),
.A2(n_30),
.B1(n_1),
.B2(n_0),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_106),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_90),
.A2(n_30),
.B1(n_14),
.B2(n_3),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_0),
.B(n_1),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_110),
.B(n_14),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_201),
.B(n_202),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_82),
.B(n_14),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_112),
.B(n_15),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_206),
.B(n_212),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_93),
.B(n_15),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_123),
.B(n_15),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_213),
.B(n_220),
.Y(n_269)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_125),
.Y(n_215)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_74),
.A2(n_30),
.B1(n_9),
.B2(n_5),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_216),
.B(n_8),
.Y(n_259)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_84),
.Y(n_219)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_92),
.B(n_18),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_100),
.Y(n_221)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_101),
.B(n_9),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_222),
.B(n_170),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_172),
.Y(n_223)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_223),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_138),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_224),
.Y(n_341)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_162),
.Y(n_225)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_225),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_228),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_147),
.A2(n_124),
.B1(n_119),
.B2(n_117),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_229),
.A2(n_231),
.B1(n_233),
.B2(n_257),
.Y(n_314)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_151),
.Y(n_232)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_232),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_183),
.A2(n_98),
.B1(n_70),
.B2(n_0),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_161),
.Y(n_234)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_234),
.Y(n_303)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_150),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_235),
.Y(n_327)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_152),
.Y(n_236)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_236),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_211),
.A2(n_9),
.B1(n_17),
.B2(n_5),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_238),
.A2(n_243),
.B1(n_270),
.B2(n_281),
.Y(n_320)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_143),
.Y(n_239)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_239),
.Y(n_346)
);

A2O1A1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_134),
.A2(n_8),
.B(n_16),
.C(n_17),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_240),
.B(n_246),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_143),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_241),
.Y(n_325)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_160),
.Y(n_245)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_245),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_172),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_165),
.Y(n_247)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_247),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_187),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_248),
.B(n_287),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_146),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_249),
.Y(n_358)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_150),
.Y(n_250)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_250),
.Y(n_307)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_163),
.Y(n_251)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_251),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_138),
.Y(n_252)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_252),
.Y(n_329)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_253),
.Y(n_337)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_166),
.Y(n_254)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_254),
.Y(n_344)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_191),
.Y(n_255)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_255),
.Y(n_336)
);

OAI22xp33_ASAP7_75t_L g257 ( 
.A1(n_131),
.A2(n_8),
.B1(n_16),
.B2(n_17),
.Y(n_257)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_199),
.Y(n_258)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_258),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_259),
.Y(n_316)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_178),
.Y(n_260)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_260),
.Y(n_348)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_140),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_261),
.Y(n_340)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_148),
.Y(n_263)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_263),
.Y(n_352)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_140),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_264),
.B(n_265),
.Y(n_313)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_218),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_158),
.Y(n_266)
);

INVx11_ASAP7_75t_L g324 ( 
.A(n_266),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_136),
.B(n_18),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_268),
.B(n_271),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_211),
.A2(n_8),
.B1(n_16),
.B2(n_155),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_192),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_208),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_272),
.B(n_273),
.Y(n_334)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_169),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_158),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_274),
.B(n_277),
.Y(n_338)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_151),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_275),
.Y(n_306)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_194),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_276),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_164),
.B(n_149),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_214),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_278),
.B(n_279),
.Y(n_347)
);

BUFx12f_ASAP7_75t_L g279 ( 
.A(n_205),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_153),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_280),
.B(n_282),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_136),
.A2(n_135),
.B1(n_144),
.B2(n_132),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_207),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_180),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_283),
.B(n_286),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_284),
.A2(n_289),
.B1(n_292),
.B2(n_295),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_189),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_285),
.Y(n_330)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_194),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_129),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_133),
.B(n_130),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_177),
.Y(n_317)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_179),
.Y(n_289)
);

A2O1A1O1Ixp25_ASAP7_75t_L g290 ( 
.A1(n_210),
.A2(n_195),
.B(n_156),
.C(n_200),
.D(n_190),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_290),
.A2(n_270),
.B(n_238),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_293),
.Y(n_305)
);

OAI22x1_ASAP7_75t_L g292 ( 
.A1(n_155),
.A2(n_196),
.B1(n_139),
.B2(n_142),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_168),
.B(n_181),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_154),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_296),
.Y(n_312)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_182),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_203),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_176),
.B(n_187),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_298),
.Y(n_321)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_185),
.Y(n_298)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_185),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_301),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_300),
.A2(n_177),
.B1(n_167),
.B2(n_157),
.Y(n_315)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_204),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_189),
.B(n_217),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_285),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_249),
.A2(n_173),
.B(n_209),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_304),
.A2(n_360),
.B(n_306),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_231),
.A2(n_217),
.B1(n_154),
.B2(n_209),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_308),
.A2(n_315),
.B1(n_326),
.B2(n_341),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_237),
.B(n_141),
.CI(n_184),
.CON(n_309),
.SN(n_309)
);

A2O1A1Ixp33_ASAP7_75t_L g369 ( 
.A1(n_309),
.A2(n_339),
.B(n_335),
.C(n_328),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_317),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_269),
.A2(n_157),
.B1(n_167),
.B2(n_184),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_326),
.A2(n_335),
.B1(n_339),
.B2(n_357),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_332),
.B(n_349),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_292),
.A2(n_259),
.B1(n_267),
.B2(n_262),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_244),
.A2(n_268),
.B1(n_242),
.B2(n_290),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_256),
.B(n_288),
.C(n_226),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_343),
.B(n_279),
.C(n_225),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_240),
.B(n_230),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_356),
.A2(n_320),
.B(n_360),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_244),
.A2(n_233),
.B1(n_257),
.B2(n_252),
.Y(n_357)
);

NAND2x1_ASAP7_75t_L g360 ( 
.A(n_244),
.B(n_239),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_357),
.A2(n_227),
.B1(n_266),
.B2(n_241),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_SL g425 ( 
.A1(n_361),
.A2(n_362),
.B1(n_390),
.B2(n_376),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_358),
.A2(n_276),
.B1(n_253),
.B2(n_258),
.Y(n_362)
);

BUFx8_ASAP7_75t_L g363 ( 
.A(n_325),
.Y(n_363)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_363),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_223),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_364),
.B(n_381),
.C(n_394),
.Y(n_416)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_312),
.Y(n_365)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_365),
.Y(n_414)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_312),
.Y(n_366)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_366),
.Y(n_418)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_322),
.Y(n_367)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_367),
.Y(n_439)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_311),
.Y(n_368)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_368),
.Y(n_441)
);

OAI21xp33_ASAP7_75t_L g428 ( 
.A1(n_369),
.A2(n_389),
.B(n_331),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_338),
.B(n_228),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_371),
.B(n_384),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_354),
.A2(n_224),
.B1(n_251),
.B2(n_286),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_372),
.A2(n_374),
.B1(n_392),
.B2(n_396),
.Y(n_419)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_322),
.Y(n_373)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_373),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_314),
.A2(n_358),
.B1(n_305),
.B2(n_304),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_332),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_375),
.B(n_379),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_314),
.A2(n_250),
.B1(n_299),
.B2(n_275),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_376),
.A2(n_324),
.B1(n_341),
.B2(n_346),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_377),
.B(n_399),
.Y(n_433)
);

A2O1A1Ixp33_ASAP7_75t_SL g378 ( 
.A1(n_360),
.A2(n_232),
.B(n_279),
.C(n_356),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_378),
.A2(n_395),
.B(n_401),
.Y(n_407)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_311),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_318),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_380),
.B(n_310),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_305),
.B(n_321),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_349),
.B(n_321),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_383),
.B(n_387),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_347),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_329),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_385),
.B(n_386),
.Y(n_412)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_324),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_317),
.B(n_309),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_318),
.B(n_333),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_388),
.B(n_398),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_309),
.B(n_319),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_391),
.B(n_400),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_316),
.A2(n_315),
.B1(n_333),
.B2(n_336),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_336),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_393),
.B(n_397),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_334),
.B(n_359),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_316),
.A2(n_353),
.B(n_355),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_330),
.A2(n_323),
.B1(n_325),
.B2(n_306),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_342),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_313),
.B(n_352),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_350),
.Y(n_400)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_352),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_402),
.B(n_310),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_323),
.B(n_303),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_403),
.B(n_404),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_346),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_303),
.B(n_348),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_405),
.B(n_379),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_401),
.A2(n_340),
.B(n_327),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_408),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_369),
.A2(n_340),
.B(n_327),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_410),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_421),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_370),
.A2(n_330),
.B1(n_341),
.B2(n_329),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_415),
.A2(n_424),
.B1(n_420),
.B2(n_429),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_417),
.B(n_396),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g460 ( 
.A1(n_420),
.A2(n_425),
.B1(n_363),
.B2(n_385),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_383),
.B(n_344),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_382),
.B(n_344),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_423),
.B(n_436),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_370),
.A2(n_331),
.B1(n_348),
.B2(n_351),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_364),
.B(n_337),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_427),
.B(n_434),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_R g457 ( 
.A(n_428),
.B(n_438),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_374),
.A2(n_351),
.B1(n_337),
.B2(n_345),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_429),
.A2(n_432),
.B1(n_380),
.B2(n_405),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_399),
.B(n_345),
.C(n_307),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_433),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_375),
.A2(n_307),
.B1(n_365),
.B2(n_366),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_381),
.B(n_382),
.Y(n_434)
);

AND2x2_ASAP7_75t_SL g438 ( 
.A(n_387),
.B(n_367),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_373),
.B(n_403),
.Y(n_440)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_440),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_444),
.A2(n_445),
.B1(n_467),
.B2(n_411),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_406),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_377),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_461),
.C(n_433),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_414),
.A2(n_378),
.B1(n_391),
.B2(n_392),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_449),
.A2(n_454),
.B1(n_460),
.B2(n_469),
.Y(n_486)
);

CKINVDCx14_ASAP7_75t_R g506 ( 
.A(n_450),
.Y(n_506)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_441),
.Y(n_451)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_451),
.Y(n_478)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_441),
.Y(n_453)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_453),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_419),
.A2(n_394),
.B1(n_378),
.B2(n_389),
.Y(n_454)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_435),
.Y(n_456)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_456),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_419),
.A2(n_378),
.B1(n_372),
.B2(n_363),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_458),
.B(n_411),
.Y(n_491)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_435),
.Y(n_459)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_459),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_416),
.B(n_395),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_436),
.Y(n_462)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_462),
.Y(n_490)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_413),
.Y(n_463)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_463),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_409),
.B(n_404),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_464),
.B(n_465),
.Y(n_505)
);

OAI21xp33_ASAP7_75t_SL g465 ( 
.A1(n_430),
.A2(n_378),
.B(n_400),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_432),
.Y(n_466)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_466),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_406),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_406),
.Y(n_468)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_468),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_409),
.A2(n_386),
.B1(n_397),
.B2(n_418),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_471),
.A2(n_472),
.B1(n_439),
.B2(n_417),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_424),
.A2(n_415),
.B1(n_418),
.B2(n_414),
.Y(n_472)
);

OAI22x1_ASAP7_75t_L g473 ( 
.A1(n_407),
.A2(n_408),
.B1(n_410),
.B2(n_430),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_473),
.Y(n_507)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_440),
.Y(n_475)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_475),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_422),
.Y(n_476)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_476),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_446),
.A2(n_442),
.B1(n_439),
.B2(n_407),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_477),
.A2(n_487),
.B1(n_489),
.B2(n_495),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_479),
.B(n_482),
.C(n_499),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_447),
.B(n_427),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_480),
.B(n_488),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_443),
.B(n_431),
.C(n_434),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_449),
.A2(n_438),
.B1(n_426),
.B2(n_442),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_483),
.A2(n_498),
.B1(n_502),
.B2(n_477),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_443),
.B(n_438),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_446),
.A2(n_423),
.B1(n_426),
.B2(n_421),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_491),
.B(n_478),
.Y(n_530)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_493),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_475),
.A2(n_412),
.B1(n_437),
.B2(n_466),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_455),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_508),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_456),
.A2(n_459),
.B1(n_462),
.B2(n_445),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_470),
.B(n_461),
.C(n_468),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_455),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_500),
.B(n_453),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_467),
.A2(n_452),
.B1(n_472),
.B2(n_471),
.Y(n_502)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_451),
.Y(n_504)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_504),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_474),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_503),
.Y(n_510)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_510),
.Y(n_546)
);

AND2x2_ASAP7_75t_SL g548 ( 
.A(n_512),
.B(n_530),
.Y(n_548)
);

XNOR2x1_ASAP7_75t_L g514 ( 
.A(n_483),
.B(n_473),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_514),
.B(n_486),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_505),
.A2(n_452),
.B(n_448),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_515),
.B(n_521),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_480),
.B(n_470),
.C(n_448),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_516),
.B(n_517),
.C(n_527),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_479),
.B(n_463),
.C(n_474),
.Y(n_517)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_518),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_506),
.A2(n_457),
.B1(n_458),
.B2(n_507),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_519),
.A2(n_491),
.B1(n_490),
.B2(n_501),
.Y(n_549)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_498),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_481),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_522),
.B(n_523),
.Y(n_542)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_481),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_496),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_524),
.B(n_525),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_497),
.B(n_457),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_496),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_526),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_482),
.B(n_499),
.C(n_488),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_508),
.B(n_489),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_529),
.B(n_532),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_492),
.B(n_495),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_503),
.B(n_501),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_533),
.B(n_534),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_502),
.Y(n_534)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_535),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_531),
.B(n_484),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_537),
.Y(n_568)
);

XNOR2x2_ASAP7_75t_L g543 ( 
.A(n_525),
.B(n_507),
.Y(n_543)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_543),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_517),
.B(n_494),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_544),
.B(n_547),
.C(n_550),
.Y(n_555)
);

FAx1_ASAP7_75t_SL g545 ( 
.A(n_516),
.B(n_484),
.CI(n_485),
.CON(n_545),
.SN(n_545)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_545),
.B(n_532),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_531),
.B(n_485),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_549),
.A2(n_512),
.B1(n_521),
.B2(n_509),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_513),
.B(n_494),
.C(n_490),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_513),
.B(n_492),
.C(n_478),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_552),
.B(n_554),
.C(n_515),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_527),
.B(n_504),
.C(n_514),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_556),
.A2(n_565),
.B1(n_567),
.B2(n_537),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_557),
.B(n_559),
.Y(n_576)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_553),
.Y(n_558)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_558),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_552),
.B(n_528),
.C(n_509),
.Y(n_559)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_560),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_SL g561 ( 
.A1(n_538),
.A2(n_511),
.B(n_529),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_SL g582 ( 
.A1(n_561),
.A2(n_530),
.B(n_524),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_550),
.B(n_554),
.C(n_541),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_563),
.B(n_566),
.Y(n_578)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_536),
.Y(n_564)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_564),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_539),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_SL g566 ( 
.A1(n_551),
.A2(n_519),
.B1(n_546),
.B2(n_526),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_540),
.Y(n_567)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_542),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_569),
.B(n_570),
.Y(n_577)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_540),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_573),
.B(n_562),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_562),
.A2(n_548),
.B1(n_511),
.B2(n_530),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_574),
.A2(n_585),
.B1(n_571),
.B2(n_567),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_559),
.B(n_544),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_575),
.A2(n_580),
.B(n_581),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_557),
.B(n_547),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_555),
.B(n_535),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_582),
.A2(n_561),
.B(n_564),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_555),
.B(n_548),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_583),
.B(n_568),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_556),
.A2(n_548),
.B1(n_545),
.B2(n_520),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_575),
.B(n_563),
.C(n_541),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_586),
.B(n_590),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_587),
.B(n_589),
.Y(n_600)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_572),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_572),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_591),
.B(n_592),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_593),
.B(n_581),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_584),
.B(n_571),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_594),
.B(n_595),
.Y(n_602)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_582),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_576),
.B(n_565),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_596),
.A2(n_578),
.B(n_583),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_SL g599 ( 
.A(n_586),
.B(n_580),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_599),
.B(n_588),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_601),
.B(n_603),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_597),
.B(n_577),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_604),
.B(n_606),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_SL g610 ( 
.A1(n_605),
.A2(n_607),
.B(n_600),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_602),
.A2(n_589),
.B1(n_587),
.B2(n_579),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_600),
.A2(n_592),
.B(n_585),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_610),
.B(n_608),
.C(n_598),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_SL g612 ( 
.A1(n_611),
.A2(n_609),
.B(n_573),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_612),
.A2(n_574),
.B(n_520),
.Y(n_613)
);

AO21x1_ASAP7_75t_L g614 ( 
.A1(n_613),
.A2(n_522),
.B(n_523),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_614),
.B(n_543),
.Y(n_615)
);


endmodule