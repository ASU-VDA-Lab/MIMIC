module fake_ariane_1710_n_1798 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1798);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1798;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1769;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_148),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_149),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_61),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_43),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_29),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_100),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_1),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_133),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_7),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_5),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_54),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_136),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_88),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_19),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_110),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_14),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_20),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_125),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_80),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_6),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_18),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_154),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_127),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_48),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_93),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_108),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_62),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_113),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_142),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_152),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_102),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_65),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g194 ( 
.A(n_58),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_27),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_3),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_121),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_109),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_7),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_63),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_10),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_60),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_26),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_66),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_44),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_98),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_9),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_27),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_33),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_25),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_39),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_40),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_87),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_0),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_77),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_1),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_116),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_151),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_24),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_6),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_99),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_155),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_31),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_106),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_10),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_55),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_76),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_128),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_33),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_105),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_101),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_147),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_56),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_39),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_42),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_120),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_26),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_146),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_75),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_51),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_74),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_20),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_72),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_14),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_2),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_44),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_140),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_94),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_15),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_25),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_22),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_67),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_112),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_138),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_157),
.Y(n_255)
);

BUFx2_ASAP7_75t_SL g256 ( 
.A(n_12),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_126),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_9),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_5),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_114),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_159),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_23),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_35),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_36),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_68),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_21),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_59),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_24),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_35),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_40),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_50),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_115),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_103),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_95),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_69),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_52),
.Y(n_276)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_11),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_18),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_38),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_85),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_32),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_47),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_111),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_131),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_23),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_15),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_79),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_83),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_53),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_2),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_0),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_82),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_45),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_47),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_84),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_22),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_141),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_11),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_37),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_123),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_96),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_97),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_129),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_73),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_16),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_48),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_21),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_122),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_36),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_135),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_119),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_130),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_46),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_8),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_78),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_86),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_8),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_117),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_28),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_4),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_256),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_169),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_264),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_169),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_169),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_169),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_242),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_169),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_178),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_178),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_242),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_266),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_167),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_212),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_184),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_178),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_178),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_212),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_198),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_240),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_178),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_254),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_196),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_234),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_196),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_196),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_249),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_199),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_201),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_203),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_196),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_170),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_163),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_250),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_208),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_282),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_209),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_196),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_312),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_211),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_306),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_223),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_229),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_164),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_164),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_306),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_306),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_306),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_181),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_190),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_182),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_306),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_194),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_177),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_177),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_235),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_210),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_170),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_210),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_172),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_172),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_222),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_222),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_233),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_244),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_205),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_233),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_243),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_243),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_271),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_245),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_271),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_245),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_194),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_245),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_246),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_285),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_285),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_345),
.B(n_174),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_352),
.B(n_188),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_346),
.B(n_176),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g402 ( 
.A(n_352),
.B(n_188),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_333),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_378),
.B(n_348),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_380),
.B(n_206),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_378),
.B(n_226),
.Y(n_406)
);

OA21x2_ASAP7_75t_L g407 ( 
.A1(n_322),
.A2(n_221),
.B(n_217),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_322),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_343),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_343),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_368),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_368),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_340),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_324),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_324),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_325),
.Y(n_416)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_380),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_344),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_323),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_325),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_326),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_327),
.B(n_226),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_326),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_328),
.Y(n_424)
);

NOR2xp67_ASAP7_75t_L g425 ( 
.A(n_381),
.B(n_276),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_328),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_329),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_329),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_381),
.B(n_224),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_364),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_330),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_382),
.B(n_227),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_330),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_336),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_382),
.B(n_230),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_336),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_337),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_337),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_341),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_332),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_364),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_341),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_351),
.Y(n_443)
);

OR2x6_ASAP7_75t_L g444 ( 
.A(n_393),
.B(n_195),
.Y(n_444)
);

OR2x6_ASAP7_75t_L g445 ( 
.A(n_397),
.B(n_207),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_351),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_359),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_358),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_358),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_361),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_361),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_383),
.B(n_238),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_366),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_366),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_367),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_383),
.B(n_239),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_367),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_331),
.B(n_194),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_372),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_372),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_384),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_384),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_387),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_387),
.Y(n_464)
);

OA21x2_ASAP7_75t_L g465 ( 
.A1(n_388),
.A2(n_247),
.B(n_241),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_342),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_373),
.A2(n_394),
.B1(n_391),
.B2(n_395),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_388),
.B(n_389),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_389),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_390),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_390),
.B(n_248),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_392),
.Y(n_472)
);

NAND3xp33_ASAP7_75t_L g473 ( 
.A(n_404),
.B(n_350),
.C(n_349),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_419),
.B(n_365),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_463),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_453),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_463),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_458),
.B(n_355),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_462),
.Y(n_479)
);

NAND2xp33_ASAP7_75t_R g480 ( 
.A(n_440),
.B(n_357),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_454),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_463),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_458),
.B(n_468),
.Y(n_483)
);

INVx8_ASAP7_75t_L g484 ( 
.A(n_422),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_422),
.B(n_360),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_462),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_408),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_458),
.B(n_362),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_422),
.B(n_363),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_463),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_422),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_445),
.Y(n_492)
);

OR2x6_ASAP7_75t_L g493 ( 
.A(n_445),
.B(n_331),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_454),
.Y(n_494)
);

NAND3xp33_ASAP7_75t_L g495 ( 
.A(n_430),
.B(n_385),
.C(n_376),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_464),
.Y(n_496)
);

BUFx4f_ASAP7_75t_L g497 ( 
.A(n_465),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_454),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_408),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_400),
.B(n_396),
.Y(n_500)
);

OAI22xp33_ASAP7_75t_L g501 ( 
.A1(n_444),
.A2(n_445),
.B1(n_430),
.B2(n_441),
.Y(n_501)
);

AND2x2_ASAP7_75t_SL g502 ( 
.A(n_440),
.B(n_273),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_418),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_454),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_414),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_453),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_414),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_414),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_420),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_415),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_417),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_463),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_400),
.B(n_321),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_400),
.B(n_392),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_415),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_415),
.Y(n_516)
);

INVx5_ASAP7_75t_L g517 ( 
.A(n_412),
.Y(n_517)
);

AO21x2_ASAP7_75t_L g518 ( 
.A1(n_399),
.A2(n_267),
.B(n_261),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_464),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_472),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_472),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_403),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_445),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_428),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_399),
.B(n_398),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_468),
.B(n_386),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_445),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_401),
.B(n_417),
.Y(n_528)
);

BUFx10_ASAP7_75t_L g529 ( 
.A(n_413),
.Y(n_529)
);

CKINVDCx6p67_ASAP7_75t_R g530 ( 
.A(n_466),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_428),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_463),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_428),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_419),
.Y(n_534)
);

INVx6_ASAP7_75t_L g535 ( 
.A(n_417),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_400),
.B(n_370),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_402),
.B(n_160),
.Y(n_537)
);

INVx5_ASAP7_75t_L g538 ( 
.A(n_412),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_431),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_468),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_468),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_470),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_431),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_420),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_402),
.B(n_353),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_431),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_L g547 ( 
.A(n_470),
.B(n_252),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_433),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_466),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_445),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_417),
.B(n_334),
.Y(n_551)
);

OAI22xp33_ASAP7_75t_L g552 ( 
.A1(n_444),
.A2(n_317),
.B1(n_258),
.B2(n_173),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_402),
.B(n_369),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_433),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_453),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_402),
.B(n_160),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_406),
.B(n_338),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_421),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_433),
.Y(n_559)
);

BUFx6f_ASAP7_75t_SL g560 ( 
.A(n_444),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_L g561 ( 
.A(n_470),
.B(n_252),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_434),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_434),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_470),
.Y(n_564)
);

NOR3xp33_ASAP7_75t_L g565 ( 
.A(n_441),
.B(n_277),
.C(n_168),
.Y(n_565)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_465),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_434),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_412),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_465),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_465),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_406),
.B(n_371),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_446),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_446),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_446),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_421),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_448),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_423),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_423),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_470),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_401),
.B(n_335),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_L g581 ( 
.A(n_470),
.B(n_252),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_406),
.B(n_425),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_416),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_424),
.Y(n_584)
);

BUFx4f_ASAP7_75t_L g585 ( 
.A(n_465),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_424),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_427),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_427),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_448),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_436),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_448),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_449),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_406),
.B(n_192),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_467),
.B(n_347),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_407),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_444),
.B(n_339),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_436),
.Y(n_597)
);

XOR2x2_ASAP7_75t_SL g598 ( 
.A(n_467),
.B(n_354),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_437),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_SL g600 ( 
.A(n_405),
.B(n_166),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_437),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_439),
.Y(n_602)
);

AND2x6_ASAP7_75t_L g603 ( 
.A(n_461),
.B(n_273),
.Y(n_603)
);

NOR2x1p5_ASAP7_75t_L g604 ( 
.A(n_444),
.B(n_166),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_425),
.B(n_161),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_412),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_412),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_407),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_449),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_412),
.Y(n_610)
);

INVx6_ASAP7_75t_L g611 ( 
.A(n_416),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_461),
.B(n_252),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_449),
.Y(n_613)
);

NOR2x1p5_ASAP7_75t_L g614 ( 
.A(n_444),
.B(n_168),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_455),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_439),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_442),
.Y(n_617)
);

INVx5_ASAP7_75t_L g618 ( 
.A(n_416),
.Y(n_618)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_447),
.B(n_356),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_405),
.B(n_161),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_442),
.Y(n_621)
);

INVx8_ASAP7_75t_L g622 ( 
.A(n_416),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_492),
.B(n_162),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_491),
.A2(n_276),
.B1(n_162),
.B2(n_297),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_492),
.B(n_165),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_491),
.B(n_461),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_525),
.B(n_469),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_505),
.Y(n_628)
);

AND2x6_ASAP7_75t_SL g629 ( 
.A(n_596),
.B(n_214),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_528),
.B(n_469),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_507),
.Y(n_631)
);

AO22x2_ASAP7_75t_L g632 ( 
.A1(n_598),
.A2(n_471),
.B1(n_429),
.B2(n_432),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_549),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_523),
.B(n_165),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_484),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_534),
.Y(n_636)
);

AND2x6_ASAP7_75t_SL g637 ( 
.A(n_522),
.B(n_216),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_476),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_484),
.B(n_469),
.Y(n_639)
);

NOR2xp67_ASAP7_75t_L g640 ( 
.A(n_549),
.B(n_429),
.Y(n_640)
);

O2A1O1Ixp5_ASAP7_75t_L g641 ( 
.A1(n_511),
.A2(n_620),
.B(n_605),
.C(n_532),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_487),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_502),
.A2(n_407),
.B1(n_452),
.B2(n_471),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_485),
.B(n_432),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_507),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_487),
.Y(n_646)
);

NAND3xp33_ASAP7_75t_L g647 ( 
.A(n_480),
.B(n_296),
.C(n_185),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_484),
.B(n_483),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_484),
.B(n_435),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_534),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_483),
.B(n_435),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_508),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_493),
.B(n_452),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_526),
.B(n_456),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_493),
.B(n_456),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_508),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_526),
.B(n_443),
.Y(n_657)
);

BUFx5_ASAP7_75t_L g658 ( 
.A(n_612),
.Y(n_658)
);

INVxp67_ASAP7_75t_SL g659 ( 
.A(n_523),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_510),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_551),
.B(n_540),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_510),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_L g663 ( 
.A1(n_527),
.A2(n_185),
.B1(n_296),
.B2(n_298),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_550),
.B(n_171),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_550),
.A2(n_175),
.B1(n_311),
.B2(n_304),
.Y(n_665)
);

INVx8_ASAP7_75t_L g666 ( 
.A(n_493),
.Y(n_666)
);

INVx8_ASAP7_75t_L g667 ( 
.A(n_493),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_L g668 ( 
.A(n_522),
.B(n_175),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_604),
.B(n_614),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_551),
.B(n_443),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_515),
.Y(n_671)
);

BUFx6f_ASAP7_75t_SL g672 ( 
.A(n_529),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_530),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_502),
.A2(n_407),
.B1(n_459),
.B2(n_457),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_541),
.B(n_450),
.Y(n_675)
);

NOR3xp33_ASAP7_75t_L g676 ( 
.A(n_478),
.B(n_220),
.C(n_219),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_617),
.B(n_179),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_518),
.A2(n_407),
.B1(n_459),
.B2(n_457),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_489),
.B(n_450),
.Y(n_679)
);

NAND2x1p5_ASAP7_75t_L g680 ( 
.A(n_476),
.B(n_460),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_475),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_500),
.B(n_251),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_529),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_580),
.B(n_460),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_515),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_474),
.B(n_374),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_479),
.B(n_200),
.Y(n_687)
);

NOR2xp67_ASAP7_75t_L g688 ( 
.A(n_473),
.B(n_455),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_486),
.B(n_283),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_499),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_474),
.B(n_557),
.Y(n_691)
);

NOR2xp67_ASAP7_75t_L g692 ( 
.A(n_495),
.B(n_455),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_496),
.B(n_289),
.Y(n_693)
);

OR2x6_ASAP7_75t_L g694 ( 
.A(n_536),
.B(n_374),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_617),
.B(n_179),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_509),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_488),
.B(n_263),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_511),
.B(n_270),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_511),
.B(n_278),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_516),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_516),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_519),
.B(n_520),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_524),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_509),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_521),
.B(n_316),
.Y(n_705)
);

NAND2x1p5_ASAP7_75t_L g706 ( 
.A(n_506),
.B(n_272),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_531),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_SL g708 ( 
.A(n_529),
.B(n_231),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_582),
.B(n_180),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_531),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_L g711 ( 
.A(n_481),
.B(n_180),
.Y(n_711)
);

CKINVDCx14_ASAP7_75t_R g712 ( 
.A(n_503),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_544),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_533),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_L g715 ( 
.A(n_481),
.B(n_183),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_533),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_593),
.B(n_183),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_557),
.B(n_186),
.Y(n_718)
);

BUFx5_ASAP7_75t_L g719 ( 
.A(n_612),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_475),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_619),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_497),
.A2(n_299),
.B(n_262),
.C(n_259),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_617),
.B(n_497),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_497),
.B(n_186),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_513),
.B(n_292),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_518),
.A2(n_225),
.B1(n_294),
.B2(n_237),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_585),
.B(n_475),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_585),
.B(n_292),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_585),
.B(n_297),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_565),
.B(n_375),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_514),
.B(n_300),
.Y(n_731)
);

O2A1O1Ixp5_ASAP7_75t_L g732 ( 
.A1(n_512),
.A2(n_308),
.B(n_295),
.C(n_310),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_535),
.A2(n_309),
.B1(n_305),
.B2(n_313),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_544),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_539),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_560),
.A2(n_303),
.B1(n_300),
.B2(n_301),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_475),
.B(n_301),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_475),
.B(n_477),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_503),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_539),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_537),
.B(n_279),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_543),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_545),
.B(n_302),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_553),
.B(n_571),
.Y(n_744)
);

NOR2xp67_ASAP7_75t_L g745 ( 
.A(n_558),
.B(n_575),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_619),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_518),
.B(n_302),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_566),
.A2(n_314),
.B1(n_268),
.B2(n_269),
.Y(n_748)
);

OAI22xp33_ASAP7_75t_L g749 ( 
.A1(n_501),
.A2(n_307),
.B1(n_281),
.B2(n_293),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_594),
.B(n_375),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_566),
.A2(n_319),
.B1(n_231),
.B2(n_411),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_558),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_506),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_556),
.B(n_286),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_477),
.B(n_303),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_535),
.B(n_304),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_535),
.B(n_290),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_535),
.B(n_311),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_477),
.B(n_275),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_543),
.Y(n_760)
);

NAND2x1_ASAP7_75t_L g761 ( 
.A(n_611),
.B(n_416),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_575),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_555),
.B(n_377),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_566),
.A2(n_231),
.B1(n_409),
.B2(n_411),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_569),
.A2(n_409),
.B1(n_410),
.B2(n_411),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_577),
.B(n_291),
.Y(n_766)
);

AOI22x1_ASAP7_75t_L g767 ( 
.A1(n_494),
.A2(n_298),
.B1(n_313),
.B2(n_305),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_587),
.B(n_320),
.Y(n_768)
);

BUFx8_ASAP7_75t_L g769 ( 
.A(n_560),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_588),
.B(n_309),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_578),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_590),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_546),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_477),
.B(n_315),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_578),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_560),
.B(n_318),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_477),
.B(n_416),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_546),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_512),
.B(n_532),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_594),
.B(n_377),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_548),
.Y(n_781)
);

A2O1A1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_584),
.A2(n_379),
.B(n_410),
.C(n_409),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_548),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_554),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_482),
.B(n_426),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_494),
.B(n_187),
.Y(n_786)
);

INVxp33_ASAP7_75t_L g787 ( 
.A(n_598),
.Y(n_787)
);

INVx5_ASAP7_75t_L g788 ( 
.A(n_635),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_632),
.A2(n_552),
.B1(n_570),
.B2(n_569),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_642),
.Y(n_790)
);

AND2x4_ASAP7_75t_SL g791 ( 
.A(n_673),
.B(n_512),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_666),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_681),
.B(n_498),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_683),
.Y(n_794)
);

NOR3xp33_ASAP7_75t_L g795 ( 
.A(n_697),
.B(n_600),
.C(n_621),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_636),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_630),
.A2(n_504),
.B(n_498),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_627),
.A2(n_504),
.B(n_621),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_646),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_644),
.B(n_586),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_644),
.B(n_586),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_672),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_632),
.A2(n_748),
.B1(n_726),
.B2(n_749),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_648),
.B(n_532),
.Y(n_804)
);

NOR2x2_ASAP7_75t_L g805 ( 
.A(n_694),
.B(n_600),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_690),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_683),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_654),
.B(n_597),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_635),
.B(n_482),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_739),
.Y(n_810)
);

CKINVDCx8_ASAP7_75t_R g811 ( 
.A(n_637),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_696),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_704),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_653),
.B(n_542),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_SL g815 ( 
.A(n_633),
.B(n_569),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_651),
.B(n_684),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_653),
.B(n_542),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_686),
.Y(n_818)
);

INVx5_ASAP7_75t_L g819 ( 
.A(n_666),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_745),
.A2(n_599),
.B(n_597),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_691),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_640),
.B(n_599),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_661),
.B(n_601),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_652),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_632),
.A2(n_570),
.B1(n_595),
.B2(n_608),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_681),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_666),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_681),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_667),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_650),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_716),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_713),
.A2(n_616),
.B(n_601),
.C(n_602),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_734),
.Y(n_833)
);

NOR3xp33_ASAP7_75t_SL g834 ( 
.A(n_733),
.B(n_602),
.C(n_616),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_750),
.B(n_379),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_752),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_744),
.B(n_570),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_723),
.B(n_482),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_655),
.A2(n_579),
.B1(n_542),
.B2(n_564),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_682),
.B(n_554),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_762),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_716),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_771),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_760),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_682),
.B(n_559),
.Y(n_845)
);

AO22x2_ASAP7_75t_L g846 ( 
.A1(n_780),
.A2(n_787),
.B1(n_749),
.B2(n_747),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_760),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_712),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_775),
.Y(n_849)
);

AND2x6_ASAP7_75t_L g850 ( 
.A(n_655),
.B(n_482),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_681),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_723),
.B(n_482),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_720),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_669),
.B(n_694),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_649),
.B(n_720),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_702),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_669),
.B(n_564),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_784),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_748),
.A2(n_595),
.B1(n_608),
.B2(n_615),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_667),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_763),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_726),
.A2(n_595),
.B1(n_608),
.B2(n_615),
.Y(n_862)
);

AO22x1_ASAP7_75t_L g863 ( 
.A1(n_787),
.A2(n_603),
.B1(n_612),
.B2(n_215),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_698),
.B(n_559),
.Y(n_864)
);

NOR2x1p5_ASAP7_75t_L g865 ( 
.A(n_647),
.B(n_564),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_720),
.B(n_490),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_763),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_772),
.Y(n_868)
);

OAI22xp33_ASAP7_75t_L g869 ( 
.A1(n_708),
.A2(n_579),
.B1(n_613),
.B2(n_576),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_730),
.B(n_562),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_698),
.B(n_562),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_675),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_699),
.B(n_563),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_784),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_628),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_699),
.B(n_563),
.Y(n_876)
);

OR2x6_ASAP7_75t_L g877 ( 
.A(n_667),
.B(n_622),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_631),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_679),
.B(n_567),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_657),
.B(n_567),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_645),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_643),
.B(n_572),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_643),
.B(n_572),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_656),
.Y(n_884)
);

INVx4_ASAP7_75t_L g885 ( 
.A(n_672),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_660),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_662),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_720),
.B(n_490),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_671),
.Y(n_889)
);

OAI22xp33_ASAP7_75t_L g890 ( 
.A1(n_670),
.A2(n_579),
.B1(n_613),
.B2(n_573),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_685),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_724),
.A2(n_583),
.B(n_622),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_638),
.Y(n_893)
);

OR2x6_ASAP7_75t_L g894 ( 
.A(n_706),
.B(n_622),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_700),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_659),
.B(n_583),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_701),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_677),
.A2(n_583),
.B1(n_611),
.B2(n_490),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_757),
.B(n_574),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_703),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_638),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_677),
.A2(n_611),
.B1(n_490),
.B2(n_622),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_779),
.A2(n_589),
.B(n_574),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_707),
.Y(n_904)
);

INVxp67_ASAP7_75t_SL g905 ( 
.A(n_639),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_710),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_714),
.Y(n_907)
);

AND2x2_ASAP7_75t_SL g908 ( 
.A(n_674),
.B(n_547),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_769),
.Y(n_909)
);

AOI221xp5_ASAP7_75t_SL g910 ( 
.A1(n_663),
.A2(n_609),
.B1(n_592),
.B2(n_591),
.C(n_589),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_753),
.B(n_490),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_SL g912 ( 
.A(n_721),
.B(n_603),
.Y(n_912)
);

OR2x6_ASAP7_75t_L g913 ( 
.A(n_706),
.B(n_576),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_753),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_676),
.B(n_606),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_735),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_695),
.B(n_606),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_757),
.B(n_591),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_695),
.A2(n_611),
.B1(n_603),
.B2(n_609),
.Y(n_919)
);

AOI211xp5_ASAP7_75t_L g920 ( 
.A1(n_697),
.A2(n_561),
.B(n_547),
.C(n_581),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_740),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_687),
.B(n_592),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_727),
.B(n_618),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_769),
.Y(n_924)
);

NOR3xp33_ASAP7_75t_SL g925 ( 
.A(n_770),
.B(n_189),
.C(n_191),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_689),
.B(n_607),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_693),
.B(n_607),
.Y(n_927)
);

NAND2xp33_ASAP7_75t_L g928 ( 
.A(n_756),
.B(n_618),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_705),
.B(n_718),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_742),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_680),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_773),
.Y(n_932)
);

BUFx12f_ASAP7_75t_L g933 ( 
.A(n_629),
.Y(n_933)
);

NAND3xp33_ASAP7_75t_SL g934 ( 
.A(n_624),
.B(n_193),
.C(n_197),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_680),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_717),
.B(n_610),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_725),
.B(n_776),
.Y(n_937)
);

NOR3xp33_ASAP7_75t_SL g938 ( 
.A(n_766),
.B(n_202),
.C(n_204),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_674),
.A2(n_603),
.B1(n_410),
.B2(n_612),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_778),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_781),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_746),
.B(n_603),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_751),
.A2(n_612),
.B1(n_561),
.B2(n_426),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_668),
.B(n_426),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_761),
.Y(n_945)
);

OAI21xp33_ASAP7_75t_L g946 ( 
.A1(n_741),
.A2(n_754),
.B(n_768),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_776),
.B(n_618),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_741),
.B(n_426),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_623),
.B(n_625),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_783),
.Y(n_950)
);

INVxp67_ASAP7_75t_L g951 ( 
.A(n_623),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_626),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_751),
.A2(n_612),
.B1(n_426),
.B2(n_438),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_743),
.B(n_618),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_731),
.B(n_618),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_727),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_709),
.B(n_517),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_782),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_754),
.B(n_517),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_665),
.B(n_517),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_782),
.Y(n_961)
);

NOR2x1p5_ASAP7_75t_L g962 ( 
.A(n_758),
.B(n_213),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_777),
.Y(n_963)
);

BUFx4f_ASAP7_75t_L g964 ( 
.A(n_625),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_779),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_692),
.B(n_517),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_634),
.A2(n_274),
.B1(n_228),
.B2(n_232),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_786),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_688),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_800),
.A2(n_738),
.B(n_729),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_837),
.A2(n_724),
.B(n_728),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_819),
.B(n_634),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_801),
.A2(n_738),
.B(n_728),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_819),
.B(n_664),
.Y(n_974)
);

AOI21x1_ASAP7_75t_L g975 ( 
.A1(n_838),
.A2(n_729),
.B(n_759),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_816),
.A2(n_871),
.B(n_864),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_790),
.Y(n_977)
);

AOI222xp33_ASAP7_75t_L g978 ( 
.A1(n_803),
.A2(n_821),
.B1(n_933),
.B2(n_846),
.C1(n_835),
.C2(n_946),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_796),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_803),
.A2(n_722),
.B1(n_764),
.B2(n_664),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_873),
.A2(n_641),
.B(n_715),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_937),
.B(n_736),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_794),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_856),
.B(n_722),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_964),
.B(n_767),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_929),
.B(n_737),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_819),
.B(n_785),
.Y(n_987)
);

NAND2xp33_ASAP7_75t_SL g988 ( 
.A(n_834),
.B(n_737),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_872),
.B(n_818),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_808),
.A2(n_764),
.B1(n_755),
.B2(n_765),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_799),
.Y(n_991)
);

NOR3xp33_ASAP7_75t_L g992 ( 
.A(n_934),
.B(n_755),
.C(n_711),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_795),
.A2(n_732),
.B(n_774),
.C(n_759),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_949),
.A2(n_774),
.B1(n_777),
.B2(n_785),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_949),
.A2(n_765),
.B(n_678),
.C(n_568),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_802),
.Y(n_996)
);

INVx4_ASAP7_75t_L g997 ( 
.A(n_819),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_792),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_876),
.A2(n_823),
.B(n_820),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_830),
.B(n_854),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_870),
.B(n_678),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_820),
.A2(n_517),
.B(n_538),
.Y(n_1002)
);

BUFx4_ASAP7_75t_SL g1003 ( 
.A(n_924),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_834),
.A2(n_568),
.B(n_538),
.C(n_426),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_840),
.A2(n_538),
.B(n_568),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_845),
.A2(n_538),
.B(n_568),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_957),
.A2(n_538),
.B(n_568),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_806),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_797),
.A2(n_265),
.B(n_236),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_797),
.A2(n_280),
.B(n_253),
.Y(n_1010)
);

INVx5_ASAP7_75t_L g1011 ( 
.A(n_877),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_846),
.A2(n_719),
.B1(n_658),
.B2(n_451),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_846),
.B(n_719),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_861),
.A2(n_719),
.B1(n_658),
.B2(n_451),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_879),
.A2(n_284),
.B(n_255),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_955),
.A2(n_287),
.B(n_257),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_795),
.A2(n_3),
.B(n_4),
.C(n_12),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_830),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_812),
.Y(n_1019)
);

OR2x6_ASAP7_75t_L g1020 ( 
.A(n_792),
.B(n_719),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_SL g1021 ( 
.A1(n_832),
.A2(n_965),
.B(n_852),
.C(n_838),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_798),
.A2(n_288),
.B(n_260),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_867),
.B(n_719),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_810),
.Y(n_1024)
);

NAND3xp33_ASAP7_75t_SL g1025 ( 
.A(n_811),
.B(n_925),
.C(n_967),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_SL g1026 ( 
.A1(n_804),
.A2(n_892),
.B(n_798),
.C(n_914),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_788),
.B(n_719),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_822),
.A2(n_13),
.B(n_16),
.C(n_17),
.Y(n_1028)
);

NAND3xp33_ASAP7_75t_L g1029 ( 
.A(n_815),
.B(n_968),
.C(n_832),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_934),
.A2(n_951),
.B(n_868),
.C(n_833),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_917),
.A2(n_451),
.B(n_438),
.C(n_218),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_952),
.B(n_658),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_827),
.B(n_438),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_892),
.A2(n_903),
.B(n_852),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_854),
.B(n_438),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_813),
.Y(n_1036)
);

AO21x1_ASAP7_75t_L g1037 ( 
.A1(n_855),
.A2(n_658),
.B(n_451),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_788),
.B(n_658),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_899),
.A2(n_252),
.B(n_451),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_942),
.B(n_13),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_807),
.Y(n_1041)
);

CKINVDCx11_ASAP7_75t_R g1042 ( 
.A(n_885),
.Y(n_1042)
);

AO21x1_ASAP7_75t_L g1043 ( 
.A1(n_855),
.A2(n_451),
.B(n_438),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_836),
.B(n_17),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_909),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_918),
.A2(n_438),
.B(n_89),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_788),
.B(n_19),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_857),
.B(n_848),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_841),
.B(n_28),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_954),
.A2(n_90),
.B(n_156),
.Y(n_1050)
);

BUFx12f_ASAP7_75t_L g1051 ( 
.A(n_885),
.Y(n_1051)
);

AO21x1_ASAP7_75t_L g1052 ( 
.A1(n_869),
.A2(n_890),
.B(n_923),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_788),
.B(n_29),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_908),
.A2(n_789),
.B1(n_891),
.B2(n_950),
.Y(n_1054)
);

OR2x6_ASAP7_75t_L g1055 ( 
.A(n_877),
.B(n_30),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_905),
.A2(n_91),
.B(n_153),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_824),
.Y(n_1057)
);

O2A1O1Ixp5_ASAP7_75t_L g1058 ( 
.A1(n_809),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_905),
.A2(n_92),
.B(n_150),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_938),
.Y(n_1060)
);

NOR2xp67_ASAP7_75t_L g1061 ( 
.A(n_829),
.B(n_860),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_831),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_793),
.A2(n_81),
.B(n_144),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_869),
.B(n_34),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_814),
.B(n_34),
.Y(n_1065)
);

NAND2x1p5_ASAP7_75t_L g1066 ( 
.A(n_931),
.B(n_935),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_843),
.B(n_37),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_849),
.B(n_38),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_880),
.A2(n_107),
.B(n_143),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_928),
.A2(n_104),
.B(n_139),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_917),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_877),
.B(n_41),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_910),
.A2(n_45),
.B(n_46),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_828),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_857),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_828),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_814),
.B(n_49),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_817),
.B(n_49),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_935),
.B(n_57),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_791),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_817),
.A2(n_64),
.B1(n_70),
.B2(n_71),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_865),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_828),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_908),
.A2(n_118),
.B1(n_124),
.B2(n_132),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_969),
.B(n_134),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_850),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_969),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_828),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_850),
.B(n_158),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_842),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_866),
.A2(n_888),
.B(n_936),
.Y(n_1091)
);

BUFx2_ASAP7_75t_R g1092 ( 
.A(n_945),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_804),
.A2(n_911),
.B(n_925),
.C(n_893),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_850),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_935),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_866),
.A2(n_888),
.B(n_890),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_915),
.B(n_922),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_959),
.A2(n_911),
.B(n_923),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_809),
.A2(n_927),
.B(n_926),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_948),
.A2(n_958),
.B(n_961),
.C(n_920),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_947),
.A2(n_882),
.B(n_883),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_850),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_875),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_960),
.A2(n_896),
.B(n_963),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_850),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_935),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_901),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_SL g1108 ( 
.A1(n_912),
.A2(n_805),
.B1(n_915),
.B2(n_913),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_844),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_SL g1110 ( 
.A1(n_826),
.A2(n_851),
.B(n_853),
.C(n_898),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_789),
.B(n_913),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_896),
.A2(n_826),
.B(n_853),
.Y(n_1112)
);

OAI21xp33_ASAP7_75t_L g1113 ( 
.A1(n_938),
.A2(n_839),
.B(n_944),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_913),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_919),
.A2(n_825),
.B(n_962),
.C(n_902),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1034),
.A2(n_825),
.B(n_874),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_976),
.A2(n_851),
.B(n_894),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1000),
.B(n_900),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_986),
.B(n_847),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_977),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_991),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_979),
.B(n_901),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1078),
.A2(n_939),
.B1(n_859),
.B2(n_953),
.Y(n_1123)
);

CKINVDCx14_ASAP7_75t_R g1124 ( 
.A(n_996),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1008),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_1018),
.B(n_901),
.Y(n_1126)
);

O2A1O1Ixp5_ASAP7_75t_L g1127 ( 
.A1(n_988),
.A2(n_863),
.B(n_966),
.C(n_858),
.Y(n_1127)
);

BUFx12f_ASAP7_75t_L g1128 ( 
.A(n_1042),
.Y(n_1128)
);

AND2x2_ASAP7_75t_SL g1129 ( 
.A(n_1086),
.B(n_939),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1043),
.A2(n_1052),
.A3(n_1037),
.B(n_1013),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1091),
.A2(n_1098),
.B(n_1099),
.Y(n_1131)
);

AO31x2_ASAP7_75t_L g1132 ( 
.A1(n_1101),
.A2(n_1115),
.A3(n_980),
.B(n_995),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1097),
.B(n_862),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1029),
.A2(n_859),
.B(n_862),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_998),
.Y(n_1135)
);

AOI21x1_ASAP7_75t_L g1136 ( 
.A1(n_999),
.A2(n_894),
.B(n_966),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1019),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1096),
.A2(n_878),
.B(n_881),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_1071),
.A2(n_894),
.B(n_886),
.C(n_887),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_R g1140 ( 
.A(n_1051),
.B(n_901),
.Y(n_1140)
);

OA21x2_ASAP7_75t_L g1141 ( 
.A1(n_971),
.A2(n_943),
.B(n_889),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1055),
.A2(n_953),
.B1(n_956),
.B2(n_897),
.Y(n_1142)
);

O2A1O1Ixp5_ASAP7_75t_SL g1143 ( 
.A1(n_985),
.A2(n_884),
.B(n_895),
.C(n_941),
.Y(n_1143)
);

O2A1O1Ixp5_ASAP7_75t_L g1144 ( 
.A1(n_1064),
.A2(n_921),
.B(n_940),
.C(n_907),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_R g1145 ( 
.A(n_1041),
.B(n_1045),
.Y(n_1145)
);

BUFx5_ASAP7_75t_L g1146 ( 
.A(n_1102),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1039),
.A2(n_930),
.B(n_932),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1011),
.B(n_956),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_978),
.B(n_904),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_998),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_978),
.B(n_906),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1104),
.A2(n_916),
.B(n_956),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1046),
.A2(n_956),
.B(n_981),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1029),
.A2(n_971),
.B(n_970),
.Y(n_1154)
);

NAND2x1p5_ASAP7_75t_L g1155 ( 
.A(n_1086),
.B(n_1094),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1021),
.A2(n_973),
.B(n_1026),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1036),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1100),
.A2(n_990),
.B(n_1073),
.Y(n_1158)
);

NAND3xp33_ASAP7_75t_L g1159 ( 
.A(n_992),
.B(n_1028),
.C(n_1022),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_989),
.B(n_1075),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1003),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1011),
.B(n_1114),
.Y(n_1162)
);

NOR2xp67_ASAP7_75t_L g1163 ( 
.A(n_983),
.B(n_1087),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1108),
.B(n_1048),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_990),
.A2(n_1007),
.B(n_1002),
.Y(n_1165)
);

NAND2x1p5_ASAP7_75t_L g1166 ( 
.A(n_1094),
.B(n_1011),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1103),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1049),
.Y(n_1168)
);

AO21x1_ASAP7_75t_L g1169 ( 
.A1(n_980),
.A2(n_1022),
.B(n_1093),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_975),
.A2(n_1006),
.B(n_1005),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_1092),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1072),
.B(n_1085),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1073),
.A2(n_993),
.B(n_1004),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1070),
.A2(n_1050),
.B(n_1056),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_984),
.B(n_1001),
.Y(n_1175)
);

AOI221x1_ASAP7_75t_L g1176 ( 
.A1(n_1113),
.A2(n_1040),
.B1(n_1111),
.B2(n_1031),
.C(n_1059),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_994),
.A2(n_1030),
.B(n_1068),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1049),
.Y(n_1178)
);

AOI211x1_ASAP7_75t_L g1179 ( 
.A1(n_1065),
.A2(n_1068),
.B(n_1044),
.C(n_1067),
.Y(n_1179)
);

NAND2x1p5_ASAP7_75t_L g1180 ( 
.A(n_1011),
.B(n_1105),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1063),
.A2(n_1069),
.B(n_1032),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1110),
.A2(n_1112),
.B(n_1032),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1084),
.A2(n_1058),
.B(n_1009),
.Y(n_1183)
);

BUFx8_ASAP7_75t_SL g1184 ( 
.A(n_1024),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_997),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1027),
.A2(n_1038),
.B(n_1016),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_997),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1047),
.A2(n_1053),
.B(n_1010),
.Y(n_1188)
);

OA21x2_ASAP7_75t_L g1189 ( 
.A1(n_1012),
.A2(n_1054),
.B(n_1023),
.Y(n_1189)
);

OAI21xp33_ASAP7_75t_L g1190 ( 
.A1(n_1025),
.A2(n_1060),
.B(n_1055),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1089),
.A2(n_1083),
.B(n_1074),
.Y(n_1191)
);

INVx4_ASAP7_75t_L g1192 ( 
.A(n_998),
.Y(n_1192)
);

INVx3_ASAP7_75t_SL g1193 ( 
.A(n_1055),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1074),
.A2(n_1083),
.B(n_1079),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_SL g1195 ( 
.A1(n_1020),
.A2(n_1072),
.B(n_974),
.Y(n_1195)
);

INVx5_ASAP7_75t_L g1196 ( 
.A(n_1020),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1057),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1035),
.B(n_1114),
.Y(n_1198)
);

INVx5_ASAP7_75t_L g1199 ( 
.A(n_1020),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1062),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1014),
.A2(n_1066),
.B(n_1090),
.Y(n_1201)
);

BUFx2_ASAP7_75t_SL g1202 ( 
.A(n_1080),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1066),
.A2(n_1109),
.B(n_1081),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1077),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1015),
.A2(n_1061),
.B(n_1076),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_972),
.B(n_974),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1076),
.A2(n_1088),
.B(n_1106),
.Y(n_1207)
);

NAND2xp33_ASAP7_75t_L g1208 ( 
.A(n_1076),
.B(n_1088),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1082),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_972),
.B(n_1088),
.Y(n_1210)
);

OR2x2_ASAP7_75t_SL g1211 ( 
.A(n_1095),
.B(n_1106),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_987),
.A2(n_1033),
.B1(n_1107),
.B2(n_1106),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1095),
.A2(n_1043),
.A3(n_1052),
.B(n_1037),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_987),
.A2(n_1034),
.B(n_1091),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1033),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1018),
.B(n_691),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1018),
.B(n_691),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1034),
.A2(n_1091),
.B(n_1098),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_976),
.A2(n_801),
.B(n_800),
.Y(n_1219)
);

AO31x2_ASAP7_75t_L g1220 ( 
.A1(n_1043),
.A2(n_1052),
.A3(n_1037),
.B(n_1013),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_998),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_986),
.B(n_800),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_986),
.B(n_549),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1000),
.B(n_821),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1034),
.A2(n_1091),
.B(n_1098),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1011),
.B(n_819),
.Y(n_1226)
);

INVxp67_ASAP7_75t_L g1227 ( 
.A(n_1000),
.Y(n_1227)
);

NOR4xp25_ASAP7_75t_L g1228 ( 
.A(n_1017),
.B(n_803),
.C(n_1071),
.D(n_749),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_998),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_986),
.B(n_549),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_986),
.B(n_800),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_979),
.B(n_522),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_998),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1000),
.B(n_691),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_976),
.A2(n_801),
.B(n_800),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1034),
.A2(n_1091),
.B(n_1098),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_986),
.A2(n_946),
.B(n_949),
.C(n_988),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1029),
.A2(n_971),
.B(n_976),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_976),
.A2(n_801),
.B(n_800),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_979),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1034),
.A2(n_1091),
.B(n_1098),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1018),
.B(n_691),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1018),
.B(n_691),
.Y(n_1243)
);

INVxp67_ASAP7_75t_SL g1244 ( 
.A(n_1018),
.Y(n_1244)
);

INVxp67_ASAP7_75t_SL g1245 ( 
.A(n_1018),
.Y(n_1245)
);

AO31x2_ASAP7_75t_L g1246 ( 
.A1(n_1043),
.A2(n_1052),
.A3(n_1037),
.B(n_1013),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1000),
.B(n_691),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1034),
.A2(n_1091),
.B(n_1098),
.Y(n_1248)
);

NAND3xp33_ASAP7_75t_L g1249 ( 
.A(n_1017),
.B(n_834),
.C(n_946),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_977),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1024),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1018),
.B(n_691),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1018),
.B(n_691),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_R g1254 ( 
.A(n_996),
.B(n_503),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1034),
.A2(n_1091),
.B(n_1098),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1034),
.A2(n_1091),
.B(n_1098),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_976),
.A2(n_801),
.B(n_800),
.Y(n_1257)
);

AOI21xp33_ASAP7_75t_L g1258 ( 
.A1(n_978),
.A2(n_632),
.B(n_980),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1034),
.A2(n_1091),
.B(n_1098),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1034),
.A2(n_1091),
.B(n_1098),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_986),
.B(n_800),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1123),
.A2(n_1190),
.B1(n_1172),
.B2(n_1232),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1223),
.B(n_1230),
.Y(n_1263)
);

NAND3xp33_ASAP7_75t_SL g1264 ( 
.A(n_1237),
.B(n_1169),
.C(n_1177),
.Y(n_1264)
);

CKINVDCx11_ASAP7_75t_R g1265 ( 
.A(n_1128),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1249),
.A2(n_1159),
.B(n_1222),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1170),
.A2(n_1153),
.B(n_1218),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_1254),
.Y(n_1268)
);

OAI221xp5_ASAP7_75t_L g1269 ( 
.A1(n_1228),
.A2(n_1249),
.B1(n_1159),
.B2(n_1177),
.C(n_1190),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1225),
.A2(n_1241),
.B(n_1236),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1222),
.A2(n_1261),
.B1(n_1231),
.B2(n_1204),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1120),
.Y(n_1272)
);

CKINVDCx11_ASAP7_75t_R g1273 ( 
.A(n_1171),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1234),
.B(n_1247),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_1145),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1248),
.A2(n_1256),
.B(n_1255),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1259),
.A2(n_1260),
.B(n_1165),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1116),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1131),
.A2(n_1181),
.B(n_1156),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1161),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1226),
.Y(n_1281)
);

NAND3xp33_ASAP7_75t_L g1282 ( 
.A(n_1179),
.B(n_1261),
.C(n_1231),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1158),
.A2(n_1243),
.B1(n_1242),
.B2(n_1252),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1136),
.A2(n_1174),
.B(n_1191),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1143),
.A2(n_1138),
.B(n_1214),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1132),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1238),
.A2(n_1154),
.B(n_1158),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1121),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1176),
.A2(n_1182),
.A3(n_1142),
.B(n_1239),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1130),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_1226),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1132),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1124),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1134),
.A2(n_1258),
.B(n_1183),
.C(n_1219),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1117),
.A2(n_1147),
.B(n_1152),
.Y(n_1295)
);

OA21x2_ASAP7_75t_L g1296 ( 
.A1(n_1238),
.A2(n_1154),
.B(n_1134),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1186),
.A2(n_1257),
.B(n_1235),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1125),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1228),
.A2(n_1178),
.B(n_1168),
.C(n_1139),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1224),
.B(n_1227),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1142),
.A2(n_1175),
.A3(n_1133),
.B(n_1119),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1203),
.A2(n_1194),
.B(n_1127),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1184),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1137),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1201),
.A2(n_1188),
.B(n_1207),
.Y(n_1305)
);

NOR2x1_ASAP7_75t_SL g1306 ( 
.A(n_1196),
.B(n_1199),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1258),
.A2(n_1149),
.B1(n_1151),
.B2(n_1133),
.Y(n_1307)
);

O2A1O1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1216),
.A2(n_1253),
.B(n_1217),
.C(n_1245),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1144),
.A2(n_1205),
.B(n_1155),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_1171),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1157),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1118),
.B(n_1160),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1250),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1132),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1193),
.B(n_1240),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1244),
.B(n_1175),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1167),
.Y(n_1317)
);

AOI21xp33_ASAP7_75t_L g1318 ( 
.A1(n_1141),
.A2(n_1198),
.B(n_1129),
.Y(n_1318)
);

NOR2x1_ASAP7_75t_SL g1319 ( 
.A(n_1196),
.B(n_1199),
.Y(n_1319)
);

NAND3xp33_ASAP7_75t_L g1320 ( 
.A(n_1126),
.B(n_1122),
.C(n_1209),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1197),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1163),
.A2(n_1208),
.B(n_1155),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1206),
.A2(n_1196),
.B(n_1199),
.C(n_1164),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1195),
.A2(n_1166),
.B(n_1189),
.Y(n_1324)
);

OR2x6_ASAP7_75t_L g1325 ( 
.A(n_1166),
.B(n_1180),
.Y(n_1325)
);

BUFx12f_ASAP7_75t_L g1326 ( 
.A(n_1135),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1189),
.A2(n_1200),
.B1(n_1206),
.B2(n_1215),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1210),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1185),
.A2(n_1187),
.B(n_1212),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1210),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1180),
.A2(n_1187),
.B(n_1185),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1212),
.A2(n_1213),
.B(n_1246),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1130),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1202),
.B(n_1140),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1211),
.B(n_1162),
.Y(n_1335)
);

OAI222xp33_ASAP7_75t_L g1336 ( 
.A1(n_1162),
.A2(n_1148),
.B1(n_1192),
.B2(n_1146),
.C1(n_1246),
.C2(n_1130),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1220),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1135),
.B(n_1221),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1213),
.A2(n_1246),
.B(n_1220),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1220),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1146),
.A2(n_1150),
.B(n_1221),
.Y(n_1341)
);

BUFx2_ASAP7_75t_R g1342 ( 
.A(n_1146),
.Y(n_1342)
);

INVx2_ASAP7_75t_R g1343 ( 
.A(n_1229),
.Y(n_1343)
);

OA21x2_ASAP7_75t_L g1344 ( 
.A1(n_1229),
.A2(n_1165),
.B(n_1156),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1233),
.B(n_1222),
.Y(n_1345)
);

CKINVDCx11_ASAP7_75t_R g1346 ( 
.A(n_1128),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1120),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1170),
.A2(n_1153),
.B(n_1218),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1120),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1237),
.A2(n_1249),
.B(n_1159),
.Y(n_1350)
);

CKINVDCx14_ASAP7_75t_R g1351 ( 
.A(n_1254),
.Y(n_1351)
);

AO21x2_ASAP7_75t_L g1352 ( 
.A1(n_1177),
.A2(n_1258),
.B(n_1013),
.Y(n_1352)
);

CKINVDCx16_ASAP7_75t_R g1353 ( 
.A(n_1254),
.Y(n_1353)
);

AND2x6_ASAP7_75t_L g1354 ( 
.A(n_1226),
.B(n_1111),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1226),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1211),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1120),
.Y(n_1357)
);

NAND2x1p5_ASAP7_75t_L g1358 ( 
.A(n_1196),
.B(n_1086),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1162),
.B(n_1215),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1254),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1120),
.Y(n_1361)
);

NAND3xp33_ASAP7_75t_L g1362 ( 
.A(n_1237),
.B(n_1249),
.C(n_708),
.Y(n_1362)
);

AO21x2_ASAP7_75t_L g1363 ( 
.A1(n_1177),
.A2(n_1258),
.B(n_1013),
.Y(n_1363)
);

NOR2xp67_ASAP7_75t_SL g1364 ( 
.A(n_1128),
.B(n_683),
.Y(n_1364)
);

OR2x6_ASAP7_75t_L g1365 ( 
.A(n_1195),
.B(n_1142),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1170),
.A2(n_1153),
.B(n_1218),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1226),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1226),
.Y(n_1368)
);

AO21x2_ASAP7_75t_L g1369 ( 
.A1(n_1177),
.A2(n_1258),
.B(n_1013),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_SL g1370 ( 
.A1(n_1123),
.A2(n_632),
.B1(n_846),
.B2(n_502),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1249),
.A2(n_1231),
.B1(n_1261),
.B2(n_1222),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1258),
.A2(n_978),
.B1(n_632),
.B2(n_846),
.Y(n_1372)
);

NAND3xp33_ASAP7_75t_L g1373 ( 
.A(n_1237),
.B(n_1249),
.C(n_708),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1258),
.A2(n_978),
.B1(n_632),
.B2(n_846),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1116),
.Y(n_1375)
);

NOR3xp33_ASAP7_75t_L g1376 ( 
.A(n_1249),
.B(n_1237),
.C(n_1159),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1251),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1234),
.B(n_1247),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1258),
.A2(n_978),
.B1(n_632),
.B2(n_846),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1237),
.A2(n_946),
.B(n_982),
.C(n_1223),
.Y(n_1380)
);

O2A1O1Ixp5_ASAP7_75t_L g1381 ( 
.A1(n_1158),
.A2(n_1169),
.B(n_988),
.C(n_1173),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1120),
.Y(n_1382)
);

OA21x2_ASAP7_75t_L g1383 ( 
.A1(n_1165),
.A2(n_1156),
.B(n_1131),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1258),
.A2(n_978),
.B1(n_632),
.B2(n_846),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1251),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1162),
.B(n_1215),
.Y(n_1386)
);

INVxp33_ASAP7_75t_L g1387 ( 
.A(n_1232),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1177),
.A2(n_1258),
.B(n_1013),
.Y(n_1388)
);

NOR2x1_ASAP7_75t_SL g1389 ( 
.A(n_1196),
.B(n_1199),
.Y(n_1389)
);

O2A1O1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1350),
.A2(n_1269),
.B(n_1376),
.C(n_1380),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_SL g1391 ( 
.A1(n_1353),
.A2(n_1351),
.B1(n_1360),
.B2(n_1268),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1356),
.B(n_1359),
.Y(n_1392)
);

NOR2x1_ASAP7_75t_SL g1393 ( 
.A(n_1365),
.B(n_1325),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1271),
.B(n_1316),
.Y(n_1394)
);

INVx4_ASAP7_75t_L g1395 ( 
.A(n_1326),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1371),
.B(n_1312),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1300),
.B(n_1274),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1378),
.B(n_1377),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1356),
.B(n_1359),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1272),
.Y(n_1400)
);

NOR3xp33_ASAP7_75t_L g1401 ( 
.A(n_1362),
.B(n_1373),
.C(n_1264),
.Y(n_1401)
);

OA21x2_ASAP7_75t_L g1402 ( 
.A1(n_1339),
.A2(n_1279),
.B(n_1297),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1280),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1345),
.B(n_1266),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1386),
.B(n_1335),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1262),
.A2(n_1370),
.B1(n_1376),
.B2(n_1387),
.Y(n_1406)
);

BUFx12f_ASAP7_75t_L g1407 ( 
.A(n_1265),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1273),
.Y(n_1408)
);

OA21x2_ASAP7_75t_L g1409 ( 
.A1(n_1277),
.A2(n_1285),
.B(n_1381),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1383),
.A2(n_1294),
.B(n_1344),
.Y(n_1410)
);

NOR2x1_ASAP7_75t_SL g1411 ( 
.A(n_1365),
.B(n_1325),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1383),
.A2(n_1344),
.B(n_1287),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1385),
.B(n_1263),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1288),
.Y(n_1414)
);

NOR2xp67_ASAP7_75t_L g1415 ( 
.A(n_1320),
.B(n_1282),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_SL g1416 ( 
.A1(n_1308),
.A2(n_1299),
.B(n_1322),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1268),
.Y(n_1417)
);

BUFx12f_ASAP7_75t_L g1418 ( 
.A(n_1265),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1298),
.Y(n_1419)
);

OAI211xp5_ASAP7_75t_L g1420 ( 
.A1(n_1370),
.A2(n_1283),
.B(n_1263),
.C(n_1384),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1328),
.B(n_1330),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1387),
.A2(n_1374),
.B1(n_1384),
.B2(n_1372),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1304),
.B(n_1311),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_1273),
.Y(n_1424)
);

O2A1O1Ixp5_ASAP7_75t_L g1425 ( 
.A1(n_1286),
.A2(n_1314),
.B(n_1292),
.C(n_1336),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1372),
.A2(n_1374),
.B1(n_1379),
.B2(n_1351),
.Y(n_1426)
);

O2A1O1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1287),
.A2(n_1296),
.B(n_1315),
.C(n_1329),
.Y(n_1427)
);

AOI221x1_ASAP7_75t_SL g1428 ( 
.A1(n_1313),
.A2(n_1361),
.B1(n_1382),
.B2(n_1347),
.C(n_1357),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1317),
.B(n_1349),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1379),
.A2(n_1360),
.B1(n_1307),
.B2(n_1287),
.Y(n_1430)
);

AOI211xp5_ASAP7_75t_L g1431 ( 
.A1(n_1315),
.A2(n_1364),
.B(n_1275),
.C(n_1334),
.Y(n_1431)
);

BUFx5_ASAP7_75t_L g1432 ( 
.A(n_1354),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1326),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1383),
.A2(n_1344),
.B(n_1267),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1301),
.B(n_1296),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1307),
.A2(n_1296),
.B1(n_1310),
.B2(n_1293),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1310),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1293),
.A2(n_1342),
.B1(n_1323),
.B2(n_1327),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1303),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1321),
.B(n_1338),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1346),
.Y(n_1441)
);

AOI211xp5_ASAP7_75t_L g1442 ( 
.A1(n_1290),
.A2(n_1336),
.B(n_1323),
.C(n_1318),
.Y(n_1442)
);

NAND3xp33_ASAP7_75t_L g1443 ( 
.A(n_1327),
.B(n_1341),
.C(n_1314),
.Y(n_1443)
);

AOI21x1_ASAP7_75t_SL g1444 ( 
.A1(n_1278),
.A2(n_1366),
.B(n_1348),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1301),
.B(n_1363),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1355),
.B(n_1368),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1343),
.B(n_1368),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1301),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1281),
.B(n_1367),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1289),
.Y(n_1450)
);

AOI221x1_ASAP7_75t_SL g1451 ( 
.A1(n_1346),
.A2(n_1333),
.B1(n_1340),
.B2(n_1337),
.C(n_1289),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1352),
.Y(n_1452)
);

A2O1A1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1324),
.A2(n_1332),
.B(n_1333),
.C(n_1340),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1291),
.B(n_1367),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1289),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1354),
.A2(n_1369),
.B1(n_1363),
.B2(n_1388),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1284),
.A2(n_1270),
.B(n_1276),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1295),
.A2(n_1302),
.B(n_1305),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1306),
.A2(n_1389),
.B(n_1319),
.Y(n_1459)
);

NOR3xp33_ASAP7_75t_L g1460 ( 
.A(n_1331),
.B(n_1309),
.C(n_1375),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1358),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1312),
.B(n_1316),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_SL g1463 ( 
.A1(n_1353),
.A2(n_1351),
.B1(n_1360),
.B2(n_1268),
.Y(n_1463)
);

O2A1O1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1350),
.A2(n_1237),
.B(n_1269),
.C(n_1376),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1271),
.B(n_1316),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1272),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1308),
.A2(n_1123),
.B(n_1172),
.Y(n_1467)
);

CKINVDCx20_ASAP7_75t_R g1468 ( 
.A(n_1293),
.Y(n_1468)
);

O2A1O1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1350),
.A2(n_1237),
.B(n_1269),
.C(n_1376),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1262),
.A2(n_1373),
.B1(n_1362),
.B2(n_1269),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1274),
.B(n_1378),
.Y(n_1471)
);

O2A1O1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1350),
.A2(n_1237),
.B(n_1269),
.C(n_1376),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_SL g1473 ( 
.A1(n_1308),
.A2(n_1123),
.B(n_1172),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1274),
.B(n_1378),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_R g1475 ( 
.A(n_1351),
.B(n_1161),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1274),
.B(n_1378),
.Y(n_1476)
);

A2O1A1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1262),
.A2(n_946),
.B(n_1373),
.C(n_1362),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1400),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1434),
.A2(n_1412),
.B(n_1410),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1466),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1423),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1435),
.B(n_1450),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1429),
.Y(n_1483)
);

OAI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1390),
.A2(n_1469),
.B(n_1464),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1448),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1414),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1394),
.B(n_1465),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1402),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1432),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1419),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1455),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1432),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1432),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1396),
.B(n_1428),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_SL g1495 ( 
.A1(n_1390),
.A2(n_1464),
.B(n_1469),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1421),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1425),
.A2(n_1456),
.B(n_1453),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1452),
.Y(n_1498)
);

INVxp67_ASAP7_75t_L g1499 ( 
.A(n_1440),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1409),
.B(n_1445),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1458),
.B(n_1427),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1427),
.B(n_1404),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1443),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1471),
.B(n_1474),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1462),
.B(n_1397),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1447),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1476),
.B(n_1413),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1460),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1457),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1457),
.B(n_1398),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_1475),
.Y(n_1511)
);

OR2x6_ASAP7_75t_L g1512 ( 
.A(n_1459),
.B(n_1438),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1436),
.B(n_1430),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1415),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1472),
.B(n_1401),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1393),
.Y(n_1516)
);

OAI21xp33_ASAP7_75t_SL g1517 ( 
.A1(n_1467),
.A2(n_1473),
.B(n_1416),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1451),
.Y(n_1518)
);

OR2x6_ASAP7_75t_L g1519 ( 
.A(n_1420),
.B(n_1392),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1487),
.B(n_1472),
.Y(n_1520)
);

AND2x2_ASAP7_75t_SL g1521 ( 
.A(n_1497),
.B(n_1392),
.Y(n_1521)
);

OAI33xp33_ASAP7_75t_L g1522 ( 
.A1(n_1515),
.A2(n_1406),
.A3(n_1470),
.B1(n_1422),
.B2(n_1426),
.B3(n_1463),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1510),
.B(n_1442),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1511),
.Y(n_1524)
);

AOI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_1484),
.A2(n_1420),
.B1(n_1477),
.B2(n_1431),
.C(n_1391),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1487),
.B(n_1437),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1489),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1510),
.B(n_1411),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1509),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1510),
.B(n_1446),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1502),
.B(n_1405),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1498),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1491),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1500),
.B(n_1501),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1489),
.B(n_1399),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1500),
.B(n_1449),
.Y(n_1536)
);

NOR4xp25_ASAP7_75t_SL g1537 ( 
.A(n_1518),
.B(n_1424),
.C(n_1408),
.D(n_1441),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1509),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1485),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1485),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1502),
.B(n_1405),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1505),
.B(n_1454),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1478),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1491),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1492),
.B(n_1399),
.Y(n_1545)
);

AOI211xp5_ASAP7_75t_SL g1546 ( 
.A1(n_1495),
.A2(n_1468),
.B(n_1461),
.C(n_1407),
.Y(n_1546)
);

BUFx4f_ASAP7_75t_SL g1547 ( 
.A(n_1511),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1488),
.B(n_1444),
.Y(n_1548)
);

AOI21xp33_ASAP7_75t_L g1549 ( 
.A1(n_1520),
.A2(n_1517),
.B(n_1484),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1539),
.Y(n_1550)
);

OR2x6_ASAP7_75t_L g1551 ( 
.A(n_1523),
.B(n_1516),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1539),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1534),
.B(n_1523),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1539),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1534),
.B(n_1507),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1522),
.A2(n_1515),
.B1(n_1517),
.B2(n_1513),
.Y(n_1556)
);

NAND5xp2_ASAP7_75t_SL g1557 ( 
.A(n_1524),
.B(n_1403),
.C(n_1504),
.D(n_1507),
.E(n_1418),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1547),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1520),
.A2(n_1514),
.B1(n_1494),
.B2(n_1512),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1540),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1527),
.B(n_1493),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1534),
.B(n_1507),
.Y(n_1562)
);

AND2x4_ASAP7_75t_SL g1563 ( 
.A(n_1535),
.B(n_1545),
.Y(n_1563)
);

OAI31xp33_ASAP7_75t_SL g1564 ( 
.A1(n_1523),
.A2(n_1504),
.A3(n_1518),
.B(n_1503),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1531),
.B(n_1514),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1529),
.Y(n_1566)
);

INVxp67_ASAP7_75t_SL g1567 ( 
.A(n_1533),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1533),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1530),
.B(n_1504),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1540),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1525),
.A2(n_1512),
.B1(n_1494),
.B2(n_1513),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1530),
.Y(n_1572)
);

INVxp67_ASAP7_75t_SL g1573 ( 
.A(n_1544),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1540),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1531),
.B(n_1499),
.Y(n_1575)
);

AOI33xp33_ASAP7_75t_L g1576 ( 
.A1(n_1525),
.A2(n_1503),
.A3(n_1486),
.B1(n_1490),
.B2(n_1483),
.B3(n_1480),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1530),
.B(n_1506),
.Y(n_1577)
);

AOI221xp5_ASAP7_75t_L g1578 ( 
.A1(n_1522),
.A2(n_1508),
.B1(n_1513),
.B2(n_1499),
.C(n_1481),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1544),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1528),
.B(n_1506),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1542),
.B(n_1505),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1529),
.Y(n_1582)
);

AOI221xp5_ASAP7_75t_L g1583 ( 
.A1(n_1548),
.A2(n_1508),
.B1(n_1481),
.B2(n_1488),
.C(n_1496),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1521),
.A2(n_1497),
.B1(n_1519),
.B2(n_1512),
.Y(n_1584)
);

INVxp67_ASAP7_75t_SL g1585 ( 
.A(n_1541),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1538),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1536),
.Y(n_1587)
);

INVx4_ASAP7_75t_L g1588 ( 
.A(n_1561),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1563),
.B(n_1527),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1568),
.Y(n_1590)
);

OA21x2_ASAP7_75t_L g1591 ( 
.A1(n_1566),
.A2(n_1479),
.B(n_1488),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1550),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1563),
.B(n_1561),
.Y(n_1593)
);

INVxp67_ASAP7_75t_SL g1594 ( 
.A(n_1556),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1553),
.B(n_1548),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1585),
.B(n_1543),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1550),
.Y(n_1597)
);

AND2x4_ASAP7_75t_SL g1598 ( 
.A(n_1555),
.B(n_1512),
.Y(n_1598)
);

INVxp67_ASAP7_75t_L g1599 ( 
.A(n_1559),
.Y(n_1599)
);

NAND3xp33_ASAP7_75t_SL g1600 ( 
.A(n_1556),
.B(n_1546),
.C(n_1537),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1552),
.Y(n_1601)
);

INVx4_ASAP7_75t_SL g1602 ( 
.A(n_1559),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1552),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1582),
.Y(n_1604)
);

BUFx2_ASAP7_75t_L g1605 ( 
.A(n_1561),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1579),
.Y(n_1606)
);

BUFx2_ASAP7_75t_L g1607 ( 
.A(n_1561),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1549),
.B(n_1526),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1554),
.Y(n_1609)
);

INVx3_ASAP7_75t_L g1610 ( 
.A(n_1553),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1554),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1582),
.Y(n_1612)
);

BUFx2_ASAP7_75t_L g1613 ( 
.A(n_1567),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1586),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1555),
.B(n_1548),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1562),
.B(n_1528),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1560),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1570),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1594),
.B(n_1581),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1591),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1591),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1610),
.B(n_1562),
.Y(n_1622)
);

AND4x1_ASAP7_75t_L g1623 ( 
.A(n_1608),
.B(n_1546),
.C(n_1564),
.D(n_1576),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1610),
.B(n_1595),
.Y(n_1624)
);

INVx2_ASAP7_75t_SL g1625 ( 
.A(n_1589),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1594),
.B(n_1581),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1610),
.B(n_1587),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1596),
.B(n_1575),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1591),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1596),
.B(n_1565),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1610),
.B(n_1595),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1610),
.B(n_1587),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1595),
.B(n_1569),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1591),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1608),
.B(n_1578),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1613),
.B(n_1583),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1600),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1613),
.B(n_1570),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1600),
.A2(n_1571),
.B1(n_1521),
.B2(n_1497),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1592),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1613),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1615),
.B(n_1569),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1609),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1615),
.B(n_1572),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1592),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1599),
.B(n_1547),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1597),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1615),
.B(n_1572),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1590),
.B(n_1573),
.Y(n_1649)
);

NAND4xp25_ASAP7_75t_L g1650 ( 
.A(n_1599),
.B(n_1558),
.C(n_1584),
.D(n_1417),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1590),
.B(n_1574),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1616),
.B(n_1580),
.Y(n_1652)
);

AOI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1609),
.A2(n_1541),
.B1(n_1557),
.B2(n_1482),
.C(n_1532),
.Y(n_1653)
);

OAI31xp33_ASAP7_75t_SL g1654 ( 
.A1(n_1602),
.A2(n_1557),
.A3(n_1528),
.B(n_1577),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1591),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1605),
.B(n_1551),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1605),
.B(n_1551),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1605),
.B(n_1551),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1607),
.B(n_1551),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1635),
.B(n_1606),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1641),
.B(n_1602),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1640),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1640),
.Y(n_1663)
);

NOR2x1_ASAP7_75t_L g1664 ( 
.A(n_1641),
.B(n_1439),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1641),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1645),
.Y(n_1666)
);

AND2x2_ASAP7_75t_SL g1667 ( 
.A(n_1623),
.B(n_1598),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1654),
.B(n_1593),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1635),
.B(n_1606),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1619),
.B(n_1597),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1645),
.Y(n_1671)
);

INVxp67_ASAP7_75t_SL g1672 ( 
.A(n_1637),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1623),
.B(n_1602),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1647),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1624),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1647),
.Y(n_1676)
);

NOR2x1p5_ASAP7_75t_L g1677 ( 
.A(n_1650),
.B(n_1524),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1625),
.B(n_1602),
.Y(n_1678)
);

OAI22xp33_ASAP7_75t_SL g1679 ( 
.A1(n_1637),
.A2(n_1607),
.B1(n_1602),
.B2(n_1512),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1654),
.B(n_1593),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1625),
.B(n_1602),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1651),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1639),
.A2(n_1521),
.B1(n_1497),
.B2(n_1512),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1619),
.B(n_1609),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1626),
.B(n_1601),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1626),
.B(n_1601),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1651),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1651),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1628),
.B(n_1603),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1643),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1638),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1638),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1633),
.B(n_1593),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1633),
.B(n_1593),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1636),
.B(n_1603),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1671),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1665),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1672),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1664),
.B(n_1625),
.Y(n_1699)
);

INVx1_ASAP7_75t_SL g1700 ( 
.A(n_1661),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1693),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1660),
.B(n_1628),
.Y(n_1702)
);

OR2x6_ASAP7_75t_L g1703 ( 
.A(n_1673),
.B(n_1395),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1671),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_1661),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1669),
.B(n_1630),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1695),
.B(n_1630),
.Y(n_1707)
);

NOR2x1_ASAP7_75t_L g1708 ( 
.A(n_1661),
.B(n_1678),
.Y(n_1708)
);

A2O1A1Ixp33_ASAP7_75t_SL g1709 ( 
.A1(n_1692),
.A2(n_1636),
.B(n_1646),
.C(n_1537),
.Y(n_1709)
);

CKINVDCx14_ASAP7_75t_R g1710 ( 
.A(n_1678),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1662),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1690),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1691),
.B(n_1633),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1667),
.A2(n_1653),
.B1(n_1521),
.B2(n_1620),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1667),
.A2(n_1653),
.B1(n_1634),
.B2(n_1629),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1675),
.B(n_1649),
.Y(n_1716)
);

INVxp67_ASAP7_75t_L g1717 ( 
.A(n_1682),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1678),
.B(n_1650),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1693),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1663),
.Y(n_1720)
);

NAND3xp33_ASAP7_75t_SL g1721 ( 
.A(n_1683),
.B(n_1680),
.C(n_1668),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1710),
.B(n_1677),
.Y(n_1722)
);

AOI21xp33_ASAP7_75t_L g1723 ( 
.A1(n_1698),
.A2(n_1679),
.B(n_1692),
.Y(n_1723)
);

AO221x1_ASAP7_75t_L g1724 ( 
.A1(n_1701),
.A2(n_1675),
.B1(n_1607),
.B2(n_1687),
.C(n_1688),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1696),
.Y(n_1725)
);

NAND2x1p5_ASAP7_75t_L g1726 ( 
.A(n_1708),
.B(n_1681),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1699),
.Y(n_1727)
);

INVxp67_ASAP7_75t_L g1728 ( 
.A(n_1703),
.Y(n_1728)
);

INVx2_ASAP7_75t_SL g1729 ( 
.A(n_1699),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1712),
.B(n_1687),
.Y(n_1730)
);

INVxp67_ASAP7_75t_L g1731 ( 
.A(n_1703),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1715),
.B(n_1681),
.Y(n_1732)
);

OAI32xp33_ASAP7_75t_L g1733 ( 
.A1(n_1714),
.A2(n_1668),
.A3(n_1680),
.B1(n_1684),
.B2(n_1685),
.Y(n_1733)
);

INVx3_ASAP7_75t_SL g1734 ( 
.A(n_1703),
.Y(n_1734)
);

NOR2x1_ASAP7_75t_L g1735 ( 
.A(n_1697),
.B(n_1681),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1705),
.B(n_1694),
.Y(n_1736)
);

NAND4xp25_ASAP7_75t_L g1737 ( 
.A(n_1712),
.B(n_1694),
.C(n_1686),
.D(n_1666),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1697),
.B(n_1642),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1702),
.B(n_1670),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1721),
.A2(n_1655),
.B1(n_1629),
.B2(n_1621),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1719),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1724),
.B(n_1706),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1735),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1736),
.B(n_1705),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1739),
.B(n_1700),
.Y(n_1745)
);

BUFx3_ASAP7_75t_L g1746 ( 
.A(n_1734),
.Y(n_1746)
);

INVxp33_ASAP7_75t_L g1747 ( 
.A(n_1726),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1726),
.Y(n_1748)
);

INVx1_ASAP7_75t_SL g1749 ( 
.A(n_1730),
.Y(n_1749)
);

INVx2_ASAP7_75t_SL g1750 ( 
.A(n_1729),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1722),
.B(n_1727),
.Y(n_1751)
);

NAND3x1_ASAP7_75t_L g1752 ( 
.A(n_1730),
.B(n_1718),
.C(n_1711),
.Y(n_1752)
);

AO21x1_ASAP7_75t_L g1753 ( 
.A1(n_1742),
.A2(n_1747),
.B(n_1732),
.Y(n_1753)
);

A2O1A1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1749),
.A2(n_1723),
.B(n_1740),
.C(n_1733),
.Y(n_1754)
);

AOI311xp33_ASAP7_75t_L g1755 ( 
.A1(n_1742),
.A2(n_1723),
.A3(n_1738),
.B(n_1709),
.C(n_1725),
.Y(n_1755)
);

AOI221xp5_ASAP7_75t_L g1756 ( 
.A1(n_1749),
.A2(n_1743),
.B1(n_1737),
.B2(n_1717),
.C(n_1748),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_SL g1757 ( 
.A1(n_1744),
.A2(n_1737),
.B(n_1731),
.Y(n_1757)
);

AOI221xp5_ASAP7_75t_L g1758 ( 
.A1(n_1745),
.A2(n_1704),
.B1(n_1720),
.B2(n_1741),
.C(n_1728),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1746),
.B(n_1707),
.Y(n_1759)
);

AOI222xp33_ASAP7_75t_L g1760 ( 
.A1(n_1750),
.A2(n_1621),
.B1(n_1629),
.B2(n_1620),
.C1(n_1655),
.C2(n_1634),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1751),
.B(n_1716),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_SL g1762 ( 
.A(n_1752),
.B(n_1649),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1746),
.B(n_1624),
.Y(n_1763)
);

OAI321xp33_ASAP7_75t_L g1764 ( 
.A1(n_1754),
.A2(n_1713),
.A3(n_1655),
.B1(n_1621),
.B2(n_1634),
.C(n_1620),
.Y(n_1764)
);

AOI322xp5_ASAP7_75t_L g1765 ( 
.A1(n_1756),
.A2(n_1676),
.A3(n_1674),
.B1(n_1657),
.B2(n_1656),
.C1(n_1658),
.C2(n_1659),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1761),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1759),
.Y(n_1767)
);

AOI31xp33_ASAP7_75t_L g1768 ( 
.A1(n_1753),
.A2(n_1685),
.A3(n_1670),
.B(n_1689),
.Y(n_1768)
);

AOI221xp5_ASAP7_75t_L g1769 ( 
.A1(n_1762),
.A2(n_1643),
.B1(n_1689),
.B2(n_1658),
.C(n_1657),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1767),
.B(n_1763),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1768),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1766),
.B(n_1763),
.Y(n_1772)
);

XOR2x2_ASAP7_75t_L g1773 ( 
.A(n_1769),
.B(n_1758),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1764),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1765),
.B(n_1755),
.Y(n_1775)
);

OAI322xp33_ASAP7_75t_L g1776 ( 
.A1(n_1771),
.A2(n_1757),
.A3(n_1760),
.B1(n_1659),
.B2(n_1658),
.C1(n_1657),
.C2(n_1656),
.Y(n_1776)
);

OAI211xp5_ASAP7_75t_L g1777 ( 
.A1(n_1775),
.A2(n_1659),
.B(n_1656),
.C(n_1624),
.Y(n_1777)
);

XNOR2x1_ASAP7_75t_L g1778 ( 
.A(n_1773),
.B(n_1631),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1770),
.B(n_1631),
.Y(n_1779)
);

XNOR2x1_ASAP7_75t_L g1780 ( 
.A(n_1773),
.B(n_1631),
.Y(n_1780)
);

NOR4xp75_ASAP7_75t_SL g1781 ( 
.A(n_1778),
.B(n_1770),
.C(n_1772),
.D(n_1774),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1780),
.B(n_1770),
.Y(n_1782)
);

XNOR2xp5_ASAP7_75t_L g1783 ( 
.A(n_1779),
.B(n_1598),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1782),
.Y(n_1784)
);

OAI322xp33_ASAP7_75t_SL g1785 ( 
.A1(n_1784),
.A2(n_1781),
.A3(n_1776),
.B1(n_1777),
.B2(n_1783),
.C1(n_1618),
.C2(n_1617),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1785),
.A2(n_1642),
.B1(n_1644),
.B2(n_1648),
.Y(n_1786)
);

OR3x1_ASAP7_75t_L g1787 ( 
.A(n_1785),
.B(n_1617),
.C(n_1611),
.Y(n_1787)
);

AO21x2_ASAP7_75t_L g1788 ( 
.A1(n_1787),
.A2(n_1642),
.B(n_1648),
.Y(n_1788)
);

AOI22x1_ASAP7_75t_L g1789 ( 
.A1(n_1786),
.A2(n_1588),
.B1(n_1632),
.B2(n_1627),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1789),
.A2(n_1788),
.B1(n_1644),
.B2(n_1648),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1788),
.A2(n_1644),
.B1(n_1622),
.B2(n_1627),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1790),
.A2(n_1622),
.B1(n_1632),
.B2(n_1627),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1791),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1793),
.A2(n_1604),
.B1(n_1612),
.B2(n_1614),
.Y(n_1794)
);

AO21x2_ASAP7_75t_L g1795 ( 
.A1(n_1794),
.A2(n_1792),
.B(n_1622),
.Y(n_1795)
);

INVxp67_ASAP7_75t_L g1796 ( 
.A(n_1795),
.Y(n_1796)
);

AOI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1796),
.A2(n_1395),
.B1(n_1433),
.B2(n_1632),
.Y(n_1797)
);

AOI211xp5_ASAP7_75t_L g1798 ( 
.A1(n_1797),
.A2(n_1433),
.B(n_1526),
.C(n_1652),
.Y(n_1798)
);


endmodule