module real_aes_7131_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_527;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g242 ( .A1(n_0), .A2(n_243), .B(n_244), .C(n_248), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_1), .B(n_184), .Y(n_249) );
INVx1_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_3), .B(n_156), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_4), .A2(n_142), .B(n_147), .C(n_513), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_5), .A2(n_137), .B(n_551), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_6), .A2(n_137), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_7), .B(n_184), .Y(n_557) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_8), .A2(n_172), .B(n_188), .Y(n_187) );
AND2x6_ASAP7_75t_L g142 ( .A(n_9), .B(n_143), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_10), .A2(n_142), .B(n_147), .C(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g495 ( .A(n_11), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_12), .B(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_12), .B(n_41), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_13), .B(n_247), .Y(n_515) );
INVx1_ASAP7_75t_L g166 ( .A(n_14), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_15), .B(n_156), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_16), .A2(n_157), .B(n_503), .C(n_505), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_17), .B(n_184), .Y(n_506) );
AOI22xp5_ASAP7_75t_SL g470 ( .A1(n_18), .A2(n_464), .B1(n_471), .B2(n_752), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_19), .A2(n_47), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_19), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_19), .B(n_221), .Y(n_594) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_20), .A2(n_147), .B(n_198), .C(n_217), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_21), .A2(n_196), .B(n_246), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_22), .B(n_247), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_23), .B(n_247), .Y(n_535) );
CKINVDCx16_ASAP7_75t_R g542 ( .A(n_24), .Y(n_542) );
INVx1_ASAP7_75t_L g534 ( .A(n_25), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_26), .A2(n_147), .B(n_191), .C(n_198), .Y(n_190) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_27), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_28), .Y(n_511) );
INVx1_ASAP7_75t_L g591 ( .A(n_29), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_30), .A2(n_137), .B(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g140 ( .A(n_31), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_32), .A2(n_145), .B(n_160), .C(n_206), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_33), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g553 ( .A1(n_34), .A2(n_246), .B(n_554), .C(n_556), .Y(n_553) );
INVxp67_ASAP7_75t_L g592 ( .A(n_35), .Y(n_592) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_36), .A2(n_46), .B1(n_128), .B2(n_129), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_36), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_37), .B(n_193), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_38), .A2(n_147), .B(n_198), .C(n_533), .Y(n_532) );
CKINVDCx14_ASAP7_75t_R g552 ( .A(n_39), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_40), .A2(n_45), .B1(n_478), .B2(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_40), .Y(n_479) );
INVx1_ASAP7_75t_L g114 ( .A(n_41), .Y(n_114) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_42), .A2(n_248), .B(n_493), .C(n_494), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_43), .B(n_215), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_44), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_45), .Y(n_478) );
INVx1_ASAP7_75t_L g129 ( .A(n_46), .Y(n_129) );
INVx1_ASAP7_75t_L g125 ( .A(n_47), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_48), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_49), .B(n_137), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_50), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_51), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_52), .A2(n_105), .B1(n_115), .B2(n_757), .Y(n_104) );
A2O1A1Ixp33_ASAP7_75t_L g144 ( .A1(n_53), .A2(n_145), .B(n_150), .C(n_160), .Y(n_144) );
INVx1_ASAP7_75t_L g245 ( .A(n_54), .Y(n_245) );
INVx1_ASAP7_75t_L g151 ( .A(n_55), .Y(n_151) );
INVx1_ASAP7_75t_L g523 ( .A(n_56), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_57), .B(n_137), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_58), .Y(n_224) );
CKINVDCx14_ASAP7_75t_R g491 ( .A(n_59), .Y(n_491) );
INVx1_ASAP7_75t_L g143 ( .A(n_60), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_61), .B(n_137), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_62), .B(n_184), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_63), .A2(n_178), .B(n_180), .C(n_182), .Y(n_177) );
INVx1_ASAP7_75t_L g165 ( .A(n_64), .Y(n_165) );
INVx1_ASAP7_75t_SL g555 ( .A(n_65), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_66), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_67), .B(n_156), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_68), .B(n_184), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_69), .B(n_157), .Y(n_259) );
INVx1_ASAP7_75t_L g545 ( .A(n_70), .Y(n_545) );
CKINVDCx16_ASAP7_75t_R g241 ( .A(n_71), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_72), .B(n_153), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_73), .A2(n_147), .B(n_160), .C(n_230), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g176 ( .A(n_74), .Y(n_176) );
INVx1_ASAP7_75t_L g112 ( .A(n_75), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_76), .A2(n_137), .B(n_490), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_77), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_78), .A2(n_137), .B(n_500), .Y(n_499) );
OAI22xp5_ASAP7_75t_SL g472 ( .A1(n_79), .A2(n_473), .B1(n_474), .B2(n_480), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_79), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_80), .A2(n_215), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g501 ( .A(n_81), .Y(n_501) );
CKINVDCx16_ASAP7_75t_R g531 ( .A(n_82), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_83), .B(n_152), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_84), .A2(n_475), .B1(n_476), .B2(n_477), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_84), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_85), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_86), .A2(n_137), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g504 ( .A(n_87), .Y(n_504) );
INVx2_ASAP7_75t_L g163 ( .A(n_88), .Y(n_163) );
INVx1_ASAP7_75t_L g514 ( .A(n_89), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_90), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_91), .B(n_247), .Y(n_260) );
INVx2_ASAP7_75t_L g109 ( .A(n_92), .Y(n_109) );
OR2x2_ASAP7_75t_L g463 ( .A(n_92), .B(n_464), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_93), .A2(n_147), .B(n_160), .C(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_94), .B(n_137), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_95), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g207 ( .A(n_96), .Y(n_207) );
INVxp67_ASAP7_75t_L g181 ( .A(n_97), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_98), .B(n_172), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g231 ( .A(n_100), .Y(n_231) );
INVx1_ASAP7_75t_L g255 ( .A(n_101), .Y(n_255) );
INVx2_ASAP7_75t_L g526 ( .A(n_102), .Y(n_526) );
AND2x2_ASAP7_75t_L g167 ( .A(n_103), .B(n_162), .Y(n_167) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_106), .Y(n_757) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_113), .Y(n_106) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .C(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g465 ( .A(n_108), .B(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g482 ( .A(n_109), .Y(n_482) );
INVx1_ASAP7_75t_L g751 ( .A(n_109), .Y(n_751) );
NOR2x2_ASAP7_75t_L g754 ( .A(n_109), .B(n_464), .Y(n_754) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_469), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_SL g756 ( .A(n_119), .Y(n_756) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_460), .B(n_467), .Y(n_121) );
XNOR2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_126), .Y(n_122) );
XOR2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_130), .Y(n_126) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_130), .A2(n_482), .B1(n_483), .B2(n_750), .Y(n_481) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OR5x1_ASAP7_75t_L g131 ( .A(n_132), .B(n_333), .C(n_411), .D(n_435), .E(n_452), .Y(n_131) );
OAI211xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_199), .B(n_250), .C(n_310), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_168), .Y(n_133) );
AND2x2_ASAP7_75t_L g264 ( .A(n_134), .B(n_170), .Y(n_264) );
INVx5_ASAP7_75t_SL g292 ( .A(n_134), .Y(n_292) );
AND2x2_ASAP7_75t_L g328 ( .A(n_134), .B(n_313), .Y(n_328) );
OR2x2_ASAP7_75t_L g367 ( .A(n_134), .B(n_169), .Y(n_367) );
OR2x2_ASAP7_75t_L g398 ( .A(n_134), .B(n_289), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_134), .B(n_302), .Y(n_434) );
AND2x2_ASAP7_75t_L g446 ( .A(n_134), .B(n_289), .Y(n_446) );
OR2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_167), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_144), .B(n_162), .Y(n_135) );
BUFx2_ASAP7_75t_L g215 ( .A(n_137), .Y(n_215) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_142), .Y(n_137) );
NAND2x1p5_ASAP7_75t_L g256 ( .A(n_138), .B(n_142), .Y(n_256) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
INVx1_ASAP7_75t_L g182 ( .A(n_139), .Y(n_182) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
INVx1_ASAP7_75t_L g197 ( .A(n_140), .Y(n_197) );
INVx1_ASAP7_75t_L g149 ( .A(n_141), .Y(n_149) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_141), .Y(n_154) );
INVx3_ASAP7_75t_L g157 ( .A(n_141), .Y(n_157) );
INVx1_ASAP7_75t_L g193 ( .A(n_141), .Y(n_193) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_141), .Y(n_247) );
INVx4_ASAP7_75t_SL g161 ( .A(n_142), .Y(n_161) );
BUFx3_ASAP7_75t_L g198 ( .A(n_142), .Y(n_198) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g175 ( .A1(n_146), .A2(n_161), .B(n_176), .C(n_177), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_SL g240 ( .A1(n_146), .A2(n_161), .B(n_241), .C(n_242), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g490 ( .A1(n_146), .A2(n_161), .B(n_491), .C(n_492), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_SL g500 ( .A1(n_146), .A2(n_161), .B(n_501), .C(n_502), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_SL g522 ( .A1(n_146), .A2(n_161), .B(n_523), .C(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g551 ( .A1(n_146), .A2(n_161), .B(n_552), .C(n_553), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_SL g587 ( .A1(n_146), .A2(n_161), .B(n_588), .C(n_589), .Y(n_587) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
BUFx3_ASAP7_75t_L g159 ( .A(n_148), .Y(n_159) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_148), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_155), .C(n_158), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_152), .A2(n_158), .B(n_207), .C(n_208), .Y(n_206) );
O2A1O1Ixp5_ASAP7_75t_L g513 ( .A1(n_152), .A2(n_514), .B(n_515), .C(n_516), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g544 ( .A1(n_152), .A2(n_516), .B(n_545), .C(n_546), .Y(n_544) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx4_ASAP7_75t_L g179 ( .A(n_154), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_156), .B(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g243 ( .A(n_156), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_156), .A2(n_220), .B(n_534), .C(n_535), .Y(n_533) );
OAI22xp33_ASAP7_75t_L g590 ( .A1(n_156), .A2(n_179), .B1(n_591), .B2(n_592), .Y(n_590) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_157), .B(n_495), .Y(n_494) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g248 ( .A(n_159), .Y(n_248) );
INVx1_ASAP7_75t_L g505 ( .A(n_159), .Y(n_505) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_162), .A2(n_204), .B(n_205), .Y(n_203) );
INVx2_ASAP7_75t_L g222 ( .A(n_162), .Y(n_222) );
INVx1_ASAP7_75t_L g225 ( .A(n_162), .Y(n_225) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_162), .A2(n_489), .B(n_496), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_162), .A2(n_256), .B(n_531), .C(n_532), .Y(n_530) );
AND2x2_ASAP7_75t_SL g162 ( .A(n_163), .B(n_164), .Y(n_162) );
AND2x2_ASAP7_75t_L g173 ( .A(n_163), .B(n_164), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
AND2x2_ASAP7_75t_L g445 ( .A(n_168), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g168 ( .A(n_169), .Y(n_168) );
OR2x2_ASAP7_75t_L g308 ( .A(n_169), .B(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_186), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_170), .B(n_289), .Y(n_288) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_170), .Y(n_301) );
INVx3_ASAP7_75t_L g316 ( .A(n_170), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_170), .B(n_186), .Y(n_340) );
OR2x2_ASAP7_75t_L g349 ( .A(n_170), .B(n_292), .Y(n_349) );
AND2x2_ASAP7_75t_L g353 ( .A(n_170), .B(n_313), .Y(n_353) );
AND2x2_ASAP7_75t_L g359 ( .A(n_170), .B(n_360), .Y(n_359) );
INVxp67_ASAP7_75t_L g396 ( .A(n_170), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_170), .B(n_253), .Y(n_410) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_174), .B(n_183), .Y(n_170) );
OA21x2_ASAP7_75t_L g498 ( .A1(n_171), .A2(n_499), .B(n_506), .Y(n_498) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_171), .A2(n_521), .B(n_527), .Y(n_520) );
OA21x2_ASAP7_75t_L g549 ( .A1(n_171), .A2(n_550), .B(n_557), .Y(n_549) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx4_ASAP7_75t_L g185 ( .A(n_172), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_172), .A2(n_189), .B(n_190), .Y(n_188) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g263 ( .A(n_173), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_178), .A2(n_231), .B(n_232), .C(n_233), .Y(n_230) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_179), .B(n_504), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_179), .B(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g220 ( .A(n_182), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_182), .B(n_590), .Y(n_589) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_184), .A2(n_239), .B(n_249), .Y(n_238) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_185), .B(n_210), .Y(n_209) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_185), .A2(n_228), .B(n_236), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_185), .B(n_237), .Y(n_236) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_185), .A2(n_254), .B(n_261), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_185), .B(n_518), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_185), .B(n_537), .Y(n_536) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_185), .A2(n_541), .B(n_547), .Y(n_540) );
OR2x2_ASAP7_75t_L g302 ( .A(n_186), .B(n_253), .Y(n_302) );
AND2x2_ASAP7_75t_L g313 ( .A(n_186), .B(n_289), .Y(n_313) );
AND2x2_ASAP7_75t_L g325 ( .A(n_186), .B(n_316), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_186), .B(n_253), .Y(n_348) );
INVx1_ASAP7_75t_SL g360 ( .A(n_186), .Y(n_360) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g252 ( .A(n_187), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_187), .B(n_292), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_194), .B(n_195), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_195), .A2(n_259), .B(n_260), .Y(n_258) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_211), .Y(n_200) );
AND2x2_ASAP7_75t_L g273 ( .A(n_201), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_201), .B(n_226), .Y(n_277) );
AND2x2_ASAP7_75t_L g280 ( .A(n_201), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_201), .B(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g305 ( .A(n_201), .B(n_296), .Y(n_305) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_201), .Y(n_324) );
AND2x2_ASAP7_75t_L g345 ( .A(n_201), .B(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g355 ( .A(n_201), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g401 ( .A(n_201), .B(n_284), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_201), .B(n_307), .Y(n_428) );
INVx5_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
BUFx2_ASAP7_75t_L g298 ( .A(n_202), .Y(n_298) );
AND2x2_ASAP7_75t_L g364 ( .A(n_202), .B(n_296), .Y(n_364) );
AND2x2_ASAP7_75t_L g448 ( .A(n_202), .B(n_316), .Y(n_448) );
OR2x6_ASAP7_75t_L g202 ( .A(n_203), .B(n_209), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_211), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g437 ( .A(n_211), .Y(n_437) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_226), .Y(n_211) );
AND2x2_ASAP7_75t_L g267 ( .A(n_212), .B(n_268), .Y(n_267) );
AND2x4_ASAP7_75t_L g276 ( .A(n_212), .B(n_274), .Y(n_276) );
INVx5_ASAP7_75t_L g284 ( .A(n_212), .Y(n_284) );
AND2x2_ASAP7_75t_L g307 ( .A(n_212), .B(n_238), .Y(n_307) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_212), .Y(n_344) );
OR2x6_ASAP7_75t_L g212 ( .A(n_213), .B(n_223), .Y(n_212) );
AOI21xp5_ASAP7_75t_SL g213 ( .A1(n_214), .A2(n_216), .B(n_221), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_220), .Y(n_217) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_222), .B(n_548), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_225), .A2(n_510), .B(n_517), .Y(n_509) );
INVx1_ASAP7_75t_L g385 ( .A(n_226), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_226), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g418 ( .A(n_226), .B(n_284), .Y(n_418) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_226), .A2(n_341), .B(n_448), .C(n_449), .Y(n_447) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_238), .Y(n_226) );
BUFx2_ASAP7_75t_L g268 ( .A(n_227), .Y(n_268) );
INVx2_ASAP7_75t_L g272 ( .A(n_227), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_235), .Y(n_228) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx3_ASAP7_75t_L g556 ( .A(n_234), .Y(n_556) );
INVx2_ASAP7_75t_L g274 ( .A(n_238), .Y(n_274) );
AND2x2_ASAP7_75t_L g281 ( .A(n_238), .B(n_272), .Y(n_281) );
AND2x2_ASAP7_75t_L g372 ( .A(n_238), .B(n_284), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_246), .B(n_555), .Y(n_554) );
INVx4_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g493 ( .A(n_247), .Y(n_493) );
INVx2_ASAP7_75t_L g516 ( .A(n_248), .Y(n_516) );
AOI211x1_ASAP7_75t_SL g250 ( .A1(n_251), .A2(n_265), .B(n_278), .C(n_303), .Y(n_250) );
INVx1_ASAP7_75t_L g369 ( .A(n_251), .Y(n_369) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_264), .Y(n_251) );
INVx5_ASAP7_75t_SL g289 ( .A(n_253), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_253), .B(n_359), .Y(n_358) );
AOI311xp33_ASAP7_75t_L g377 ( .A1(n_253), .A2(n_378), .A3(n_380), .B(n_381), .C(n_387), .Y(n_377) );
A2O1A1Ixp33_ASAP7_75t_L g412 ( .A1(n_253), .A2(n_325), .B(n_413), .C(n_416), .Y(n_412) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_257), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_256), .A2(n_511), .B(n_512), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g541 ( .A1(n_256), .A2(n_542), .B(n_543), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g584 ( .A(n_263), .Y(n_584) );
INVxp67_ASAP7_75t_L g332 ( .A(n_264), .Y(n_332) );
NAND4xp25_ASAP7_75t_SL g265 ( .A(n_266), .B(n_269), .C(n_275), .D(n_277), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_266), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g323 ( .A(n_267), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_273), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_270), .B(n_276), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_270), .B(n_283), .Y(n_403) );
BUFx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_271), .B(n_284), .Y(n_421) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g296 ( .A(n_272), .Y(n_296) );
INVxp67_ASAP7_75t_L g331 ( .A(n_273), .Y(n_331) );
AND2x4_ASAP7_75t_L g283 ( .A(n_274), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g357 ( .A(n_274), .B(n_296), .Y(n_357) );
INVx1_ASAP7_75t_L g384 ( .A(n_274), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_274), .B(n_371), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_275), .B(n_345), .Y(n_365) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_276), .B(n_298), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_276), .B(n_345), .Y(n_444) );
INVx1_ASAP7_75t_L g455 ( .A(n_277), .Y(n_455) );
A2O1A1Ixp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_282), .B(n_285), .C(n_293), .Y(n_278) );
INVx1_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g297 ( .A(n_281), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g335 ( .A(n_281), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g317 ( .A(n_282), .Y(n_317) );
AND2x2_ASAP7_75t_L g294 ( .A(n_283), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_283), .B(n_345), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_283), .B(n_364), .Y(n_388) );
OR2x2_ASAP7_75t_L g304 ( .A(n_284), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g336 ( .A(n_284), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_284), .B(n_296), .Y(n_351) );
AND2x2_ASAP7_75t_L g408 ( .A(n_284), .B(n_364), .Y(n_408) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_284), .Y(n_415) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_286), .A2(n_298), .B1(n_420), .B2(n_422), .C(n_425), .Y(n_419) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g309 ( .A(n_289), .B(n_292), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_289), .B(n_359), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_289), .B(n_316), .Y(n_424) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g409 ( .A(n_291), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g423 ( .A(n_291), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_292), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g320 ( .A(n_292), .B(n_313), .Y(n_320) );
AND2x2_ASAP7_75t_L g390 ( .A(n_292), .B(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_292), .B(n_339), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_292), .B(n_440), .Y(n_439) );
OAI21xp5_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_297), .B(n_299), .Y(n_293) );
INVx2_ASAP7_75t_L g326 ( .A(n_294), .Y(n_326) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g346 ( .A(n_296), .Y(n_346) );
OR2x2_ASAP7_75t_L g350 ( .A(n_298), .B(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g453 ( .A(n_298), .B(n_421), .Y(n_453) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AOI21xp33_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_306), .B(n_308), .Y(n_303) );
INVx1_ASAP7_75t_L g457 ( .A(n_304), .Y(n_457) );
INVx2_ASAP7_75t_SL g371 ( .A(n_305), .Y(n_371) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
A2O1A1Ixp33_ASAP7_75t_L g452 ( .A1(n_308), .A2(n_389), .B(n_453), .C(n_454), .Y(n_452) );
OAI322xp33_ASAP7_75t_SL g321 ( .A1(n_309), .A2(n_322), .A3(n_325), .B1(n_326), .B2(n_327), .C1(n_329), .C2(n_332), .Y(n_321) );
INVx2_ASAP7_75t_L g341 ( .A(n_309), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_317), .B1(n_318), .B2(n_320), .C(n_321), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OAI22xp33_ASAP7_75t_SL g387 ( .A1(n_312), .A2(n_388), .B1(n_389), .B2(n_392), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_313), .B(n_316), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_313), .B(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g386 ( .A(n_315), .B(n_348), .Y(n_386) );
INVx1_ASAP7_75t_L g376 ( .A(n_316), .Y(n_376) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_320), .A2(n_430), .B(n_432), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g354 ( .A1(n_322), .A2(n_355), .B(n_358), .Y(n_354) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NOR2xp67_ASAP7_75t_SL g383 ( .A(n_324), .B(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_324), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g440 ( .A(n_325), .Y(n_440) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND4xp25_ASAP7_75t_L g333 ( .A(n_334), .B(n_361), .C(n_377), .D(n_393), .Y(n_333) );
AOI211xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_337), .B(n_342), .C(n_354), .Y(n_334) );
INVx1_ASAP7_75t_L g426 ( .A(n_335), .Y(n_426) );
AND2x2_ASAP7_75t_L g374 ( .A(n_336), .B(n_357), .Y(n_374) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_341), .B(n_376), .Y(n_375) );
OAI22xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_347), .B1(n_350), .B2(n_352), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_344), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g392 ( .A(n_345), .Y(n_392) );
O2A1O1Ixp33_ASAP7_75t_L g406 ( .A1(n_345), .A2(n_384), .B(n_407), .C(n_409), .Y(n_406) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g391 ( .A(n_348), .Y(n_391) );
INVx1_ASAP7_75t_L g451 ( .A(n_349), .Y(n_451) );
NAND2xp33_ASAP7_75t_SL g441 ( .A(n_350), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g380 ( .A(n_359), .Y(n_380) );
O2A1O1Ixp33_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B(n_366), .C(n_368), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B1(n_373), .B2(n_375), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_371), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_376), .B(n_397), .Y(n_459) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI21xp33_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_385), .B(n_386), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_399), .B1(n_402), .B2(n_404), .C(n_406), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_409), .A2(n_426), .B1(n_427), .B2(n_428), .Y(n_425) );
NAND3xp33_ASAP7_75t_SL g411 ( .A(n_412), .B(n_419), .C(n_429), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
CKINVDCx16_ASAP7_75t_R g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI211xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_437), .B(n_438), .C(n_447), .Y(n_435) );
INVx1_ASAP7_75t_L g456 ( .A(n_436), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_441), .B1(n_443), .B2(n_445), .Y(n_438) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B1(n_457), .B2(n_458), .Y(n_454) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g468 ( .A(n_463), .Y(n_468) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND3xp33_ASAP7_75t_L g469 ( .A(n_467), .B(n_470), .C(n_755), .Y(n_469) );
XNOR2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_481), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_474), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_680), .Y(n_483) );
NAND5xp2_ASAP7_75t_L g484 ( .A(n_485), .B(n_595), .C(n_627), .D(n_644), .E(n_667), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_528), .B1(n_558), .B2(n_562), .C(n_566), .Y(n_485) );
INVx1_ASAP7_75t_L g707 ( .A(n_486), .Y(n_707) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_507), .Y(n_486) );
AND3x2_ASAP7_75t_L g682 ( .A(n_487), .B(n_509), .C(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_497), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_488), .B(n_564), .Y(n_563) );
BUFx3_ASAP7_75t_L g573 ( .A(n_488), .Y(n_573) );
AND2x2_ASAP7_75t_L g577 ( .A(n_488), .B(n_519), .Y(n_577) );
INVx2_ASAP7_75t_L g604 ( .A(n_488), .Y(n_604) );
OR2x2_ASAP7_75t_L g615 ( .A(n_488), .B(n_520), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_488), .B(n_508), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_488), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g694 ( .A(n_488), .B(n_520), .Y(n_694) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_497), .Y(n_576) );
AND2x2_ASAP7_75t_L g635 ( .A(n_497), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_497), .B(n_508), .Y(n_654) );
INVx1_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g565 ( .A(n_498), .B(n_508), .Y(n_565) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_498), .Y(n_572) );
AND2x2_ASAP7_75t_L g621 ( .A(n_498), .B(n_520), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g646 ( .A(n_498), .B(n_507), .C(n_604), .Y(n_646) );
AND2x2_ASAP7_75t_L g711 ( .A(n_498), .B(n_509), .Y(n_711) );
AND2x2_ASAP7_75t_L g745 ( .A(n_498), .B(n_508), .Y(n_745) );
INVxp67_ASAP7_75t_L g574 ( .A(n_507), .Y(n_574) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_519), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_508), .B(n_604), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_508), .B(n_635), .Y(n_643) );
AND2x2_ASAP7_75t_L g693 ( .A(n_508), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g721 ( .A(n_508), .Y(n_721) );
INVx4_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g628 ( .A(n_509), .B(n_621), .Y(n_628) );
BUFx3_ASAP7_75t_L g660 ( .A(n_509), .Y(n_660) );
INVx2_ASAP7_75t_L g636 ( .A(n_519), .Y(n_636) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_520), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_528), .A2(n_696), .B1(n_698), .B2(n_699), .Y(n_695) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_538), .Y(n_528) );
AND2x2_ASAP7_75t_L g558 ( .A(n_529), .B(n_559), .Y(n_558) );
INVx3_ASAP7_75t_SL g569 ( .A(n_529), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_529), .B(n_599), .Y(n_631) );
OR2x2_ASAP7_75t_L g650 ( .A(n_529), .B(n_539), .Y(n_650) );
AND2x2_ASAP7_75t_L g655 ( .A(n_529), .B(n_607), .Y(n_655) );
AND2x2_ASAP7_75t_L g658 ( .A(n_529), .B(n_600), .Y(n_658) );
AND2x2_ASAP7_75t_L g670 ( .A(n_529), .B(n_549), .Y(n_670) );
AND2x2_ASAP7_75t_L g686 ( .A(n_529), .B(n_540), .Y(n_686) );
AND2x4_ASAP7_75t_L g689 ( .A(n_529), .B(n_560), .Y(n_689) );
OR2x2_ASAP7_75t_L g706 ( .A(n_529), .B(n_642), .Y(n_706) );
OR2x2_ASAP7_75t_L g737 ( .A(n_529), .B(n_582), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g739 ( .A(n_529), .B(n_665), .Y(n_739) );
OR2x6_ASAP7_75t_L g529 ( .A(n_530), .B(n_536), .Y(n_529) );
AND2x2_ASAP7_75t_L g613 ( .A(n_538), .B(n_580), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_538), .B(n_600), .Y(n_732) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_549), .Y(n_538) );
AND2x2_ASAP7_75t_L g568 ( .A(n_539), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g599 ( .A(n_539), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g607 ( .A(n_539), .B(n_582), .Y(n_607) );
AND2x2_ASAP7_75t_L g625 ( .A(n_539), .B(n_560), .Y(n_625) );
OR2x2_ASAP7_75t_L g642 ( .A(n_539), .B(n_600), .Y(n_642) );
INVx2_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
BUFx2_ASAP7_75t_L g561 ( .A(n_540), .Y(n_561) );
AND2x2_ASAP7_75t_L g665 ( .A(n_540), .B(n_549), .Y(n_665) );
INVx2_ASAP7_75t_L g560 ( .A(n_549), .Y(n_560) );
INVx1_ASAP7_75t_L g677 ( .A(n_549), .Y(n_677) );
AND2x2_ASAP7_75t_L g727 ( .A(n_549), .B(n_569), .Y(n_727) );
AND2x2_ASAP7_75t_L g579 ( .A(n_559), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g611 ( .A(n_559), .B(n_569), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_559), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
AND2x2_ASAP7_75t_L g598 ( .A(n_560), .B(n_569), .Y(n_598) );
OR2x2_ASAP7_75t_L g714 ( .A(n_561), .B(n_688), .Y(n_714) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_564), .B(n_694), .Y(n_700) );
INVx2_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
OAI32xp33_ASAP7_75t_L g656 ( .A1(n_565), .A2(n_657), .A3(n_659), .B1(n_661), .B2(n_662), .Y(n_656) );
OR2x2_ASAP7_75t_L g673 ( .A(n_565), .B(n_615), .Y(n_673) );
OAI21xp33_ASAP7_75t_SL g698 ( .A1(n_565), .A2(n_575), .B(n_603), .Y(n_698) );
OAI22xp33_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_570), .B1(n_575), .B2(n_578), .Y(n_566) );
INVxp33_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_568), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_569), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g624 ( .A(n_569), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g724 ( .A(n_569), .B(n_665), .Y(n_724) );
OR2x2_ASAP7_75t_L g748 ( .A(n_569), .B(n_642), .Y(n_748) );
AOI21xp33_ASAP7_75t_L g731 ( .A1(n_570), .A2(n_630), .B(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_574), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
INVx1_ASAP7_75t_L g608 ( .A(n_572), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_572), .B(n_577), .Y(n_626) );
AND2x2_ASAP7_75t_L g648 ( .A(n_573), .B(n_621), .Y(n_648) );
INVx1_ASAP7_75t_L g661 ( .A(n_573), .Y(n_661) );
OR2x2_ASAP7_75t_L g666 ( .A(n_573), .B(n_600), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_576), .B(n_615), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g596 ( .A1(n_577), .A2(n_597), .B1(n_602), .B2(n_606), .Y(n_596) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_580), .A2(n_639), .B1(n_646), .B2(n_647), .Y(n_645) );
AND2x2_ASAP7_75t_L g723 ( .A(n_580), .B(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_582), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g742 ( .A(n_582), .B(n_625), .Y(n_742) );
AO21x2_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_585), .B(n_593), .Y(n_582) );
INVx1_ASAP7_75t_L g601 ( .A(n_583), .Y(n_601) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OA21x2_ASAP7_75t_L g600 ( .A1(n_586), .A2(n_594), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_608), .B1(n_609), .B2(n_614), .C(n_616), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_598), .B(n_600), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_598), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g617 ( .A(n_599), .Y(n_617) );
O2A1O1Ixp33_ASAP7_75t_L g704 ( .A1(n_599), .A2(n_705), .B(n_706), .C(n_707), .Y(n_704) );
AND2x2_ASAP7_75t_L g709 ( .A(n_599), .B(n_689), .Y(n_709) );
O2A1O1Ixp33_ASAP7_75t_SL g747 ( .A1(n_599), .A2(n_688), .B(n_748), .C(n_749), .Y(n_747) );
BUFx3_ASAP7_75t_L g639 ( .A(n_600), .Y(n_639) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_603), .B(n_660), .Y(n_703) );
AOI211xp5_ASAP7_75t_L g722 ( .A1(n_603), .A2(n_723), .B(n_725), .C(n_731), .Y(n_722) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVxp67_ASAP7_75t_L g683 ( .A(n_605), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_607), .B(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_610), .B(n_612), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
AOI211xp5_ASAP7_75t_L g627 ( .A1(n_611), .A2(n_628), .B(n_629), .C(n_637), .Y(n_627) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g712 ( .A(n_615), .Y(n_712) );
OR2x2_ASAP7_75t_L g729 ( .A(n_615), .B(n_659), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B1(n_623), .B2(n_626), .Y(n_616) );
OAI22xp33_ASAP7_75t_L g629 ( .A1(n_618), .A2(n_630), .B1(n_631), .B2(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
OR2x2_ASAP7_75t_L g716 ( .A(n_620), .B(n_660), .Y(n_716) );
INVx1_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g671 ( .A(n_621), .B(n_661), .Y(n_671) );
INVx1_ASAP7_75t_L g679 ( .A(n_622), .Y(n_679) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_625), .B(n_639), .Y(n_687) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_635), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g744 ( .A(n_636), .Y(n_744) );
AOI21xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .B(n_643), .Y(n_637) );
INVx1_ASAP7_75t_L g674 ( .A(n_638), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_639), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_639), .B(n_670), .Y(n_669) );
NAND2x1p5_ASAP7_75t_L g690 ( .A(n_639), .B(n_665), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_639), .B(n_686), .Y(n_697) );
OAI211xp5_ASAP7_75t_L g701 ( .A1(n_639), .A2(n_649), .B(n_689), .C(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
AOI221xp5_ASAP7_75t_SL g644 ( .A1(n_645), .A2(n_649), .B1(n_651), .B2(n_655), .C(n_656), .Y(n_644) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVxp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_653), .B(n_661), .Y(n_735) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g746 ( .A1(n_655), .A2(n_670), .B(n_672), .C(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_658), .B(n_665), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g749 ( .A(n_659), .B(n_712), .Y(n_749) );
CKINVDCx16_ASAP7_75t_R g659 ( .A(n_660), .Y(n_659) );
INVxp33_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
AOI21xp33_ASAP7_75t_SL g675 ( .A1(n_664), .A2(n_676), .B(n_678), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_664), .B(n_737), .Y(n_736) );
INVx2_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_665), .B(n_719), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_671), .B1(n_672), .B2(n_674), .C(n_675), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_671), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g705 ( .A(n_677), .Y(n_705) );
NAND5xp2_ASAP7_75t_L g680 ( .A(n_681), .B(n_708), .C(n_722), .D(n_733), .E(n_746), .Y(n_680) );
AOI211xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_684), .B(n_691), .C(n_704), .Y(n_681) );
INVx2_ASAP7_75t_SL g728 ( .A(n_682), .Y(n_728) );
NAND4xp25_ASAP7_75t_SL g684 ( .A(n_685), .B(n_687), .C(n_688), .D(n_690), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx3_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI211xp5_ASAP7_75t_SL g691 ( .A1(n_690), .A2(n_692), .B(n_695), .C(n_701), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_693), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g733 ( .A1(n_693), .A2(n_734), .B1(n_736), .B2(n_738), .C(n_740), .Y(n_733) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI221xp5_ASAP7_75t_SL g708 ( .A1(n_709), .A2(n_710), .B1(n_713), .B2(n_715), .C(n_717), .Y(n_708) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_716), .A2(n_739), .B1(n_741), .B2(n_743), .Y(n_740) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_725) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
endmodule