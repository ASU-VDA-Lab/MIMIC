module fake_jpeg_10862_n_88 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_10),
.B(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_39),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_36),
.B1(n_39),
.B2(n_32),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_36),
.A2(n_13),
.B1(n_27),
.B2(n_25),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_42),
.B1(n_32),
.B2(n_31),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_34),
.B(n_37),
.C(n_29),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_46),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_2),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_62)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_3),
.Y(n_61)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_6),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_6),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_58),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_33),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_43),
.B1(n_34),
.B2(n_5),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_50),
.B1(n_48),
.B2(n_8),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_64),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_50),
.B1(n_48),
.B2(n_7),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_15),
.C(n_21),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_12),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_4),
.Y(n_64)
);

NOR2x1_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_8),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_62),
.B1(n_63),
.B2(n_60),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_71),
.Y(n_78)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_16),
.B1(n_17),
.B2(n_20),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_28),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_80),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_68),
.B1(n_73),
.B2(n_69),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_73),
.C(n_74),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_76),
.Y(n_83)
);

NOR3xp33_ASAP7_75t_SL g84 ( 
.A(n_83),
.B(n_78),
.C(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_79),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_82),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_77),
.Y(n_88)
);


endmodule