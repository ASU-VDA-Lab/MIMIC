module fake_netlist_1_4845_n_501 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_501);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_501;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g71 ( .A(n_52), .Y(n_71) );
CKINVDCx16_ASAP7_75t_R g72 ( .A(n_37), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_64), .Y(n_73) );
BUFx6f_ASAP7_75t_L g74 ( .A(n_25), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_31), .Y(n_75) );
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_44), .Y(n_76) );
HB1xp67_ASAP7_75t_L g77 ( .A(n_27), .Y(n_77) );
CKINVDCx16_ASAP7_75t_R g78 ( .A(n_47), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_49), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_36), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_11), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_69), .Y(n_82) );
BUFx5_ASAP7_75t_L g83 ( .A(n_19), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_43), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_16), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_6), .Y(n_86) );
BUFx6f_ASAP7_75t_L g87 ( .A(n_21), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_59), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_20), .Y(n_89) );
BUFx10_ASAP7_75t_L g90 ( .A(n_10), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_56), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_10), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_55), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_51), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_3), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_62), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_34), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_38), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_45), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_66), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_24), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_48), .Y(n_102) );
INVxp33_ASAP7_75t_L g103 ( .A(n_61), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_65), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_70), .Y(n_105) );
AND2x2_ASAP7_75t_L g106 ( .A(n_103), .B(n_0), .Y(n_106) );
INVx3_ASAP7_75t_L g107 ( .A(n_74), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_77), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_77), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_71), .Y(n_110) );
INVx1_ASAP7_75t_SL g111 ( .A(n_81), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_72), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_73), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_74), .Y(n_114) );
BUFx8_ASAP7_75t_L g115 ( .A(n_83), .Y(n_115) );
AND2x4_ASAP7_75t_L g116 ( .A(n_85), .B(n_0), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_75), .Y(n_117) );
AND2x4_ASAP7_75t_L g118 ( .A(n_86), .B(n_1), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_78), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_103), .B(n_1), .Y(n_120) );
AND2x4_ASAP7_75t_L g121 ( .A(n_92), .B(n_2), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_83), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_79), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_74), .Y(n_124) );
INVxp67_ASAP7_75t_L g125 ( .A(n_90), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_80), .Y(n_126) );
AND2x6_ASAP7_75t_L g127 ( .A(n_82), .B(n_29), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_83), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_83), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_108), .B(n_84), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_122), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_122), .Y(n_132) );
BUFx3_ASAP7_75t_L g133 ( .A(n_115), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_122), .Y(n_134) );
BUFx3_ASAP7_75t_L g135 ( .A(n_115), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_108), .B(n_76), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_109), .B(n_76), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_114), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_109), .B(n_90), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_128), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_114), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_128), .Y(n_142) );
NAND2x1p5_ASAP7_75t_L g143 ( .A(n_116), .B(n_105), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_119), .B(n_104), .Y(n_144) );
BUFx6f_ASAP7_75t_SL g145 ( .A(n_127), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_119), .B(n_102), .Y(n_146) );
INVx4_ASAP7_75t_L g147 ( .A(n_127), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_128), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_116), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_129), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_125), .B(n_101), .Y(n_151) );
AND2x6_ASAP7_75t_L g152 ( .A(n_116), .B(n_100), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_129), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_114), .Y(n_154) );
NAND2xp33_ASAP7_75t_R g155 ( .A(n_112), .B(n_99), .Y(n_155) );
AOI22xp5_ASAP7_75t_L g156 ( .A1(n_139), .A2(n_146), .B1(n_144), .B2(n_152), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_136), .B(n_111), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_135), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_139), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
INVxp67_ASAP7_75t_L g161 ( .A(n_155), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_135), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_152), .B(n_116), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g165 ( .A1(n_131), .A2(n_127), .B(n_129), .Y(n_165) );
OR2x2_ASAP7_75t_L g166 ( .A(n_137), .B(n_106), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_152), .A2(n_106), .B1(n_120), .B2(n_118), .Y(n_167) );
INVx2_ASAP7_75t_SL g168 ( .A(n_133), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_130), .B(n_115), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_149), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_143), .B(n_115), .Y(n_172) );
INVx5_ASAP7_75t_L g173 ( .A(n_152), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_133), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_143), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_149), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_149), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_142), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_142), .Y(n_181) );
INVx1_ASAP7_75t_SL g182 ( .A(n_152), .Y(n_182) );
BUFx2_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
BUFx4f_ASAP7_75t_L g184 ( .A(n_131), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_132), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_151), .B(n_110), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_132), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_134), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_134), .Y(n_189) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_171), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_175), .B(n_118), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_189), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_158), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_189), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_185), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_178), .Y(n_196) );
BUFx2_ASAP7_75t_L g197 ( .A(n_159), .Y(n_197) );
NOR2x1_ASAP7_75t_L g198 ( .A(n_172), .B(n_147), .Y(n_198) );
BUFx12f_ASAP7_75t_L g199 ( .A(n_164), .Y(n_199) );
BUFx10_ASAP7_75t_L g200 ( .A(n_164), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_179), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_178), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_159), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_185), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_162), .Y(n_205) );
BUFx2_ASAP7_75t_L g206 ( .A(n_158), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_160), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_179), .Y(n_208) );
INVx5_ASAP7_75t_L g209 ( .A(n_160), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_162), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_160), .Y(n_211) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_165), .A2(n_97), .B(n_88), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_160), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_170), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_164), .B(n_118), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_180), .B(n_118), .Y(n_216) );
INVx2_ASAP7_75t_SL g217 ( .A(n_160), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_181), .Y(n_218) );
NAND3xp33_ASAP7_75t_L g219 ( .A(n_156), .B(n_121), .C(n_113), .Y(n_219) );
BUFx4f_ASAP7_75t_L g220 ( .A(n_163), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_170), .A2(n_147), .B(n_153), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_196), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_215), .A2(n_157), .B1(n_166), .B2(n_186), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_190), .B(n_166), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_215), .A2(n_167), .B1(n_161), .B2(n_176), .Y(n_225) );
OR2x2_ASAP7_75t_L g226 ( .A(n_197), .B(n_187), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_190), .B(n_173), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_219), .A2(n_184), .B1(n_188), .B2(n_169), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_215), .A2(n_176), .B1(n_95), .B2(n_177), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_195), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_192), .B(n_184), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_197), .B(n_184), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_196), .Y(n_233) );
OAI22xp33_ASAP7_75t_L g234 ( .A1(n_203), .A2(n_182), .B1(n_173), .B2(n_168), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_195), .Y(n_235) );
BUFx2_ASAP7_75t_R g236 ( .A(n_212), .Y(n_236) );
BUFx2_ASAP7_75t_L g237 ( .A(n_199), .Y(n_237) );
OAI222xp33_ASAP7_75t_L g238 ( .A1(n_204), .A2(n_121), .B1(n_99), .B2(n_110), .C1(n_113), .C2(n_117), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_219), .A2(n_121), .B1(n_117), .B2(n_126), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_199), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_204), .Y(n_241) );
AOI22xp33_ASAP7_75t_SL g242 ( .A1(n_199), .A2(n_168), .B1(n_127), .B2(n_173), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_221), .A2(n_183), .B(n_126), .C(n_123), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_200), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_215), .A2(n_147), .B1(n_173), .B2(n_127), .Y(n_245) );
AOI221xp5_ASAP7_75t_L g246 ( .A1(n_191), .A2(n_123), .B1(n_140), .B2(n_148), .C(n_150), .Y(n_246) );
OAI21xp5_ASAP7_75t_SL g247 ( .A1(n_191), .A2(n_163), .B(n_96), .Y(n_247) );
BUFx2_ASAP7_75t_L g248 ( .A(n_222), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_224), .B(n_192), .Y(n_249) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_243), .A2(n_221), .B(n_194), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_223), .A2(n_192), .B1(n_194), .B2(n_191), .Y(n_251) );
AOI221xp5_ASAP7_75t_L g252 ( .A1(n_224), .A2(n_191), .B1(n_205), .B2(n_214), .C(n_210), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_247), .A2(n_194), .B1(n_191), .B2(n_218), .Y(n_253) );
INVx3_ASAP7_75t_L g254 ( .A(n_244), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_222), .Y(n_255) );
AOI222xp33_ASAP7_75t_L g256 ( .A1(n_229), .A2(n_205), .B1(n_214), .B2(n_210), .C1(n_216), .C2(n_127), .Y(n_256) );
NOR2x1_ASAP7_75t_SL g257 ( .A(n_247), .B(n_209), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_230), .B(n_196), .Y(n_258) );
OAI22xp33_ASAP7_75t_L g259 ( .A1(n_226), .A2(n_202), .B1(n_218), .B2(n_206), .Y(n_259) );
INVx3_ASAP7_75t_L g260 ( .A(n_244), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_230), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_235), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_244), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_244), .B(n_209), .Y(n_264) );
AOI221xp5_ASAP7_75t_L g265 ( .A1(n_239), .A2(n_216), .B1(n_153), .B2(n_212), .C(n_89), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_237), .Y(n_266) );
NOR2x1p5_ASAP7_75t_L g267 ( .A(n_266), .B(n_235), .Y(n_267) );
AOI221xp5_ASAP7_75t_L g268 ( .A1(n_252), .A2(n_238), .B1(n_232), .B2(n_225), .C(n_241), .Y(n_268) );
OAI31xp33_ASAP7_75t_L g269 ( .A1(n_259), .A2(n_228), .A3(n_237), .B(n_231), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_249), .B(n_222), .Y(n_270) );
OA21x2_ASAP7_75t_L g271 ( .A1(n_250), .A2(n_228), .B(n_241), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_249), .B(n_233), .Y(n_272) );
OA222x2_ASAP7_75t_L g273 ( .A1(n_266), .A2(n_236), .B1(n_233), .B2(n_193), .C1(n_211), .C2(n_212), .Y(n_273) );
NAND3xp33_ASAP7_75t_L g274 ( .A(n_265), .B(n_233), .C(n_114), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_261), .Y(n_275) );
OAI221xp5_ASAP7_75t_SL g276 ( .A1(n_256), .A2(n_246), .B1(n_93), .B2(n_98), .C(n_91), .Y(n_276) );
AOI31xp33_ASAP7_75t_L g277 ( .A1(n_253), .A2(n_240), .A3(n_242), .B(n_227), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_258), .B(n_231), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_255), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_255), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_248), .Y(n_281) );
NAND3xp33_ASAP7_75t_L g282 ( .A(n_256), .B(n_114), .C(n_87), .Y(n_282) );
AND2x4_ASAP7_75t_L g283 ( .A(n_248), .B(n_227), .Y(n_283) );
AOI221xp5_ASAP7_75t_L g284 ( .A1(n_251), .A2(n_216), .B1(n_94), .B2(n_234), .C(n_227), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_257), .B(n_227), .Y(n_285) );
OAI221xp5_ASAP7_75t_L g286 ( .A1(n_268), .A2(n_262), .B1(n_250), .B2(n_260), .C(n_254), .Y(n_286) );
INVx2_ASAP7_75t_SL g287 ( .A(n_267), .Y(n_287) );
OR2x2_ASAP7_75t_L g288 ( .A(n_272), .B(n_254), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_272), .B(n_254), .Y(n_289) );
NAND3xp33_ASAP7_75t_L g290 ( .A(n_269), .B(n_74), .C(n_87), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_279), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_281), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_278), .B(n_260), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_277), .B(n_264), .Y(n_294) );
INVxp67_ASAP7_75t_L g295 ( .A(n_270), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_270), .B(n_257), .Y(n_296) );
OAI221xp5_ASAP7_75t_L g297 ( .A1(n_269), .A2(n_260), .B1(n_263), .B2(n_245), .C(n_87), .Y(n_297) );
INVx4_ASAP7_75t_L g298 ( .A(n_285), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_282), .A2(n_264), .B1(n_263), .B2(n_127), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_275), .B(n_264), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_278), .B(n_263), .Y(n_301) );
AO21x2_ASAP7_75t_L g302 ( .A1(n_282), .A2(n_264), .B(n_181), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_275), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_267), .B(n_2), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_284), .A2(n_127), .B1(n_200), .B2(n_198), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_279), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_285), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_279), .B(n_83), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_280), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_280), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_280), .B(n_83), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_283), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_283), .Y(n_313) );
OAI22xp5_ASAP7_75t_SL g314 ( .A1(n_285), .A2(n_4), .B1(n_5), .B2(n_7), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_298), .B(n_271), .Y(n_315) );
OAI221xp5_ASAP7_75t_L g316 ( .A1(n_314), .A2(n_277), .B1(n_276), .B2(n_274), .C(n_271), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_303), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_292), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_292), .Y(n_319) );
NOR3xp33_ASAP7_75t_L g320 ( .A(n_304), .B(n_107), .C(n_124), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_295), .B(n_283), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_296), .B(n_283), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_298), .B(n_285), .Y(n_323) );
INVx4_ASAP7_75t_L g324 ( .A(n_298), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_300), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_296), .B(n_271), .Y(n_326) );
INVx1_ASAP7_75t_SL g327 ( .A(n_307), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_307), .B(n_271), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_306), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_307), .B(n_273), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_312), .B(n_273), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_287), .B(n_4), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_293), .B(n_5), .Y(n_333) );
NAND3xp33_ASAP7_75t_L g334 ( .A(n_290), .B(n_114), .C(n_107), .Y(n_334) );
NAND4xp25_ASAP7_75t_SL g335 ( .A(n_299), .B(n_297), .C(n_286), .D(n_301), .Y(n_335) );
OAI211xp5_ASAP7_75t_L g336 ( .A1(n_294), .A2(n_107), .B(n_124), .C(n_209), .Y(n_336) );
NOR3xp33_ASAP7_75t_SL g337 ( .A(n_294), .B(n_8), .C(n_9), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_287), .B(n_8), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_288), .B(n_9), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_291), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_308), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_309), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_313), .B(n_54), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_289), .B(n_11), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_310), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_310), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_308), .B(n_311), .Y(n_347) );
INVx2_ASAP7_75t_SL g348 ( .A(n_311), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_302), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_302), .B(n_12), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_305), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_298), .B(n_12), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_291), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_291), .Y(n_354) );
OAI33xp33_ASAP7_75t_L g355 ( .A1(n_314), .A2(n_13), .A3(n_14), .B1(n_15), .B2(n_16), .B3(n_17), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_318), .B(n_124), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_319), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_322), .B(n_14), .Y(n_358) );
NOR2xp67_ASAP7_75t_SL g359 ( .A(n_324), .B(n_209), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_317), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_323), .B(n_15), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_325), .B(n_17), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_329), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_347), .B(n_18), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_342), .Y(n_365) );
A2O1A1Ixp33_ASAP7_75t_L g366 ( .A1(n_337), .A2(n_220), .B(n_209), .C(n_211), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_352), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_323), .B(n_330), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_352), .B(n_22), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_323), .B(n_23), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_327), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_332), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_321), .B(n_326), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_324), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_346), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_316), .A2(n_220), .B1(n_209), .B2(n_207), .Y(n_376) );
INVx1_ASAP7_75t_SL g377 ( .A(n_324), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_344), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_331), .B(n_26), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_331), .B(n_207), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_340), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_330), .B(n_28), .Y(n_382) );
NAND2x1_ASAP7_75t_L g383 ( .A(n_315), .B(n_207), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_315), .B(n_30), .Y(n_384) );
INVxp67_ASAP7_75t_SL g385 ( .A(n_340), .Y(n_385) );
OAI22xp5_ASAP7_75t_SL g386 ( .A1(n_338), .A2(n_209), .B1(n_201), .B2(n_208), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_348), .B(n_32), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_345), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_341), .B(n_33), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_353), .B(n_207), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_354), .Y(n_391) );
XOR2x2_ASAP7_75t_L g392 ( .A(n_338), .B(n_35), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_354), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_339), .B(n_39), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_328), .B(n_40), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_333), .Y(n_396) );
OR2x6_ASAP7_75t_L g397 ( .A(n_336), .B(n_217), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_355), .B(n_41), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_368), .B(n_349), .Y(n_399) );
XNOR2x1_ASAP7_75t_L g400 ( .A(n_392), .B(n_351), .Y(n_400) );
OAI31xp33_ASAP7_75t_L g401 ( .A1(n_376), .A2(n_335), .A3(n_320), .B(n_350), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_360), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_372), .B(n_343), .Y(n_403) );
OAI21xp5_ASAP7_75t_SL g404 ( .A1(n_377), .A2(n_334), .B(n_343), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_363), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_365), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_373), .B(n_349), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_367), .B(n_343), .Y(n_408) );
INVxp67_ASAP7_75t_L g409 ( .A(n_371), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_396), .B(n_42), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_357), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_371), .B(n_46), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_378), .B(n_50), .Y(n_413) );
INVxp67_ASAP7_75t_SL g414 ( .A(n_385), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_375), .B(n_53), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_380), .B(n_57), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_356), .Y(n_417) );
O2A1O1Ixp33_ASAP7_75t_L g418 ( .A1(n_376), .A2(n_217), .B(n_201), .C(n_208), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_380), .B(n_383), .Y(n_419) );
INVx1_ASAP7_75t_SL g420 ( .A(n_377), .Y(n_420) );
BUFx2_ASAP7_75t_SL g421 ( .A(n_374), .Y(n_421) );
XNOR2xp5_ASAP7_75t_L g422 ( .A(n_361), .B(n_198), .Y(n_422) );
XNOR2xp5_ASAP7_75t_L g423 ( .A(n_382), .B(n_58), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_356), .Y(n_424) );
NAND2xp33_ASAP7_75t_SL g425 ( .A(n_359), .B(n_213), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_381), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_388), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_374), .B(n_209), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_391), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_393), .Y(n_430) );
CKINVDCx16_ASAP7_75t_R g431 ( .A(n_358), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_362), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_362), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_379), .B(n_60), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_395), .B(n_63), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_370), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_390), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_384), .B(n_67), .Y(n_438) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_384), .B(n_220), .Y(n_439) );
OAI31xp33_ASAP7_75t_SL g440 ( .A1(n_398), .A2(n_68), .A3(n_220), .B(n_200), .Y(n_440) );
XOR2xp5_ASAP7_75t_L g441 ( .A(n_364), .B(n_213), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_390), .B(n_138), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_387), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_389), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_369), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_394), .Y(n_446) );
AOI32xp33_ASAP7_75t_L g447 ( .A1(n_366), .A2(n_208), .A3(n_201), .B1(n_200), .B2(n_213), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_397), .B(n_141), .Y(n_448) );
INVxp67_ASAP7_75t_L g449 ( .A(n_386), .Y(n_449) );
XNOR2x1_ASAP7_75t_L g450 ( .A(n_397), .B(n_174), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_397), .Y(n_451) );
OAI31xp33_ASAP7_75t_SL g452 ( .A1(n_377), .A2(n_200), .A3(n_173), .B(n_145), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_373), .B(n_141), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_368), .B(n_154), .Y(n_454) );
XNOR2xp5_ASAP7_75t_L g455 ( .A(n_392), .B(n_145), .Y(n_455) );
OAI221xp5_ASAP7_75t_L g456 ( .A1(n_376), .A2(n_163), .B1(n_174), .B2(n_337), .C(n_377), .Y(n_456) );
OAI21xp33_ASAP7_75t_L g457 ( .A1(n_368), .A2(n_174), .B(n_330), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_371), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_357), .B(n_318), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_360), .Y(n_460) );
NOR2x1_ASAP7_75t_L g461 ( .A(n_456), .B(n_404), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_432), .A2(n_433), .B1(n_401), .B2(n_445), .C(n_460), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_456), .A2(n_409), .B(n_449), .C(n_428), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_406), .A2(n_405), .B1(n_402), .B2(n_411), .C(n_424), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_427), .Y(n_465) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_428), .A2(n_409), .B(n_423), .Y(n_466) );
NAND3xp33_ASAP7_75t_SL g467 ( .A(n_420), .B(n_447), .C(n_425), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_414), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_457), .A2(n_451), .B1(n_403), .B2(n_436), .Y(n_469) );
NOR2x1_ASAP7_75t_L g470 ( .A(n_421), .B(n_413), .Y(n_470) );
NOR2x1_ASAP7_75t_SL g471 ( .A(n_458), .B(n_419), .Y(n_471) );
OAI22xp33_ASAP7_75t_L g472 ( .A1(n_414), .A2(n_431), .B1(n_439), .B2(n_446), .Y(n_472) );
OAI21xp5_ASAP7_75t_SL g473 ( .A1(n_440), .A2(n_452), .B(n_439), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_403), .A2(n_400), .B1(n_399), .B2(n_444), .Y(n_474) );
OAI211xp5_ASAP7_75t_SL g475 ( .A1(n_417), .A2(n_459), .B(n_407), .C(n_434), .Y(n_475) );
OAI211xp5_ASAP7_75t_L g476 ( .A1(n_425), .A2(n_441), .B(n_454), .C(n_408), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_427), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_471), .Y(n_478) );
NOR2x1_ASAP7_75t_L g479 ( .A(n_461), .B(n_438), .Y(n_479) );
OAI221xp5_ASAP7_75t_L g480 ( .A1(n_462), .A2(n_459), .B1(n_422), .B2(n_410), .C(n_412), .Y(n_480) );
AOI221xp5_ASAP7_75t_L g481 ( .A1(n_472), .A2(n_429), .B1(n_430), .B2(n_426), .C(n_437), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_468), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_466), .A2(n_450), .B1(n_443), .B2(n_418), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_465), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_477), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_463), .Y(n_486) );
NOR4xp25_ASAP7_75t_L g487 ( .A(n_486), .B(n_467), .C(n_466), .D(n_473), .Y(n_487) );
OAI222xp33_ASAP7_75t_L g488 ( .A1(n_479), .A2(n_474), .B1(n_470), .B2(n_469), .C1(n_453), .C2(n_476), .Y(n_488) );
NOR3xp33_ASAP7_75t_L g489 ( .A(n_483), .B(n_475), .C(n_464), .Y(n_489) );
INVxp67_ASAP7_75t_SL g490 ( .A(n_478), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_483), .B(n_481), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_490), .A2(n_480), .B1(n_485), .B2(n_482), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_489), .B(n_484), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_491), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_494), .A2(n_487), .B1(n_488), .B2(n_437), .Y(n_495) );
XNOR2x1_ASAP7_75t_L g496 ( .A(n_493), .B(n_455), .Y(n_496) );
XNOR2xp5_ASAP7_75t_L g497 ( .A(n_496), .B(n_492), .Y(n_497) );
OAI22xp5_ASAP7_75t_SL g498 ( .A1(n_495), .A2(n_435), .B1(n_416), .B2(n_415), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_497), .A2(n_448), .B(n_442), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_499), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_500), .A2(n_498), .B(n_448), .Y(n_501) );
endmodule