module fake_jpeg_14748_n_315 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_16),
.B1(n_32),
.B2(n_29),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_45),
.A2(n_51),
.B1(n_27),
.B2(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_32),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_63),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_16),
.B1(n_29),
.B2(n_33),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_22),
.Y(n_56)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_42),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_33),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_18),
.B(n_27),
.C(n_22),
.Y(n_61)
);

FAx1_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_18),
.CI(n_26),
.CON(n_71),
.SN(n_71)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_16),
.B1(n_29),
.B2(n_18),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_30),
.B1(n_39),
.B2(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_30),
.Y(n_64)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_26),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_30),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_18),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_61),
.Y(n_92)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_73),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_81),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_72),
.A2(n_59),
.B1(n_56),
.B2(n_28),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_53),
.B1(n_52),
.B2(n_58),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_79),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_82),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_42),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_36),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_90),
.Y(n_117)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_61),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_55),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_66),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_0),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_95),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_96),
.B(n_19),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_45),
.B1(n_44),
.B2(n_67),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_100),
.B1(n_106),
.B2(n_111),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_58),
.B1(n_39),
.B2(n_38),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_120),
.B1(n_123),
.B2(n_69),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_71),
.B1(n_92),
.B2(n_87),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_50),
.C(n_36),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_109),
.C(n_114),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_66),
.C(n_36),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_44),
.B1(n_39),
.B2(n_59),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_65),
.C(n_64),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_23),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_59),
.B1(n_42),
.B2(n_44),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_42),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_79),
.B(n_85),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_72),
.A2(n_57),
.B1(n_54),
.B2(n_31),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_57),
.B1(n_54),
.B2(n_31),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_57),
.B1(n_31),
.B2(n_20),
.Y(n_123)
);

AO22x1_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_94),
.B1(n_69),
.B2(n_70),
.Y(n_124)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

NOR2x1_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_94),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_125),
.A2(n_140),
.B(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_73),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_130),
.B(n_138),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_101),
.Y(n_131)
);

XNOR2x1_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_146),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_133),
.A2(n_135),
.B1(n_137),
.B2(n_119),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_112),
.A2(n_85),
.B1(n_80),
.B2(n_95),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_118),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_136),
.B(n_149),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_82),
.B1(n_78),
.B2(n_77),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_89),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

NAND2x1p5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_70),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_112),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_143),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_145),
.B1(n_123),
.B2(n_120),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_100),
.A2(n_31),
.B1(n_20),
.B2(n_28),
.Y(n_145)
);

OR2x4_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_17),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_93),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_97),
.B(n_93),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_154),
.B(n_158),
.Y(n_187)
);

CKINVDCx10_ASAP7_75t_R g157 ( 
.A(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_157),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_138),
.Y(n_158)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_164),
.B1(n_174),
.B2(n_105),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_110),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_166),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_143),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_118),
.B(n_116),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_169),
.A2(n_132),
.B(n_129),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_109),
.C(n_114),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_136),
.C(n_109),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_141),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_175),
.A2(n_169),
.B(n_173),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_134),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_179),
.C(n_191),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_151),
.A2(n_131),
.B1(n_125),
.B2(n_146),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_178),
.A2(n_181),
.B1(n_188),
.B2(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_161),
.A2(n_125),
.B1(n_144),
.B2(n_128),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_159),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_183),
.B(n_185),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_168),
.B(n_153),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_159),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_127),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_196),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_151),
.A2(n_133),
.B1(n_128),
.B2(n_137),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_190),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_107),
.C(n_149),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_124),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_195),
.C(n_199),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_99),
.C(n_124),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_124),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_160),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_198),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_160),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_115),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_152),
.B(n_103),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_166),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_177),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_180),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_205),
.B(n_219),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_208),
.B(n_213),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_175),
.A2(n_173),
.B(n_172),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_172),
.C(n_152),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_215),
.C(n_221),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_167),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_214),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_156),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_175),
.A2(n_167),
.B1(n_174),
.B2(n_153),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_217),
.A2(n_177),
.B1(n_196),
.B2(n_195),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_181),
.A2(n_154),
.B(n_157),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g220 ( 
.A(n_192),
.B(n_164),
.CI(n_150),
.CON(n_220),
.SN(n_220)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_220),
.B(n_189),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_98),
.C(n_102),
.Y(n_221)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_184),
.C(n_178),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_220),
.Y(n_233)
);

INVx11_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_216),
.Y(n_245)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_233),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_231),
.A2(n_206),
.B(n_223),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_217),
.A2(n_190),
.B1(n_186),
.B2(n_194),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_232),
.A2(n_235),
.B1(n_242),
.B2(n_243),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_182),
.B1(n_200),
.B2(n_98),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_239),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_121),
.C(n_113),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_240),
.C(n_212),
.Y(n_247)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_121),
.C(n_25),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_0),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_208),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_209),
.A2(n_24),
.B1(n_17),
.B2(n_20),
.Y(n_243)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_227),
.A2(n_216),
.B1(n_210),
.B2(n_219),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_246),
.A2(n_243),
.B1(n_2),
.B2(n_4),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_248),
.C(n_249),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_221),
.C(n_215),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_202),
.C(n_213),
.Y(n_249)
);

OAI321xp33_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_233),
.A3(n_236),
.B1(n_235),
.B2(n_234),
.C(n_225),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_202),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_259),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_220),
.B1(n_218),
.B2(n_222),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_222),
.C(n_20),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_255),
.C(n_241),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_25),
.C(n_19),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_234),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_19),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_15),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_260),
.B(n_0),
.Y(n_271)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_269),
.B(n_270),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_1),
.C(n_4),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_239),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_266),
.B(n_267),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_242),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_226),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_249),
.A2(n_236),
.B(n_226),
.Y(n_270)
);

OAI321xp33_ASAP7_75t_L g279 ( 
.A1(n_271),
.A2(n_272),
.A3(n_12),
.B1(n_13),
.B2(n_11),
.C(n_10),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_256),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_273),
.A2(n_246),
.B1(n_255),
.B2(n_254),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_1),
.C(n_2),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_4),
.C(n_5),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_6),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_247),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_279),
.B(n_281),
.Y(n_290)
);

NOR2xp67_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_256),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_5),
.C(n_6),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_263),
.A2(n_13),
.B(n_11),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_274),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_9),
.B(n_10),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_9),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_286),
.B(n_4),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_268),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_287),
.B(n_291),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_276),
.B(n_265),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_292),
.A2(n_277),
.B(n_284),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_9),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_294),
.Y(n_298)
);

OAI211xp5_ASAP7_75t_L g301 ( 
.A1(n_295),
.A2(n_290),
.B(n_291),
.C(n_296),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_296),
.Y(n_299)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_303),
.B(n_299),
.Y(n_307)
);

AOI31xp67_ASAP7_75t_L g303 ( 
.A1(n_288),
.A2(n_286),
.A3(n_10),
.B(n_8),
.Y(n_303)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_6),
.B(n_7),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_7),
.C(n_8),
.Y(n_306)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_306),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_308),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_301),
.A2(n_7),
.B(n_8),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_300),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_8),
.Y(n_310)
);

OA21x2_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_310),
.B(n_309),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_305),
.B(n_312),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_298),
.Y(n_315)
);


endmodule