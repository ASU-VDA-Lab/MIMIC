module fake_jpeg_24924_n_185 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_185);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_36),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_0),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_30),
.C(n_26),
.Y(n_51)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_17),
.Y(n_37)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_15),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_15),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_40)
);

NOR2x1_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_17),
.Y(n_41)
);

OR2x2_ASAP7_75t_SL g80 ( 
.A(n_41),
.B(n_49),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_23),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_51),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_32),
.A2(n_24),
.B1(n_29),
.B2(n_22),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_53),
.B1(n_38),
.B2(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_28),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_29),
.B1(n_28),
.B2(n_25),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_38),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_51),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_SL g91 ( 
.A(n_58),
.B(n_73),
.C(n_35),
.Y(n_91)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_63),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_33),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_26),
.C(n_23),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_65),
.Y(n_95)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_66),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_67),
.B(n_27),
.Y(n_98)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_70),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_72),
.Y(n_101)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_35),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_76),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_25),
.B(n_39),
.C(n_40),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_36),
.Y(n_93)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_34),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_78),
.B(n_79),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_36),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_45),
.B(n_18),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_82),
.B(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_27),
.Y(n_83)
);

INVxp33_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_105),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_SL g86 ( 
.A(n_80),
.B(n_25),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_89),
.B(n_65),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_91),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_79),
.A2(n_36),
.B(n_22),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_35),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_67),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_16),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_60),
.B(n_2),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_58),
.B(n_57),
.Y(n_118)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_78),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_124),
.C(n_125),
.Y(n_128)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_114),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_55),
.B1(n_62),
.B2(n_75),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_109),
.A2(n_121),
.B1(n_122),
.B2(n_104),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_110),
.A2(n_118),
.B(n_103),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_58),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_117),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_90),
.B(n_86),
.Y(n_129)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_115),
.B(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_57),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_123),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_68),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_57),
.B1(n_70),
.B2(n_71),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_93),
.A2(n_73),
.B1(n_66),
.B2(n_31),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_73),
.C(n_64),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_63),
.C(n_59),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_21),
.Y(n_126)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_141),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_90),
.B(n_98),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_136),
.B(n_142),
.Y(n_157)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_114),
.Y(n_134)
);

OAI322xp33_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_108),
.A3(n_21),
.B1(n_19),
.B2(n_20),
.C1(n_31),
.C2(n_14),
.Y(n_150)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_102),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_100),
.C(n_94),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_113),
.C(n_125),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_104),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_109),
.A2(n_94),
.B1(n_100),
.B2(n_96),
.Y(n_142)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

BUFx12_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_135),
.A2(n_117),
.B1(n_111),
.B2(n_124),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_151),
.C(n_156),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_19),
.B(n_131),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_108),
.C(n_92),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_152),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_142),
.A2(n_139),
.B1(n_136),
.B2(n_140),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_154),
.B(n_155),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_143),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_92),
.C(n_84),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_157),
.A2(n_132),
.B(n_129),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_161),
.B(n_146),
.Y(n_170)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_139),
.C(n_141),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_84),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_156),
.C(n_149),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_165),
.C(n_148),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_127),
.C(n_133),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_169),
.B(n_170),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_147),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_171),
.B(n_174),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_146),
.C(n_152),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_173),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_166),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_170),
.A2(n_160),
.B(n_161),
.Y(n_175)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_173),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_179),
.A2(n_181),
.B(n_7),
.Y(n_183)
);

AOI21x1_ASAP7_75t_SL g181 ( 
.A1(n_177),
.A2(n_4),
.B(n_6),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_178),
.C(n_8),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_183),
.B(n_181),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_184),
.B(n_7),
.Y(n_185)
);


endmodule