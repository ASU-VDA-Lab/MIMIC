module fake_jpeg_10578_n_313 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_28),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_17),
.B1(n_31),
.B2(n_24),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_37),
.B1(n_22),
.B2(n_30),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_17),
.B1(n_31),
.B2(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_51),
.B1(n_42),
.B2(n_28),
.Y(n_76)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_58),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_17),
.B1(n_31),
.B2(n_29),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_28),
.B1(n_33),
.B2(n_32),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_53),
.A2(n_33),
.B1(n_39),
.B2(n_35),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_31),
.B1(n_24),
.B2(n_21),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_70),
.B1(n_18),
.B2(n_26),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_66),
.B(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_27),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_69),
.Y(n_85)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_68),
.B(n_27),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_20),
.C(n_21),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_24),
.B1(n_21),
.B2(n_30),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_82),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_73),
.A2(n_80),
.B1(n_84),
.B2(n_57),
.Y(n_118)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_53),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_76),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_77),
.B(n_106),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_78),
.A2(n_105),
.B1(n_53),
.B2(n_63),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_39),
.B1(n_36),
.B2(n_45),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_86),
.B(n_53),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_18),
.B1(n_26),
.B2(n_25),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_62),
.A2(n_25),
.B1(n_22),
.B2(n_45),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_81),
.A2(n_95),
.B1(n_102),
.B2(n_104),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_62),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_39),
.B1(n_36),
.B2(n_45),
.Y(n_84)
);

OR2x2_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_23),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_41),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_41),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_91),
.Y(n_112)
);

INVx6_ASAP7_75t_SL g91 ( 
.A(n_48),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_28),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_86),
.B(n_96),
.C(n_88),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_56),
.A2(n_19),
.B1(n_28),
.B2(n_12),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_39),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_99),
.Y(n_131)
);

CKINVDCx6p67_ASAP7_75t_R g98 ( 
.A(n_61),
.Y(n_98)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_19),
.B1(n_12),
.B2(n_16),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_103),
.Y(n_123)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_49),
.B(n_16),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_114),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_109),
.A2(n_115),
.B(n_121),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_34),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_57),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_120),
.C(n_133),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_127),
.B1(n_83),
.B2(n_104),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_94),
.C(n_84),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_50),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_132),
.Y(n_142)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_9),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_125),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_97),
.A2(n_33),
.B1(n_35),
.B2(n_32),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_82),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_73),
.B(n_50),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_76),
.B(n_50),
.C(n_67),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_35),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_32),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_126),
.B(n_105),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_157),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_105),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_136),
.B(n_143),
.C(n_148),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_124),
.A2(n_99),
.B1(n_82),
.B2(n_83),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_139),
.A2(n_156),
.B1(n_158),
.B2(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_141),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_91),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_79),
.B(n_92),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_128),
.B(n_125),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_74),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_146),
.A2(n_150),
.B1(n_151),
.B2(n_165),
.Y(n_191)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_149),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_98),
.C(n_79),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_103),
.B1(n_101),
.B2(n_98),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_98),
.B1(n_33),
.B2(n_32),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_93),
.Y(n_154)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_93),
.Y(n_155)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_32),
.B1(n_72),
.B2(n_34),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_133),
.A2(n_72),
.B1(n_34),
.B2(n_2),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_108),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_160),
.A2(n_126),
.B(n_119),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_112),
.B(n_34),
.C(n_1),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_166),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_112),
.A2(n_34),
.B1(n_1),
.B2(n_2),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_14),
.Y(n_164)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_13),
.B1(n_9),
.B2(n_3),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_116),
.B(n_0),
.C(n_1),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_167),
.A2(n_192),
.B(n_194),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_107),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_169),
.B(n_172),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_116),
.B(n_109),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_171),
.A2(n_173),
.B(n_178),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_143),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_116),
.B(n_121),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_139),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_175),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_150),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_159),
.A2(n_121),
.B(n_107),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_121),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_181),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_114),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_119),
.Y(n_184)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_157),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_186),
.A2(n_197),
.B1(n_194),
.B2(n_168),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_188),
.A2(n_146),
.B1(n_144),
.B2(n_166),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_190),
.A2(n_158),
.B(n_163),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_141),
.A2(n_114),
.B(n_123),
.Y(n_192)
);

XNOR2x2_ASAP7_75t_SL g193 ( 
.A(n_142),
.B(n_111),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_193),
.A2(n_198),
.B(n_123),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_147),
.B(n_0),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_142),
.B(n_113),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_156),
.Y(n_209)
);

A2O1A1O1Ixp25_ASAP7_75t_L g198 ( 
.A1(n_159),
.A2(n_111),
.B(n_110),
.C(n_9),
.D(n_113),
.Y(n_198)
);

NOR2x1_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_160),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_199),
.A2(n_213),
.B(n_219),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_180),
.B(n_153),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_206),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_205),
.A2(n_113),
.B1(n_3),
.B2(n_4),
.Y(n_245)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_144),
.B1(n_151),
.B2(n_149),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_207),
.A2(n_188),
.B1(n_212),
.B2(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_211),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_189),
.C(n_179),
.Y(n_227)
);

NAND3xp33_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_165),
.C(n_135),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_L g241 ( 
.A1(n_210),
.A2(n_185),
.B(n_176),
.Y(n_241)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_167),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_212),
.B(n_217),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_183),
.B(n_161),
.Y(n_215)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_197),
.B(n_144),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_216),
.B(n_221),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_194),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_218),
.A2(n_196),
.B1(n_110),
.B2(n_113),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_178),
.B(n_113),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_171),
.A2(n_111),
.B(n_1),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_223),
.A2(n_224),
.B(n_191),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_192),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_189),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_237),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_231),
.C(n_234),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_203),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_232),
.Y(n_253)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_230),
.A2(n_241),
.B(n_226),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_172),
.C(n_169),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_214),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_233),
.A2(n_208),
.B1(n_202),
.B2(n_207),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_181),
.C(n_176),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_198),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_224),
.A2(n_170),
.B1(n_191),
.B2(n_187),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_245),
.B1(n_200),
.B2(n_240),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_182),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_246),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_223),
.B(n_218),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_0),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_233),
.A2(n_205),
.B1(n_221),
.B2(n_216),
.Y(n_248)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_199),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_255),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_251),
.B(n_237),
.Y(n_272)
);

AOI21x1_ASAP7_75t_SL g252 ( 
.A1(n_230),
.A2(n_199),
.B(n_210),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_242),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_219),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_257),
.C(n_231),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_206),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_204),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_217),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_261),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_260),
.Y(n_265)
);

OAI321xp33_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_200),
.A3(n_213),
.B1(n_202),
.B2(n_215),
.C(n_211),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_243),
.B(n_229),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_263),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_238),
.B(n_226),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_264),
.A2(n_270),
.B(n_274),
.Y(n_284)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_272),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_234),
.C(n_236),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_277),
.C(n_256),
.Y(n_288)
);

AOI21x1_ASAP7_75t_L g274 ( 
.A1(n_251),
.A2(n_243),
.B(n_229),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_258),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_263),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_246),
.C(n_3),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_267),
.B(n_253),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_278),
.B(n_279),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_277),
.B(n_249),
.Y(n_279)
);

INVx11_ASAP7_75t_L g280 ( 
.A(n_275),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_0),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_285),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_268),
.B(n_248),
.Y(n_285)
);

AND2x6_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_257),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_286),
.A2(n_4),
.B(n_5),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_249),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_287),
.B(n_4),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_288),
.B(n_269),
.C(n_272),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_256),
.C(n_254),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_265),
.C(n_3),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_296),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_284),
.A2(n_264),
.B(n_271),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_294),
.B(n_298),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_295),
.Y(n_304)
);

XNOR2x1_ASAP7_75t_SL g297 ( 
.A(n_286),
.B(n_4),
.Y(n_297)
);

NAND3xp33_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_5),
.C(n_6),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_299),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_281),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_301),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_283),
.C1(n_304),
.C2(n_300),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_297),
.A2(n_280),
.B1(n_284),
.B2(n_288),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_302),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_308)
);

OAI221xp5_ASAP7_75t_L g305 ( 
.A1(n_303),
.A2(n_291),
.B1(n_294),
.B2(n_283),
.C(n_289),
.Y(n_305)
);

AO21x2_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_306),
.B(n_8),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_6),
.C(n_7),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_309),
.Y(n_311)
);

AO21x2_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_310),
.B(n_307),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_8),
.Y(n_313)
);


endmodule