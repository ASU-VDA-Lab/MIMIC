module fake_jpeg_25110_n_149 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_149);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx11_ASAP7_75t_SL g48 ( 
.A(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_10),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_0),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_12),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_27),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_1),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_63),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_74),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_52),
.B1(n_49),
.B2(n_59),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_83),
.B1(n_56),
.B2(n_50),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_86),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_52),
.B1(n_60),
.B2(n_69),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_54),
.C(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_47),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_92),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_53),
.B1(n_56),
.B2(n_62),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_50),
.B1(n_67),
.B2(n_64),
.Y(n_107)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_97),
.Y(n_102)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_79),
.B1(n_3),
.B2(n_4),
.Y(n_112)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_79),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_53),
.C(n_47),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_22),
.C(n_37),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_2),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_93),
.B1(n_7),
.B2(n_8),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_46),
.B1(n_58),
.B2(n_55),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_108),
.A2(n_112),
.B1(n_90),
.B2(n_96),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_20),
.C(n_45),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_0),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_124),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_117),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_25),
.B1(n_41),
.B2(n_38),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

AND2x4_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_13),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_123),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_19),
.B(n_35),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_6),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_9),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_122),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_11),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_132),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_127),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_137),
.C(n_138),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_122),
.B1(n_113),
.B2(n_110),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_103),
.C(n_15),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_128),
.C(n_129),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_135),
.C(n_133),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_140),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_14),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_26),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_145),
.B(n_31),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_32),
.B(n_34),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_147),
.B(n_43),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_113),
.Y(n_149)
);


endmodule