module real_jpeg_25857_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_2),
.A2(n_25),
.B1(n_35),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_2),
.A2(n_56),
.B1(n_57),
.B2(n_65),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_65),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_3),
.A2(n_24),
.B1(n_68),
.B2(n_71),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_3),
.A2(n_25),
.B1(n_35),
.B2(n_71),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_3),
.A2(n_56),
.B1(n_57),
.B2(n_71),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_71),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_4),
.A2(n_25),
.B1(n_35),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_4),
.A2(n_39),
.B1(n_40),
.B2(n_62),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_4),
.A2(n_56),
.B1(n_57),
.B2(n_62),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_5),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_5),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_5),
.A2(n_25),
.B1(n_35),
.B2(n_82),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_5),
.A2(n_56),
.B1(n_57),
.B2(n_82),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_82),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_6),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx8_ASAP7_75t_SL g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_9),
.B(n_77),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_9),
.A2(n_33),
.B1(n_56),
.B2(n_57),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_9),
.A2(n_40),
.B(n_97),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_9),
.B(n_114),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_9),
.A2(n_87),
.B1(n_173),
.B2(n_176),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_9),
.A2(n_35),
.B(n_188),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_10),
.A2(n_46),
.B1(n_56),
.B2(n_57),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_11),
.A2(n_39),
.B1(n_40),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_11),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_11),
.A2(n_56),
.B1(n_57),
.B2(n_94),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_15),
.Y(n_159)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_15),
.Y(n_176)
);

HAxp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_132),
.CON(n_16),
.SN(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_116),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_20),
.B(n_116),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_83),
.B1(n_84),
.B2(n_115),
.Y(n_20)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_21),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_51),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_23),
.A2(n_36),
.B1(n_37),
.B2(n_120),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_23),
.Y(n_120)
);

OAI32xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.A3(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_23)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_25),
.A2(n_35),
.B1(n_55),
.B2(n_59),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_25),
.A2(n_28),
.B1(n_29),
.B2(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_25),
.B(n_33),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_28),
.A2(n_29),
.B1(n_69),
.B2(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_31),
.A2(n_33),
.B(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_33),
.A2(n_57),
.B(n_99),
.C(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_33),
.B(n_96),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_33),
.B(n_176),
.Y(n_178)
);

OAI32xp33_ASAP7_75t_L g196 ( 
.A1(n_35),
.A2(n_55),
.A3(n_57),
.B1(n_189),
.B2(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_37)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_38),
.B(n_93),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_38),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_39),
.A2(n_40),
.B1(n_97),
.B2(n_99),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_39),
.B(n_178),
.Y(n_177)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_45),
.A2(n_48),
.B(n_129),
.Y(n_128)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g166 ( 
.A(n_48),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_66),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_61),
.B(n_63),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_53),
.A2(n_61),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_53),
.A2(n_113),
.B1(n_114),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_53),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_54),
.A2(n_125),
.B1(n_187),
.B2(n_190),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_54)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_56),
.A2(n_57),
.B1(n_97),
.B2(n_99),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_56),
.B(n_59),
.Y(n_197)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_67),
.A2(n_72),
.B1(n_77),
.B2(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_74),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_106),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_95),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B(n_89),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_87),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_87),
.A2(n_159),
.B1(n_164),
.B2(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_87),
.A2(n_89),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B(n_101),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_103),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_96),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_139)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

BUFx24_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_108),
.B(n_109),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_104),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_104),
.A2(n_143),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_104),
.A2(n_151),
.B1(n_152),
.B2(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.C(n_112),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_112),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_108),
.B(n_151),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.C(n_121),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_117),
.B(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_119),
.A2(n_121),
.B1(n_122),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_119),
.Y(n_223)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.C(n_127),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_123),
.B(n_208),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_126),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_219),
.B(n_224),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_203),
.B(n_218),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_182),
.B(n_202),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_160),
.B(n_181),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_146),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_137),
.B(n_146),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_144),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_138),
.A2(n_139),
.B1(n_144),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_141),
.A2(n_214),
.B(n_215),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_144),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_154),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_153),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_153),
.C(n_154),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_155),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_169),
.B(n_180),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_167),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_162),
.B(n_167),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_174),
.B(n_179),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_171),
.B(n_172),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_183),
.B(n_184),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_195),
.B1(n_200),
.B2(n_201),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_185),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_185)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_191),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_194),
.C(n_200),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_192),
.Y(n_214)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_195),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_198),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_204),
.B(n_205),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_213),
.C(n_216),
.Y(n_220)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_216),
.B2(n_217),
.Y(n_211)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_213),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_220),
.B(n_221),
.Y(n_224)
);


endmodule