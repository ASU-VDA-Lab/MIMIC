module fake_netlist_5_203_n_1675 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1675);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1675;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_117),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_77),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_33),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_119),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_23),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_34),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_95),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_88),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_18),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_152),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_30),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_93),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_135),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_11),
.Y(n_172)
);

BUFx10_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_8),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_116),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_51),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_16),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_98),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_59),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_63),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_58),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_87),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_104),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_2),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_127),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_12),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_68),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_90),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_113),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_85),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_99),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_24),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_109),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_35),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_149),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_72),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_31),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_81),
.Y(n_202)
);

BUFx2_ASAP7_75t_R g203 ( 
.A(n_79),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_144),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_52),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_51),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_19),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_52),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_25),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_29),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_89),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_153),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_91),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_20),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_130),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_36),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_22),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_114),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_31),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_125),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_49),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_138),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_12),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_74),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_151),
.Y(n_227)
);

HB1xp67_ASAP7_75t_SL g228 ( 
.A(n_96),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_24),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_5),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_5),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_10),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_101),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_115),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_38),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_129),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_42),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_110),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_66),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_22),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_56),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_120),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_28),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_124),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_100),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_29),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_73),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_75),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_25),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_4),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_123),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_40),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_54),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_147),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_118),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_76),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_126),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_44),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_13),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_112),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_38),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_132),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_92),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_26),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_23),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_40),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_60),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_47),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_86),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_16),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_13),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_150),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_33),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_106),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_78),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_108),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_71),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_37),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_80),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_70),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_64),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_19),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_26),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_49),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_27),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_18),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_20),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_3),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_21),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_69),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_45),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_105),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_46),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_3),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_54),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_8),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_11),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_57),
.Y(n_298)
);

BUFx5_ASAP7_75t_L g299 ( 
.A(n_15),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_140),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_47),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_65),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_122),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_7),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_97),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_44),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_145),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_55),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_32),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_271),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_158),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_169),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_184),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_155),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_156),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_161),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_166),
.B(n_0),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_271),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_190),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_163),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_299),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_225),
.B(n_0),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_299),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_165),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_299),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_218),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_235),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_168),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_217),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_299),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_308),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_299),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_175),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_274),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_292),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_178),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_299),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_235),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_299),
.Y(n_339)
);

NOR2xp67_ASAP7_75t_L g340 ( 
.A(n_235),
.B(n_1),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_236),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_218),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_309),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_299),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_166),
.B(n_1),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_159),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_225),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_179),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_185),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_232),
.B(n_2),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_187),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_299),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_309),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_191),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_236),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_309),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_192),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_309),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_280),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_228),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_197),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_249),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_309),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_199),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_232),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_157),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_180),
.B(n_260),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_157),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_170),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_200),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_224),
.B(n_4),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_204),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_211),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_224),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_282),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_215),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_222),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_282),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_283),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_283),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_226),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_177),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_177),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_233),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_234),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_343),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_311),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_312),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_313),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_314),
.B(n_170),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_315),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_316),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_320),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_343),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_324),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_319),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_337),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_337),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_360),
.B(n_173),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_328),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_360),
.Y(n_401)
);

OA21x2_ASAP7_75t_L g402 ( 
.A1(n_321),
.A2(n_171),
.B(n_162),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_340),
.B(n_343),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_333),
.B(n_269),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_336),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_181),
.Y(n_406)
);

INVx6_ASAP7_75t_L g407 ( 
.A(n_369),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_329),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_337),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_334),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_348),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_327),
.B(n_269),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_352),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_353),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_353),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_356),
.Y(n_416)
);

BUFx8_ASAP7_75t_L g417 ( 
.A(n_322),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_349),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_356),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_351),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_335),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_362),
.B(n_173),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_359),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_352),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_367),
.B(n_180),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_354),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_362),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_358),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_357),
.B(n_303),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_352),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_361),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_358),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_370),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_321),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_372),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_369),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_373),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_381),
.B(n_303),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_346),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_363),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_323),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_363),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_382),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_364),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_327),
.B(n_186),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_347),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_338),
.B(n_186),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_384),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_385),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_376),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g452 ( 
.A1(n_323),
.A2(n_171),
.B(n_162),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_338),
.B(n_260),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_325),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_383),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_377),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_325),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_386),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_390),
.B(n_367),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_403),
.B(n_436),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_397),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_403),
.B(n_369),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_427),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_403),
.B(n_330),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_386),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_397),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_394),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_427),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_409),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_397),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_407),
.Y(n_472)
);

BUFx10_ASAP7_75t_L g473 ( 
.A(n_406),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_403),
.B(n_193),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_412),
.B(n_368),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_434),
.Y(n_476)
);

INVx4_ASAP7_75t_SL g477 ( 
.A(n_454),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_434),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_434),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_436),
.B(n_330),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_L g481 ( 
.A(n_425),
.B(n_345),
.C(n_317),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_412),
.B(n_368),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_404),
.B(n_429),
.Y(n_484)
);

INVx4_ASAP7_75t_SL g485 ( 
.A(n_454),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_446),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_436),
.B(n_340),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_445),
.A2(n_371),
.B1(n_322),
.B2(n_318),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_441),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_386),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_417),
.B(n_445),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_456),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_407),
.B(n_332),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_386),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_417),
.B(n_193),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_413),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_417),
.B(n_447),
.Y(n_497)
);

OR2x6_ASAP7_75t_L g498 ( 
.A(n_399),
.B(n_366),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_407),
.B(n_332),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_423),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_444),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_417),
.B(n_195),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_447),
.A2(n_310),
.B1(n_318),
.B2(n_350),
.Y(n_503)
);

BUFx10_ASAP7_75t_L g504 ( 
.A(n_391),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_413),
.Y(n_505)
);

AND2x6_ASAP7_75t_L g506 ( 
.A(n_441),
.B(n_195),
.Y(n_506)
);

BUFx4f_ASAP7_75t_L g507 ( 
.A(n_402),
.Y(n_507)
);

BUFx10_ASAP7_75t_L g508 ( 
.A(n_392),
.Y(n_508)
);

INVx5_ASAP7_75t_L g509 ( 
.A(n_457),
.Y(n_509)
);

AND2x6_ASAP7_75t_L g510 ( 
.A(n_441),
.B(n_202),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_439),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_438),
.B(n_202),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_430),
.Y(n_513)
);

BUFx10_ASAP7_75t_L g514 ( 
.A(n_393),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_407),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_409),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_407),
.B(n_339),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_386),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_430),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_453),
.B(n_310),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_402),
.A2(n_350),
.B1(n_331),
.B2(n_188),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_454),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_422),
.B(n_347),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_402),
.A2(n_452),
.B1(n_450),
.B2(n_443),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_454),
.Y(n_525)
);

INVxp33_ASAP7_75t_L g526 ( 
.A(n_443),
.Y(n_526)
);

OR2x6_ASAP7_75t_L g527 ( 
.A(n_450),
.B(n_366),
.Y(n_527)
);

AO22x2_ASAP7_75t_L g528 ( 
.A1(n_455),
.A2(n_221),
.B1(n_231),
.B2(n_188),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_430),
.Y(n_529)
);

BUFx4f_ASAP7_75t_L g530 ( 
.A(n_402),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_457),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_395),
.B(n_341),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_409),
.Y(n_533)
);

BUFx10_ASAP7_75t_L g534 ( 
.A(n_400),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_401),
.Y(n_535)
);

BUFx8_ASAP7_75t_SL g536 ( 
.A(n_387),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_398),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_401),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_457),
.B(n_339),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_409),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_457),
.B(n_344),
.Y(n_541)
);

OAI22xp33_ASAP7_75t_L g542 ( 
.A1(n_405),
.A2(n_265),
.B1(n_219),
.B2(n_252),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_455),
.B(n_365),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_398),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_414),
.B(n_365),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_457),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_409),
.B(n_182),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_414),
.Y(n_548)
);

NAND3xp33_ASAP7_75t_L g549 ( 
.A(n_411),
.B(n_326),
.C(n_342),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_418),
.B(n_183),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_420),
.B(n_355),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_415),
.Y(n_552)
);

INVx6_ASAP7_75t_L g553 ( 
.A(n_426),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_416),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_452),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_416),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_451),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_452),
.B(n_326),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_419),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_419),
.B(n_182),
.Y(n_560)
);

AND2x2_ASAP7_75t_SL g561 ( 
.A(n_452),
.B(n_189),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_431),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_398),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_424),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_428),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_428),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_424),
.B(n_189),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_424),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_424),
.B(n_344),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_433),
.B(n_342),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_432),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_432),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_388),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_440),
.Y(n_574)
);

INVx5_ASAP7_75t_L g575 ( 
.A(n_440),
.Y(n_575)
);

INVxp33_ASAP7_75t_L g576 ( 
.A(n_442),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_442),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_435),
.B(n_238),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_437),
.B(n_375),
.Y(n_579)
);

NAND2xp33_ASAP7_75t_L g580 ( 
.A(n_448),
.B(n_183),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_449),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_389),
.B(n_160),
.Y(n_582)
);

AND2x2_ASAP7_75t_SL g583 ( 
.A(n_396),
.B(n_194),
.Y(n_583)
);

INVx5_ASAP7_75t_L g584 ( 
.A(n_408),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_410),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_421),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_427),
.B(n_383),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_394),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_409),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_390),
.B(n_164),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_409),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_407),
.Y(n_592)
);

OR2x6_ASAP7_75t_L g593 ( 
.A(n_399),
.B(n_209),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_407),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_390),
.B(n_167),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_427),
.B(n_375),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_409),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_397),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_397),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_390),
.B(n_172),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_561),
.A2(n_231),
.B1(n_237),
.B2(n_221),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_577),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_463),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_543),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_577),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_484),
.B(n_194),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_461),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_553),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_472),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_459),
.B(n_174),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_461),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_553),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_475),
.B(n_212),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_475),
.B(n_212),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_568),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_543),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_481),
.A2(n_272),
.B1(n_307),
.B2(n_251),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_507),
.B(n_183),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_561),
.A2(n_253),
.B1(n_259),
.B2(n_261),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_545),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_587),
.B(n_176),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_467),
.Y(n_622)
);

NOR3xp33_ASAP7_75t_L g623 ( 
.A(n_468),
.B(n_230),
.C(n_306),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_483),
.B(n_213),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_564),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_488),
.A2(n_248),
.B1(n_247),
.B2(n_245),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_L g627 ( 
.A(n_558),
.B(n_239),
.Y(n_627)
);

NOR2x1p5_ASAP7_75t_L g628 ( 
.A(n_587),
.B(n_196),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_590),
.B(n_214),
.Y(n_629)
);

OR2x6_ASAP7_75t_L g630 ( 
.A(n_553),
.B(n_203),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_520),
.B(n_198),
.Y(n_631)
);

BUFx5_ASAP7_75t_L g632 ( 
.A(n_567),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_595),
.B(n_214),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_471),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_600),
.B(n_220),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_472),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_536),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_536),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_462),
.B(n_220),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_SL g640 ( 
.A1(n_583),
.A2(n_207),
.B1(n_206),
.B2(n_205),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_593),
.A2(n_241),
.B1(n_242),
.B2(n_244),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_507),
.B(n_183),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_530),
.B(n_558),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_SL g644 ( 
.A1(n_492),
.A2(n_201),
.B1(n_243),
.B2(n_304),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_487),
.B(n_245),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_584),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_480),
.B(n_247),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_460),
.B(n_248),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_464),
.B(n_255),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_537),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_593),
.A2(n_290),
.B1(n_305),
.B2(n_277),
.Y(n_651)
);

AOI221xp5_ASAP7_75t_L g652 ( 
.A1(n_542),
.A2(n_237),
.B1(n_210),
.B2(n_209),
.C(n_253),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_588),
.B(n_255),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_520),
.B(n_208),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_548),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_555),
.A2(n_287),
.B1(n_288),
.B2(n_210),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_526),
.B(n_216),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_555),
.A2(n_287),
.B1(n_288),
.B2(n_266),
.Y(n_658)
);

BUFx5_ASAP7_75t_L g659 ( 
.A(n_567),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_584),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_596),
.B(n_378),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_596),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_512),
.B(n_552),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_486),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_593),
.A2(n_257),
.B1(n_281),
.B2(n_254),
.Y(n_665)
);

BUFx6f_ASAP7_75t_SL g666 ( 
.A(n_504),
.Y(n_666)
);

NOR2x1p5_ASAP7_75t_L g667 ( 
.A(n_523),
.B(n_549),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_554),
.B(n_262),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_556),
.B(n_559),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_565),
.B(n_263),
.Y(n_670)
);

NOR2xp67_ASAP7_75t_L g671 ( 
.A(n_562),
.B(n_256),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_526),
.B(n_223),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_515),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_466),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_466),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_566),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_571),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_572),
.B(n_263),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_574),
.B(n_302),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_564),
.B(n_302),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_570),
.B(n_380),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_530),
.B(n_227),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_576),
.B(n_267),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_555),
.A2(n_259),
.B1(n_261),
.B2(n_266),
.Y(n_684)
);

NOR2xp67_ASAP7_75t_L g685 ( 
.A(n_562),
.B(n_275),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_470),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_530),
.B(n_227),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_524),
.B(n_227),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_576),
.B(n_276),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_579),
.B(n_380),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_528),
.A2(n_293),
.B1(n_296),
.B2(n_227),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_593),
.A2(n_497),
.B1(n_491),
.B2(n_579),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_521),
.B(n_279),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_540),
.B(n_298),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_544),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_578),
.B(n_300),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_503),
.A2(n_293),
.B(n_296),
.C(n_379),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_560),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_523),
.B(n_229),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_491),
.A2(n_173),
.B1(n_227),
.B2(n_301),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_511),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_582),
.Y(n_702)
);

INVx8_ASAP7_75t_L g703 ( 
.A(n_584),
.Y(n_703)
);

AOI21x1_ASAP7_75t_L g704 ( 
.A1(n_493),
.A2(n_379),
.B(n_378),
.Y(n_704)
);

NOR3xp33_ASAP7_75t_L g705 ( 
.A(n_497),
.B(n_297),
.C(n_295),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_560),
.B(n_82),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_563),
.Y(n_707)
);

NOR2xp67_ASAP7_75t_L g708 ( 
.A(n_584),
.B(n_83),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_495),
.A2(n_173),
.B1(n_291),
.B2(n_289),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_499),
.B(n_294),
.Y(n_710)
);

A2O1A1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_495),
.A2(n_268),
.B(n_285),
.C(n_284),
.Y(n_711)
);

OAI221xp5_ASAP7_75t_L g712 ( 
.A1(n_498),
.A2(n_286),
.B1(n_278),
.B2(n_273),
.C(n_270),
.Y(n_712)
);

AOI221xp5_ASAP7_75t_L g713 ( 
.A1(n_528),
.A2(n_264),
.B1(n_258),
.B2(n_250),
.C(n_246),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_474),
.B(n_240),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_515),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_538),
.Y(n_716)
);

AND2x6_ASAP7_75t_SL g717 ( 
.A(n_586),
.B(n_6),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_SL g718 ( 
.A(n_504),
.B(n_6),
.Y(n_718)
);

NOR3xp33_ASAP7_75t_L g719 ( 
.A(n_532),
.B(n_7),
.C(n_9),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_592),
.B(n_154),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_527),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_496),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_528),
.A2(n_9),
.B1(n_10),
.B2(n_14),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_594),
.B(n_141),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_469),
.B(n_136),
.Y(n_725)
);

OAI22x1_ASAP7_75t_L g726 ( 
.A1(n_535),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_563),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_502),
.A2(n_133),
.B1(n_131),
.B2(n_128),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_551),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_517),
.B(n_102),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_469),
.B(n_94),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_539),
.B(n_84),
.Y(n_732)
);

NOR3xp33_ASAP7_75t_L g733 ( 
.A(n_550),
.B(n_17),
.C(n_21),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_550),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_L g735 ( 
.A(n_567),
.B(n_547),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_505),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_527),
.B(n_28),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_527),
.B(n_30),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_527),
.B(n_32),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_473),
.B(n_34),
.Y(n_740)
);

AOI22x1_ASAP7_75t_L g741 ( 
.A1(n_528),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_498),
.B(n_39),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_505),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_473),
.B(n_39),
.Y(n_744)
);

A2O1A1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_502),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_745)
);

CKINVDCx16_ASAP7_75t_R g746 ( 
.A(n_504),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_602),
.Y(n_747)
);

NOR2xp67_ASAP7_75t_SL g748 ( 
.A(n_625),
.B(n_584),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_610),
.B(n_580),
.Y(n_749)
);

OAI21xp5_ASAP7_75t_L g750 ( 
.A1(n_643),
.A2(n_541),
.B(n_531),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_702),
.B(n_581),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_602),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_610),
.B(n_606),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_662),
.B(n_473),
.Y(n_754)
);

NOR3xp33_ASAP7_75t_L g755 ( 
.A(n_712),
.B(n_729),
.C(n_640),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_603),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_681),
.B(n_580),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_605),
.Y(n_758)
);

AOI21x1_ASAP7_75t_L g759 ( 
.A1(n_688),
.A2(n_546),
.B(n_525),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_643),
.A2(n_476),
.B(n_489),
.Y(n_760)
);

NOR2x1_ASAP7_75t_L g761 ( 
.A(n_608),
.B(n_498),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_609),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_629),
.B(n_498),
.Y(n_763)
);

OAI21xp5_ASAP7_75t_L g764 ( 
.A1(n_618),
.A2(n_478),
.B(n_479),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_633),
.B(n_516),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_635),
.B(n_516),
.Y(n_766)
);

NOR2x1_ASAP7_75t_L g767 ( 
.A(n_608),
.B(n_612),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_613),
.A2(n_569),
.B(n_598),
.C(n_599),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_601),
.B(n_533),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_601),
.B(n_533),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_618),
.A2(n_522),
.B(n_465),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_619),
.B(n_533),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_664),
.Y(n_773)
);

OAI21xp5_ASAP7_75t_L g774 ( 
.A1(n_642),
.A2(n_589),
.B(n_591),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_619),
.B(n_589),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_642),
.A2(n_522),
.B(n_458),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_605),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_661),
.B(n_690),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_607),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_655),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_734),
.A2(n_583),
.B1(n_597),
.B2(n_591),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_607),
.Y(n_782)
);

AOI21x1_ASAP7_75t_L g783 ( 
.A1(n_682),
.A2(n_599),
.B(n_598),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_L g784 ( 
.A1(n_682),
.A2(n_519),
.B(n_513),
.Y(n_784)
);

OAI21xp5_ASAP7_75t_L g785 ( 
.A1(n_687),
.A2(n_627),
.B(n_624),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_621),
.B(n_513),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_621),
.B(n_557),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_676),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_716),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_657),
.B(n_519),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_611),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_657),
.B(n_529),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_699),
.B(n_514),
.Y(n_793)
);

OAI22xp33_ASAP7_75t_L g794 ( 
.A1(n_718),
.A2(n_535),
.B1(n_492),
.B2(n_501),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_611),
.Y(n_795)
);

INVx11_ASAP7_75t_L g796 ( 
.A(n_666),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_715),
.A2(n_490),
.B(n_482),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_677),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_694),
.A2(n_494),
.B(n_518),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_672),
.B(n_529),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_701),
.B(n_573),
.Y(n_801)
);

NAND2xp33_ASAP7_75t_L g802 ( 
.A(n_632),
.B(n_567),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_692),
.B(n_534),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_672),
.B(n_614),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_609),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_622),
.Y(n_806)
);

A2O1A1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_699),
.A2(n_585),
.B(n_500),
.C(n_575),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_631),
.B(n_654),
.Y(n_808)
);

INVx1_ASAP7_75t_SL g809 ( 
.A(n_742),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_696),
.B(n_534),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_634),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_698),
.B(n_567),
.Y(n_812)
);

BUFx4f_ASAP7_75t_L g813 ( 
.A(n_703),
.Y(n_813)
);

NOR2x1p5_ASAP7_75t_SL g814 ( 
.A(n_632),
.B(n_477),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_721),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_612),
.B(n_585),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_663),
.A2(n_482),
.B(n_465),
.Y(n_817)
);

AO32x2_ASAP7_75t_L g818 ( 
.A1(n_626),
.A2(n_547),
.A3(n_506),
.B1(n_510),
.B2(n_48),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_648),
.A2(n_465),
.B(n_458),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_669),
.A2(n_509),
.B(n_575),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_693),
.A2(n_500),
.B1(n_575),
.B2(n_509),
.Y(n_821)
);

OAI21x1_ASAP7_75t_L g822 ( 
.A1(n_725),
.A2(n_477),
.B(n_485),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_609),
.Y(n_823)
);

O2A1O1Ixp5_ASAP7_75t_L g824 ( 
.A1(n_649),
.A2(n_510),
.B(n_506),
.C(n_547),
.Y(n_824)
);

NAND3xp33_ASAP7_75t_L g825 ( 
.A(n_631),
.B(n_654),
.C(n_713),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_700),
.A2(n_575),
.B(n_509),
.C(n_534),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_604),
.B(n_477),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_616),
.B(n_477),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_609),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_656),
.A2(n_684),
.B1(n_658),
.B2(n_620),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_738),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_645),
.A2(n_509),
.B(n_575),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_745),
.A2(n_547),
.B(n_510),
.C(n_506),
.Y(n_833)
);

O2A1O1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_745),
.A2(n_547),
.B(n_510),
.C(n_506),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_706),
.B(n_485),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_706),
.B(n_485),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_636),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_656),
.B(n_547),
.Y(n_838)
);

O2A1O1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_697),
.A2(n_506),
.B(n_510),
.C(n_46),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_680),
.A2(n_509),
.B(n_510),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_628),
.B(n_514),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_683),
.B(n_508),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_615),
.A2(n_506),
.B(n_67),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_658),
.B(n_508),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_707),
.Y(n_845)
);

O2A1O1Ixp5_ASAP7_75t_L g846 ( 
.A1(n_639),
.A2(n_41),
.B(n_43),
.C(n_48),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_684),
.B(n_508),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_636),
.A2(n_61),
.B(n_62),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_636),
.A2(n_50),
.B(n_53),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_689),
.B(n_50),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_674),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_697),
.A2(n_53),
.B(n_55),
.C(n_711),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_705),
.A2(n_667),
.B1(n_710),
.B2(n_714),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_636),
.A2(n_673),
.B(n_720),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_637),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_740),
.B(n_744),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_671),
.B(n_685),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_644),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_674),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_673),
.A2(n_724),
.B(n_735),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_646),
.B(n_660),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_740),
.B(n_744),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_675),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_617),
.B(n_737),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_668),
.B(n_679),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_691),
.A2(n_723),
.B1(n_711),
.B2(n_660),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_670),
.B(n_678),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_675),
.Y(n_868)
);

NOR2x1p5_ASAP7_75t_SL g869 ( 
.A(n_632),
.B(n_659),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_647),
.A2(n_653),
.B(n_732),
.C(n_710),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_737),
.B(n_739),
.Y(n_871)
);

NOR3xp33_ASAP7_75t_L g872 ( 
.A(n_739),
.B(n_652),
.C(n_719),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_646),
.B(n_708),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_733),
.A2(n_665),
.B(n_651),
.C(n_641),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_623),
.A2(n_727),
.B1(n_650),
.B2(n_695),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_746),
.B(n_709),
.Y(n_876)
);

CKINVDCx10_ASAP7_75t_R g877 ( 
.A(n_630),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_630),
.B(n_703),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_R g879 ( 
.A(n_638),
.B(n_703),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_686),
.B(n_743),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_630),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_731),
.A2(n_732),
.B(n_730),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_726),
.Y(n_883)
);

AO21x1_ASAP7_75t_L g884 ( 
.A1(n_730),
.A2(n_728),
.B(n_722),
.Y(n_884)
);

NOR3xp33_ASAP7_75t_L g885 ( 
.A(n_704),
.B(n_736),
.C(n_722),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_741),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_691),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_723),
.B(n_717),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_632),
.A2(n_625),
.B(n_530),
.Y(n_889)
);

NAND2x1p5_ASAP7_75t_L g890 ( 
.A(n_632),
.B(n_659),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_659),
.B(n_702),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_659),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_609),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_625),
.A2(n_530),
.B(n_507),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_625),
.A2(n_530),
.B(n_507),
.Y(n_895)
);

BUFx12f_ASAP7_75t_L g896 ( 
.A(n_603),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_601),
.A2(n_619),
.B1(n_606),
.B2(n_734),
.Y(n_897)
);

OAI321xp33_ASAP7_75t_L g898 ( 
.A1(n_626),
.A2(n_723),
.A3(n_610),
.B1(n_481),
.B2(n_317),
.C(n_371),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_662),
.B(n_427),
.Y(n_899)
);

NOR2x1_ASAP7_75t_L g900 ( 
.A(n_608),
.B(n_612),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_610),
.B(n_484),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_610),
.B(n_484),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_625),
.A2(n_530),
.B(n_507),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_610),
.B(n_484),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_610),
.B(n_484),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_609),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_610),
.A2(n_484),
.B1(n_692),
.B2(n_459),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_610),
.B(n_484),
.Y(n_908)
);

O2A1O1Ixp5_ASAP7_75t_SL g909 ( 
.A1(n_629),
.A2(n_633),
.B(n_635),
.C(n_606),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_625),
.A2(n_530),
.B(n_507),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_901),
.B(n_902),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_904),
.B(n_905),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_907),
.B(n_808),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_908),
.A2(n_753),
.B1(n_825),
.B2(n_897),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_889),
.A2(n_895),
.B(n_894),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_903),
.A2(n_910),
.B(n_802),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_909),
.A2(n_804),
.B(n_749),
.Y(n_917)
);

OAI21x1_ASAP7_75t_L g918 ( 
.A1(n_799),
.A2(n_759),
.B(n_854),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_838),
.A2(n_770),
.B(n_769),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_SL g920 ( 
.A1(n_890),
.A2(n_830),
.B(n_873),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_823),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_864),
.A2(n_871),
.B1(n_862),
.B2(n_856),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_899),
.B(n_787),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_778),
.B(n_871),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_780),
.Y(n_925)
);

CKINVDCx14_ASAP7_75t_R g926 ( 
.A(n_879),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_823),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_788),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_773),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_793),
.B(n_757),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_793),
.B(n_763),
.Y(n_931)
);

AOI21x1_ASAP7_75t_L g932 ( 
.A1(n_790),
.A2(n_800),
.B(n_792),
.Y(n_932)
);

O2A1O1Ixp5_ASAP7_75t_L g933 ( 
.A1(n_886),
.A2(n_884),
.B(n_882),
.C(n_764),
.Y(n_933)
);

OAI21x1_ASAP7_75t_L g934 ( 
.A1(n_824),
.A2(n_750),
.B(n_784),
.Y(n_934)
);

AO31x2_ASAP7_75t_L g935 ( 
.A1(n_866),
.A2(n_826),
.A3(n_807),
.B(n_772),
.Y(n_935)
);

INVx6_ASAP7_75t_SL g936 ( 
.A(n_816),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_751),
.B(n_865),
.Y(n_937)
);

AO31x2_ASAP7_75t_L g938 ( 
.A1(n_775),
.A2(n_786),
.A3(n_781),
.B(n_850),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_870),
.A2(n_898),
.B(n_768),
.Y(n_939)
);

AOI21x1_ASAP7_75t_L g940 ( 
.A1(n_771),
.A2(n_776),
.B(n_819),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_867),
.B(n_891),
.Y(n_941)
);

INVx4_ASAP7_75t_L g942 ( 
.A(n_823),
.Y(n_942)
);

OAI21x1_ASAP7_75t_L g943 ( 
.A1(n_817),
.A2(n_774),
.B(n_797),
.Y(n_943)
);

AO31x2_ASAP7_75t_L g944 ( 
.A1(n_765),
.A2(n_766),
.A3(n_887),
.B(n_891),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_831),
.B(n_809),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_870),
.A2(n_768),
.B(n_760),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_SL g947 ( 
.A1(n_873),
.A2(n_892),
.B(n_906),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_773),
.Y(n_948)
);

AOI21xp33_ASAP7_75t_L g949 ( 
.A1(n_844),
.A2(n_847),
.B(n_801),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_798),
.B(n_806),
.Y(n_950)
);

AO31x2_ASAP7_75t_L g951 ( 
.A1(n_874),
.A2(n_821),
.A3(n_747),
.B(n_752),
.Y(n_951)
);

NAND2xp33_ASAP7_75t_L g952 ( 
.A(n_823),
.B(n_829),
.Y(n_952)
);

OAI21x1_ASAP7_75t_L g953 ( 
.A1(n_824),
.A2(n_834),
.B(n_833),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_811),
.B(n_853),
.Y(n_954)
);

AOI21x1_ASAP7_75t_SL g955 ( 
.A1(n_827),
.A2(n_828),
.B(n_812),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_779),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_835),
.A2(n_836),
.B(n_892),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_831),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_872),
.A2(n_852),
.B(n_888),
.C(n_755),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_782),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_791),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_833),
.A2(n_834),
.B(n_880),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_795),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_861),
.A2(n_857),
.B(n_805),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_829),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_762),
.A2(n_893),
.B(n_813),
.Y(n_966)
);

AND3x4_ASAP7_75t_L g967 ( 
.A(n_755),
.B(n_872),
.C(n_761),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_789),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_813),
.A2(n_803),
.B(n_840),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_754),
.B(n_756),
.Y(n_970)
);

OAI21x1_ASAP7_75t_SL g971 ( 
.A1(n_839),
.A2(n_852),
.B(n_849),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_758),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_832),
.A2(n_820),
.B(n_843),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_794),
.B(n_842),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_885),
.A2(n_777),
.B(n_851),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_885),
.A2(n_868),
.B(n_859),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_L g977 ( 
.A(n_883),
.B(n_815),
.C(n_876),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_863),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_845),
.A2(n_875),
.B(n_848),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_896),
.Y(n_980)
);

OAI21x1_ASAP7_75t_L g981 ( 
.A1(n_839),
.A2(n_900),
.B(n_767),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_846),
.A2(n_883),
.B(n_869),
.C(n_878),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_816),
.B(n_815),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_829),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_748),
.B(n_810),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_846),
.A2(n_858),
.B(n_841),
.C(n_814),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_818),
.A2(n_881),
.B(n_906),
.C(n_829),
.Y(n_987)
);

OAI21x1_ASAP7_75t_L g988 ( 
.A1(n_837),
.A2(n_906),
.B(n_818),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_837),
.B(n_855),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_818),
.A2(n_837),
.B(n_877),
.C(n_796),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_901),
.A2(n_904),
.B(n_905),
.C(n_902),
.Y(n_991)
);

OAI21x1_ASAP7_75t_L g992 ( 
.A1(n_822),
.A2(n_783),
.B(n_860),
.Y(n_992)
);

O2A1O1Ixp5_ASAP7_75t_L g993 ( 
.A1(n_808),
.A2(n_753),
.B(n_902),
.C(n_901),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_901),
.A2(n_904),
.B(n_905),
.C(n_902),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_899),
.B(n_427),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_901),
.B(n_902),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_773),
.Y(n_997)
);

OAI21x1_ASAP7_75t_L g998 ( 
.A1(n_822),
.A2(n_783),
.B(n_860),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_780),
.Y(n_999)
);

OR2x6_ASAP7_75t_L g1000 ( 
.A(n_896),
.B(n_703),
.Y(n_1000)
);

OAI21x1_ASAP7_75t_L g1001 ( 
.A1(n_822),
.A2(n_783),
.B(n_860),
.Y(n_1001)
);

AOI21x1_ASAP7_75t_L g1002 ( 
.A1(n_759),
.A2(n_642),
.B(n_618),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_822),
.A2(n_783),
.B(n_860),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_779),
.Y(n_1004)
);

BUFx4f_ASAP7_75t_L g1005 ( 
.A(n_896),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_901),
.A2(n_904),
.B(n_902),
.Y(n_1006)
);

OA21x2_ASAP7_75t_L g1007 ( 
.A1(n_785),
.A2(n_764),
.B(n_760),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_780),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_808),
.A2(n_901),
.B1(n_904),
.B2(n_902),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_780),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_896),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_SL g1012 ( 
.A(n_808),
.B(n_902),
.C(n_901),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_901),
.B(n_902),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_901),
.B(n_902),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_901),
.A2(n_904),
.B(n_905),
.C(n_902),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_901),
.A2(n_904),
.B(n_905),
.C(n_902),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_901),
.B(n_902),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_780),
.Y(n_1018)
);

INVxp67_ASAP7_75t_L g1019 ( 
.A(n_773),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_822),
.A2(n_783),
.B(n_860),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_901),
.A2(n_904),
.B(n_902),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_SL g1022 ( 
.A1(n_833),
.A2(n_834),
.B(n_839),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_901),
.B(n_902),
.Y(n_1023)
);

OR2x6_ASAP7_75t_L g1024 ( 
.A(n_896),
.B(n_703),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_808),
.B(n_901),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_901),
.B(n_902),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_901),
.A2(n_904),
.B(n_902),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_822),
.A2(n_783),
.B(n_860),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_901),
.A2(n_904),
.B(n_902),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_901),
.B(n_902),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_779),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_901),
.A2(n_902),
.B1(n_905),
.B2(n_904),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_823),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_901),
.B(n_902),
.Y(n_1034)
);

AOI221xp5_ASAP7_75t_SL g1035 ( 
.A1(n_901),
.A2(n_626),
.B1(n_902),
.B2(n_905),
.C(n_904),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_SL g1036 ( 
.A(n_816),
.Y(n_1036)
);

AO31x2_ASAP7_75t_L g1037 ( 
.A1(n_884),
.A2(n_886),
.A3(n_866),
.B(n_897),
.Y(n_1037)
);

AO21x2_ASAP7_75t_L g1038 ( 
.A1(n_785),
.A2(n_885),
.B(n_882),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_956),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_925),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_1025),
.A2(n_922),
.B(n_1009),
.C(n_1006),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_1025),
.A2(n_911),
.B1(n_912),
.B2(n_996),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_1021),
.A2(n_1029),
.B(n_1027),
.C(n_959),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_989),
.B(n_983),
.Y(n_1044)
);

O2A1O1Ixp5_ASAP7_75t_L g1045 ( 
.A1(n_939),
.A2(n_913),
.B(n_917),
.C(n_914),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_945),
.B(n_970),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1013),
.A2(n_1017),
.B1(n_1034),
.B2(n_1014),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_948),
.Y(n_1048)
);

AND2x6_ASAP7_75t_L g1049 ( 
.A(n_921),
.B(n_965),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_913),
.A2(n_967),
.B1(n_1012),
.B2(n_974),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_929),
.Y(n_1051)
);

CKINVDCx8_ASAP7_75t_R g1052 ( 
.A(n_980),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1023),
.A2(n_1026),
.B1(n_1030),
.B2(n_937),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_923),
.B(n_995),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_929),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_991),
.A2(n_1015),
.B(n_1016),
.C(n_994),
.Y(n_1056)
);

INVx3_ASAP7_75t_SL g1057 ( 
.A(n_968),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_959),
.A2(n_993),
.B(n_994),
.C(n_991),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_958),
.B(n_928),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1032),
.B(n_924),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1015),
.B(n_1016),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_997),
.Y(n_1062)
);

AO21x1_ASAP7_75t_L g1063 ( 
.A1(n_930),
.A2(n_931),
.B(n_941),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_967),
.A2(n_1012),
.B1(n_974),
.B2(n_949),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_960),
.Y(n_1065)
);

INVxp67_ASAP7_75t_SL g1066 ( 
.A(n_1019),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_999),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_954),
.B(n_1035),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_919),
.B(n_987),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1008),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_987),
.A2(n_990),
.B1(n_950),
.B2(n_1010),
.Y(n_1071)
);

O2A1O1Ixp5_ASAP7_75t_L g1072 ( 
.A1(n_993),
.A2(n_933),
.B(n_915),
.C(n_932),
.Y(n_1072)
);

NOR2x1_ASAP7_75t_L g1073 ( 
.A(n_942),
.B(n_984),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1018),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_972),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_990),
.A2(n_982),
.B1(n_986),
.B2(n_962),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_921),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_1019),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_961),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_986),
.A2(n_982),
.B(n_971),
.C(n_1022),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_958),
.B(n_1000),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_961),
.B(n_963),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_977),
.B(n_963),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_1000),
.B(n_1024),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_978),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1036),
.A2(n_926),
.B1(n_985),
.B2(n_1011),
.Y(n_1086)
);

CKINVDCx6p67_ASAP7_75t_R g1087 ( 
.A(n_1011),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1036),
.A2(n_926),
.B1(n_1005),
.B2(n_1024),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_1000),
.B(n_1024),
.Y(n_1089)
);

CKINVDCx6p67_ASAP7_75t_R g1090 ( 
.A(n_921),
.Y(n_1090)
);

INVxp67_ASAP7_75t_SL g1091 ( 
.A(n_952),
.Y(n_1091)
);

O2A1O1Ixp5_ASAP7_75t_L g1092 ( 
.A1(n_933),
.A2(n_916),
.B(n_940),
.C(n_1002),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_1004),
.B(n_1031),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1004),
.B(n_1031),
.Y(n_1094)
);

CKINVDCx16_ASAP7_75t_R g1095 ( 
.A(n_942),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1037),
.B(n_944),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1037),
.B(n_944),
.Y(n_1097)
);

NAND2xp33_ASAP7_75t_L g1098 ( 
.A(n_965),
.B(n_966),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_936),
.B(n_920),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1037),
.B(n_944),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_927),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_979),
.A2(n_964),
.B(n_969),
.C(n_981),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_965),
.Y(n_1103)
);

INVxp33_ASAP7_75t_L g1104 ( 
.A(n_1005),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_965),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_927),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_951),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_936),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_SL g1109 ( 
.A1(n_952),
.A2(n_1007),
.B1(n_1038),
.B2(n_984),
.Y(n_1109)
);

BUFx12f_ASAP7_75t_L g1110 ( 
.A(n_936),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_951),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1033),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1033),
.B(n_951),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1038),
.A2(n_957),
.B1(n_976),
.B2(n_975),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_938),
.B(n_935),
.Y(n_1115)
);

INVx3_ASAP7_75t_SL g1116 ( 
.A(n_1007),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_988),
.Y(n_1117)
);

CKINVDCx11_ASAP7_75t_R g1118 ( 
.A(n_947),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_938),
.B(n_935),
.Y(n_1119)
);

INVxp67_ASAP7_75t_L g1120 ( 
.A(n_953),
.Y(n_1120)
);

INVx3_ASAP7_75t_SL g1121 ( 
.A(n_1007),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_938),
.B(n_935),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_944),
.B(n_938),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_935),
.B(n_934),
.Y(n_1124)
);

OR2x2_ASAP7_75t_SL g1125 ( 
.A(n_955),
.B(n_918),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_943),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_934),
.Y(n_1127)
);

OR2x6_ASAP7_75t_SL g1128 ( 
.A(n_973),
.B(n_992),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_998),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_1001),
.B(n_1003),
.Y(n_1130)
);

INVx5_ASAP7_75t_L g1131 ( 
.A(n_1020),
.Y(n_1131)
);

INVxp67_ASAP7_75t_L g1132 ( 
.A(n_1028),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1025),
.B(n_911),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_925),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1025),
.B(n_911),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_956),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_948),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_921),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_995),
.B(n_463),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_925),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_926),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_923),
.B(n_995),
.Y(n_1142)
);

OR2x2_ASAP7_75t_L g1143 ( 
.A(n_995),
.B(n_463),
.Y(n_1143)
);

OR2x2_ASAP7_75t_L g1144 ( 
.A(n_995),
.B(n_463),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_956),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_922),
.A2(n_1025),
.B1(n_902),
.B2(n_904),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_925),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_922),
.A2(n_808),
.B1(n_864),
.B2(n_1025),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_921),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_926),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_913),
.A2(n_808),
.B1(n_864),
.B2(n_825),
.Y(n_1151)
);

INVx3_ASAP7_75t_SL g1152 ( 
.A(n_968),
.Y(n_1152)
);

AOI221x1_ASAP7_75t_L g1153 ( 
.A1(n_939),
.A2(n_808),
.B1(n_862),
.B2(n_856),
.C(n_914),
.Y(n_1153)
);

AOI221xp5_ASAP7_75t_L g1154 ( 
.A1(n_1025),
.A2(n_808),
.B1(n_922),
.B2(n_898),
.C(n_1032),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_929),
.Y(n_1155)
);

BUFx8_ASAP7_75t_L g1156 ( 
.A(n_1036),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1025),
.B(n_911),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_989),
.B(n_767),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_989),
.B(n_767),
.Y(n_1159)
);

NOR2x1_ASAP7_75t_SL g1160 ( 
.A(n_921),
.B(n_965),
.Y(n_1160)
);

OR2x2_ASAP7_75t_SL g1161 ( 
.A(n_977),
.B(n_746),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1025),
.B(n_911),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_921),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_922),
.B(n_808),
.Y(n_1164)
);

OAI22x1_ASAP7_75t_L g1165 ( 
.A1(n_922),
.A2(n_967),
.B1(n_862),
.B2(n_856),
.Y(n_1165)
);

OA21x2_ASAP7_75t_L g1166 ( 
.A1(n_946),
.A2(n_939),
.B(n_933),
.Y(n_1166)
);

INVx6_ASAP7_75t_SL g1167 ( 
.A(n_1000),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_956),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1025),
.B(n_911),
.Y(n_1169)
);

BUFx12f_ASAP7_75t_L g1170 ( 
.A(n_980),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_921),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_956),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_921),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1164),
.A2(n_1154),
.B1(n_1151),
.B2(n_1165),
.Y(n_1174)
);

OA21x2_ASAP7_75t_L g1175 ( 
.A1(n_1072),
.A2(n_1092),
.B(n_1045),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1044),
.B(n_1084),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_1156),
.Y(n_1177)
);

AND2x2_ASAP7_75t_SL g1178 ( 
.A(n_1154),
.B(n_1064),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1113),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1067),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1070),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1050),
.B(n_1041),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1148),
.B(n_1043),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1062),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1074),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1146),
.A2(n_1076),
.B1(n_1042),
.B2(n_1142),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1134),
.Y(n_1187)
);

INVxp67_ASAP7_75t_L g1188 ( 
.A(n_1139),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_1099),
.B(n_1131),
.Y(n_1189)
);

BUFx2_ASAP7_75t_L g1190 ( 
.A(n_1137),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1140),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1147),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1075),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1079),
.Y(n_1194)
);

AO21x1_ASAP7_75t_L g1195 ( 
.A1(n_1076),
.A2(n_1056),
.B(n_1080),
.Y(n_1195)
);

BUFx10_ASAP7_75t_L g1196 ( 
.A(n_1141),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1065),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1085),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1133),
.A2(n_1135),
.B1(n_1169),
.B2(n_1157),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1136),
.Y(n_1200)
);

BUFx12f_ASAP7_75t_L g1201 ( 
.A(n_1156),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_1059),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1062),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_SL g1204 ( 
.A1(n_1091),
.A2(n_1080),
.B(n_1153),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1145),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1168),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_1046),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1172),
.Y(n_1208)
);

AO21x1_ASAP7_75t_L g1209 ( 
.A1(n_1056),
.A2(n_1061),
.B(n_1060),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1044),
.B(n_1084),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1046),
.Y(n_1211)
);

OAI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1146),
.A2(n_1162),
.B1(n_1133),
.B2(n_1157),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1135),
.A2(n_1169),
.B1(n_1162),
.B2(n_1042),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1059),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1054),
.A2(n_1053),
.B1(n_1047),
.B2(n_1060),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1143),
.A2(n_1144),
.B1(n_1161),
.B2(n_1066),
.Y(n_1216)
);

NOR2x1_ASAP7_75t_L g1217 ( 
.A(n_1073),
.B(n_1048),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1071),
.A2(n_1069),
.B1(n_1083),
.B2(n_1118),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1093),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1150),
.Y(n_1220)
);

INVx3_ASAP7_75t_SL g1221 ( 
.A(n_1057),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1152),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1082),
.Y(n_1223)
);

AO21x1_ASAP7_75t_L g1224 ( 
.A1(n_1068),
.A2(n_1069),
.B(n_1114),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1051),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_SL g1226 ( 
.A1(n_1089),
.A2(n_1081),
.B1(n_1166),
.B2(n_1158),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1115),
.B(n_1119),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1052),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_1087),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1094),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1055),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1049),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1101),
.Y(n_1233)
);

OAI21xp33_ASAP7_75t_L g1234 ( 
.A1(n_1058),
.A2(n_1068),
.B(n_1104),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1122),
.B(n_1063),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1166),
.B(n_1045),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1106),
.Y(n_1237)
);

AO21x1_ASAP7_75t_L g1238 ( 
.A1(n_1123),
.A2(n_1100),
.B(n_1097),
.Y(n_1238)
);

INVx4_ASAP7_75t_L g1239 ( 
.A(n_1049),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1107),
.B(n_1111),
.Y(n_1240)
);

BUFx2_ASAP7_75t_R g1241 ( 
.A(n_1108),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_SL g1242 ( 
.A1(n_1081),
.A2(n_1089),
.B1(n_1159),
.B2(n_1158),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1049),
.Y(n_1243)
);

AO21x1_ASAP7_75t_L g1244 ( 
.A1(n_1123),
.A2(n_1100),
.B(n_1097),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1112),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1155),
.A2(n_1086),
.B1(n_1078),
.B2(n_1095),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_SL g1247 ( 
.A1(n_1159),
.A2(n_1170),
.B1(n_1110),
.B2(n_1098),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1088),
.A2(n_1109),
.B1(n_1167),
.B2(n_1102),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1096),
.B(n_1121),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1117),
.Y(n_1250)
);

NAND2x1p5_ASAP7_75t_L g1251 ( 
.A(n_1131),
.B(n_1117),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1116),
.B(n_1096),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1090),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1167),
.A2(n_1126),
.B1(n_1124),
.B2(n_1127),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1120),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1124),
.B(n_1173),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1103),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1125),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1149),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1129),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_1103),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1160),
.A2(n_1126),
.B1(n_1105),
.B2(n_1103),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1129),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1138),
.Y(n_1264)
);

INVx11_ASAP7_75t_L g1265 ( 
.A(n_1163),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1130),
.A2(n_1163),
.B1(n_1171),
.B2(n_1132),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1171),
.B(n_1128),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1040),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1113),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1113),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1040),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1044),
.B(n_1084),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1062),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1040),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1040),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1040),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1050),
.B(n_1041),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1039),
.Y(n_1278)
);

NAND2x1p5_ASAP7_75t_L g1279 ( 
.A(n_1099),
.B(n_1113),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1040),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1039),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1040),
.Y(n_1282)
);

INVx6_ASAP7_75t_L g1283 ( 
.A(n_1077),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1184),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1203),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1256),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1227),
.B(n_1179),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1273),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1238),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1227),
.B(n_1179),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1238),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1244),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1250),
.B(n_1258),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1199),
.B(n_1212),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1244),
.Y(n_1295)
);

OR2x2_ASAP7_75t_L g1296 ( 
.A(n_1249),
.B(n_1269),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_SL g1297 ( 
.A(n_1241),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1269),
.B(n_1270),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1255),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1255),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1190),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1240),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1213),
.B(n_1215),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1270),
.B(n_1235),
.Y(n_1304)
);

AO31x2_ASAP7_75t_L g1305 ( 
.A1(n_1224),
.A2(n_1195),
.A3(n_1209),
.B(n_1258),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1174),
.B(n_1183),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1190),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1236),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1250),
.B(n_1256),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1235),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1224),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1236),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1183),
.B(n_1252),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1195),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1252),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1194),
.Y(n_1316)
);

AOI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1178),
.A2(n_1277),
.B1(n_1182),
.B2(n_1216),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1182),
.B(n_1277),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1175),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1207),
.B(n_1211),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1279),
.B(n_1186),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1180),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1181),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1188),
.B(n_1178),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1231),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1279),
.B(n_1219),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_SL g1327 ( 
.A(n_1222),
.B(n_1228),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1234),
.B(n_1176),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1185),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1187),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1191),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1279),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1204),
.A2(n_1218),
.B(n_1248),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1202),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1192),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1193),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1242),
.A2(n_1246),
.B1(n_1272),
.B2(n_1176),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1225),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1268),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1189),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1271),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1274),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1267),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1251),
.Y(n_1344)
);

AO21x2_ASAP7_75t_L g1345 ( 
.A1(n_1204),
.A2(n_1263),
.B(n_1260),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1275),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1276),
.B(n_1280),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1282),
.Y(n_1348)
);

INVx2_ASAP7_75t_SL g1349 ( 
.A(n_1283),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1176),
.B(n_1210),
.Y(n_1350)
);

AOI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1263),
.A2(n_1237),
.B(n_1245),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1254),
.B(n_1226),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1210),
.B(n_1272),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1239),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1210),
.B(n_1272),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1223),
.B(n_1230),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1202),
.Y(n_1357)
);

BUFx6f_ASAP7_75t_L g1358 ( 
.A(n_1239),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1286),
.B(n_1233),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1347),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_1284),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1285),
.B(n_1214),
.Y(n_1362)
);

AOI222xp33_ASAP7_75t_L g1363 ( 
.A1(n_1333),
.A2(n_1201),
.B1(n_1177),
.B2(n_1221),
.C1(n_1228),
.C2(n_1222),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1309),
.B(n_1239),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1308),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1308),
.B(n_1266),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1304),
.B(n_1259),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1288),
.B(n_1313),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1351),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1308),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1312),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1313),
.B(n_1208),
.Y(n_1372)
);

NAND3xp33_ASAP7_75t_L g1373 ( 
.A(n_1317),
.B(n_1247),
.C(n_1217),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1351),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1316),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1310),
.B(n_1315),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1296),
.B(n_1200),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1324),
.B(n_1221),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1319),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1296),
.B(n_1206),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1327),
.B(n_1220),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1294),
.B(n_1281),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1301),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1287),
.B(n_1278),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1319),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1290),
.B(n_1309),
.Y(n_1386)
);

AOI221xp5_ASAP7_75t_L g1387 ( 
.A1(n_1306),
.A2(n_1198),
.B1(n_1205),
.B2(n_1197),
.C(n_1220),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1298),
.B(n_1205),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1298),
.B(n_1197),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1307),
.B(n_1264),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1303),
.A2(n_1201),
.B1(n_1196),
.B2(n_1177),
.Y(n_1391)
);

OAI221xp5_ASAP7_75t_L g1392 ( 
.A1(n_1317),
.A2(n_1262),
.B1(n_1253),
.B2(n_1243),
.C(n_1232),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1326),
.B(n_1302),
.Y(n_1393)
);

INVxp67_ASAP7_75t_SL g1394 ( 
.A(n_1325),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1334),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1289),
.B(n_1257),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1365),
.B(n_1291),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1386),
.B(n_1291),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1386),
.B(n_1292),
.Y(n_1399)
);

OAI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1363),
.A2(n_1337),
.B1(n_1328),
.B2(n_1343),
.C(n_1338),
.Y(n_1400)
);

NAND3xp33_ASAP7_75t_SL g1401 ( 
.A(n_1363),
.B(n_1343),
.C(n_1352),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1373),
.A2(n_1297),
.B1(n_1318),
.B2(n_1352),
.Y(n_1402)
);

NAND3xp33_ASAP7_75t_L g1403 ( 
.A(n_1373),
.B(n_1311),
.C(n_1314),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1361),
.B(n_1326),
.Y(n_1404)
);

AOI221xp5_ASAP7_75t_L g1405 ( 
.A1(n_1387),
.A2(n_1318),
.B1(n_1320),
.B2(n_1311),
.C(n_1314),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1368),
.B(n_1299),
.Y(n_1406)
);

AND2x2_ASAP7_75t_SL g1407 ( 
.A(n_1364),
.B(n_1332),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1394),
.B(n_1383),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1393),
.B(n_1295),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1365),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1365),
.B(n_1295),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1375),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1388),
.B(n_1300),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1388),
.B(n_1300),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1378),
.B(n_1321),
.C(n_1340),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1370),
.B(n_1332),
.Y(n_1416)
);

NAND3xp33_ASAP7_75t_L g1417 ( 
.A(n_1382),
.B(n_1340),
.C(n_1336),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1389),
.B(n_1322),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1389),
.B(n_1323),
.Y(n_1419)
);

AOI221xp5_ASAP7_75t_L g1420 ( 
.A1(n_1362),
.A2(n_1323),
.B1(n_1329),
.B2(n_1330),
.C(n_1348),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1370),
.B(n_1345),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_1381),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1391),
.B(n_1350),
.Y(n_1423)
);

OAI21xp33_ASAP7_75t_L g1424 ( 
.A1(n_1372),
.A2(n_1347),
.B(n_1356),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1359),
.B(n_1329),
.Y(n_1425)
);

OAI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1392),
.A2(n_1358),
.B1(n_1354),
.B2(n_1349),
.Y(n_1426)
);

OAI221xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1366),
.A2(n_1357),
.B1(n_1335),
.B2(n_1330),
.C(n_1346),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1359),
.B(n_1331),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1364),
.B(n_1353),
.Y(n_1429)
);

NAND3xp33_ASAP7_75t_L g1430 ( 
.A(n_1390),
.B(n_1342),
.C(n_1335),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1371),
.B(n_1345),
.Y(n_1431)
);

NOR2x1_ASAP7_75t_L g1432 ( 
.A(n_1369),
.B(n_1344),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1371),
.B(n_1345),
.Y(n_1433)
);

NAND3xp33_ASAP7_75t_L g1434 ( 
.A(n_1395),
.B(n_1341),
.C(n_1331),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1377),
.A2(n_1261),
.B1(n_1354),
.B2(n_1358),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1364),
.A2(n_1353),
.B1(n_1355),
.B2(n_1293),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1377),
.B(n_1336),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1380),
.A2(n_1261),
.B1(n_1354),
.B2(n_1229),
.Y(n_1438)
);

NAND3xp33_ASAP7_75t_L g1439 ( 
.A(n_1396),
.B(n_1342),
.C(n_1339),
.Y(n_1439)
);

OAI221xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1380),
.A2(n_1357),
.B1(n_1341),
.B2(n_1339),
.C(n_1348),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1384),
.B(n_1346),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1412),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1412),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1411),
.B(n_1305),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1397),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1432),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1410),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1409),
.B(n_1305),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1398),
.B(n_1399),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1410),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1421),
.B(n_1379),
.Y(n_1451)
);

NOR2x1_ASAP7_75t_L g1452 ( 
.A(n_1403),
.B(n_1374),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1425),
.B(n_1305),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1416),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1431),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1433),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1437),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1432),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1428),
.B(n_1305),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1406),
.B(n_1441),
.Y(n_1460)
);

INVx4_ASAP7_75t_L g1461 ( 
.A(n_1407),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1418),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1424),
.B(n_1305),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1419),
.B(n_1385),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1413),
.Y(n_1465)
);

NAND3xp33_ASAP7_75t_L g1466 ( 
.A(n_1452),
.B(n_1403),
.C(n_1405),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1442),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1442),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1442),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1444),
.B(n_1408),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1443),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1443),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_SL g1473 ( 
.A(n_1461),
.B(n_1422),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1458),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1461),
.B(n_1429),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_1460),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1461),
.B(n_1439),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1443),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1445),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1451),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1457),
.B(n_1424),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1445),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1460),
.B(n_1422),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1461),
.B(n_1404),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1451),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1445),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1447),
.Y(n_1487)
);

AOI33xp33_ASAP7_75t_L g1488 ( 
.A1(n_1457),
.A2(n_1426),
.A3(n_1420),
.B1(n_1360),
.B2(n_1376),
.B3(n_1367),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1444),
.B(n_1448),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1457),
.B(n_1414),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1458),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1447),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1461),
.B(n_1360),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1465),
.B(n_1415),
.Y(n_1494)
);

INVx3_ASAP7_75t_L g1495 ( 
.A(n_1451),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1465),
.B(n_1430),
.Y(n_1496)
);

INVxp67_ASAP7_75t_SL g1497 ( 
.A(n_1452),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1450),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1465),
.B(n_1423),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1450),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1496),
.B(n_1453),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1475),
.B(n_1446),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1467),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1499),
.B(n_1462),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1476),
.B(n_1462),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1475),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1475),
.B(n_1449),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1467),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1468),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1468),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_R g1511 ( 
.A(n_1473),
.B(n_1229),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1469),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1488),
.B(n_1462),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1494),
.B(n_1453),
.Y(n_1514)
);

INVxp67_ASAP7_75t_L g1515 ( 
.A(n_1483),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1481),
.B(n_1462),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1471),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1471),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1484),
.B(n_1449),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1493),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1484),
.B(n_1449),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1466),
.B(n_1465),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1470),
.B(n_1459),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1472),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1479),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1477),
.A2(n_1401),
.B1(n_1402),
.B2(n_1400),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1469),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1490),
.B(n_1459),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1472),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1478),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1477),
.A2(n_1364),
.B1(n_1463),
.B2(n_1435),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1479),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1477),
.B(n_1493),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1470),
.B(n_1448),
.Y(n_1534)
);

NAND2xp67_ASAP7_75t_L g1535 ( 
.A(n_1480),
.B(n_1458),
.Y(n_1535)
);

OAI32xp33_ASAP7_75t_L g1536 ( 
.A1(n_1489),
.A2(n_1463),
.A3(n_1458),
.B1(n_1456),
.B2(n_1455),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1477),
.B(n_1455),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1497),
.B(n_1464),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1482),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1489),
.B(n_1464),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1482),
.B(n_1454),
.Y(n_1541)
);

NAND2x1p5_ASAP7_75t_L g1542 ( 
.A(n_1495),
.B(n_1446),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1486),
.B(n_1196),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1525),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1532),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1526),
.A2(n_1427),
.B1(n_1440),
.B2(n_1430),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1502),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1539),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1512),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1503),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1507),
.B(n_1495),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1507),
.B(n_1533),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_1511),
.Y(n_1553)
);

OR2x6_ASAP7_75t_L g1554 ( 
.A(n_1506),
.B(n_1446),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1522),
.B(n_1486),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1513),
.B(n_1478),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1511),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1508),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1506),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1512),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1504),
.B(n_1498),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1516),
.B(n_1498),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1509),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1533),
.B(n_1495),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1510),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1517),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1519),
.B(n_1480),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1527),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1515),
.B(n_1543),
.Y(n_1569)
);

INVx2_ASAP7_75t_SL g1570 ( 
.A(n_1502),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1543),
.B(n_1464),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1518),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1519),
.B(n_1521),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1521),
.B(n_1485),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1524),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1528),
.B(n_1454),
.Y(n_1576)
);

INVxp67_ASAP7_75t_R g1577 ( 
.A(n_1537),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1502),
.B(n_1485),
.Y(n_1578)
);

AND3x1_ASAP7_75t_L g1579 ( 
.A(n_1531),
.B(n_1491),
.C(n_1474),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1553),
.B(n_1528),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1556),
.B(n_1514),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1553),
.B(n_1514),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1544),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1550),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1559),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1577),
.B(n_1520),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1557),
.B(n_1520),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1569),
.B(n_1552),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1550),
.Y(n_1589)
);

AOI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1546),
.A2(n_1536),
.B1(n_1538),
.B2(n_1501),
.C(n_1537),
.Y(n_1590)
);

OAI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1546),
.A2(n_1542),
.B(n_1501),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1558),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1559),
.Y(n_1593)
);

OAI322xp33_ASAP7_75t_L g1594 ( 
.A1(n_1556),
.A2(n_1542),
.A3(n_1523),
.B1(n_1534),
.B2(n_1505),
.C1(n_1529),
.C2(n_1530),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1552),
.B(n_1540),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1577),
.B(n_1534),
.Y(n_1596)
);

INVx2_ASAP7_75t_SL g1597 ( 
.A(n_1559),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1547),
.B(n_1196),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1547),
.B(n_1523),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1554),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1573),
.B(n_1527),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1558),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1563),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1579),
.A2(n_1436),
.B1(n_1541),
.B2(n_1417),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1563),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1580),
.B(n_1570),
.Y(n_1606)
);

NOR3xp33_ASAP7_75t_SL g1607 ( 
.A(n_1587),
.B(n_1548),
.C(n_1545),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1593),
.B(n_1570),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1584),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1586),
.B(n_1573),
.Y(n_1610)
);

INVxp67_ASAP7_75t_L g1611 ( 
.A(n_1597),
.Y(n_1611)
);

INVx2_ASAP7_75t_SL g1612 ( 
.A(n_1597),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1585),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1588),
.B(n_1583),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1585),
.B(n_1545),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1584),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1582),
.B(n_1571),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1602),
.Y(n_1618)
);

OAI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1591),
.A2(n_1554),
.B1(n_1548),
.B2(n_1555),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1596),
.B(n_1555),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1596),
.B(n_1565),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1595),
.B(n_1576),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1602),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1601),
.B(n_1565),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1601),
.B(n_1566),
.Y(n_1625)
);

AOI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1607),
.A2(n_1594),
.B1(n_1590),
.B2(n_1579),
.C(n_1604),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1607),
.A2(n_1619),
.B1(n_1611),
.B2(n_1606),
.Y(n_1627)
);

AOI211x1_ASAP7_75t_L g1628 ( 
.A1(n_1619),
.A2(n_1586),
.B(n_1599),
.C(n_1603),
.Y(n_1628)
);

OAI211xp5_ASAP7_75t_SL g1629 ( 
.A1(n_1614),
.A2(n_1592),
.B(n_1589),
.C(n_1605),
.Y(n_1629)
);

AOI21xp33_ASAP7_75t_L g1630 ( 
.A1(n_1611),
.A2(n_1600),
.B(n_1598),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1620),
.A2(n_1600),
.B(n_1605),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1610),
.A2(n_1578),
.B1(n_1564),
.B2(n_1581),
.Y(n_1632)
);

NAND2xp33_ASAP7_75t_R g1633 ( 
.A(n_1608),
.B(n_1581),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1617),
.B(n_1561),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1612),
.Y(n_1635)
);

INVxp67_ASAP7_75t_L g1636 ( 
.A(n_1633),
.Y(n_1636)
);

NAND2x1_ASAP7_75t_SL g1637 ( 
.A(n_1635),
.B(n_1613),
.Y(n_1637)
);

NAND3xp33_ASAP7_75t_SL g1638 ( 
.A(n_1626),
.B(n_1621),
.C(n_1615),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1628),
.B(n_1624),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1627),
.B(n_1625),
.Y(n_1640)
);

NOR2x1_ASAP7_75t_L g1641 ( 
.A(n_1629),
.B(n_1609),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1632),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1634),
.B(n_1622),
.Y(n_1643)
);

NOR2x1_ASAP7_75t_L g1644 ( 
.A(n_1631),
.B(n_1616),
.Y(n_1644)
);

NAND4xp25_ASAP7_75t_SL g1645 ( 
.A(n_1639),
.B(n_1630),
.C(n_1623),
.D(n_1618),
.Y(n_1645)
);

O2A1O1Ixp33_ASAP7_75t_L g1646 ( 
.A1(n_1636),
.A2(n_1554),
.B(n_1575),
.C(n_1572),
.Y(n_1646)
);

O2A1O1Ixp33_ASAP7_75t_L g1647 ( 
.A1(n_1638),
.A2(n_1640),
.B(n_1644),
.C(n_1641),
.Y(n_1647)
);

NOR4xp75_ASAP7_75t_L g1648 ( 
.A(n_1637),
.B(n_1564),
.C(n_1578),
.D(n_1551),
.Y(n_1648)
);

NAND4xp25_ASAP7_75t_L g1649 ( 
.A(n_1642),
.B(n_1575),
.C(n_1566),
.D(n_1572),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1646),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1649),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1648),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1645),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1647),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1648),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1651),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1654),
.Y(n_1657)
);

NOR3xp33_ASAP7_75t_L g1658 ( 
.A(n_1653),
.B(n_1643),
.C(n_1560),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1652),
.Y(n_1659)
);

NAND4xp25_ASAP7_75t_L g1660 ( 
.A(n_1655),
.B(n_1560),
.C(n_1549),
.D(n_1568),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1657),
.A2(n_1654),
.B(n_1650),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1659),
.Y(n_1662)
);

NOR3xp33_ASAP7_75t_L g1663 ( 
.A(n_1656),
.B(n_1652),
.C(n_1560),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1662),
.A2(n_1658),
.B1(n_1554),
.B2(n_1549),
.Y(n_1664)
);

OAI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1664),
.A2(n_1660),
.B1(n_1661),
.B2(n_1554),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1665),
.A2(n_1663),
.B1(n_1549),
.B2(n_1568),
.Y(n_1666)
);

AO21x2_ASAP7_75t_L g1667 ( 
.A1(n_1665),
.A2(n_1568),
.B(n_1551),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1667),
.A2(n_1561),
.B1(n_1562),
.B2(n_1567),
.Y(n_1668)
);

OAI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1666),
.A2(n_1562),
.B(n_1567),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1668),
.B(n_1574),
.Y(n_1670)
);

AOI21xp33_ASAP7_75t_L g1671 ( 
.A1(n_1669),
.A2(n_1253),
.B(n_1574),
.Y(n_1671)
);

OAI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1670),
.A2(n_1491),
.B(n_1474),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1672),
.A2(n_1671),
.B1(n_1492),
.B2(n_1487),
.Y(n_1673)
);

OAI221xp5_ASAP7_75t_R g1674 ( 
.A1(n_1673),
.A2(n_1535),
.B1(n_1265),
.B2(n_1500),
.C(n_1492),
.Y(n_1674)
);

AOI211xp5_ASAP7_75t_L g1675 ( 
.A1(n_1674),
.A2(n_1434),
.B(n_1500),
.C(n_1438),
.Y(n_1675)
);


endmodule