module fake_jpeg_19113_n_148 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_SL g48 ( 
.A(n_5),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_21),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_26),
.Y(n_64)
);

INVx8_ASAP7_75t_SL g65 ( 
.A(n_47),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_6),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_6),
.Y(n_71)
);

INVx11_ASAP7_75t_SL g72 ( 
.A(n_2),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_31),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_0),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_28),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_76),
.B(n_82),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_80),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_1),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_30),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_82),
.A2(n_73),
.B1(n_49),
.B2(n_66),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_89),
.B1(n_63),
.B2(n_69),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_52),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_73),
.B1(n_49),
.B2(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_91),
.B(n_93),
.Y(n_98)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_90),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_100),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_72),
.B1(n_58),
.B2(n_65),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_71),
.B1(n_74),
.B2(n_54),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_96),
.A2(n_97),
.B1(n_105),
.B2(n_57),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_50),
.B1(n_53),
.B2(n_64),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_69),
.B1(n_62),
.B2(n_60),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_70),
.B1(n_55),
.B2(n_83),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_62),
.B1(n_59),
.B2(n_56),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_59),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_3),
.Y(n_113)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_111),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_114),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_35),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_123),
.Y(n_124)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_117),
.B(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_10),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_11),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_108),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_37),
.B1(n_14),
.B2(n_16),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_36),
.B(n_38),
.C(n_40),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_39),
.B1(n_20),
.B2(n_25),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_11),
.B(n_33),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_131),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_123),
.Y(n_134)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_133),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_126),
.B(n_112),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_124),
.C(n_115),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_139),
.A2(n_124),
.B1(n_138),
.B2(n_135),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_136),
.B1(n_129),
.B2(n_128),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_141),
.A2(n_128),
.B1(n_131),
.B2(n_132),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_116),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_121),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_122),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_122),
.C(n_42),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_41),
.C(n_43),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_45),
.Y(n_148)
);


endmodule