module fake_jpeg_3168_n_43 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_43);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_15;

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_10),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_12),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_18),
.Y(n_22)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

NAND2x1_ASAP7_75t_SL g19 ( 
.A(n_15),
.B(n_0),
.Y(n_19)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_12),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_15),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_22),
.A2(n_15),
.B1(n_14),
.B2(n_16),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_26),
.B1(n_19),
.B2(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_18),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_18),
.B1(n_19),
.B2(n_14),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_19),
.C(n_16),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_30),
.C(n_11),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_26),
.B1(n_13),
.B2(n_16),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_14),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_13),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_35),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_13),
.B(n_4),
.Y(n_33)
);

OAI21x1_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_34),
.B(n_3),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_7),
.Y(n_40)
);

A2O1A1O1Ixp25_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_9),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_3),
.B(n_5),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_40),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_41),
.B(n_38),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_7),
.B1(n_8),
.B2(n_25),
.Y(n_43)
);


endmodule