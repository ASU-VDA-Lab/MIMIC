module real_jpeg_26834_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_80;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_244;
wire n_128;
wire n_213;
wire n_202;
wire n_179;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_SL g60 ( 
.A(n_0),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_1),
.Y(n_119)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_1),
.Y(n_136)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_4),
.A2(n_9),
.B1(n_24),
.B2(n_28),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_4),
.A2(n_28),
.B1(n_58),
.B2(n_59),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_4),
.A2(n_28),
.B1(n_41),
.B2(n_43),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_6),
.A2(n_41),
.B1(n_43),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_6),
.A2(n_9),
.B1(n_24),
.B2(n_62),
.Y(n_100)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_8),
.A2(n_9),
.B1(n_24),
.B2(n_31),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_8),
.A2(n_31),
.B1(n_41),
.B2(n_43),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_SL g115 ( 
.A1(n_8),
.A2(n_9),
.B(n_23),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_8),
.A2(n_31),
.B1(n_58),
.B2(n_59),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_8),
.B(n_21),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_SL g160 ( 
.A1(n_8),
.A2(n_10),
.B(n_41),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_8),
.A2(n_55),
.B(n_59),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_8),
.B(n_40),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_9),
.A2(n_11),
.B1(n_24),
.B2(n_39),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_9),
.A2(n_10),
.B1(n_24),
.B2(n_42),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_9),
.A2(n_31),
.B(n_159),
.C(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_10),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_11),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_11),
.A2(n_39),
.B1(n_58),
.B2(n_59),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_103),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_102),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_89),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_16),
.B(n_89),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_63),
.C(n_71),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_17),
.B(n_63),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_34),
.B2(n_35),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_18),
.A2(n_19),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_18),
.A2(n_19),
.B1(n_143),
.B2(n_145),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_18),
.A2(n_19),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_18),
.B(n_223),
.C(n_225),
.Y(n_243)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_19),
.B(n_37),
.C(n_49),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_19),
.B(n_123),
.C(n_124),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_25),
.B(n_29),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_21),
.B(n_32),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_21),
.A2(n_30),
.B1(n_32),
.B2(n_95),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_22),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_22),
.A2(n_27),
.B(n_31),
.C(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_30),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_31),
.A2(n_41),
.B(n_56),
.C(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_31),
.B(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_31),
.B(n_57),
.Y(n_198)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_49),
.B2(n_50),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_40),
.B(n_44),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_38),
.A2(n_40),
.B1(n_47),
.B2(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_40),
.B(n_47),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_45),
.A2(n_68),
.B(n_70),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_49),
.A2(n_50),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_61),
.Y(n_50)
);

INVxp33_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_52),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_53),
.A2(n_57),
.B1(n_61),
.B2(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_53),
.A2(n_57),
.B1(n_84),
.B2(n_132),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_65),
.B(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_58),
.B(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_78),
.Y(n_77)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_63),
.A2(n_64),
.B(n_66),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_66),
.A2(n_93),
.B1(n_94),
.B2(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_66),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_66),
.B(n_149),
.C(n_150),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_66),
.A2(n_111),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_69),
.B(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_71),
.A2(n_72),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_80),
.B(n_85),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_73),
.A2(n_81),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_73),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_73),
.A2(n_85),
.B1(n_86),
.B2(n_241),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_74),
.A2(n_77),
.B1(n_119),
.B2(n_137),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_76),
.B(n_140),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_77),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_80),
.B(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_81),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_83),
.A2(n_131),
.B(n_133),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_101),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_93),
.A2(n_94),
.B1(n_123),
.B2(n_144),
.Y(n_238)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_94),
.B(n_111),
.C(n_112),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_94),
.B(n_144),
.C(n_237),
.Y(n_253)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_256),
.B(n_261),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_245),
.B(n_255),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_231),
.B(n_244),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_152),
.B(n_214),
.C(n_230),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_141),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_108),
.B(n_141),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_120),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_109),
.B(n_121),
.C(n_128),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_116),
.A2(n_147),
.B1(n_183),
.B2(n_186),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_116),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_116),
.B(n_198),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_116),
.B(n_173),
.C(n_185),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_117),
.A2(n_119),
.B(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

INVx11_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_127),
.B2(n_128),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_123),
.A2(n_129),
.B1(n_130),
.B2(n_144),
.Y(n_205)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_134),
.B2(n_135),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_129),
.A2(n_130),
.B1(n_180),
.B2(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_129),
.B(n_135),
.Y(n_223)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_144),
.C(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_130),
.B(n_180),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B(n_138),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.C(n_148),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_142),
.B(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_143),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_146),
.B(n_148),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_149),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_213),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_208),
.B(n_212),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_176),
.B(n_207),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_164),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_156),
.B(n_164),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_158),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_163),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_170),
.B2(n_171),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_173),
.C(n_174),
.Y(n_209)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_167),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_168),
.B(n_189),
.Y(n_200)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_172),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_175),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_173),
.A2(n_175),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_173),
.B(n_220),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_202),
.B(n_206),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_187),
.B(n_201),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_182),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_180),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_183),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_184),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_191),
.B(n_200),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_197),
.B(n_199),
.Y(n_191)
);

INVx5_ASAP7_75t_SL g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_204),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_210),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_215),
.B(n_216),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_228),
.B2(n_229),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_222),
.C(n_229),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_220),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_228),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_232),
.B(n_233),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_243),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_240),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_240),
.C(n_243),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_246),
.B(n_247),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_253),
.B2(n_254),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_251),
.C(n_254),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_253),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_257),
.B(n_258),
.Y(n_261)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_259),
.Y(n_260)
);


endmodule