module fake_jpeg_25943_n_229 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_41),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_0),
.C(n_1),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_26),
.B1(n_22),
.B2(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_28),
.B1(n_27),
.B2(n_30),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_54),
.B1(n_41),
.B2(n_16),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_55),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_28),
.B1(n_18),
.B2(n_27),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_43),
.B1(n_24),
.B2(n_32),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_28),
.B1(n_30),
.B2(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_22),
.Y(n_64)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_66),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_61),
.A2(n_68),
.B1(n_26),
.B2(n_22),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_42),
.C(n_35),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_71),
.C(n_75),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_64),
.A2(n_38),
.B(n_34),
.C(n_19),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_76),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_23),
.C(n_31),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_21),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_73),
.B(n_77),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_31),
.C(n_20),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_21),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_78),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_79),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_45),
.C(n_58),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_71),
.C(n_68),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_51),
.B(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_82),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_17),
.B(n_16),
.C(n_32),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_26),
.B(n_1),
.Y(n_113)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_22),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_94),
.B(n_113),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_31),
.B1(n_20),
.B2(n_24),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_96),
.A2(n_104),
.B1(n_107),
.B2(n_29),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_31),
.B1(n_20),
.B2(n_38),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_87),
.B1(n_69),
.B2(n_82),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_92),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_60),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_111),
.Y(n_115)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_38),
.B1(n_19),
.B2(n_29),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_72),
.B1(n_86),
.B2(n_84),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_111),
.A2(n_84),
.B1(n_65),
.B2(n_105),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_116),
.A2(n_137),
.B1(n_132),
.B2(n_118),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_130),
.B1(n_135),
.B2(n_107),
.Y(n_146)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_119),
.B(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_126),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_103),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_123),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_88),
.C(n_67),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_136),
.C(n_96),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_102),
.B(n_14),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_131),
.B(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_134),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_78),
.B1(n_74),
.B2(n_19),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_93),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_138),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_92),
.B(n_29),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_108),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_154),
.C(n_2),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_142),
.B(n_151),
.Y(n_174)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_158),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_2),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_113),
.B(n_104),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_115),
.A2(n_98),
.B(n_106),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_153),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_98),
.B(n_110),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_114),
.C(n_110),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_93),
.B1(n_112),
.B2(n_3),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_122),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_0),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_130),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_161),
.Y(n_172)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_165),
.B(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_125),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_169),
.B(n_170),
.Y(n_189)
);

AO22x1_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_153),
.B1(n_146),
.B2(n_137),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_147),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_171),
.A2(n_176),
.B1(n_177),
.B2(n_149),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_178),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_160),
.C(n_142),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_156),
.B(n_10),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_3),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_172),
.A2(n_154),
.B1(n_159),
.B2(n_143),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_180),
.A2(n_192),
.B1(n_179),
.B2(n_164),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_175),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_185),
.Y(n_196)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_147),
.B1(n_143),
.B2(n_145),
.Y(n_187)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_170),
.A2(n_157),
.B1(n_158),
.B2(n_152),
.Y(n_190)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_191)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

OAI22x1_ASAP7_75t_L g192 ( 
.A1(n_163),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_188),
.A2(n_174),
.B1(n_192),
.B2(n_189),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_182),
.Y(n_211)
);

XOR2x2_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_168),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_183),
.B(n_200),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_181),
.A2(n_166),
.B(n_168),
.C(n_167),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_200),
.Y(n_209)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_202),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_180),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_178),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_211),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_207),
.A2(n_208),
.B(n_197),
.Y(n_217)
);

NOR3xp33_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_186),
.C(n_173),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_203),
.B(n_179),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_210),
.B(n_209),
.Y(n_214)
);

AOI21x1_ASAP7_75t_SL g213 ( 
.A1(n_205),
.A2(n_202),
.B(n_195),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_217),
.B(n_6),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_215),
.Y(n_221)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_194),
.C(n_196),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

NOR2x1_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_198),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_9),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_220),
.A2(n_215),
.B1(n_212),
.B2(n_8),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_223),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_212),
.C(n_7),
.Y(n_223)
);

OAI21x1_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_6),
.B(n_7),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_226),
.C(n_223),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_219),
.Y(n_229)
);


endmodule