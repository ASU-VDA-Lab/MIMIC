module fake_jpeg_9497_n_64 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_64);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_64;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_5),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_0),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_28),
.B(n_9),
.C(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_18),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_25),
.A2(n_14),
.B1(n_24),
.B2(n_3),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_7),
.B1(n_12),
.B2(n_13),
.Y(n_48)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_30),
.Y(n_47)
);

NOR2x1_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_1),
.C(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_55)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_22),
.Y(n_53)
);

MAJx2_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_16),
.C(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_51),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.B(n_56),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_55),
.C(n_54),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_53),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_SL g64 ( 
.A1(n_63),
.A2(n_57),
.B(n_42),
.C(n_41),
.Y(n_64)
);


endmodule