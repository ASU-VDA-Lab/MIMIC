module fake_jpeg_15908_n_47 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx11_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx12_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

HAxp5_ASAP7_75t_SL g15 ( 
.A(n_10),
.B(n_0),
.CON(n_15),
.SN(n_15)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_15),
.A2(n_18),
.B1(n_7),
.B2(n_4),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_22),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_11),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_11),
.A2(n_7),
.B1(n_9),
.B2(n_14),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_19),
.A2(n_13),
.B1(n_23),
.B2(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_15),
.B(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_21),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_30),
.C(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_34),
.B(n_38),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_37),
.B(n_24),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_32),
.C(n_29),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_40),
.C(n_34),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_43),
.B(n_44),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

AOI221xp5_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_28),
.B1(n_33),
.B2(n_41),
.C(n_45),
.Y(n_47)
);


endmodule