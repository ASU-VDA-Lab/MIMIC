module fake_jpeg_22978_n_346 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_41),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

CKINVDCx6p67_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_44),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_46),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_37),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_31),
.B1(n_35),
.B2(n_47),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_65),
.B1(n_22),
.B2(n_23),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_31),
.B1(n_47),
.B2(n_35),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_31),
.B1(n_35),
.B2(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_60),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_31),
.B1(n_35),
.B2(n_47),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

OR2x2_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_40),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_71),
.A2(n_26),
.B1(n_17),
.B2(n_32),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_72),
.A2(n_21),
.B1(n_36),
.B2(n_19),
.Y(n_112)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_76),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_26),
.B1(n_25),
.B2(n_22),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_75),
.A2(n_90),
.B(n_103),
.Y(n_117)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_84),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_85),
.B1(n_87),
.B2(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_46),
.B(n_44),
.C(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_81),
.B(n_93),
.Y(n_123)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_25),
.B1(n_46),
.B2(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_86),
.B(n_92),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_54),
.A2(n_40),
.B1(n_45),
.B2(n_38),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_96),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_26),
.B1(n_25),
.B2(n_19),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_40),
.B1(n_45),
.B2(n_38),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_53),
.B(n_41),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_42),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_102),
.Y(n_116)
);

AO22x1_ASAP7_75t_SL g98 ( 
.A1(n_59),
.A2(n_38),
.B1(n_48),
.B2(n_42),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_51),
.B1(n_45),
.B2(n_64),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_42),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_60),
.A2(n_26),
.B1(n_36),
.B2(n_22),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_0),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_105),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_0),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_122),
.B1(n_126),
.B2(n_128),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_112),
.A2(n_121),
.B1(n_135),
.B2(n_77),
.Y(n_136)
);

FAx1_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_42),
.CI(n_39),
.CON(n_113),
.SN(n_113)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_113),
.B(n_82),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_44),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_34),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_39),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_131),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_79),
.A2(n_91),
.B1(n_87),
.B2(n_71),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_81),
.A2(n_98),
.B1(n_102),
.B2(n_96),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_36),
.B(n_23),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_124),
.A2(n_125),
.B(n_134),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_19),
.B(n_23),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_84),
.A2(n_41),
.B1(n_28),
.B2(n_21),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_92),
.A2(n_28),
.B1(n_33),
.B2(n_29),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g145 ( 
.A1(n_130),
.A2(n_17),
.B(n_32),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_28),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_1),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_97),
.A2(n_26),
.B1(n_21),
.B2(n_28),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_141),
.B1(n_145),
.B2(n_159),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_20),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_140),
.Y(n_170)
);

O2A1O1Ixp33_ASAP7_75t_SL g178 ( 
.A1(n_138),
.A2(n_166),
.B(n_115),
.C(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_117),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_139),
.B(n_152),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_109),
.B(n_99),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_121),
.A2(n_74),
.B1(n_73),
.B2(n_101),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_74),
.A3(n_21),
.B1(n_34),
.B2(n_83),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_126),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_143),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_108),
.A2(n_117),
.B1(n_118),
.B2(n_113),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_147),
.A2(n_132),
.B1(n_94),
.B2(n_114),
.Y(n_200)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_148),
.B(n_150),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_95),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_124),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_116),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_151),
.Y(n_185)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_154),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_17),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_106),
.B(n_101),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_160),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_100),
.Y(n_156)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_15),
.B(n_14),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_163),
.C(n_125),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_108),
.A2(n_86),
.B1(n_78),
.B2(n_18),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_158),
.A2(n_146),
.B1(n_135),
.B2(n_166),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_113),
.A2(n_33),
.B1(n_18),
.B2(n_32),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_119),
.B(n_18),
.Y(n_161)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_83),
.C(n_34),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_34),
.Y(n_164)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_131),
.C(n_123),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_167),
.B(n_179),
.C(n_198),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_168),
.A2(n_180),
.B1(n_142),
.B2(n_152),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_169),
.A2(n_165),
.B(n_163),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_111),
.B1(n_123),
.B2(n_113),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_200),
.B1(n_173),
.B2(n_196),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_176),
.B(n_187),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_178),
.A2(n_183),
.B(n_197),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_144),
.C(n_151),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_146),
.A2(n_130),
.B1(n_115),
.B2(n_107),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_139),
.A2(n_110),
.B(n_107),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_184),
.B(n_190),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_134),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_134),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_2),
.Y(n_224)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_192),
.Y(n_202)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_194),
.Y(n_207)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_137),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_195),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_153),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_144),
.B(n_128),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_129),
.Y(n_198)
);

NOR2x1_ASAP7_75t_L g199 ( 
.A(n_154),
.B(n_129),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_20),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_200),
.B(n_136),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_159),
.Y(n_203)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_206),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_226),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_181),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_208),
.B(n_225),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_150),
.B(n_160),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_209),
.A2(n_230),
.B(n_231),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_211),
.A2(n_222),
.B1(n_8),
.B2(n_14),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_212),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_114),
.Y(n_213)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_214),
.B(n_211),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_20),
.Y(n_215)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_168),
.A2(n_24),
.B1(n_33),
.B2(n_88),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_217),
.A2(n_199),
.B1(n_172),
.B2(n_170),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_182),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_218),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_24),
.Y(n_219)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_175),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_220),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_188),
.A2(n_24),
.B1(n_9),
.B2(n_11),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_189),
.B(n_174),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_224),
.Y(n_243)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_171),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_167),
.C(n_186),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_187),
.C(n_176),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_175),
.A2(n_2),
.B(n_3),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_180),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_234),
.B(n_237),
.C(n_251),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_244),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_213),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_236),
.B(n_245),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_184),
.C(n_173),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_240),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_178),
.B1(n_197),
.B2(n_169),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_242),
.A2(n_246),
.B1(n_247),
.B2(n_203),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_197),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_214),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_210),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_253),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_9),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_3),
.C(n_5),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_256),
.Y(n_260)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_261),
.B(n_266),
.Y(n_291)
);

XNOR2x1_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_206),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_278),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_248),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_264),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_216),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_267),
.A2(n_269),
.B(n_270),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_208),
.B1(n_220),
.B2(n_204),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_268),
.A2(n_277),
.B1(n_252),
.B2(n_222),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_257),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_274),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_218),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_247),
.C(n_244),
.Y(n_282)
);

AOI211xp5_ASAP7_75t_L g276 ( 
.A1(n_255),
.A2(n_228),
.B(n_209),
.C(n_216),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_243),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_255),
.A2(n_228),
.B(n_230),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_242),
.B(n_224),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_SL g280 ( 
.A1(n_269),
.A2(n_254),
.B(n_235),
.C(n_238),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_280),
.A2(n_293),
.B1(n_295),
.B2(n_13),
.Y(n_310)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_282),
.Y(n_304)
);

OAI21xp33_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_239),
.B(n_237),
.Y(n_283)
);

XNOR2x1_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_265),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_259),
.B(n_207),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_284),
.B(n_294),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_234),
.C(n_227),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_287),
.C(n_288),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_286),
.B(n_276),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_227),
.C(n_229),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_267),
.C(n_278),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_268),
.A2(n_217),
.B1(n_251),
.B2(n_240),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_258),
.B(n_233),
.Y(n_294)
);

OAI322xp33_ASAP7_75t_L g296 ( 
.A1(n_262),
.A2(n_243),
.A3(n_205),
.B1(n_12),
.B2(n_8),
.C1(n_11),
.C2(n_13),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_263),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_271),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_299),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_277),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_272),
.C(n_265),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_308),
.Y(n_312)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_302),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_303),
.A2(n_310),
.B1(n_286),
.B2(n_293),
.Y(n_314)
);

NOR2x1_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_270),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_305),
.A2(n_307),
.B(n_283),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_275),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_282),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_205),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_8),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_311),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_287),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_289),
.Y(n_313)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_313),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_316),
.Y(n_324)
);

NOR2xp67_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_280),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_317),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_303),
.A2(n_281),
.B(n_280),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_316),
.A2(n_320),
.B(n_321),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_291),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_299),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_SL g321 ( 
.A(n_298),
.B(n_16),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_325),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_317),
.B(n_304),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_328),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_297),
.Y(n_327)
);

AOI21x1_ASAP7_75t_SL g335 ( 
.A1(n_327),
.A2(n_319),
.B(n_16),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_311),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_322),
.A2(n_16),
.B1(n_6),
.B2(n_7),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_330),
.B(n_323),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_335),
.Y(n_340)
);

AO21x1_ASAP7_75t_L g337 ( 
.A1(n_329),
.A2(n_5),
.B(n_6),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_337),
.A2(n_332),
.B(n_7),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_331),
.A2(n_5),
.B1(n_7),
.B2(n_329),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_338),
.Y(n_339)
);

AOI21xp33_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_337),
.B(n_7),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_339),
.C(n_335),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_343),
.A2(n_334),
.B(n_336),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_327),
.C(n_340),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_5),
.Y(n_346)
);


endmodule