module fake_netlist_6_69_n_1668 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1668);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1668;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx8_ASAP7_75t_SL g159 ( 
.A(n_93),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_22),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_49),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_49),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_109),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_32),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_53),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_146),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_85),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g171 ( 
.A(n_37),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_23),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_132),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_92),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_82),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_39),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_105),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_69),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_71),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_8),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_1),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_37),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_137),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_46),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_61),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_5),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_39),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_150),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_51),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_11),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_84),
.Y(n_193)
);

INVxp33_ASAP7_75t_R g194 ( 
.A(n_10),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_149),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_47),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_87),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_112),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_54),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_151),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_7),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_73),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_89),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_142),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_147),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_94),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_79),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_77),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_13),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_2),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_7),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_126),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_128),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_52),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_50),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_111),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_24),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_95),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_43),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_8),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_108),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_80),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_40),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_46),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_17),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_113),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_138),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_97),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_72),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_125),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_134),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_131),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_102),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_5),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_34),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_91),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_6),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_62),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_4),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_106),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_28),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_21),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_16),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_107),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_0),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_153),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_13),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_155),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_103),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_33),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_15),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_98),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_58),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_123),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_139),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_144),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_52),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_17),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_157),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_18),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_41),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_35),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_130),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_121),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_110),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_63),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_65),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_12),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_36),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_25),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_56),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_35),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_16),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_0),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_152),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_143),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_68),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_75),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_47),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_20),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_145),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_64),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_14),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_41),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_31),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_148),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_70),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_100),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_28),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_43),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_83),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_27),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_90),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_25),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_60),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_78),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_81),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_40),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_1),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_11),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_23),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_9),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_24),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_38),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_30),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_66),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_59),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_50),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_156),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_76),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_33),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_34),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_30),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_26),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_14),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_104),
.Y(n_316)
);

BUFx2_ASAP7_75t_SL g317 ( 
.A(n_198),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_172),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_159),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_L g320 ( 
.A(n_196),
.B(n_2),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_200),
.Y(n_321)
);

OAI21x1_ASAP7_75t_L g322 ( 
.A1(n_168),
.A2(n_3),
.B(n_4),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_204),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_275),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_R g325 ( 
.A(n_228),
.B(n_173),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_172),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_172),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_205),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_196),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_188),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_208),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_172),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_240),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_196),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_201),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_201),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_201),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_215),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_209),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_188),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_209),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_282),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_220),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_220),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_273),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_192),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_206),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_192),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_207),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_161),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_273),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_280),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_280),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_160),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_181),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_185),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_212),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_211),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_217),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_213),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_224),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_216),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_287),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_222),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_295),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_227),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_235),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_230),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_198),
.B(n_3),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_231),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_221),
.B(n_6),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_233),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_239),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_161),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_242),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_243),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_247),
.Y(n_377)
);

INVxp33_ASAP7_75t_SL g378 ( 
.A(n_166),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_244),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_249),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_293),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_251),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_258),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_221),
.B(n_9),
.Y(n_384)
);

INVxp33_ASAP7_75t_SL g385 ( 
.A(n_166),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_188),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_296),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_262),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_269),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_270),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_234),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_325),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_366),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_318),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_318),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_381),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_326),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_387),
.Y(n_398)
);

AND2x6_ASAP7_75t_L g399 ( 
.A(n_329),
.B(n_162),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_331),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_326),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_338),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_321),
.Y(n_403)
);

NAND3xp33_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_171),
.C(n_225),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_327),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_337),
.B(n_300),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_327),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_332),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_323),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_328),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_347),
.B(n_165),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_332),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_330),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_349),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_333),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_357),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_329),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_360),
.B(n_165),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_342),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_363),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_350),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_365),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_362),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_334),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_324),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_364),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_335),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_352),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_368),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_352),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_370),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_372),
.B(n_229),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_378),
.B(n_237),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_322),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_322),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_379),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_380),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_335),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_319),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g440 ( 
.A(n_371),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_336),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_336),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_317),
.Y(n_443)
);

AND2x6_ASAP7_75t_L g444 ( 
.A(n_384),
.B(n_162),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_317),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_339),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_340),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_339),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_341),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_374),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g452 ( 
.A1(n_341),
.A2(n_344),
.B(n_343),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_356),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_385),
.B(n_310),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_386),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_343),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_344),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_345),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_345),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_391),
.B(n_310),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_445),
.B(n_402),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_395),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_407),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_453),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_394),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_395),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_395),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_397),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_413),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_407),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_440),
.B(n_346),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_440),
.B(n_168),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_451),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_454),
.B(n_348),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_408),
.Y(n_475)
);

BUFx10_ASAP7_75t_L g476 ( 
.A(n_392),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_401),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_456),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_452),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_434),
.B(n_199),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_405),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_411),
.B(n_358),
.Y(n_482)
);

BUFx10_ASAP7_75t_L g483 ( 
.A(n_392),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_395),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_456),
.Y(n_485)
);

NAND2xp33_ASAP7_75t_L g486 ( 
.A(n_444),
.B(n_162),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_443),
.B(n_199),
.Y(n_487)
);

AND2x2_ASAP7_75t_SL g488 ( 
.A(n_460),
.B(n_238),
.Y(n_488)
);

AND2x6_ASAP7_75t_L g489 ( 
.A(n_434),
.B(n_238),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_444),
.A2(n_320),
.B1(n_300),
.B2(n_259),
.Y(n_490)
);

AND3x2_ASAP7_75t_L g491 ( 
.A(n_413),
.B(n_259),
.C(n_254),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_424),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_427),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_444),
.B(n_229),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_438),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_406),
.B(n_232),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_418),
.B(n_359),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_432),
.B(n_421),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_444),
.B(n_232),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_443),
.B(n_354),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_425),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_441),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_444),
.B(n_167),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_412),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_446),
.B(n_254),
.Y(n_505)
);

INVx4_ASAP7_75t_SL g506 ( 
.A(n_399),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_446),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_434),
.B(n_288),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_444),
.A2(n_316),
.B1(n_288),
.B2(n_290),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_412),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_L g511 ( 
.A(n_444),
.B(n_162),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_406),
.Y(n_512)
);

NAND3xp33_ASAP7_75t_L g513 ( 
.A(n_404),
.B(n_214),
.C(n_210),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_434),
.A2(n_316),
.B1(n_289),
.B2(n_294),
.Y(n_514)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_412),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_456),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_434),
.A2(n_304),
.B1(n_308),
.B2(n_312),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_426),
.B(n_354),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_456),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_417),
.B(n_203),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_435),
.A2(n_279),
.B1(n_314),
.B2(n_388),
.Y(n_521)
);

AND2x6_ASAP7_75t_L g522 ( 
.A(n_435),
.B(n_162),
.Y(n_522)
);

OR2x6_ASAP7_75t_L g523 ( 
.A(n_436),
.B(n_194),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_435),
.B(n_187),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_442),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_452),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_452),
.Y(n_527)
);

BUFx4f_ASAP7_75t_L g528 ( 
.A(n_452),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_456),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_403),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_458),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_458),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_417),
.B(n_264),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_458),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_435),
.B(n_187),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_435),
.A2(n_375),
.B1(n_389),
.B2(n_388),
.Y(n_536)
);

BUFx8_ASAP7_75t_SL g537 ( 
.A(n_448),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_403),
.B(n_355),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_433),
.Y(n_539)
);

INVxp33_ASAP7_75t_L g540 ( 
.A(n_433),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_430),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_409),
.B(n_261),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_430),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_458),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_458),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_428),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_428),
.Y(n_547)
);

OR2x6_ASAP7_75t_L g548 ( 
.A(n_447),
.B(n_355),
.Y(n_548)
);

NOR2x1p5_ASAP7_75t_L g549 ( 
.A(n_409),
.B(n_410),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_410),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_414),
.B(n_187),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_399),
.A2(n_390),
.B1(n_389),
.B2(n_383),
.Y(n_552)
);

INVx5_ASAP7_75t_L g553 ( 
.A(n_399),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_428),
.B(n_170),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_447),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_449),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_449),
.B(n_180),
.Y(n_557)
);

BUFx8_ASAP7_75t_SL g558 ( 
.A(n_400),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_414),
.B(n_390),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_L g560 ( 
.A(n_416),
.B(n_219),
.C(n_223),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_416),
.B(n_361),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_423),
.B(n_361),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_450),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_450),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_423),
.B(n_187),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_457),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_457),
.B(n_383),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_459),
.Y(n_568)
);

INVx4_ASAP7_75t_SL g569 ( 
.A(n_399),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_399),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_459),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_399),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_399),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_431),
.B(n_186),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_431),
.A2(n_373),
.B1(n_377),
.B2(n_376),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_393),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_429),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_437),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_455),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_439),
.A2(n_373),
.B1(n_377),
.B2(n_376),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_SL g581 ( 
.A1(n_393),
.A2(n_234),
.B1(n_245),
.B2(n_226),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_396),
.B(n_197),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_396),
.B(n_202),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_419),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_398),
.B(n_367),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_398),
.A2(n_382),
.B1(n_375),
.B2(n_367),
.Y(n_586)
);

BUFx10_ASAP7_75t_L g587 ( 
.A(n_415),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_420),
.B(n_187),
.Y(n_588)
);

OR2x6_ASAP7_75t_L g589 ( 
.A(n_422),
.B(n_382),
.Y(n_589)
);

OR2x6_ASAP7_75t_L g590 ( 
.A(n_402),
.B(n_218),
.Y(n_590)
);

BUFx4f_ASAP7_75t_L g591 ( 
.A(n_444),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_453),
.Y(n_592)
);

INVxp67_ASAP7_75t_SL g593 ( 
.A(n_395),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_407),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_395),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_392),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_407),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_395),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_440),
.B(n_306),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_399),
.Y(n_600)
);

BUFx10_ASAP7_75t_L g601 ( 
.A(n_392),
.Y(n_601)
);

AND2x6_ASAP7_75t_L g602 ( 
.A(n_434),
.B(n_306),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_406),
.B(n_351),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_440),
.B(n_306),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_488),
.A2(n_163),
.B1(n_284),
.B2(n_306),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_464),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_461),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_592),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_488),
.B(n_236),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_492),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_482),
.B(n_246),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_547),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_518),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_603),
.B(n_351),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_493),
.Y(n_615)
);

BUFx5_ASAP7_75t_L g616 ( 
.A(n_479),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_482),
.B(n_248),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_547),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_564),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_498),
.B(n_164),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_479),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_495),
.Y(n_622)
);

A2O1A1Ixp33_ASAP7_75t_L g623 ( 
.A1(n_528),
.A2(n_252),
.B(n_253),
.C(n_307),
.Y(n_623)
);

A2O1A1Ixp33_ASAP7_75t_L g624 ( 
.A1(n_528),
.A2(n_265),
.B(n_266),
.C(n_297),
.Y(n_624)
);

NOR2x1p5_ASAP7_75t_L g625 ( 
.A(n_530),
.B(n_574),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_497),
.B(n_512),
.Y(n_626)
);

AND3x1_ASAP7_75t_L g627 ( 
.A(n_585),
.B(n_353),
.C(n_286),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_564),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_526),
.A2(n_306),
.B1(n_276),
.B2(n_278),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_497),
.B(n_164),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_498),
.B(n_169),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_536),
.B(n_174),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_514),
.A2(n_175),
.B1(n_174),
.B2(n_177),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_538),
.B(n_175),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_527),
.A2(n_176),
.B1(n_315),
.B2(n_313),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_538),
.B(n_178),
.Y(n_636)
);

AND2x4_ASAP7_75t_SL g637 ( 
.A(n_587),
.B(n_226),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_471),
.B(n_178),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_471),
.B(n_179),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_502),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_525),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_568),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_559),
.B(n_234),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_500),
.B(n_179),
.Y(n_644)
);

INVx5_ASAP7_75t_L g645 ( 
.A(n_522),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_561),
.B(n_562),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_561),
.B(n_184),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_514),
.B(n_184),
.Y(n_648)
);

NAND2x1p5_ASAP7_75t_L g649 ( 
.A(n_591),
.B(n_353),
.Y(n_649)
);

AND2x6_ASAP7_75t_L g650 ( 
.A(n_572),
.B(n_226),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_474),
.B(n_190),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_562),
.B(n_193),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_469),
.B(n_473),
.Y(n_653)
);

OAI221xp5_ASAP7_75t_L g654 ( 
.A1(n_472),
.A2(n_241),
.B1(n_298),
.B2(n_299),
.C(n_301),
.Y(n_654)
);

NOR3xp33_ASAP7_75t_L g655 ( 
.A(n_588),
.B(n_271),
.C(n_195),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_558),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_474),
.B(n_255),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_599),
.B(n_255),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_548),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_585),
.B(n_256),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_580),
.B(n_245),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_509),
.A2(n_315),
.B1(n_313),
.B2(n_311),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_603),
.B(n_256),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_521),
.A2(n_271),
.B1(n_309),
.B2(n_281),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_603),
.B(n_263),
.Y(n_665)
);

AND2x6_ASAP7_75t_L g666 ( 
.A(n_494),
.B(n_245),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_586),
.B(n_263),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_521),
.B(n_267),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_568),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_599),
.B(n_267),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_604),
.B(n_277),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_465),
.B(n_277),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_571),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_571),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_604),
.A2(n_291),
.B1(n_309),
.B2(n_305),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_487),
.B(n_302),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_468),
.B(n_303),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_477),
.B(n_311),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_588),
.A2(n_292),
.B1(n_285),
.B2(n_283),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_L g680 ( 
.A(n_522),
.B(n_292),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_496),
.A2(n_285),
.B1(n_283),
.B2(n_274),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_487),
.B(n_274),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_481),
.B(n_272),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_558),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_505),
.B(n_272),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_463),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_509),
.A2(n_268),
.B1(n_260),
.B2(n_257),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_505),
.B(n_582),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_463),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_496),
.B(n_268),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_496),
.A2(n_260),
.B1(n_257),
.B2(n_250),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_583),
.B(n_250),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_524),
.B(n_191),
.Y(n_693)
);

OAI22xp33_ASAP7_75t_L g694 ( 
.A1(n_542),
.A2(n_191),
.B1(n_189),
.B2(n_183),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_501),
.B(n_189),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_470),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_551),
.B(n_183),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_SL g698 ( 
.A(n_517),
.B(n_182),
.C(n_176),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_524),
.B(n_182),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_551),
.B(n_10),
.Y(n_700)
);

NOR2xp67_ASAP7_75t_SL g701 ( 
.A(n_553),
.B(n_12),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_586),
.B(n_15),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_535),
.B(n_67),
.Y(n_703)
);

OR2x6_ASAP7_75t_L g704 ( 
.A(n_589),
.B(n_18),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_517),
.B(n_74),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_503),
.A2(n_86),
.B1(n_154),
.B2(n_140),
.Y(n_706)
);

BUFx6f_ASAP7_75t_SL g707 ( 
.A(n_476),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_475),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_575),
.B(n_19),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_575),
.B(n_580),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_490),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_SL g712 ( 
.A(n_476),
.B(n_22),
.Y(n_712)
);

A2O1A1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_508),
.A2(n_26),
.B(n_27),
.C(n_29),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_589),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_490),
.B(n_96),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_508),
.B(n_99),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_594),
.B(n_88),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_594),
.B(n_101),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_597),
.Y(n_719)
);

OR2x6_ASAP7_75t_L g720 ( 
.A(n_589),
.B(n_29),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_597),
.B(n_115),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_507),
.B(n_31),
.Y(n_722)
);

AND2x6_ASAP7_75t_L g723 ( 
.A(n_499),
.B(n_116),
.Y(n_723)
);

AO22x1_ASAP7_75t_L g724 ( 
.A1(n_480),
.A2(n_489),
.B1(n_602),
.B2(n_522),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_565),
.B(n_32),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_491),
.Y(n_726)
);

O2A1O1Ixp5_ASAP7_75t_L g727 ( 
.A1(n_591),
.A2(n_36),
.B(n_38),
.C(n_42),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_565),
.B(n_42),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_546),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_520),
.B(n_118),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_567),
.B(n_119),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_L g732 ( 
.A(n_522),
.B(n_117),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_560),
.B(n_44),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_567),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_567),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_539),
.B(n_44),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_480),
.A2(n_122),
.B1(n_135),
.B2(n_133),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_533),
.B(n_57),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_550),
.B(n_45),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_601),
.B(n_45),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_541),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_SL g742 ( 
.A(n_483),
.B(n_48),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_555),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_513),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_543),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_556),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_576),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_563),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_522),
.B(n_55),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_601),
.B(n_48),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_566),
.B(n_127),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_576),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_601),
.B(n_596),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_602),
.B(n_129),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_478),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_480),
.A2(n_51),
.B1(n_158),
.B2(n_489),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_480),
.A2(n_489),
.B1(n_602),
.B2(n_511),
.Y(n_757)
);

AND2x2_ASAP7_75t_SL g758 ( 
.A(n_486),
.B(n_552),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_576),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_602),
.B(n_593),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_602),
.B(n_489),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_480),
.B(n_489),
.Y(n_762)
);

NOR3xp33_ASAP7_75t_L g763 ( 
.A(n_581),
.B(n_557),
.C(n_584),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_478),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_760),
.A2(n_573),
.B(n_570),
.Y(n_765)
);

A2O1A1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_620),
.A2(n_544),
.B(n_531),
.C(n_529),
.Y(n_766)
);

OAI21xp33_ASAP7_75t_SL g767 ( 
.A1(n_710),
.A2(n_552),
.B(n_549),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_724),
.A2(n_573),
.B(n_570),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_645),
.A2(n_515),
.B(n_504),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_621),
.Y(n_770)
);

A2O1A1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_620),
.A2(n_631),
.B(n_688),
.C(n_639),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_707),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_688),
.B(n_631),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_734),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_621),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_643),
.B(n_613),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_626),
.B(n_462),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_747),
.B(n_590),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_646),
.B(n_540),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_752),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_711),
.A2(n_590),
.B1(n_540),
.B2(n_576),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_661),
.B(n_590),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_616),
.B(n_621),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_645),
.A2(n_484),
.B(n_515),
.Y(n_784)
);

AND2x6_ASAP7_75t_SL g785 ( 
.A(n_704),
.B(n_523),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_636),
.B(n_462),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_702),
.A2(n_554),
.B(n_534),
.C(n_545),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_638),
.B(n_596),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_645),
.A2(n_484),
.B(n_504),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_652),
.B(n_579),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_645),
.A2(n_598),
.B(n_595),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_761),
.A2(n_598),
.B(n_595),
.Y(n_792)
);

INVx5_ASAP7_75t_L g793 ( 
.A(n_723),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_762),
.A2(n_598),
.B(n_595),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_716),
.A2(n_598),
.B(n_595),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_629),
.A2(n_510),
.B(n_600),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_711),
.A2(n_577),
.B1(n_584),
.B2(n_523),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_629),
.A2(n_510),
.B(n_600),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_639),
.B(n_483),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_703),
.A2(n_510),
.B(n_600),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_651),
.B(n_466),
.Y(n_801)
);

AOI21xp33_ASAP7_75t_L g802 ( 
.A1(n_692),
.A2(n_577),
.B(n_578),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_616),
.B(n_600),
.Y(n_803)
);

OR2x6_ASAP7_75t_L g804 ( 
.A(n_704),
.B(n_523),
.Y(n_804)
);

INVx5_ASAP7_75t_L g805 ( 
.A(n_723),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_695),
.Y(n_806)
);

O2A1O1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_709),
.A2(n_531),
.B(n_545),
.C(n_485),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_649),
.A2(n_510),
.B(n_553),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_758),
.A2(n_532),
.B(n_544),
.Y(n_809)
);

AOI21x1_ASAP7_75t_L g810 ( 
.A1(n_686),
.A2(n_532),
.B(n_519),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_657),
.B(n_467),
.Y(n_811)
);

OAI321xp33_ASAP7_75t_L g812 ( 
.A1(n_635),
.A2(n_516),
.A3(n_587),
.B1(n_537),
.B2(n_467),
.C(n_569),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_635),
.A2(n_553),
.B1(n_506),
.B2(n_569),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_605),
.A2(n_758),
.B1(n_756),
.B2(n_609),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_623),
.A2(n_553),
.B(n_506),
.Y(n_815)
);

AOI21x1_ASAP7_75t_L g816 ( 
.A1(n_689),
.A2(n_506),
.B(n_569),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_649),
.A2(n_587),
.B(n_537),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_630),
.B(n_692),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_611),
.B(n_617),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_759),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_757),
.A2(n_612),
.B(n_738),
.Y(n_821)
);

NOR3xp33_ASAP7_75t_L g822 ( 
.A(n_694),
.B(n_660),
.C(n_634),
.Y(n_822)
);

AOI22x1_ASAP7_75t_L g823 ( 
.A1(n_755),
.A2(n_764),
.B1(n_618),
.B2(n_622),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_757),
.A2(n_612),
.B(n_730),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_715),
.A2(n_731),
.B(n_735),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_731),
.A2(n_732),
.B(n_708),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_719),
.A2(n_705),
.B(n_729),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_717),
.A2(n_718),
.B(n_721),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_644),
.B(n_658),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_658),
.B(n_670),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_763),
.A2(n_655),
.B1(n_676),
.B2(n_616),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_607),
.B(n_647),
.Y(n_832)
);

NOR2xp67_ASAP7_75t_L g833 ( 
.A(n_653),
.B(n_753),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_619),
.A2(n_669),
.B(n_642),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_628),
.A2(n_673),
.B(n_674),
.Y(n_835)
);

AO21x1_ASAP7_75t_L g836 ( 
.A1(n_700),
.A2(n_728),
.B(n_671),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_670),
.B(n_671),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_616),
.B(n_676),
.Y(n_838)
);

AO21x1_ASAP7_75t_L g839 ( 
.A1(n_700),
.A2(n_728),
.B(n_697),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_606),
.A2(n_608),
.B(n_640),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_751),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_690),
.B(n_663),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_741),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_610),
.A2(n_641),
.B(n_615),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_616),
.B(n_763),
.Y(n_845)
);

NOR2xp67_ASAP7_75t_L g846 ( 
.A(n_654),
.B(n_675),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_749),
.A2(n_754),
.B(n_665),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_614),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_698),
.A2(n_685),
.B1(n_682),
.B2(n_655),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_614),
.B(n_743),
.Y(n_850)
);

CKINVDCx10_ASAP7_75t_R g851 ( 
.A(n_707),
.Y(n_851)
);

NAND3xp33_ASAP7_75t_L g852 ( 
.A(n_605),
.B(n_627),
.C(n_667),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_746),
.B(n_748),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_751),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_745),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_693),
.B(n_699),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_672),
.A2(n_677),
.B(n_632),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_659),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_756),
.A2(n_624),
.B(n_648),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_727),
.A2(n_698),
.B(n_713),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_678),
.A2(n_683),
.B(n_668),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_725),
.B(n_666),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_666),
.B(n_650),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_666),
.B(n_650),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_666),
.B(n_650),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_727),
.A2(n_680),
.B(n_691),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_681),
.A2(n_733),
.B(n_706),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_736),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_737),
.A2(n_726),
.B(n_739),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_666),
.B(n_650),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_722),
.A2(n_750),
.B(n_740),
.Y(n_871)
);

NOR3xp33_ASAP7_75t_SL g872 ( 
.A(n_694),
.B(n_664),
.C(n_633),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_662),
.A2(n_687),
.B(n_742),
.C(n_712),
.Y(n_873)
);

INVx3_ASAP7_75t_SL g874 ( 
.A(n_704),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_714),
.A2(n_637),
.B(n_650),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_679),
.B(n_687),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_662),
.B(n_625),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_723),
.A2(n_720),
.B(n_701),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_656),
.A2(n_684),
.B(n_723),
.C(n_720),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_720),
.A2(n_591),
.B(n_528),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_688),
.B(n_620),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_646),
.B(n_620),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_760),
.A2(n_591),
.B(n_528),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_696),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_710),
.A2(n_488),
.B1(n_698),
.B2(n_700),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_688),
.B(n_620),
.Y(n_886)
);

AOI21x1_ASAP7_75t_L g887 ( 
.A1(n_724),
.A2(n_535),
.B(n_524),
.Y(n_887)
);

O2A1O1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_710),
.A2(n_646),
.B(n_702),
.C(n_709),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_758),
.A2(n_528),
.B(n_527),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_688),
.B(n_620),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_760),
.A2(n_591),
.B(n_528),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_758),
.A2(n_528),
.B(n_527),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_688),
.A2(n_631),
.B1(n_620),
.B2(n_744),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_688),
.B(n_620),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_688),
.B(n_620),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_760),
.A2(n_591),
.B(n_528),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_760),
.A2(n_591),
.B(n_528),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_643),
.B(n_559),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_621),
.Y(n_899)
);

NAND2xp33_ASAP7_75t_L g900 ( 
.A(n_616),
.B(n_621),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_688),
.B(n_620),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_688),
.B(n_620),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_646),
.B(n_620),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_710),
.A2(n_711),
.B1(n_629),
.B2(n_635),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_688),
.A2(n_631),
.B1(n_620),
.B2(n_744),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_688),
.A2(n_631),
.B1(n_620),
.B2(n_744),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_747),
.B(n_752),
.Y(n_907)
);

AOI21x1_ASAP7_75t_L g908 ( 
.A1(n_724),
.A2(n_535),
.B(n_524),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_760),
.A2(n_591),
.B(n_528),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_760),
.A2(n_591),
.B(n_528),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_621),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_688),
.A2(n_631),
.B1(n_620),
.B2(n_744),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_760),
.A2(n_591),
.B(n_528),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_760),
.A2(n_591),
.B(n_528),
.Y(n_914)
);

AOI21x1_ASAP7_75t_L g915 ( 
.A1(n_724),
.A2(n_535),
.B(n_524),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_758),
.A2(n_528),
.B(n_527),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_734),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_710),
.A2(n_646),
.B(n_702),
.C(n_709),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_643),
.B(n_559),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_688),
.B(n_620),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_760),
.A2(n_591),
.B(n_528),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_688),
.B(n_620),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_688),
.B(n_620),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_621),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_760),
.A2(n_591),
.B(n_528),
.Y(n_925)
);

AOI21x1_ASAP7_75t_L g926 ( 
.A1(n_724),
.A2(n_535),
.B(n_524),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_621),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_760),
.A2(n_591),
.B(n_528),
.Y(n_928)
);

OAI21xp33_ASAP7_75t_L g929 ( 
.A1(n_620),
.A2(n_631),
.B(n_638),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_760),
.A2(n_591),
.B(n_528),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_760),
.A2(n_591),
.B(n_528),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_688),
.B(n_620),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_688),
.B(n_620),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_760),
.A2(n_591),
.B(n_528),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_760),
.A2(n_591),
.B(n_528),
.Y(n_935)
);

AOI21xp33_ASAP7_75t_L g936 ( 
.A1(n_929),
.A2(n_903),
.B(n_882),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_900),
.A2(n_825),
.B(n_838),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_774),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_773),
.B(n_881),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_886),
.B(n_890),
.Y(n_940)
);

OAI21x1_ASAP7_75t_L g941 ( 
.A1(n_794),
.A2(n_908),
.B(n_887),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_893),
.B(n_905),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_894),
.B(n_895),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_906),
.B(n_912),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_899),
.Y(n_945)
);

NAND2x1_ASAP7_75t_L g946 ( 
.A(n_899),
.B(n_911),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_771),
.A2(n_892),
.B(n_889),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_901),
.B(n_902),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_920),
.B(n_922),
.Y(n_949)
);

AO31x2_ASAP7_75t_L g950 ( 
.A1(n_836),
.A2(n_839),
.A3(n_766),
.B(n_814),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_915),
.A2(n_926),
.B(n_792),
.Y(n_951)
);

AO21x2_ASAP7_75t_L g952 ( 
.A1(n_831),
.A2(n_860),
.B(n_845),
.Y(n_952)
);

OAI21x1_ASAP7_75t_L g953 ( 
.A1(n_823),
.A2(n_891),
.B(n_883),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_896),
.A2(n_909),
.B(n_897),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_780),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_910),
.A2(n_935),
.B(n_914),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_923),
.B(n_932),
.Y(n_957)
);

NAND2x1p5_ASAP7_75t_L g958 ( 
.A(n_899),
.B(n_911),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_913),
.A2(n_925),
.B(n_921),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_889),
.A2(n_916),
.B(n_892),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_928),
.A2(n_931),
.B(n_930),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_788),
.B(n_790),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_933),
.B(n_818),
.Y(n_963)
);

AO21x1_ASAP7_75t_L g964 ( 
.A1(n_830),
.A2(n_837),
.B(n_814),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_934),
.A2(n_826),
.B(n_847),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_898),
.Y(n_966)
);

OAI21x1_ASAP7_75t_L g967 ( 
.A1(n_809),
.A2(n_824),
.B(n_821),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_765),
.A2(n_828),
.B(n_783),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_819),
.B(n_829),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_904),
.A2(n_885),
.B1(n_849),
.B2(n_876),
.Y(n_970)
);

NOR3xp33_ASAP7_75t_L g971 ( 
.A(n_799),
.B(n_873),
.C(n_781),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_809),
.A2(n_807),
.B(n_800),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_842),
.B(n_919),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_856),
.B(n_861),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_859),
.A2(n_786),
.B(n_801),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_917),
.Y(n_976)
);

AOI21xp33_ASAP7_75t_L g977 ( 
.A1(n_888),
.A2(n_918),
.B(n_852),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_853),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_841),
.B(n_854),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_806),
.B(n_779),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_841),
.B(n_854),
.Y(n_981)
);

AO21x2_ASAP7_75t_L g982 ( 
.A1(n_866),
.A2(n_865),
.B(n_864),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_911),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_916),
.A2(n_767),
.B(n_857),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_822),
.A2(n_846),
.B(n_867),
.C(n_872),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_811),
.A2(n_803),
.B(n_768),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_816),
.A2(n_787),
.B(n_834),
.Y(n_987)
);

O2A1O1Ixp5_ASAP7_75t_L g988 ( 
.A1(n_862),
.A2(n_863),
.B(n_870),
.C(n_869),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_924),
.Y(n_989)
);

OAI21x1_ASAP7_75t_L g990 ( 
.A1(n_835),
.A2(n_791),
.B(n_808),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_769),
.A2(n_789),
.B(n_784),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_777),
.A2(n_796),
.B(n_798),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_880),
.A2(n_877),
.B(n_844),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_813),
.A2(n_850),
.B(n_815),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_813),
.A2(n_815),
.B(n_840),
.Y(n_995)
);

AO31x2_ASAP7_75t_L g996 ( 
.A1(n_878),
.A2(n_879),
.A3(n_871),
.B(n_797),
.Y(n_996)
);

AOI221x1_ASAP7_75t_L g997 ( 
.A1(n_802),
.A2(n_797),
.B1(n_875),
.B2(n_782),
.C(n_832),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_855),
.B(n_843),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_770),
.A2(n_927),
.B(n_775),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_855),
.B(n_848),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_884),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_778),
.A2(n_907),
.B1(n_833),
.B2(n_858),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_812),
.A2(n_793),
.B(n_805),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_868),
.B(n_778),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_924),
.A2(n_793),
.B(n_805),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_812),
.A2(n_793),
.B(n_805),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_924),
.B(n_820),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_820),
.B(n_793),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_874),
.B(n_817),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_SL g1010 ( 
.A1(n_805),
.A2(n_804),
.B(n_772),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_804),
.B(n_785),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_851),
.A2(n_591),
.B(n_900),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_773),
.B(n_881),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_900),
.A2(n_591),
.B(n_528),
.Y(n_1014)
);

AO31x2_ASAP7_75t_L g1015 ( 
.A1(n_836),
.A2(n_839),
.A3(n_771),
.B(n_766),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_929),
.A2(n_771),
.B(n_903),
.C(n_882),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_929),
.A2(n_771),
.B(n_903),
.C(n_882),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_929),
.A2(n_771),
.B(n_903),
.C(n_882),
.Y(n_1018)
);

AOI21xp33_ASAP7_75t_L g1019 ( 
.A1(n_929),
.A2(n_903),
.B(n_882),
.Y(n_1019)
);

AOI21xp33_ASAP7_75t_L g1020 ( 
.A1(n_929),
.A2(n_903),
.B(n_882),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_907),
.B(n_759),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_907),
.B(n_759),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_898),
.B(n_919),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_771),
.A2(n_892),
.B(n_889),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_899),
.Y(n_1025)
);

AOI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_929),
.A2(n_903),
.B(n_882),
.Y(n_1026)
);

INVx8_ASAP7_75t_L g1027 ( 
.A(n_907),
.Y(n_1027)
);

AND2x6_ASAP7_75t_L g1028 ( 
.A(n_841),
.B(n_621),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_907),
.B(n_759),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_773),
.B(n_881),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_773),
.B(n_881),
.Y(n_1031)
);

BUFx12f_ASAP7_75t_L g1032 ( 
.A(n_772),
.Y(n_1032)
);

INVxp67_ASAP7_75t_L g1033 ( 
.A(n_776),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_771),
.A2(n_892),
.B(n_889),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_773),
.B(n_881),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_898),
.B(n_919),
.Y(n_1036)
);

INVx6_ASAP7_75t_SL g1037 ( 
.A(n_804),
.Y(n_1037)
);

NOR3xp33_ASAP7_75t_L g1038 ( 
.A(n_929),
.B(n_419),
.C(n_799),
.Y(n_1038)
);

INVx1_ASAP7_75t_SL g1039 ( 
.A(n_898),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_773),
.B(n_881),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_771),
.A2(n_892),
.B(n_889),
.Y(n_1041)
);

OA22x2_ASAP7_75t_L g1042 ( 
.A1(n_893),
.A2(n_710),
.B1(n_906),
.B2(n_905),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_773),
.B(n_881),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_771),
.A2(n_892),
.B(n_889),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_899),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_898),
.B(n_919),
.Y(n_1046)
);

OAI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_893),
.A2(n_906),
.B1(n_912),
.B2(n_905),
.Y(n_1047)
);

NAND2x1p5_ASAP7_75t_L g1048 ( 
.A(n_899),
.B(n_911),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_899),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_773),
.B(n_881),
.Y(n_1050)
);

AOI21xp33_ASAP7_75t_L g1051 ( 
.A1(n_929),
.A2(n_903),
.B(n_882),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_773),
.B(n_881),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_898),
.B(n_473),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_773),
.B(n_881),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_900),
.A2(n_591),
.B(n_528),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_810),
.A2(n_795),
.B(n_827),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_1027),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_1016),
.A2(n_1017),
.B(n_1018),
.C(n_985),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_955),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_969),
.A2(n_963),
.B1(n_940),
.B2(n_1040),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_1004),
.Y(n_1061)
);

INVx5_ASAP7_75t_L g1062 ( 
.A(n_1028),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_938),
.Y(n_1063)
);

NAND3xp33_ASAP7_75t_L g1064 ( 
.A(n_971),
.B(n_944),
.C(n_942),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_940),
.B(n_1040),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_966),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1023),
.B(n_1036),
.Y(n_1067)
);

OR2x2_ASAP7_75t_SL g1068 ( 
.A(n_1011),
.B(n_980),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_1053),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_1046),
.B(n_966),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_962),
.B(n_936),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_974),
.A2(n_965),
.B(n_937),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_939),
.B(n_943),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_936),
.B(n_1019),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_948),
.B(n_949),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_1039),
.B(n_973),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_957),
.B(n_1013),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1030),
.B(n_1031),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1039),
.B(n_978),
.Y(n_1079)
);

OR2x6_ASAP7_75t_L g1080 ( 
.A(n_1010),
.B(n_1027),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_976),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_1028),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_1021),
.B(n_1022),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_1033),
.Y(n_1084)
);

INVx4_ASAP7_75t_SL g1085 ( 
.A(n_1028),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1035),
.B(n_1043),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1050),
.B(n_1052),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_1021),
.B(n_1022),
.Y(n_1088)
);

NOR2x1_ASAP7_75t_L g1089 ( 
.A(n_1007),
.B(n_1008),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_1054),
.A2(n_1047),
.B1(n_1042),
.B2(n_970),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_1032),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1038),
.B(n_1029),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_1027),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_1037),
.Y(n_1094)
);

NOR2xp67_ASAP7_75t_L g1095 ( 
.A(n_1002),
.B(n_1001),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_945),
.Y(n_1096)
);

BUFx8_ASAP7_75t_SL g1097 ( 
.A(n_1009),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1019),
.B(n_1020),
.Y(n_1098)
);

NAND2xp33_ASAP7_75t_L g1099 ( 
.A(n_970),
.B(n_979),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_1037),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_1020),
.B(n_1026),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1042),
.A2(n_1026),
.B1(n_1051),
.B2(n_1044),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_996),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_998),
.Y(n_1104)
);

BUFx12f_ASAP7_75t_L g1105 ( 
.A(n_945),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_1000),
.B(n_977),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_984),
.A2(n_947),
.B(n_1034),
.C(n_1024),
.Y(n_1107)
);

BUFx12f_ASAP7_75t_L g1108 ( 
.A(n_945),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_952),
.B(n_947),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_996),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_981),
.B(n_1049),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_983),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1049),
.B(n_1015),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1024),
.B(n_1041),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1015),
.B(n_950),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_983),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_975),
.A2(n_968),
.B(n_984),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1034),
.B(n_1041),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1044),
.B(n_964),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_983),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_958),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_997),
.B(n_993),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_995),
.A2(n_959),
.B(n_961),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_960),
.B(n_950),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_989),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_989),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_958),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_1012),
.B(n_1025),
.Y(n_1128)
);

NAND2x1p5_ASAP7_75t_L g1129 ( 
.A(n_989),
.B(n_1025),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_960),
.A2(n_994),
.B1(n_1003),
.B2(n_1006),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_1025),
.Y(n_1131)
);

INVx4_ASAP7_75t_SL g1132 ( 
.A(n_1045),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_954),
.A2(n_1014),
.B(n_1055),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1045),
.Y(n_1134)
);

NAND2x1p5_ASAP7_75t_L g1135 ( 
.A(n_1045),
.B(n_946),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_993),
.Y(n_1136)
);

BUFx12f_ASAP7_75t_L g1137 ( 
.A(n_1048),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_1048),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_982),
.B(n_967),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1003),
.A2(n_1006),
.B1(n_1005),
.B2(n_992),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_999),
.B(n_988),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_986),
.A2(n_953),
.B(n_956),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_972),
.B(n_990),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_951),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_941),
.B(n_991),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_987),
.B(n_1056),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_940),
.B(n_1040),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_962),
.B(n_790),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_1021),
.B(n_1022),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_955),
.Y(n_1150)
);

INVx8_ASAP7_75t_L g1151 ( 
.A(n_1028),
.Y(n_1151)
);

OR2x6_ASAP7_75t_L g1152 ( 
.A(n_1010),
.B(n_1027),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_955),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_1053),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_1028),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_974),
.A2(n_965),
.B(n_937),
.Y(n_1156)
);

NAND3xp33_ASAP7_75t_L g1157 ( 
.A(n_971),
.B(n_929),
.C(n_771),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_966),
.Y(n_1158)
);

AND2x6_ASAP7_75t_L g1159 ( 
.A(n_974),
.B(n_831),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_974),
.A2(n_965),
.B(n_937),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1016),
.A2(n_904),
.B1(n_814),
.B2(n_771),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_1028),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_1027),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_974),
.A2(n_965),
.B(n_937),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_1027),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_940),
.B(n_1040),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1016),
.A2(n_904),
.B1(n_814),
.B2(n_771),
.Y(n_1167)
);

BUFx12f_ASAP7_75t_L g1168 ( 
.A(n_1032),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1023),
.B(n_1036),
.Y(n_1169)
);

BUFx2_ASAP7_75t_SL g1170 ( 
.A(n_955),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_966),
.B(n_576),
.Y(n_1171)
);

OR2x6_ASAP7_75t_SL g1172 ( 
.A(n_1011),
.B(n_393),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_940),
.B(n_1040),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_940),
.B(n_1040),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_955),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_955),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_974),
.A2(n_965),
.B(n_937),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_973),
.B(n_1053),
.Y(n_1178)
);

BUFx5_ASAP7_75t_L g1179 ( 
.A(n_1028),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1062),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1074),
.B(n_1101),
.Y(n_1181)
);

OAI22xp33_ASAP7_75t_SL g1182 ( 
.A1(n_1148),
.A2(n_1060),
.B1(n_1075),
.B2(n_1086),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_1069),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1065),
.B(n_1147),
.Y(n_1184)
);

BUFx12f_ASAP7_75t_L g1185 ( 
.A(n_1091),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_SL g1186 ( 
.A1(n_1136),
.A2(n_1064),
.B1(n_1090),
.B2(n_1157),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1113),
.Y(n_1187)
);

OAI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1073),
.A2(n_1075),
.B1(n_1077),
.B2(n_1078),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1081),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_SL g1190 ( 
.A1(n_1090),
.A2(n_1161),
.B1(n_1167),
.B2(n_1071),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1104),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1063),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1065),
.B(n_1147),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_SL g1194 ( 
.A(n_1097),
.B(n_1168),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1110),
.Y(n_1195)
);

OAI22xp33_ASAP7_75t_SL g1196 ( 
.A1(n_1060),
.A2(n_1078),
.B1(n_1077),
.B2(n_1073),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1106),
.A2(n_1058),
.B(n_1102),
.Y(n_1197)
);

NAND2x1p5_ASAP7_75t_L g1198 ( 
.A(n_1062),
.B(n_1128),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1092),
.A2(n_1169),
.B1(n_1067),
.B2(n_1095),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1066),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1161),
.A2(n_1167),
.B1(n_1102),
.B2(n_1159),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_1158),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1151),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1086),
.B(n_1087),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1080),
.B(n_1152),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_1154),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1079),
.Y(n_1207)
);

BUFx5_ASAP7_75t_L g1208 ( 
.A(n_1146),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1151),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1159),
.A2(n_1098),
.B1(n_1122),
.B2(n_1070),
.Y(n_1210)
);

INVx4_ASAP7_75t_L g1211 ( 
.A(n_1085),
.Y(n_1211)
);

BUFx2_ASAP7_75t_R g1212 ( 
.A(n_1172),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1076),
.Y(n_1213)
);

BUFx12f_ASAP7_75t_L g1214 ( 
.A(n_1094),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1111),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1121),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1059),
.Y(n_1217)
);

OA21x2_ASAP7_75t_L g1218 ( 
.A1(n_1123),
.A2(n_1160),
.B(n_1164),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1141),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1127),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1089),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1166),
.B(n_1173),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1084),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1166),
.B(n_1173),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1174),
.Y(n_1225)
);

OAI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1087),
.A2(n_1174),
.B1(n_1178),
.B2(n_1098),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1171),
.A2(n_1159),
.B1(n_1099),
.B2(n_1061),
.Y(n_1227)
);

OA21x2_ASAP7_75t_L g1228 ( 
.A1(n_1123),
.A2(n_1164),
.B(n_1177),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1120),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_SL g1230 ( 
.A1(n_1159),
.A2(n_1130),
.B1(n_1114),
.B2(n_1118),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1083),
.B(n_1088),
.Y(n_1231)
);

BUFx8_ASAP7_75t_SL g1232 ( 
.A(n_1105),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1125),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1080),
.B(n_1152),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1115),
.B(n_1119),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1131),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1150),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1108),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1103),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1133),
.A2(n_1142),
.B(n_1160),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1144),
.Y(n_1241)
);

INVxp67_ASAP7_75t_L g1242 ( 
.A(n_1170),
.Y(n_1242)
);

BUFx4f_ASAP7_75t_SL g1243 ( 
.A(n_1175),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1116),
.Y(n_1244)
);

BUFx8_ASAP7_75t_L g1245 ( 
.A(n_1100),
.Y(n_1245)
);

NAND2x1p5_ASAP7_75t_L g1246 ( 
.A(n_1128),
.B(n_1139),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_SL g1247 ( 
.A1(n_1140),
.A2(n_1119),
.B1(n_1152),
.B2(n_1080),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1085),
.Y(n_1248)
);

INVx3_ASAP7_75t_SL g1249 ( 
.A(n_1083),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1109),
.A2(n_1149),
.B1(n_1088),
.B2(n_1140),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1068),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1129),
.Y(n_1252)
);

BUFx4f_ASAP7_75t_SL g1253 ( 
.A(n_1176),
.Y(n_1253)
);

AND2x4_ASAP7_75t_SL g1254 ( 
.A(n_1163),
.B(n_1057),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1109),
.A2(n_1149),
.B1(n_1124),
.B2(n_1143),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1153),
.A2(n_1163),
.B1(n_1093),
.B2(n_1165),
.Y(n_1256)
);

NAND2x1p5_ASAP7_75t_L g1257 ( 
.A(n_1143),
.B(n_1145),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1138),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1135),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1132),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1124),
.A2(n_1057),
.B1(n_1165),
.B2(n_1093),
.Y(n_1261)
);

OA21x2_ASAP7_75t_L g1262 ( 
.A1(n_1072),
.A2(n_1156),
.B(n_1177),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1107),
.B(n_1162),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1135),
.Y(n_1264)
);

BUFx4f_ASAP7_75t_SL g1265 ( 
.A(n_1137),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_SL g1266 ( 
.A1(n_1179),
.A2(n_1057),
.B1(n_1165),
.B2(n_1093),
.Y(n_1266)
);

INVx8_ASAP7_75t_L g1267 ( 
.A(n_1126),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1117),
.A2(n_1145),
.B1(n_1096),
.B2(n_1162),
.Y(n_1268)
);

BUFx2_ASAP7_75t_R g1269 ( 
.A(n_1082),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1126),
.Y(n_1270)
);

INVx5_ASAP7_75t_L g1271 ( 
.A(n_1155),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1126),
.Y(n_1272)
);

AO21x2_ASAP7_75t_L g1273 ( 
.A1(n_1132),
.A2(n_1134),
.B(n_1112),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1134),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1132),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1064),
.A2(n_929),
.B1(n_971),
.B2(n_822),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1074),
.B(n_1042),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1073),
.B(n_1075),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1186),
.A2(n_1190),
.B1(n_1276),
.B2(n_1197),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1239),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1195),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1205),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1240),
.A2(n_1262),
.B(n_1228),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1235),
.B(n_1219),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1235),
.B(n_1219),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1208),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1208),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1230),
.B(n_1201),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1257),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1241),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1187),
.B(n_1277),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1262),
.A2(n_1228),
.B(n_1218),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1217),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1246),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1187),
.B(n_1277),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1181),
.B(n_1263),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1205),
.B(n_1234),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1208),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1205),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1181),
.B(n_1263),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1246),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1208),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1246),
.Y(n_1303)
);

AO21x2_ASAP7_75t_L g1304 ( 
.A1(n_1226),
.A2(n_1188),
.B(n_1227),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1182),
.A2(n_1251),
.B1(n_1196),
.B2(n_1224),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1234),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1210),
.B(n_1184),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1200),
.Y(n_1308)
);

OA21x2_ASAP7_75t_L g1309 ( 
.A1(n_1255),
.A2(n_1250),
.B(n_1268),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1208),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1184),
.B(n_1193),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1193),
.B(n_1222),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1222),
.B(n_1224),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1200),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1202),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1225),
.B(n_1204),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1202),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1234),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1251),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1198),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1247),
.B(n_1191),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1189),
.Y(n_1322)
);

AOI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1221),
.A2(n_1216),
.B(n_1220),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1223),
.Y(n_1324)
);

AO21x2_ASAP7_75t_L g1325 ( 
.A1(n_1199),
.A2(n_1278),
.B(n_1215),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1185),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1213),
.B(n_1207),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1192),
.Y(n_1328)
);

CKINVDCx11_ASAP7_75t_R g1329 ( 
.A(n_1185),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1261),
.B(n_1244),
.Y(n_1330)
);

AO21x1_ASAP7_75t_SL g1331 ( 
.A1(n_1259),
.A2(n_1264),
.B(n_1252),
.Y(n_1331)
);

AO21x2_ASAP7_75t_L g1332 ( 
.A1(n_1229),
.A2(n_1233),
.B(n_1236),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1206),
.B(n_1183),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1302),
.B(n_1274),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1299),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1299),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1279),
.A2(n_1249),
.B1(n_1194),
.B2(n_1231),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1296),
.B(n_1266),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1281),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1279),
.A2(n_1242),
.B1(n_1249),
.B2(n_1217),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1281),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1302),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1302),
.B(n_1272),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1296),
.B(n_1258),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1284),
.B(n_1272),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1296),
.B(n_1180),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1284),
.B(n_1272),
.Y(n_1347)
);

AOI221xp5_ASAP7_75t_L g1348 ( 
.A1(n_1288),
.A2(n_1305),
.B1(n_1304),
.B2(n_1324),
.C(n_1307),
.Y(n_1348)
);

NOR2x1p5_ASAP7_75t_L g1349 ( 
.A(n_1282),
.B(n_1248),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1290),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1298),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1285),
.B(n_1298),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1285),
.B(n_1271),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1290),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1288),
.A2(n_1245),
.B1(n_1214),
.B2(n_1237),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1323),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_1308),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1299),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1323),
.Y(n_1359)
);

NOR2x1_ASAP7_75t_L g1360 ( 
.A(n_1332),
.B(n_1304),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1323),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1280),
.B(n_1256),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1286),
.B(n_1209),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1286),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1289),
.B(n_1209),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1299),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1286),
.B(n_1209),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1344),
.B(n_1308),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1344),
.B(n_1315),
.Y(n_1369)
);

NAND2xp33_ASAP7_75t_SL g1370 ( 
.A(n_1349),
.B(n_1293),
.Y(n_1370)
);

AOI211xp5_ASAP7_75t_L g1371 ( 
.A1(n_1348),
.A2(n_1288),
.B(n_1333),
.C(n_1330),
.Y(n_1371)
);

NAND3xp33_ASAP7_75t_L g1372 ( 
.A(n_1348),
.B(n_1305),
.C(n_1330),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1357),
.B(n_1315),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1357),
.B(n_1324),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1339),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1352),
.B(n_1300),
.Y(n_1376)
);

NOR3xp33_ASAP7_75t_L g1377 ( 
.A(n_1340),
.B(n_1314),
.C(n_1320),
.Y(n_1377)
);

OAI21xp33_ASAP7_75t_L g1378 ( 
.A1(n_1340),
.A2(n_1316),
.B(n_1212),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1355),
.B(n_1297),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1356),
.A2(n_1292),
.B(n_1283),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1352),
.B(n_1291),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1352),
.B(n_1317),
.Y(n_1382)
);

OAI21xp5_ASAP7_75t_SL g1383 ( 
.A1(n_1337),
.A2(n_1297),
.B(n_1307),
.Y(n_1383)
);

OA211x2_ASAP7_75t_L g1384 ( 
.A1(n_1355),
.A2(n_1314),
.B(n_1316),
.C(n_1329),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1345),
.B(n_1317),
.Y(n_1385)
);

OAI221xp5_ASAP7_75t_SL g1386 ( 
.A1(n_1337),
.A2(n_1319),
.B1(n_1333),
.B2(n_1307),
.C(n_1321),
.Y(n_1386)
);

OAI221xp5_ASAP7_75t_L g1387 ( 
.A1(n_1360),
.A2(n_1319),
.B1(n_1333),
.B2(n_1303),
.C(n_1301),
.Y(n_1387)
);

AOI221xp5_ASAP7_75t_L g1388 ( 
.A1(n_1338),
.A2(n_1319),
.B1(n_1317),
.B2(n_1321),
.C(n_1295),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1338),
.A2(n_1304),
.B1(n_1297),
.B2(n_1309),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1342),
.B(n_1291),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1342),
.B(n_1291),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1342),
.B(n_1295),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1351),
.B(n_1295),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1339),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1351),
.B(n_1287),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1351),
.B(n_1287),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1346),
.B(n_1293),
.Y(n_1397)
);

OAI21xp33_ASAP7_75t_L g1398 ( 
.A1(n_1360),
.A2(n_1321),
.B(n_1312),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1345),
.B(n_1311),
.Y(n_1399)
);

OAI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1362),
.A2(n_1303),
.B1(n_1301),
.B2(n_1238),
.C(n_1327),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1345),
.B(n_1311),
.Y(n_1401)
);

OAI21xp33_ASAP7_75t_L g1402 ( 
.A1(n_1362),
.A2(n_1312),
.B(n_1327),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1347),
.B(n_1311),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1362),
.A2(n_1269),
.B1(n_1297),
.B2(n_1306),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_SL g1405 ( 
.A(n_1365),
.B(n_1297),
.Y(n_1405)
);

NAND3xp33_ASAP7_75t_L g1406 ( 
.A(n_1359),
.B(n_1328),
.C(n_1322),
.Y(n_1406)
);

OAI221xp5_ASAP7_75t_L g1407 ( 
.A1(n_1346),
.A2(n_1238),
.B1(n_1327),
.B2(n_1294),
.C(n_1237),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1349),
.A2(n_1306),
.B1(n_1318),
.B2(n_1282),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1363),
.B(n_1310),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1363),
.B(n_1310),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1347),
.B(n_1313),
.Y(n_1411)
);

NAND2xp33_ASAP7_75t_SL g1412 ( 
.A(n_1353),
.B(n_1326),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1367),
.B(n_1343),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1347),
.B(n_1313),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1334),
.B(n_1313),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1413),
.B(n_1335),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1375),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1402),
.B(n_1350),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1375),
.Y(n_1419)
);

NAND3xp33_ASAP7_75t_L g1420 ( 
.A(n_1371),
.B(n_1322),
.C(n_1328),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1394),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1394),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1381),
.B(n_1335),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1406),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1402),
.B(n_1350),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1395),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1382),
.B(n_1364),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1406),
.Y(n_1428)
);

NOR2xp67_ASAP7_75t_L g1429 ( 
.A(n_1387),
.B(n_1361),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1398),
.B(n_1354),
.Y(n_1430)
);

NOR2xp67_ASAP7_75t_L g1431 ( 
.A(n_1407),
.B(n_1361),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1390),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1405),
.B(n_1335),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1390),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1391),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1398),
.B(n_1354),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1409),
.B(n_1410),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1380),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1385),
.B(n_1415),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1368),
.B(n_1339),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1380),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1380),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1395),
.Y(n_1443)
);

INVxp67_ASAP7_75t_L g1444 ( 
.A(n_1373),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1376),
.B(n_1364),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1409),
.B(n_1336),
.Y(n_1446)
);

INVx1_ASAP7_75t_SL g1447 ( 
.A(n_1396),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1374),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1396),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1369),
.B(n_1339),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1380),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1393),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1414),
.B(n_1341),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1424),
.B(n_1399),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1424),
.B(n_1401),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1443),
.B(n_1392),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1448),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1417),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1417),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1428),
.B(n_1403),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_1448),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1419),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1419),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1421),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1433),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1444),
.B(n_1411),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1443),
.B(n_1393),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1444),
.B(n_1371),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1443),
.B(n_1358),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1448),
.B(n_1388),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1421),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1421),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1416),
.B(n_1358),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1422),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1453),
.B(n_1397),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1422),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1422),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1432),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1438),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1432),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1433),
.B(n_1358),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1453),
.B(n_1377),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1438),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1428),
.B(n_1427),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1434),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1434),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1433),
.B(n_1366),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1420),
.B(n_1372),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1416),
.B(n_1366),
.Y(n_1489)
);

AOI32xp33_ASAP7_75t_L g1490 ( 
.A1(n_1430),
.A2(n_1378),
.A3(n_1389),
.B1(n_1370),
.B2(n_1412),
.Y(n_1490)
);

OR2x6_ASAP7_75t_L g1491 ( 
.A(n_1420),
.B(n_1379),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1488),
.B(n_1431),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1458),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1468),
.B(n_1431),
.Y(n_1494)
);

OAI31xp33_ASAP7_75t_L g1495 ( 
.A1(n_1470),
.A2(n_1378),
.A3(n_1372),
.B(n_1386),
.Y(n_1495)
);

INVx2_ASAP7_75t_SL g1496 ( 
.A(n_1465),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1465),
.B(n_1437),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1458),
.Y(n_1498)
);

NAND2x1p5_ASAP7_75t_L g1499 ( 
.A(n_1457),
.B(n_1429),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1481),
.B(n_1437),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1481),
.B(n_1429),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1454),
.B(n_1439),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1459),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1459),
.Y(n_1504)
);

NAND4xp25_ASAP7_75t_L g1505 ( 
.A(n_1490),
.B(n_1384),
.C(n_1400),
.D(n_1383),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1479),
.Y(n_1506)
);

INVx1_ASAP7_75t_SL g1507 ( 
.A(n_1484),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1462),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1481),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1481),
.B(n_1437),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1484),
.B(n_1430),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1482),
.B(n_1329),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1461),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1462),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1463),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1454),
.B(n_1455),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1463),
.Y(n_1517)
);

OAI32xp33_ASAP7_75t_L g1518 ( 
.A1(n_1455),
.A2(n_1460),
.A3(n_1436),
.B1(n_1491),
.B2(n_1466),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1478),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1479),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1460),
.B(n_1436),
.Y(n_1521)
);

NOR3xp33_ASAP7_75t_L g1522 ( 
.A(n_1490),
.B(n_1404),
.C(n_1418),
.Y(n_1522)
);

NOR3xp33_ASAP7_75t_L g1523 ( 
.A(n_1475),
.B(n_1425),
.C(n_1418),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1478),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1487),
.B(n_1433),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1487),
.B(n_1433),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1491),
.B(n_1439),
.Y(n_1527)
);

AND2x6_ASAP7_75t_SL g1528 ( 
.A(n_1491),
.B(n_1214),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1491),
.B(n_1440),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1487),
.B(n_1491),
.Y(n_1530)
);

NOR3xp33_ASAP7_75t_L g1531 ( 
.A(n_1483),
.B(n_1425),
.C(n_1408),
.Y(n_1531)
);

INVxp67_ASAP7_75t_L g1532 ( 
.A(n_1480),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1480),
.B(n_1445),
.Y(n_1533)
);

NOR2xp67_ASAP7_75t_L g1534 ( 
.A(n_1487),
.B(n_1426),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1500),
.B(n_1510),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1495),
.A2(n_1450),
.B(n_1440),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1493),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1500),
.B(n_1473),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1522),
.A2(n_1384),
.B1(n_1452),
.B2(n_1447),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1505),
.A2(n_1304),
.B1(n_1325),
.B2(n_1309),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1496),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1510),
.B(n_1473),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1513),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1498),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1523),
.B(n_1467),
.Y(n_1545)
);

INVx3_ASAP7_75t_L g1546 ( 
.A(n_1501),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1525),
.B(n_1467),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1503),
.Y(n_1548)
);

INVx1_ASAP7_75t_SL g1549 ( 
.A(n_1507),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1516),
.B(n_1485),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1504),
.Y(n_1551)
);

INVx1_ASAP7_75t_SL g1552 ( 
.A(n_1492),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1494),
.B(n_1456),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1508),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1514),
.Y(n_1555)
);

NAND3xp33_ASAP7_75t_L g1556 ( 
.A(n_1529),
.B(n_1483),
.C(n_1476),
.Y(n_1556)
);

INVxp67_ASAP7_75t_L g1557 ( 
.A(n_1512),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1525),
.B(n_1456),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1529),
.B(n_1485),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1516),
.Y(n_1560)
);

BUFx12f_ASAP7_75t_L g1561 ( 
.A(n_1528),
.Y(n_1561)
);

INVx4_ASAP7_75t_L g1562 ( 
.A(n_1499),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1515),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1517),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1526),
.B(n_1469),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1519),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1524),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1532),
.Y(n_1568)
);

INVx1_ASAP7_75t_SL g1569 ( 
.A(n_1527),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1526),
.B(n_1469),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_1543),
.B(n_1512),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1549),
.B(n_1545),
.Y(n_1572)
);

O2A1O1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1557),
.A2(n_1518),
.B(n_1499),
.C(n_1501),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1540),
.A2(n_1530),
.B1(n_1509),
.B2(n_1531),
.Y(n_1574)
);

AOI31xp33_ASAP7_75t_L g1575 ( 
.A1(n_1539),
.A2(n_1530),
.A3(n_1511),
.B(n_1509),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1543),
.Y(n_1576)
);

OAI21xp5_ASAP7_75t_SL g1577 ( 
.A1(n_1540),
.A2(n_1501),
.B(n_1511),
.Y(n_1577)
);

AOI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1561),
.A2(n_1534),
.B1(n_1521),
.B2(n_1496),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1552),
.B(n_1502),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1560),
.B(n_1497),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1568),
.B(n_1497),
.Y(n_1581)
);

NAND2x1_ASAP7_75t_SL g1582 ( 
.A(n_1562),
.B(n_1506),
.Y(n_1582)
);

AOI21xp33_ASAP7_75t_SL g1583 ( 
.A1(n_1546),
.A2(n_1533),
.B(n_1520),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1546),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1561),
.A2(n_1304),
.B1(n_1533),
.B2(n_1365),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1537),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1569),
.B(n_1243),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1546),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_SL g1589 ( 
.A1(n_1562),
.A2(n_1299),
.B1(n_1306),
.B2(n_1282),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1535),
.B(n_1489),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1568),
.B(n_1486),
.Y(n_1591)
);

OAI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1536),
.A2(n_1520),
.B1(n_1506),
.B2(n_1486),
.C(n_1474),
.Y(n_1592)
);

AOI222xp33_ASAP7_75t_L g1593 ( 
.A1(n_1556),
.A2(n_1452),
.B1(n_1447),
.B2(n_1449),
.C1(n_1426),
.C2(n_1245),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1562),
.A2(n_1449),
.B1(n_1445),
.B2(n_1427),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1553),
.A2(n_1299),
.B1(n_1282),
.B2(n_1306),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_1571),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1576),
.B(n_1562),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1586),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1580),
.B(n_1581),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1582),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1581),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1584),
.B(n_1588),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1572),
.B(n_1535),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1580),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1587),
.B(n_1541),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1573),
.B(n_1575),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1593),
.A2(n_1570),
.B1(n_1565),
.B2(n_1559),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1579),
.B(n_1538),
.Y(n_1608)
);

OAI222xp33_ASAP7_75t_L g1609 ( 
.A1(n_1574),
.A2(n_1541),
.B1(n_1550),
.B2(n_1542),
.C1(n_1538),
.C2(n_1547),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1578),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1583),
.B(n_1547),
.Y(n_1611)
);

OAI222xp33_ASAP7_75t_L g1612 ( 
.A1(n_1592),
.A2(n_1550),
.B1(n_1542),
.B2(n_1558),
.C1(n_1570),
.C2(n_1565),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1591),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1590),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1606),
.A2(n_1577),
.B1(n_1594),
.B2(n_1585),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_L g1616 ( 
.A(n_1606),
.B(n_1589),
.C(n_1594),
.Y(n_1616)
);

AOI221x1_ASAP7_75t_L g1617 ( 
.A1(n_1597),
.A2(n_1548),
.B1(n_1567),
.B2(n_1537),
.C(n_1544),
.Y(n_1617)
);

AOI311xp33_ASAP7_75t_L g1618 ( 
.A1(n_1609),
.A2(n_1564),
.A3(n_1567),
.B(n_1566),
.C(n_1554),
.Y(n_1618)
);

NAND3xp33_ASAP7_75t_L g1619 ( 
.A(n_1596),
.B(n_1548),
.C(n_1544),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1596),
.A2(n_1595),
.B1(n_1558),
.B2(n_1564),
.Y(n_1620)
);

AOI221xp5_ASAP7_75t_L g1621 ( 
.A1(n_1610),
.A2(n_1566),
.B1(n_1563),
.B2(n_1555),
.C(n_1554),
.Y(n_1621)
);

OAI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1607),
.A2(n_1563),
.B1(n_1551),
.B2(n_1555),
.C(n_1474),
.Y(n_1622)
);

AOI222xp33_ASAP7_75t_L g1623 ( 
.A1(n_1612),
.A2(n_1551),
.B1(n_1442),
.B2(n_1441),
.C1(n_1451),
.C2(n_1438),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1603),
.B(n_1599),
.Y(n_1624)
);

NAND3xp33_ASAP7_75t_L g1625 ( 
.A(n_1604),
.B(n_1245),
.C(n_1476),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1605),
.B(n_1253),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_L g1627 ( 
.A(n_1618),
.B(n_1600),
.C(n_1604),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1615),
.A2(n_1611),
.B1(n_1608),
.B2(n_1600),
.Y(n_1628)
);

NAND2x1p5_ASAP7_75t_L g1629 ( 
.A(n_1626),
.B(n_1602),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1616),
.B(n_1599),
.Y(n_1630)
);

NOR2x1_ASAP7_75t_L g1631 ( 
.A(n_1619),
.B(n_1602),
.Y(n_1631)
);

NAND4xp25_ASAP7_75t_L g1632 ( 
.A(n_1621),
.B(n_1624),
.C(n_1622),
.D(n_1625),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1620),
.B(n_1601),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1623),
.B(n_1602),
.Y(n_1634)
);

AOI211xp5_ASAP7_75t_L g1635 ( 
.A1(n_1617),
.A2(n_1613),
.B(n_1614),
.C(n_1598),
.Y(n_1635)
);

AOI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1616),
.A2(n_1471),
.B(n_1464),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1626),
.B(n_1489),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1631),
.B(n_1265),
.Y(n_1638)
);

NAND3xp33_ASAP7_75t_L g1639 ( 
.A(n_1627),
.B(n_1270),
.C(n_1441),
.Y(n_1639)
);

AOI211xp5_ASAP7_75t_L g1640 ( 
.A1(n_1630),
.A2(n_1232),
.B(n_1260),
.C(n_1275),
.Y(n_1640)
);

AOI221xp5_ASAP7_75t_L g1641 ( 
.A1(n_1628),
.A2(n_1451),
.B1(n_1442),
.B2(n_1441),
.C(n_1464),
.Y(n_1641)
);

AOI222xp33_ASAP7_75t_L g1642 ( 
.A1(n_1633),
.A2(n_1451),
.B1(n_1442),
.B2(n_1477),
.C1(n_1471),
.C2(n_1472),
.Y(n_1642)
);

NOR2x1_ASAP7_75t_L g1643 ( 
.A(n_1638),
.B(n_1632),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1640),
.A2(n_1634),
.B1(n_1637),
.B2(n_1629),
.Y(n_1644)
);

AND3x4_ASAP7_75t_L g1645 ( 
.A(n_1639),
.B(n_1635),
.C(n_1232),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1641),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1642),
.B(n_1636),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1639),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1648),
.Y(n_1649)
);

NOR2x1_ASAP7_75t_L g1650 ( 
.A(n_1643),
.B(n_1211),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1644),
.B(n_1646),
.Y(n_1651)
);

NOR2x1_ASAP7_75t_L g1652 ( 
.A(n_1645),
.B(n_1211),
.Y(n_1652)
);

OAI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1647),
.A2(n_1248),
.B1(n_1211),
.B2(n_1203),
.C(n_1477),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1650),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1651),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1652),
.B(n_1423),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1655),
.Y(n_1657)
);

NAND3xp33_ASAP7_75t_L g1658 ( 
.A(n_1657),
.B(n_1654),
.C(n_1649),
.Y(n_1658)
);

OAI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1658),
.A2(n_1653),
.B1(n_1654),
.B2(n_1656),
.C(n_1248),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1658),
.Y(n_1660)
);

OR2x6_ASAP7_75t_L g1661 ( 
.A(n_1660),
.B(n_1267),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_SL g1662 ( 
.A1(n_1659),
.A2(n_1254),
.B(n_1203),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1661),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1662),
.B(n_1472),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1663),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1665),
.A2(n_1664),
.B1(n_1270),
.B2(n_1254),
.Y(n_1666)
);

OAI221xp5_ASAP7_75t_R g1667 ( 
.A1(n_1666),
.A2(n_1267),
.B1(n_1273),
.B2(n_1331),
.C(n_1435),
.Y(n_1667)
);

AOI211xp5_ASAP7_75t_L g1668 ( 
.A1(n_1667),
.A2(n_1180),
.B(n_1450),
.C(n_1446),
.Y(n_1668)
);


endmodule