module real_aes_7908_n_350 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_350);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_350;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_635;
wire n_792;
wire n_386;
wire n_673;
wire n_503;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_991;
wire n_667;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_979;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1016;
wire n_908;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_963;
wire n_865;
wire n_666;
wire n_551;
wire n_884;
wire n_537;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_994;
wire n_578;
wire n_495;
wire n_892;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_774;
wire n_992;
wire n_813;
wire n_981;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_726;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_755;
wire n_532;
wire n_656;
wire n_746;
wire n_1025;
wire n_409;
wire n_781;
wire n_748;
wire n_909;
wire n_996;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_725;
wire n_455;
wire n_960;
wire n_671;
wire n_973;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_501;
wire n_488;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_756;
wire n_713;
wire n_735;
wire n_598;
wire n_728;
wire n_997;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_366;
wire n_727;
wire n_1014;
wire n_397;
wire n_749;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_831;
wire n_487;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_789;
wire n_544;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_721;
wire n_446;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_639;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_1039;
wire n_802;
wire n_877;
wire n_868;
wire n_574;
wire n_1024;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
wire n_869;
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_0), .A2(n_144), .B1(n_532), .B2(n_535), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_1), .A2(n_148), .B1(n_518), .B2(n_716), .Y(n_924) );
INVx1_ASAP7_75t_L g959 ( .A(n_2), .Y(n_959) );
AOI22xp33_ASAP7_75t_SL g565 ( .A1(n_3), .A2(n_317), .B1(n_368), .B2(n_513), .Y(n_565) );
AOI22xp33_ASAP7_75t_SL g891 ( .A1(n_4), .A2(n_116), .B1(n_535), .B2(n_789), .Y(n_891) );
AOI222xp33_ASAP7_75t_L g1040 ( .A1(n_5), .A2(n_158), .B1(n_305), .B2(n_444), .C1(n_450), .C2(n_865), .Y(n_1040) );
AOI222xp33_ASAP7_75t_L g503 ( .A1(n_6), .A2(n_172), .B1(n_269), .B2(n_444), .C1(n_449), .C2(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_7), .A2(n_84), .B1(n_531), .B2(n_551), .Y(n_594) );
AO22x2_ASAP7_75t_L g381 ( .A1(n_8), .A2(n_200), .B1(n_373), .B2(n_378), .Y(n_381) );
INVx1_ASAP7_75t_L g992 ( .A(n_8), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_9), .A2(n_152), .B1(n_884), .B2(n_951), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_10), .A2(n_133), .B1(n_417), .B2(n_485), .Y(n_816) );
AOI222xp33_ASAP7_75t_L g895 ( .A1(n_11), .A2(n_295), .B1(n_306), .B2(n_583), .C1(n_627), .C2(n_652), .Y(n_895) );
CKINVDCx20_ASAP7_75t_R g973 ( .A(n_12), .Y(n_973) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_13), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_14), .A2(n_41), .B1(n_839), .B2(n_972), .Y(n_971) );
AOI22xp33_ASAP7_75t_SL g668 ( .A1(n_15), .A2(n_105), .B1(n_491), .B2(n_669), .Y(n_668) );
AOI22xp33_ASAP7_75t_SL g651 ( .A1(n_16), .A2(n_257), .B1(n_627), .B2(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g954 ( .A(n_17), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_18), .A2(n_286), .B1(n_483), .B2(n_620), .Y(n_619) );
AOI22xp5_ASAP7_75t_SL g515 ( .A1(n_19), .A2(n_175), .B1(n_516), .B2(n_518), .Y(n_515) );
AOI22xp33_ASAP7_75t_SL g665 ( .A1(n_20), .A2(n_237), .B1(n_420), .B2(n_666), .Y(n_665) );
AOI22xp33_ASAP7_75t_SL g600 ( .A1(n_21), .A2(n_187), .B1(n_416), .B2(n_420), .Y(n_600) );
AOI22xp33_ASAP7_75t_SL g960 ( .A1(n_22), .A2(n_176), .B1(n_437), .B2(n_450), .Y(n_960) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_23), .A2(n_94), .B1(n_473), .B2(n_474), .C(n_476), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_24), .A2(n_136), .B1(n_599), .B2(n_721), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_25), .A2(n_289), .B1(n_837), .B2(n_839), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_26), .A2(n_96), .B1(n_676), .B2(n_884), .Y(n_947) );
AOI22xp33_ASAP7_75t_SL g596 ( .A1(n_27), .A2(n_118), .B1(n_524), .B2(n_597), .Y(n_596) );
AO22x2_ASAP7_75t_L g383 ( .A1(n_28), .A2(n_102), .B1(n_373), .B2(n_374), .Y(n_383) );
AOI22xp33_ASAP7_75t_SL g559 ( .A1(n_29), .A2(n_245), .B1(n_417), .B2(n_560), .Y(n_559) );
AOI222xp33_ASAP7_75t_L g824 ( .A1(n_30), .A2(n_174), .B1(n_268), .B2(n_450), .C1(n_790), .C2(n_825), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_31), .B(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_32), .A2(n_59), .B1(n_483), .B2(n_560), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_33), .A2(n_236), .B1(n_599), .B2(n_869), .Y(n_868) );
CKINVDCx20_ASAP7_75t_R g934 ( .A(n_34), .Y(n_934) );
AOI221xp5_ASAP7_75t_L g492 ( .A1(n_35), .A2(n_183), .B1(n_493), .B2(n_496), .C(n_499), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_36), .Y(n_442) );
AOI22xp33_ASAP7_75t_SL g663 ( .A1(n_37), .A2(n_104), .B1(n_474), .B2(n_664), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g995 ( .A1(n_38), .A2(n_996), .B1(n_997), .B2(n_1019), .Y(n_995) );
CKINVDCx20_ASAP7_75t_R g1019 ( .A(n_38), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_39), .A2(n_80), .B1(n_560), .B2(n_567), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_40), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_42), .A2(n_126), .B1(n_676), .B2(n_1000), .Y(n_999) );
INVx1_ASAP7_75t_L g1011 ( .A(n_43), .Y(n_1011) );
AOI22x1_ASAP7_75t_L g363 ( .A1(n_44), .A2(n_364), .B1(n_467), .B2(n_468), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_44), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_45), .A2(n_90), .B1(n_398), .B2(n_749), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_46), .A2(n_206), .B1(n_560), .B2(n_951), .Y(n_970) );
CKINVDCx20_ASAP7_75t_R g1027 ( .A(n_47), .Y(n_1027) );
AOI222xp33_ASAP7_75t_L g791 ( .A1(n_48), .A2(n_156), .B1(n_314), .B2(n_445), .C1(n_541), .C2(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_49), .A2(n_78), .B1(n_841), .B2(n_886), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_50), .A2(n_281), .B1(n_482), .B2(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g489 ( .A(n_51), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_52), .A2(n_167), .B1(n_551), .B2(n_659), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_53), .A2(n_65), .B1(n_657), .B2(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g568 ( .A(n_54), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_55), .B(n_657), .Y(n_890) );
AOI22xp33_ASAP7_75t_SL g602 ( .A1(n_56), .A2(n_348), .B1(n_473), .B2(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_SL g566 ( .A1(n_57), .A2(n_204), .B1(n_398), .B2(n_567), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_58), .A2(n_308), .B1(n_778), .B2(n_781), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_60), .A2(n_344), .B1(n_659), .B2(n_790), .Y(n_1006) );
CKINVDCx20_ASAP7_75t_R g943 ( .A(n_61), .Y(n_943) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_62), .Y(n_624) );
AOI22xp33_ASAP7_75t_SL g562 ( .A1(n_63), .A2(n_232), .B1(n_474), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_64), .A2(n_252), .B1(n_535), .B2(n_846), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g909 ( .A(n_66), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_67), .A2(n_180), .B1(n_416), .B2(n_420), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_68), .A2(n_228), .B1(n_560), .B2(n_721), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g481 ( .A1(n_69), .A2(n_92), .B1(n_482), .B2(n_483), .C(n_486), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_70), .Y(n_769) );
AO22x2_ASAP7_75t_L g377 ( .A1(n_71), .A2(n_235), .B1(n_373), .B2(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g989 ( .A(n_71), .Y(n_989) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_72), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_73), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_74), .A2(n_89), .B1(n_483), .B2(n_686), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_75), .A2(n_213), .B1(n_474), .B2(n_620), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_76), .A2(n_128), .B1(n_531), .B2(n_865), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_77), .A2(n_195), .B1(n_531), .B2(n_534), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_79), .Y(n_431) );
AOI22xp33_ASAP7_75t_SL g556 ( .A1(n_81), .A2(n_247), .B1(n_437), .B2(n_532), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_82), .A2(n_168), .B1(n_529), .B2(n_681), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_83), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_85), .A2(n_765), .B1(n_793), .B2(n_794), .Y(n_764) );
CKINVDCx16_ASAP7_75t_R g793 ( .A(n_85), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_86), .Y(n_736) );
AOI222xp33_ASAP7_75t_L g809 ( .A1(n_87), .A2(n_98), .B1(n_160), .B2(n_444), .C1(n_652), .C2(n_661), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_88), .A2(n_342), .B1(n_504), .B2(n_789), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_91), .A2(n_240), .B1(n_398), .B2(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g500 ( .A(n_93), .Y(n_500) );
XOR2x2_ASAP7_75t_L g850 ( .A(n_95), .B(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g539 ( .A(n_97), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_99), .A2(n_251), .B1(n_664), .B2(n_775), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_100), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_101), .A2(n_244), .B1(n_406), .B2(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g993 ( .A(n_102), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_103), .A2(n_238), .B1(n_392), .B2(n_397), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_106), .A2(n_271), .B1(n_392), .B2(n_473), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_107), .Y(n_447) );
XOR2x2_ASAP7_75t_L g645 ( .A(n_108), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_109), .B(n_863), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_110), .Y(n_786) );
AO22x1_ASAP7_75t_L g829 ( .A1(n_111), .A2(n_830), .B1(n_831), .B2(n_848), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_111), .Y(n_848) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_112), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_113), .A2(n_130), .B1(n_421), .B2(n_783), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_114), .B(n_861), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_115), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_117), .A2(n_320), .B1(n_368), .B2(n_394), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_119), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_120), .A2(n_471), .B1(n_505), .B2(n_506), .Y(n_470) );
INVx1_ASAP7_75t_L g505 ( .A(n_120), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_121), .A2(n_163), .B1(n_417), .B2(n_421), .Y(n_1032) );
INVx1_ASAP7_75t_L g487 ( .A(n_122), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_123), .A2(n_143), .B1(n_386), .B2(n_923), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_124), .A2(n_315), .B1(n_666), .B2(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_125), .A2(n_203), .B1(n_671), .B2(n_920), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_127), .A2(n_140), .B1(n_518), .B2(n_841), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_129), .A2(n_329), .B1(n_781), .B2(n_871), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_131), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_132), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_134), .A2(n_186), .B1(n_789), .B2(n_790), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_135), .A2(n_273), .B1(n_686), .B2(n_884), .Y(n_883) );
AND2x6_ASAP7_75t_L g353 ( .A(n_137), .B(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g986 ( .A(n_137), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_138), .A2(n_256), .B1(n_678), .B2(n_716), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_139), .A2(n_302), .B1(n_450), .B2(n_504), .Y(n_941) );
AOI22xp33_ASAP7_75t_SL g585 ( .A1(n_141), .A2(n_241), .B1(n_586), .B2(n_589), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_142), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_145), .A2(n_294), .B1(n_716), .B2(n_718), .Y(n_715) );
AOI222xp33_ASAP7_75t_L g1018 ( .A1(n_146), .A2(n_218), .B1(n_234), .B2(n_445), .C1(n_504), .C2(n_589), .Y(n_1018) );
CKINVDCx20_ASAP7_75t_R g896 ( .A(n_147), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_149), .A2(n_280), .B1(n_522), .B2(n_676), .Y(n_675) );
AOI22xp33_ASAP7_75t_SL g605 ( .A1(n_150), .A2(n_311), .B1(n_404), .B2(n_525), .Y(n_605) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_151), .Y(n_408) );
AOI22xp33_ASAP7_75t_SL g968 ( .A1(n_153), .A2(n_331), .B1(n_563), .B2(n_783), .Y(n_968) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_154), .A2(n_284), .B1(n_522), .B2(n_525), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_155), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_157), .A2(n_229), .B1(n_416), .B2(n_420), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g874 ( .A1(n_159), .A2(n_223), .B1(n_689), .B2(n_716), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_161), .A2(n_316), .B1(n_775), .B2(n_953), .Y(n_952) );
AO22x2_ASAP7_75t_L g372 ( .A1(n_162), .A2(n_224), .B1(n_373), .B2(n_374), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g990 ( .A(n_162), .B(n_991), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_164), .A2(n_192), .B1(n_387), .B2(n_678), .Y(n_875) );
CKINVDCx20_ASAP7_75t_R g888 ( .A(n_165), .Y(n_888) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_166), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_169), .A2(n_339), .B1(n_688), .B2(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g584 ( .A(n_170), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_171), .A2(n_225), .B1(n_780), .B2(n_972), .Y(n_1031) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_173), .Y(n_650) );
AOI222xp33_ASAP7_75t_L g847 ( .A1(n_177), .A2(n_301), .B1(n_310), .B2(n_437), .C1(n_444), .C2(n_449), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_178), .B(n_550), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_179), .A2(n_227), .B1(n_685), .B2(n_686), .Y(n_684) );
XOR2x2_ASAP7_75t_L g796 ( .A(n_181), .B(n_797), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_182), .A2(n_276), .B1(n_528), .B2(n_529), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_184), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_185), .Y(n_787) );
INVx1_ASAP7_75t_L g1013 ( .A(n_188), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_189), .B(n_593), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_190), .A2(n_272), .B1(n_528), .B2(n_555), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_191), .B(n_528), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_193), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_194), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_196), .A2(n_243), .B1(n_368), .B2(n_783), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_197), .B(n_529), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_198), .A2(n_263), .B1(n_474), .B2(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_SL g549 ( .A1(n_199), .A2(n_221), .B1(n_550), .B2(n_551), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_201), .A2(n_255), .B1(n_524), .B2(n_563), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_202), .A2(n_265), .B1(n_659), .B2(n_661), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_205), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_207), .A2(n_338), .B1(n_421), .B2(n_513), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_208), .A2(n_340), .B1(n_686), .B2(n_839), .Y(n_1035) );
CKINVDCx20_ASAP7_75t_R g390 ( .A(n_209), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_210), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g904 ( .A(n_211), .Y(n_904) );
INVx1_ASAP7_75t_L g1009 ( .A(n_212), .Y(n_1009) );
INVx1_ASAP7_75t_L g502 ( .A(n_214), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_215), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_216), .A2(n_304), .B1(n_504), .B2(n_789), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_217), .A2(n_239), .B1(n_421), .B2(n_783), .Y(n_782) );
AOI222xp33_ASAP7_75t_L g690 ( .A1(n_219), .A2(n_319), .B1(n_332), .B2(n_437), .C1(n_445), .C2(n_449), .Y(n_690) );
AND2x2_ASAP7_75t_L g357 ( .A(n_220), .B(n_358), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_222), .A2(n_253), .B1(n_550), .B2(n_857), .Y(n_856) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_226), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_230), .A2(n_270), .B1(n_450), .B2(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_231), .A2(n_336), .B1(n_620), .B2(n_749), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_233), .Y(n_738) );
INVx1_ASAP7_75t_L g944 ( .A(n_242), .Y(n_944) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_246), .A2(n_732), .B1(n_755), .B2(n_756), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_246), .Y(n_755) );
AOI22xp33_ASAP7_75t_SL g670 ( .A1(n_248), .A2(n_347), .B1(n_485), .B2(n_671), .Y(n_670) );
XOR2x2_ASAP7_75t_L g578 ( .A(n_249), .B(n_579), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_250), .Y(n_706) );
INVx1_ASAP7_75t_L g373 ( .A(n_254), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_254), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_258), .A2(n_337), .B1(n_416), .B2(n_420), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_259), .B(n_657), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g905 ( .A(n_260), .Y(n_905) );
INVx1_ASAP7_75t_L g480 ( .A(n_261), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_262), .B(n_555), .Y(n_962) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_264), .A2(n_608), .B1(n_636), .B2(n_637), .Y(n_607) );
INVx1_ASAP7_75t_L g636 ( .A(n_264), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_266), .Y(n_704) );
AOI211xp5_ASAP7_75t_L g350 ( .A1(n_267), .A2(n_351), .B(n_359), .C(n_994), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_274), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g912 ( .A(n_275), .Y(n_912) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_277), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_278), .A2(n_312), .B1(n_534), .B2(n_789), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_279), .B(n_493), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_282), .A2(n_346), .B1(n_498), .B2(n_657), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_283), .A2(n_321), .B1(n_723), .B2(n_725), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_285), .Y(n_714) );
INVx1_ASAP7_75t_L g358 ( .A(n_287), .Y(n_358) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_288), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_290), .B(n_741), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g908 ( .A(n_291), .Y(n_908) );
INVx1_ASAP7_75t_L g354 ( .A(n_292), .Y(n_354) );
INVx1_ASAP7_75t_L g542 ( .A(n_293), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_296), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g855 ( .A(n_297), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_298), .A2(n_303), .B1(n_398), .B2(n_513), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g939 ( .A(n_299), .Y(n_939) );
INVx1_ASAP7_75t_L g1016 ( .A(n_300), .Y(n_1016) );
CKINVDCx20_ASAP7_75t_R g914 ( .A(n_307), .Y(n_914) );
INVx1_ASAP7_75t_L g477 ( .A(n_309), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g414 ( .A(n_313), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_318), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g1037 ( .A(n_322), .Y(n_1037) );
INVx1_ASAP7_75t_L g1003 ( .A(n_323), .Y(n_1003) );
CKINVDCx20_ASAP7_75t_R g634 ( .A(n_324), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_325), .B(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_SL g967 ( .A1(n_326), .A2(n_343), .B1(n_685), .B2(n_953), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_327), .B(n_529), .Y(n_655) );
XOR2x2_ASAP7_75t_L g672 ( .A(n_328), .B(n_673), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_330), .A2(n_692), .B1(n_726), .B2(n_727), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_330), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_333), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_334), .B(n_1005), .Y(n_1004) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_335), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_341), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g900 ( .A1(n_345), .A2(n_901), .B1(n_925), .B2(n_926), .Y(n_900) );
INVx1_ASAP7_75t_L g925 ( .A(n_345), .Y(n_925) );
CKINVDCx20_ASAP7_75t_R g936 ( .A(n_349), .Y(n_936) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
HB1xp67_ASAP7_75t_L g985 ( .A(n_354), .Y(n_985) );
OAI21xp5_ASAP7_75t_L g1025 ( .A1(n_355), .A2(n_984), .B(n_1026), .Y(n_1025) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_760), .B1(n_979), .B2(n_980), .C(n_981), .Y(n_359) );
INVx1_ASAP7_75t_L g979 ( .A(n_360), .Y(n_979) );
XOR2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_573), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_363), .B1(n_469), .B2(n_572), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g468 ( .A(n_364), .Y(n_468) );
AND2x2_ASAP7_75t_SL g364 ( .A(n_365), .B(n_424), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_366), .B(n_402), .Y(n_365) );
OAI221xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_384), .B1(n_385), .B2(n_390), .C(n_391), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_368), .Y(n_473) );
BUFx3_ASAP7_75t_L g620 ( .A(n_368), .Y(n_620) );
BUFx3_ASAP7_75t_L g923 ( .A(n_368), .Y(n_923) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_SL g664 ( .A(n_369), .Y(n_664) );
BUFx2_ASAP7_75t_SL g676 ( .A(n_369), .Y(n_676) );
INVx2_ASAP7_75t_L g872 ( .A(n_369), .Y(n_872) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_379), .Y(n_369) );
AND2x6_ASAP7_75t_L g394 ( .A(n_370), .B(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g406 ( .A(n_370), .B(n_407), .Y(n_406) );
AND2x6_ASAP7_75t_L g445 ( .A(n_370), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_376), .Y(n_370) );
AND2x2_ASAP7_75t_L g389 ( .A(n_371), .B(n_377), .Y(n_389) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_372), .B(n_377), .Y(n_401) );
AND2x2_ASAP7_75t_L g412 ( .A(n_372), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g441 ( .A(n_372), .B(n_381), .Y(n_441) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g378 ( .A(n_375), .Y(n_378) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g413 ( .A(n_377), .Y(n_413) );
INVx1_ASAP7_75t_L g440 ( .A(n_377), .Y(n_440) );
AND2x4_ASAP7_75t_L g388 ( .A(n_379), .B(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g399 ( .A(n_379), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_379), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g514 ( .A(n_379), .B(n_412), .Y(n_514) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
OR2x2_ASAP7_75t_L g396 ( .A(n_380), .B(n_383), .Y(n_396) );
AND2x2_ASAP7_75t_L g407 ( .A(n_380), .B(n_383), .Y(n_407) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g446 ( .A(n_381), .B(n_383), .Y(n_446) );
AND2x2_ASAP7_75t_L g439 ( .A(n_382), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g459 ( .A(n_382), .Y(n_459) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g423 ( .A(n_383), .Y(n_423) );
OAI221xp5_ASAP7_75t_SL g615 ( .A1(n_385), .A2(n_616), .B1(n_617), .B2(n_618), .C(n_619), .Y(n_615) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g475 ( .A(n_388), .Y(n_475) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_388), .Y(n_524) );
BUFx3_ASAP7_75t_L g775 ( .A(n_388), .Y(n_775) );
BUFx3_ASAP7_75t_L g839 ( .A(n_388), .Y(n_839) );
INVx1_ASAP7_75t_L g430 ( .A(n_389), .Y(n_430) );
NAND2x1p5_ASAP7_75t_L g434 ( .A(n_389), .B(n_407), .Y(n_434) );
AND2x4_ASAP7_75t_L g495 ( .A(n_389), .B(n_395), .Y(n_495) );
AND2x6_ASAP7_75t_L g498 ( .A(n_389), .B(n_407), .Y(n_498) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx4_ASAP7_75t_L g482 ( .A(n_393), .Y(n_482) );
INVx2_ASAP7_75t_SL g599 ( .A(n_393), .Y(n_599) );
INVx1_ASAP7_75t_L g688 ( .A(n_393), .Y(n_688) );
INVx5_ASAP7_75t_SL g780 ( .A(n_393), .Y(n_780) );
HB1xp67_ASAP7_75t_L g838 ( .A(n_393), .Y(n_838) );
INVx11_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx11_ASAP7_75t_L g561 ( .A(n_394), .Y(n_561) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g429 ( .A(n_396), .B(n_430), .Y(n_429) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g612 ( .A(n_398), .Y(n_612) );
BUFx3_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_SL g491 ( .A(n_399), .Y(n_491) );
BUFx2_ASAP7_75t_SL g525 ( .A(n_399), .Y(n_525) );
BUFx3_ASAP7_75t_L g686 ( .A(n_399), .Y(n_686) );
BUFx3_ASAP7_75t_L g725 ( .A(n_399), .Y(n_725) );
BUFx3_ASAP7_75t_L g781 ( .A(n_399), .Y(n_781) );
INVx1_ASAP7_75t_L g805 ( .A(n_399), .Y(n_805) );
BUFx2_ASAP7_75t_L g953 ( .A(n_399), .Y(n_953) );
AND2x2_ASAP7_75t_L g563 ( .A(n_400), .B(n_459), .Y(n_563) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OR2x6_ASAP7_75t_L g422 ( .A(n_401), .B(n_423), .Y(n_422) );
OAI221xp5_ASAP7_75t_SL g402 ( .A1(n_403), .A2(n_408), .B1(n_409), .B2(n_414), .C(n_415), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_403), .A2(n_409), .B1(n_768), .B2(n_769), .Y(n_767) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g689 ( .A(n_405), .Y(n_689) );
INVx2_ASAP7_75t_L g920 ( .A(n_405), .Y(n_920) );
INVx3_ASAP7_75t_L g951 ( .A(n_405), .Y(n_951) );
INVx6_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx3_ASAP7_75t_L g485 ( .A(n_406), .Y(n_485) );
BUFx3_ASAP7_75t_L g567 ( .A(n_406), .Y(n_567) );
BUFx3_ASAP7_75t_L g721 ( .A(n_406), .Y(n_721) );
AND2x2_ASAP7_75t_L g419 ( .A(n_407), .B(n_412), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_407), .B(n_412), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g1008 ( .A1(n_409), .A2(n_1009), .B1(n_1010), .B2(n_1011), .Y(n_1008) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g488 ( .A(n_410), .Y(n_488) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g466 ( .A(n_413), .Y(n_466) );
BUFx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_417), .Y(n_666) );
INVx5_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx4_ASAP7_75t_L g517 ( .A(n_418), .Y(n_517) );
BUFx3_ASAP7_75t_L g717 ( .A(n_418), .Y(n_717) );
INVx2_ASAP7_75t_L g783 ( .A(n_418), .Y(n_783) );
INVx3_ASAP7_75t_L g841 ( .A(n_418), .Y(n_841) );
INVx8_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx2_ASAP7_75t_L g518 ( .A(n_421), .Y(n_518) );
BUFx2_ASAP7_75t_L g678 ( .A(n_421), .Y(n_678) );
BUFx2_ASAP7_75t_L g886 ( .A(n_421), .Y(n_886) );
INVx6_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_422), .A2(n_477), .B1(n_478), .B2(n_480), .Y(n_476) );
INVx1_ASAP7_75t_SL g718 ( .A(n_422), .Y(n_718) );
INVx1_ASAP7_75t_L g533 ( .A(n_423), .Y(n_533) );
NOR3xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_435), .C(n_454), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B1(n_431), .B2(n_432), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_427), .A2(n_432), .B1(n_623), .B2(n_624), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_427), .A2(n_698), .B1(n_735), .B2(n_736), .Y(n_734) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_429), .Y(n_696) );
BUFx3_ASAP7_75t_L g935 ( .A(n_429), .Y(n_935) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_SL g906 ( .A(n_433), .Y(n_906) );
INVx1_ASAP7_75t_L g937 ( .A(n_433), .Y(n_937) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx3_ASAP7_75t_L g700 ( .A(n_434), .Y(n_700) );
OAI222xp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_442), .B1(n_443), .B2(n_447), .C1(n_448), .C2(n_453), .Y(n_435) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_436), .A2(n_649), .B1(n_738), .B2(n_739), .C(n_740), .Y(n_737) );
OAI221xp5_ASAP7_75t_SL g907 ( .A1(n_436), .A2(n_537), .B1(n_908), .B2(n_909), .C(n_910), .Y(n_907) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g702 ( .A(n_437), .Y(n_702) );
BUFx4f_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_438), .Y(n_504) );
BUFx2_ASAP7_75t_L g541 ( .A(n_438), .Y(n_541) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_438), .Y(n_588) );
BUFx6f_ASAP7_75t_L g865 ( .A(n_438), .Y(n_865) );
AND2x4_ASAP7_75t_L g438 ( .A(n_439), .B(n_441), .Y(n_438) );
INVx1_ASAP7_75t_L g452 ( .A(n_440), .Y(n_452) );
AND2x4_ASAP7_75t_L g451 ( .A(n_441), .B(n_452), .Y(n_451) );
NAND2x1p5_ASAP7_75t_L g458 ( .A(n_441), .B(n_459), .Y(n_458) );
AND2x4_ASAP7_75t_L g532 ( .A(n_441), .B(n_533), .Y(n_532) );
OAI222xp33_ASAP7_75t_L g625 ( .A1(n_443), .A2(n_626), .B1(n_628), .B2(n_629), .C1(n_630), .C2(n_632), .Y(n_625) );
OAI222xp33_ASAP7_75t_L g701 ( .A1(n_443), .A2(n_702), .B1(n_703), .B2(n_704), .C1(n_705), .C2(n_706), .Y(n_701) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_SL g649 ( .A(n_444), .Y(n_649) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx4_ASAP7_75t_L g538 ( .A(n_445), .Y(n_538) );
INVx2_ASAP7_75t_L g547 ( .A(n_445), .Y(n_547) );
BUFx3_ASAP7_75t_L g825 ( .A(n_445), .Y(n_825) );
INVx2_ASAP7_75t_SL g854 ( .A(n_445), .Y(n_854) );
INVx1_ASAP7_75t_L g464 ( .A(n_446), .Y(n_464) );
AND2x4_ASAP7_75t_L g535 ( .A(n_446), .B(n_466), .Y(n_535) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx4f_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g653 ( .A(n_450), .Y(n_653) );
BUFx12f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_451), .Y(n_550) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_451), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B1(n_460), .B2(n_461), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_456), .A2(n_461), .B1(n_634), .B2(n_635), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_456), .A2(n_461), .B1(n_708), .B2(n_709), .Y(n_707) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx3_ASAP7_75t_SL g913 ( .A(n_457), .Y(n_913) );
INVx4_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx3_ASAP7_75t_L g501 ( .A(n_458), .Y(n_501) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_458), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_461), .A2(n_743), .B1(n_744), .B2(n_745), .Y(n_742) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
CKINVDCx16_ASAP7_75t_R g462 ( .A(n_463), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_463), .A2(n_500), .B1(n_501), .B2(n_502), .Y(n_499) );
BUFx2_ASAP7_75t_L g915 ( .A(n_463), .Y(n_915) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_463), .A2(n_501), .B1(n_943), .B2(n_944), .Y(n_942) );
OR2x6_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_SL g572 ( .A(n_469), .Y(n_572) );
OA22x2_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_507), .B1(n_508), .B2(n_571), .Y(n_469) );
INVx1_ASAP7_75t_L g571 ( .A(n_470), .Y(n_571) );
INVx1_ASAP7_75t_L g506 ( .A(n_471), .Y(n_506) );
AND4x1_ASAP7_75t_L g471 ( .A(n_472), .B(n_481), .C(n_492), .D(n_503), .Y(n_471) );
INVx1_ASAP7_75t_SL g772 ( .A(n_473), .Y(n_772) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx2_ASAP7_75t_R g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_SL g616 ( .A(n_482), .Y(n_616) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B1(n_489), .B2(n_490), .Y(n_486) );
OAI221xp5_ASAP7_75t_SL g610 ( .A1(n_488), .A2(n_611), .B1(n_612), .B2(n_613), .C(n_614), .Y(n_610) );
INVx1_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g1005 ( .A(n_493), .Y(n_1005) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g528 ( .A(n_494), .Y(n_528) );
INVx2_ASAP7_75t_L g593 ( .A(n_494), .Y(n_593) );
INVx5_ASAP7_75t_L g657 ( .A(n_494), .Y(n_657) );
INVx4_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_SL g529 ( .A(n_497), .Y(n_529) );
INVx1_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
BUFx4f_ASAP7_75t_L g555 ( .A(n_498), .Y(n_555) );
BUFx2_ASAP7_75t_L g844 ( .A(n_498), .Y(n_844) );
BUFx2_ASAP7_75t_L g863 ( .A(n_498), .Y(n_863) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_504), .Y(n_627) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_543), .B1(n_569), .B2(n_570), .Y(n_508) );
INVx2_ASAP7_75t_SL g569 ( .A(n_509), .Y(n_569) );
XOR2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_542), .Y(n_509) );
NOR4xp75_ASAP7_75t_L g510 ( .A(n_511), .B(n_519), .C(n_526), .D(n_536), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_512), .B(n_515), .Y(n_511) );
INVx1_ASAP7_75t_L g604 ( .A(n_513), .Y(n_604) );
BUFx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx3_ASAP7_75t_L g669 ( .A(n_514), .Y(n_669) );
BUFx3_ASAP7_75t_L g685 ( .A(n_514), .Y(n_685) );
BUFx3_ASAP7_75t_L g884 ( .A(n_514), .Y(n_884) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2x1_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
INVx4_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
OAI221xp5_ASAP7_75t_SL g711 ( .A1(n_523), .A2(n_712), .B1(n_713), .B2(n_714), .C(n_715), .Y(n_711) );
INVx3_ASAP7_75t_L g1000 ( .A(n_523), .Y(n_1000) );
INVx4_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_527), .B(n_530), .Y(n_526) );
BUFx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g660 ( .A(n_532), .Y(n_660) );
BUFx3_ASAP7_75t_L g789 ( .A(n_532), .Y(n_789) );
BUFx2_ASAP7_75t_L g846 ( .A(n_532), .Y(n_846) );
INVx1_ASAP7_75t_SL g858 ( .A(n_534), .Y(n_858) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx2_ASAP7_75t_SL g551 ( .A(n_535), .Y(n_551) );
BUFx2_ASAP7_75t_SL g661 ( .A(n_535), .Y(n_661) );
BUFx3_ASAP7_75t_L g790 ( .A(n_535), .Y(n_790) );
OAI21xp5_ASAP7_75t_SL g536 ( .A1(n_537), .A2(n_539), .B(n_540), .Y(n_536) );
BUFx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx4_ASAP7_75t_L g583 ( .A(n_538), .Y(n_583) );
INVx1_ASAP7_75t_L g570 ( .A(n_543), .Y(n_570) );
XOR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_568), .Y(n_543) );
NAND2x1_ASAP7_75t_L g544 ( .A(n_545), .B(n_557), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_552), .Y(n_545) );
OAI21xp5_ASAP7_75t_SL g546 ( .A1(n_547), .A2(n_548), .B(n_549), .Y(n_546) );
BUFx3_ASAP7_75t_L g631 ( .A(n_550), .Y(n_631) );
INVx2_ASAP7_75t_L g705 ( .A(n_550), .Y(n_705) );
BUFx2_ASAP7_75t_L g792 ( .A(n_550), .Y(n_792) );
NAND3xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .C(n_556), .Y(n_552) );
NOR2x1_ASAP7_75t_L g557 ( .A(n_558), .B(n_564), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_562), .Y(n_558) );
INVx4_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_SL g671 ( .A(n_561), .Y(n_671) );
INVx3_ASAP7_75t_L g1015 ( .A(n_561), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_639), .B1(n_640), .B2(n_759), .Y(n_573) );
INVx1_ASAP7_75t_L g759 ( .A(n_574), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B1(n_606), .B2(n_638), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND3x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_595), .C(n_601), .Y(n_579) );
NOR2x1_ASAP7_75t_SL g580 ( .A(n_581), .B(n_590), .Y(n_580) );
OAI21xp5_ASAP7_75t_SL g581 ( .A1(n_582), .A2(n_584), .B(n_585), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx4_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
BUFx4f_ASAP7_75t_L g741 ( .A(n_589), .Y(n_741) );
NAND3xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .C(n_594), .Y(n_590) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_600), .Y(n_595) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_605), .Y(n_601) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g638 ( .A(n_606), .Y(n_638) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g637 ( .A(n_608), .Y(n_637) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_621), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_615), .Y(n_609) );
NOR3xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_625), .C(n_633), .Y(n_621) );
INVx2_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_729), .B2(n_730), .Y(n_640) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_644), .B1(n_691), .B2(n_728), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
XNOR2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_672), .Y(n_644) );
NAND3xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_662), .C(n_667), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_654), .Y(n_647) );
OAI21xp5_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_650), .B(n_651), .Y(n_648) );
INVx3_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .C(n_658), .Y(n_654) );
BUFx6f_ASAP7_75t_L g681 ( .A(n_657), .Y(n_681) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_657), .Y(n_861) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g724 ( .A(n_669), .Y(n_724) );
BUFx4f_ASAP7_75t_SL g869 ( .A(n_669), .Y(n_869) );
OA22x2_ASAP7_75t_L g730 ( .A1(n_672), .A2(n_731), .B1(n_757), .B2(n_758), .Y(n_730) );
INVx1_ASAP7_75t_L g758 ( .A(n_672), .Y(n_758) );
NAND4xp75_ASAP7_75t_L g673 ( .A(n_674), .B(n_679), .C(n_683), .D(n_690), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
INVx1_ASAP7_75t_L g712 ( .A(n_676), .Y(n_712) );
AND2x2_ASAP7_75t_SL g679 ( .A(n_680), .B(n_682), .Y(n_679) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_687), .Y(n_683) );
INVx1_ASAP7_75t_L g750 ( .A(n_685), .Y(n_750) );
INVxp67_ASAP7_75t_L g1010 ( .A(n_686), .Y(n_1010) );
INVx1_ASAP7_75t_L g728 ( .A(n_691), .Y(n_728) );
INVx1_ASAP7_75t_L g727 ( .A(n_692), .Y(n_727) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_710), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_701), .C(n_707), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_697), .B2(n_698), .Y(n_694) );
OAI221xp5_ASAP7_75t_SL g785 ( .A1(n_696), .A2(n_698), .B1(n_786), .B2(n_787), .C(n_788), .Y(n_785) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_696), .A2(n_904), .B1(n_905), .B2(n_906), .Y(n_903) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
BUFx3_ASAP7_75t_L g889 ( .A(n_700), .Y(n_889) );
OA211x2_ASAP7_75t_L g1036 ( .A1(n_700), .A2(n_1037), .B(n_1038), .C(n_1039), .Y(n_1036) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_719), .Y(n_710) );
INVx3_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_720), .B(n_722), .Y(n_719) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx3_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g757 ( .A(n_731), .Y(n_757) );
INVx2_ASAP7_75t_L g756 ( .A(n_732), .Y(n_756) );
AND2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_746), .Y(n_732) );
NOR3xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_737), .C(n_742), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_752), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_751), .Y(n_747) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g980 ( .A(n_760), .Y(n_980) );
AOI22xp5_ASAP7_75t_SL g760 ( .A1(n_761), .A2(n_879), .B1(n_977), .B2(n_978), .Y(n_760) );
INVx1_ASAP7_75t_L g977 ( .A(n_761), .Y(n_977) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_763), .B1(n_812), .B2(n_878), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_795), .B1(n_810), .B2(n_811), .Y(n_763) );
INVx1_ASAP7_75t_L g810 ( .A(n_764), .Y(n_810) );
INVx2_ASAP7_75t_SL g794 ( .A(n_765), .Y(n_794) );
AND4x1_ASAP7_75t_L g765 ( .A(n_766), .B(n_776), .C(n_784), .D(n_791), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_770), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_770) );
INVxp67_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
AND2x2_ASAP7_75t_L g776 ( .A(n_777), .B(n_782), .Y(n_776) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVxp67_ASAP7_75t_L g811 ( .A(n_795), .Y(n_811) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
XOR2x2_ASAP7_75t_L g849 ( .A(n_796), .B(n_850), .Y(n_849) );
NAND4xp75_ASAP7_75t_L g797 ( .A(n_798), .B(n_801), .C(n_806), .D(n_809), .Y(n_797) );
AND2x2_ASAP7_75t_SL g798 ( .A(n_799), .B(n_800), .Y(n_798) );
AND2x2_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
INVx1_ASAP7_75t_L g878 ( .A(n_812), .Y(n_878) );
AOI22xp5_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_827), .B1(n_876), .B2(n_877), .Y(n_812) );
INVx2_ASAP7_75t_SL g876 ( .A(n_813), .Y(n_876) );
XOR2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_826), .Y(n_813) );
NAND4xp75_ASAP7_75t_L g814 ( .A(n_815), .B(n_818), .C(n_821), .D(n_824), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
AND2x2_ASAP7_75t_SL g818 ( .A(n_819), .B(n_820), .Y(n_818) );
AND2x2_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
INVx3_ASAP7_75t_L g940 ( .A(n_825), .Y(n_940) );
INVx2_ASAP7_75t_L g877 ( .A(n_827), .Y(n_877) );
XNOR2x1_ASAP7_75t_L g827 ( .A(n_828), .B(n_849), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_SL g830 ( .A(n_831), .Y(n_830) );
NAND4xp75_ASAP7_75t_SL g831 ( .A(n_832), .B(n_835), .C(n_842), .D(n_847), .Y(n_831) );
AND2x2_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
AND2x2_ASAP7_75t_L g835 ( .A(n_836), .B(n_840), .Y(n_835) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
AND2x2_ASAP7_75t_SL g842 ( .A(n_843), .B(n_845), .Y(n_842) );
NAND2xp5_ASAP7_75t_SL g851 ( .A(n_852), .B(n_866), .Y(n_851) );
NOR2xp33_ASAP7_75t_SL g852 ( .A(n_853), .B(n_859), .Y(n_852) );
OAI21xp5_ASAP7_75t_SL g853 ( .A1(n_854), .A2(n_855), .B(n_856), .Y(n_853) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
NAND3xp33_ASAP7_75t_L g859 ( .A(n_860), .B(n_862), .C(n_864), .Y(n_859) );
NOR2x1_ASAP7_75t_L g866 ( .A(n_867), .B(n_873), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_870), .Y(n_867) );
INVx3_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx3_ASAP7_75t_L g972 ( .A(n_872), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_874), .B(n_875), .Y(n_873) );
INVx1_ASAP7_75t_L g978 ( .A(n_879), .Y(n_978) );
AOI22xp5_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_897), .B1(n_975), .B2(n_976), .Y(n_879) );
INVx3_ASAP7_75t_SL g975 ( .A(n_880), .Y(n_975) );
XOR2x2_ASAP7_75t_L g880 ( .A(n_881), .B(n_896), .Y(n_880) );
NAND4xp75_ASAP7_75t_L g881 ( .A(n_882), .B(n_887), .C(n_892), .D(n_895), .Y(n_881) );
AND2x2_ASAP7_75t_L g882 ( .A(n_883), .B(n_885), .Y(n_882) );
OA211x2_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_889), .B(n_890), .C(n_891), .Y(n_887) );
OA211x2_ASAP7_75t_L g1002 ( .A1(n_889), .A2(n_1003), .B(n_1004), .C(n_1006), .Y(n_1002) );
AND2x2_ASAP7_75t_L g892 ( .A(n_893), .B(n_894), .Y(n_892) );
INVx1_ASAP7_75t_L g976 ( .A(n_897), .Y(n_976) );
HB1xp67_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
AOI22xp5_ASAP7_75t_L g898 ( .A1(n_899), .A2(n_900), .B1(n_927), .B2(n_928), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx2_ASAP7_75t_L g926 ( .A(n_901), .Y(n_926) );
AND2x2_ASAP7_75t_SL g901 ( .A(n_902), .B(n_916), .Y(n_901) );
NOR3xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_907), .C(n_911), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_912), .A2(n_913), .B1(n_914), .B2(n_915), .Y(n_911) );
NOR2xp33_ASAP7_75t_L g916 ( .A(n_917), .B(n_921), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_918), .B(n_919), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_922), .B(n_924), .Y(n_921) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
AO22x1_ASAP7_75t_L g928 ( .A1(n_929), .A2(n_930), .B1(n_955), .B2(n_974), .Y(n_928) );
INVx2_ASAP7_75t_SL g929 ( .A(n_930), .Y(n_929) );
XOR2x2_ASAP7_75t_L g930 ( .A(n_931), .B(n_954), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_932), .B(n_945), .Y(n_931) );
NOR3xp33_ASAP7_75t_L g932 ( .A(n_933), .B(n_938), .C(n_942), .Y(n_932) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_934), .A2(n_935), .B1(n_936), .B2(n_937), .Y(n_933) );
OAI21xp33_ASAP7_75t_L g938 ( .A1(n_939), .A2(n_940), .B(n_941), .Y(n_938) );
OAI21xp5_ASAP7_75t_SL g958 ( .A1(n_940), .A2(n_959), .B(n_960), .Y(n_958) );
NOR2xp33_ASAP7_75t_L g945 ( .A(n_946), .B(n_949), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_947), .B(n_948), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_950), .B(n_952), .Y(n_949) );
INVx1_ASAP7_75t_L g1017 ( .A(n_951), .Y(n_1017) );
INVx3_ASAP7_75t_SL g974 ( .A(n_955), .Y(n_974) );
XOR2x2_ASAP7_75t_L g955 ( .A(n_956), .B(n_973), .Y(n_955) );
NAND2xp5_ASAP7_75t_SL g956 ( .A(n_957), .B(n_965), .Y(n_956) );
NOR2xp33_ASAP7_75t_L g957 ( .A(n_958), .B(n_961), .Y(n_957) );
NAND3xp33_ASAP7_75t_L g961 ( .A(n_962), .B(n_963), .C(n_964), .Y(n_961) );
NOR2xp33_ASAP7_75t_L g965 ( .A(n_966), .B(n_969), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_967), .B(n_968), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_970), .B(n_971), .Y(n_969) );
INVx2_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
NOR2x1_ASAP7_75t_L g982 ( .A(n_983), .B(n_987), .Y(n_982) );
OR2x2_ASAP7_75t_SL g1043 ( .A(n_983), .B(n_988), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_984), .B(n_986), .Y(n_983) );
CKINVDCx20_ASAP7_75t_R g1021 ( .A(n_984), .Y(n_1021) );
INVx1_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_985), .B(n_1023), .Y(n_1026) );
CKINVDCx16_ASAP7_75t_R g1023 ( .A(n_986), .Y(n_1023) );
CKINVDCx20_ASAP7_75t_R g987 ( .A(n_988), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_989), .B(n_990), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_992), .B(n_993), .Y(n_991) );
OAI322xp33_ASAP7_75t_L g994 ( .A1(n_995), .A2(n_1020), .A3(n_1022), .B1(n_1024), .B2(n_1027), .C1(n_1028), .C2(n_1041), .Y(n_994) );
INVx1_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
NAND4xp75_ASAP7_75t_L g997 ( .A(n_998), .B(n_1002), .C(n_1007), .D(n_1018), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_999), .B(n_1001), .Y(n_998) );
NOR2xp33_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1012), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_1013), .A2(n_1014), .B1(n_1016), .B2(n_1017), .Y(n_1012) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
HB1xp67_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
CKINVDCx16_ASAP7_75t_R g1024 ( .A(n_1025), .Y(n_1024) );
XOR2x2_ASAP7_75t_L g1028 ( .A(n_1027), .B(n_1029), .Y(n_1028) );
NAND4xp75_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1033), .C(n_1036), .D(n_1040), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1032), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1035), .Y(n_1033) );
CKINVDCx20_ASAP7_75t_R g1041 ( .A(n_1042), .Y(n_1041) );
CKINVDCx20_ASAP7_75t_R g1042 ( .A(n_1043), .Y(n_1042) );
endmodule