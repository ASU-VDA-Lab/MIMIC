module real_jpeg_3030_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_70;
wire n_74;
wire n_41;
wire n_32;
wire n_20;
wire n_228;
wire n_80;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_244;
wire n_179;
wire n_213;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_1),
.A2(n_74),
.B1(n_75),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_1),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_1),
.A2(n_59),
.B1(n_61),
.B2(n_85),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_1),
.A2(n_43),
.B1(n_44),
.B2(n_85),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_1),
.A2(n_28),
.B1(n_35),
.B2(n_85),
.Y(n_180)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_3),
.A2(n_74),
.B1(n_75),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_3),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_3),
.A2(n_59),
.B1(n_61),
.B2(n_83),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_83),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_3),
.A2(n_28),
.B1(n_35),
.B2(n_83),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_4),
.A2(n_28),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_4),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_5),
.B(n_74),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_5),
.B(n_129),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_5),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_5),
.A2(n_74),
.B(n_140),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_5),
.B(n_63),
.Y(n_202)
);

AOI21xp33_ASAP7_75t_L g209 ( 
.A1(n_5),
.A2(n_61),
.B(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_5),
.B(n_28),
.C(n_49),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_176),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_5),
.B(n_31),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_5),
.B(n_54),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_6),
.A2(n_28),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_6),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_94)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_8),
.Y(n_76)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_10),
.A2(n_58),
.B1(n_74),
.B2(n_75),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_58),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g167 ( 
.A1(n_10),
.A2(n_28),
.B1(n_35),
.B2(n_58),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_11),
.A2(n_53),
.B1(n_59),
.B2(n_61),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_11),
.A2(n_28),
.B1(n_35),
.B2(n_53),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_13),
.A2(n_74),
.B1(n_75),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_13),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_13),
.A2(n_59),
.B1(n_61),
.B2(n_150),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_150),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_13),
.A2(n_28),
.B1(n_35),
.B2(n_150),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_14),
.A2(n_74),
.B1(n_75),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_14),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_14),
.A2(n_59),
.B1(n_61),
.B2(n_128),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_128),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_14),
.A2(n_28),
.B1(n_35),
.B2(n_128),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_16),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_16),
.A2(n_46),
.B1(n_59),
.B2(n_61),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_16),
.A2(n_28),
.B1(n_35),
.B2(n_46),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_132),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_130),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_112),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_21),
.B(n_112),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_86),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_55),
.C(n_70),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_23),
.A2(n_24),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_25),
.A2(n_26),
.B1(n_39),
.B2(n_40),
.Y(n_152)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_31),
.B1(n_33),
.B2(n_37),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_27),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_27),
.A2(n_31),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_27),
.A2(n_31),
.B1(n_143),
.B2(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_27),
.A2(n_31),
.B1(n_180),
.B2(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_27),
.A2(n_31),
.B1(n_176),
.B2(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_27),
.A2(n_31),
.B1(n_230),
.B2(n_234),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_28),
.A2(n_35),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_28),
.B(n_228),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_30),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_30),
.A2(n_34),
.B1(n_100),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_30),
.A2(n_100),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_30),
.A2(n_100),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B1(n_52),
.B2(n_54),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_42),
.A2(n_51),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

AO22x2_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_44),
.B1(n_64),
.B2(n_66),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_43),
.B(n_66),
.Y(n_177)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_44),
.A2(n_61),
.A3(n_64),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_44),
.B(n_218),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_47),
.A2(n_54),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_47),
.A2(n_52),
.B1(n_54),
.B2(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_47),
.A2(n_54),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_47),
.A2(n_54),
.B1(n_172),
.B2(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_47),
.A2(n_54),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_47),
.A2(n_54),
.B1(n_200),
.B2(n_221),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_51),
.A2(n_121),
.B1(n_171),
.B2(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_55),
.B(n_70),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_62),
.B1(n_68),
.B2(n_69),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_57),
.A2(n_63),
.B1(n_90),
.B2(n_125),
.Y(n_124)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_61),
.B1(n_64),
.B2(n_66),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_61),
.B1(n_77),
.B2(n_78),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g141 ( 
.A(n_59),
.B(n_77),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_59),
.B(n_176),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI32xp33_ASAP7_75t_L g139 ( 
.A1(n_61),
.A2(n_75),
.A3(n_78),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_62),
.A2(n_69),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_62),
.A2(n_69),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_62),
.A2(n_69),
.B1(n_146),
.B2(n_162),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_62),
.A2(n_69),
.B1(n_161),
.B2(n_209),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_88)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_80),
.B1(n_81),
.B2(n_84),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_80),
.B1(n_84),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_71),
.A2(n_80),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_71),
.A2(n_80),
.B1(n_149),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_72),
.A2(n_82),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_80),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_78),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_96),
.B1(n_97),
.B2(n_111),
.Y(n_86)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_92),
.B(n_95),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_92),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_104),
.B1(n_105),
.B2(n_110),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_106),
.Y(n_116)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.C(n_117),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_116),
.Y(n_154)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_114),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_124),
.C(n_126),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_119),
.B(n_122),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_126),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_125),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_155),
.B(n_266),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_153),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_134),
.B(n_153),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.C(n_152),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_135),
.B(n_152),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_137),
.B(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_145),
.C(n_148),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_138),
.B(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_142),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_145),
.B(n_148),
.Y(n_256)
);

AOI31xp33_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_250),
.A3(n_259),
.B(n_263),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_195),
.B(n_249),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_182),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_158),
.B(n_182),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_169),
.C(n_173),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_159),
.B(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_164),
.C(n_168),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_168),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_169),
.B(n_173),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_184),
.B(n_185),
.C(n_186),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_187),
.B(n_190),
.C(n_194),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_244),
.B(n_248),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_213),
.B(n_243),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_205),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_205),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.C(n_203),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_202),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_206),
.B(n_208),
.C(n_211),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_224),
.B(n_242),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_222),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_222),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_236),
.B(n_241),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_231),
.B(n_235),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_233),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_234),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_240),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_240),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_247),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_264),
.B(n_265),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_254),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.C(n_258),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_258),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_261),
.Y(n_264)
);


endmodule