module real_aes_15023_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_139;
wire n_552;
wire n_402;
wire n_733;
wire n_602;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_679;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
OA21x2_ASAP7_75t_L g92 ( .A1(n_0), .A2(n_44), .B(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g209 ( .A(n_0), .Y(n_209) );
INVxp67_ASAP7_75t_SL g576 ( .A(n_1), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_1), .A2(n_31), .B1(n_612), .B2(n_617), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_2), .A2(n_683), .B1(n_684), .B2(n_685), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_2), .Y(n_685) );
AND2x2_ASAP7_75t_L g128 ( .A(n_3), .B(n_114), .Y(n_128) );
AOI221xp5_ASAP7_75t_L g255 ( .A1(n_4), .A2(n_72), .B1(n_152), .B2(n_182), .C(n_205), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_4), .A2(n_695), .B1(n_696), .B2(n_697), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_4), .Y(n_697) );
BUFx3_ASAP7_75t_L g503 ( .A(n_5), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_6), .B(n_91), .Y(n_121) );
INVx3_ASAP7_75t_L g549 ( .A(n_7), .Y(n_549) );
INVx2_ASAP7_75t_L g508 ( .A(n_8), .Y(n_508) );
INVx1_ASAP7_75t_L g525 ( .A(n_8), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_9), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g96 ( .A(n_10), .B(n_97), .Y(n_96) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_11), .Y(n_696) );
BUFx3_ASAP7_75t_L g102 ( .A(n_12), .Y(n_102) );
INVx1_ASAP7_75t_L g108 ( .A(n_12), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_13), .B(n_136), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_14), .Y(n_194) );
BUFx10_ASAP7_75t_L g709 ( .A(n_15), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g551 ( .A1(n_16), .A2(n_53), .B1(n_552), .B2(n_555), .C(n_557), .Y(n_551) );
INVx1_ASAP7_75t_L g610 ( .A(n_16), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_17), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_18), .B(n_187), .Y(n_191) );
OAI21xp33_ASAP7_75t_L g288 ( .A1(n_18), .A2(n_55), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g585 ( .A(n_19), .Y(n_585) );
OAI222xp33_ASAP7_75t_L g639 ( .A1(n_19), .A2(n_47), .B1(n_53), .B2(n_640), .C1(n_643), .C2(n_646), .Y(n_639) );
O2A1O1Ixp5_ASAP7_75t_L g256 ( .A1(n_20), .A2(n_116), .B(n_162), .C(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g560 ( .A(n_21), .Y(n_560) );
INVxp33_ASAP7_75t_L g595 ( .A(n_22), .Y(n_595) );
INVx1_ASAP7_75t_L g623 ( .A(n_22), .Y(n_623) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_22), .Y(n_667) );
INVx1_ASAP7_75t_L g120 ( .A(n_23), .Y(n_120) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_24), .Y(n_688) );
INVx2_ASAP7_75t_L g603 ( .A(n_25), .Y(n_603) );
OAI222xp33_ASAP7_75t_L g520 ( .A1(n_26), .A2(n_35), .B1(n_70), .B2(n_521), .C1(n_526), .C2(n_530), .Y(n_520) );
INVxp67_ASAP7_75t_SL g659 ( .A(n_26), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_27), .B(n_112), .Y(n_197) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_28), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_29), .A2(n_60), .B1(n_535), .B2(n_538), .Y(n_534) );
INVx1_ASAP7_75t_L g629 ( .A(n_29), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_30), .B(n_149), .Y(n_148) );
AOI221xp5_ASAP7_75t_L g568 ( .A1(n_31), .A2(n_47), .B1(n_569), .B2(n_572), .C(n_575), .Y(n_568) );
INVx2_ASAP7_75t_L g594 ( .A(n_32), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_32), .B(n_623), .Y(n_622) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_32), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_33), .B(n_136), .Y(n_247) );
OAI221xp5_ASAP7_75t_L g497 ( .A1(n_34), .A2(n_76), .B1(n_498), .B2(n_509), .C(n_516), .Y(n_497) );
OAI211xp5_ASAP7_75t_L g650 ( .A1(n_34), .A2(n_651), .B(n_652), .C(n_662), .Y(n_650) );
INVxp67_ASAP7_75t_SL g656 ( .A(n_35), .Y(n_656) );
AND2x4_ASAP7_75t_L g119 ( .A(n_36), .B(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_36), .Y(n_678) );
NAND2x1_ASAP7_75t_L g113 ( .A(n_37), .B(n_114), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_38), .Y(n_201) );
INVx1_ASAP7_75t_L g105 ( .A(n_39), .Y(n_105) );
INVx1_ASAP7_75t_L g507 ( .A(n_40), .Y(n_507) );
INVx1_ASAP7_75t_L g514 ( .A(n_40), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_41), .Y(n_219) );
AND2x2_ASAP7_75t_L g126 ( .A(n_42), .B(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_43), .B(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g210 ( .A(n_44), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_45), .B(n_91), .Y(n_229) );
INVx1_ASAP7_75t_L g93 ( .A(n_46), .Y(n_93) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_48), .B(n_127), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_49), .B(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_50), .B(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_51), .B(n_175), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_52), .B(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g132 ( .A(n_54), .B(n_91), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_55), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_56), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_57), .B(n_159), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_58), .B(n_175), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_59), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_60), .A2(n_76), .B1(n_633), .B2(n_635), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_61), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_62), .B(n_187), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_63), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_64), .B(n_127), .Y(n_246) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_64), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_65), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_66), .B(n_151), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_67), .B(n_177), .Y(n_176) );
BUFx3_ASAP7_75t_L g98 ( .A(n_68), .Y(n_98) );
INVx1_ASAP7_75t_L g117 ( .A(n_68), .Y(n_117) );
INVx1_ASAP7_75t_L g156 ( .A(n_68), .Y(n_156) );
INVx1_ASAP7_75t_L g692 ( .A(n_69), .Y(n_692) );
INVxp67_ASAP7_75t_SL g631 ( .A(n_70), .Y(n_631) );
INVx2_ASAP7_75t_L g604 ( .A(n_71), .Y(n_604) );
INVxp67_ASAP7_75t_SL g615 ( .A(n_71), .Y(n_615) );
AND2x2_ASAP7_75t_L g619 ( .A(n_71), .B(n_603), .Y(n_619) );
INVx1_ASAP7_75t_L g558 ( .A(n_73), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_74), .B(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g546 ( .A(n_75), .Y(n_546) );
AOI22xp33_ASAP7_75t_SL g492 ( .A1(n_77), .A2(n_493), .B1(n_494), .B2(n_495), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_77), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_479), .B(n_491), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_414), .Y(n_80) );
NOR4xp25_ASAP7_75t_L g81 ( .A(n_82), .B(n_302), .C(n_355), .D(n_396), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g82 ( .A(n_83), .B(n_276), .Y(n_82) );
AOI21xp5_ASAP7_75t_L g83 ( .A1(n_84), .A2(n_165), .B(n_230), .Y(n_83) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_84), .A2(n_334), .B1(n_381), .B2(n_383), .Y(n_380) );
AND2x2_ASAP7_75t_L g84 ( .A(n_85), .B(n_122), .Y(n_84) );
HB1xp67_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_86), .B(n_124), .Y(n_409) );
INVx1_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx2_ASAP7_75t_L g274 ( .A(n_87), .Y(n_274) );
AND2x2_ASAP7_75t_L g283 ( .A(n_87), .B(n_275), .Y(n_283) );
AND2x2_ASAP7_75t_L g309 ( .A(n_87), .B(n_236), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_87), .B(n_124), .Y(n_317) );
INVxp67_ASAP7_75t_L g325 ( .A(n_87), .Y(n_325) );
AND2x4_ASAP7_75t_SL g341 ( .A(n_87), .B(n_267), .Y(n_341) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_87), .Y(n_361) );
INVx1_ASAP7_75t_L g377 ( .A(n_87), .Y(n_377) );
BUFx6f_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
OAI21x1_ASAP7_75t_L g88 ( .A1(n_89), .A2(n_94), .B(n_121), .Y(n_88) );
INVx1_ASAP7_75t_SL g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVxp33_ASAP7_75t_L g139 ( .A(n_91), .Y(n_139) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_91), .Y(n_171) );
INVx1_ASAP7_75t_L g262 ( .A(n_91), .Y(n_262) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g145 ( .A(n_92), .Y(n_145) );
BUFx2_ASAP7_75t_L g240 ( .A(n_92), .Y(n_240) );
INVx1_ASAP7_75t_L g211 ( .A(n_93), .Y(n_211) );
OAI21x1_ASAP7_75t_L g94 ( .A1(n_95), .A2(n_109), .B(n_118), .Y(n_94) );
OAI21xp5_ASAP7_75t_L g95 ( .A1(n_96), .A2(n_99), .B(n_103), .Y(n_95) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_98), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g198 ( .A(n_98), .Y(n_198) );
INVx2_ASAP7_75t_L g248 ( .A(n_98), .Y(n_248) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx3_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx3_ASAP7_75t_L g114 ( .A(n_101), .Y(n_114) );
INVx2_ASAP7_75t_L g136 ( .A(n_101), .Y(n_136) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g112 ( .A(n_102), .Y(n_112) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_102), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
INVx1_ASAP7_75t_L g490 ( .A(n_106), .Y(n_490) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g127 ( .A(n_107), .Y(n_127) );
INVx2_ASAP7_75t_L g162 ( .A(n_107), .Y(n_162) );
INVx2_ASAP7_75t_L g200 ( .A(n_107), .Y(n_200) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g153 ( .A(n_108), .Y(n_153) );
AOI21x1_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_113), .B(n_115), .Y(n_109) );
INVx1_ASAP7_75t_L g177 ( .A(n_111), .Y(n_177) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g149 ( .A(n_112), .Y(n_149) );
INVx2_ASAP7_75t_L g175 ( .A(n_112), .Y(n_175) );
INVx2_ASAP7_75t_L g196 ( .A(n_112), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_115), .A2(n_158), .B(n_161), .Y(n_157) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g178 ( .A(n_116), .Y(n_178) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx3_ASAP7_75t_L g130 ( .A(n_117), .Y(n_130) );
INVx1_ASAP7_75t_L g164 ( .A(n_118), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_118), .A2(n_242), .B(n_245), .Y(n_241) );
BUFx6f_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx3_ASAP7_75t_L g141 ( .A(n_119), .Y(n_141) );
INVx2_ASAP7_75t_L g185 ( .A(n_119), .Y(n_185) );
INVx1_ASAP7_75t_L g207 ( .A(n_119), .Y(n_207) );
INVx1_ASAP7_75t_L g486 ( .A(n_119), .Y(n_486) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_120), .Y(n_676) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g279 ( .A(n_123), .Y(n_279) );
INVxp67_ASAP7_75t_L g391 ( .A(n_123), .Y(n_391) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_142), .Y(n_123) );
INVx2_ASAP7_75t_L g267 ( .A(n_124), .Y(n_267) );
AND2x2_ASAP7_75t_L g362 ( .A(n_124), .B(n_301), .Y(n_362) );
INVx1_ASAP7_75t_L g370 ( .A(n_124), .Y(n_370) );
AO21x2_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_131), .B(n_138), .Y(n_124) );
OAI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_128), .B(n_129), .Y(n_125) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g137 ( .A(n_130), .Y(n_137) );
NOR2xp67_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AOI21xp33_ASAP7_75t_L g138 ( .A1(n_132), .A2(n_139), .B(n_140), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_135), .B(n_137), .Y(n_133) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NOR3xp33_ASAP7_75t_L g254 ( .A(n_141), .B(n_255), .C(n_256), .Y(n_254) );
AND2x2_ASAP7_75t_L g266 ( .A(n_142), .B(n_267), .Y(n_266) );
INVx3_ASAP7_75t_L g301 ( .A(n_142), .Y(n_301) );
INVx1_ASAP7_75t_L g308 ( .A(n_142), .Y(n_308) );
AND2x2_ASAP7_75t_L g324 ( .A(n_142), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g330 ( .A(n_142), .Y(n_330) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_142), .Y(n_358) );
AND2x2_ASAP7_75t_L g417 ( .A(n_142), .B(n_333), .Y(n_417) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_146), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_144), .B(n_164), .Y(n_163) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_144), .Y(n_187) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OAI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_157), .B(n_163), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_150), .B(n_154), .Y(n_147) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_154), .A2(n_180), .B(n_183), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_154), .A2(n_223), .B(n_226), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_154), .A2(n_243), .B(n_244), .Y(n_242) );
BUFx10_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx3_ASAP7_75t_L g205 ( .A(n_156), .Y(n_205) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g202 ( .A(n_160), .Y(n_202) );
INVx1_ASAP7_75t_L g216 ( .A(n_160), .Y(n_216) );
INVx2_ASAP7_75t_L g225 ( .A(n_160), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_160), .B(n_258), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_165), .A2(n_388), .B1(n_422), .B2(n_424), .Y(n_421) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_188), .Y(n_165) );
OR2x2_ASAP7_75t_L g285 ( .A(n_166), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g420 ( .A(n_166), .B(n_379), .Y(n_420) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g306 ( .A(n_168), .B(n_271), .Y(n_306) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g343 ( .A(n_169), .B(n_253), .Y(n_343) );
OAI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_172), .B(n_186), .Y(n_169) );
OAI21x1_ASAP7_75t_L g212 ( .A1(n_170), .A2(n_213), .B(n_229), .Y(n_212) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_170), .A2(n_172), .B(n_186), .Y(n_264) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_170), .A2(n_213), .B(n_229), .Y(n_294) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OAI21x1_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_179), .B(n_184), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_176), .B(n_178), .Y(n_173) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_SL g228 ( .A(n_185), .Y(n_228) );
AND2x4_ASAP7_75t_SL g268 ( .A(n_188), .B(n_269), .Y(n_268) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_188), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g450 ( .A(n_188), .B(n_252), .Y(n_450) );
AND2x4_ASAP7_75t_L g188 ( .A(n_189), .B(n_212), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g233 ( .A(n_190), .Y(n_233) );
AND2x2_ASAP7_75t_L g336 ( .A(n_190), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g354 ( .A(n_190), .Y(n_354) );
AND2x2_ASAP7_75t_L g379 ( .A(n_190), .B(n_212), .Y(n_379) );
AND2x4_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
NAND3xp33_ASAP7_75t_L g287 ( .A(n_192), .B(n_288), .C(n_290), .Y(n_287) );
NAND3xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_199), .C(n_206), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_197), .C(n_198), .Y(n_193) );
INVx2_ASAP7_75t_SL g195 ( .A(n_196), .Y(n_195) );
OAI221xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B1(n_202), .B2(n_203), .C(n_204), .Y(n_199) );
INVx2_ASAP7_75t_L g227 ( .A(n_200), .Y(n_227) );
INVx1_ASAP7_75t_L g733 ( .A(n_201), .Y(n_733) );
INVx1_ASAP7_75t_L g722 ( .A(n_203), .Y(n_722) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_205), .A2(n_215), .B1(n_217), .B2(n_221), .Y(n_214) );
INVx2_ASAP7_75t_SL g220 ( .A(n_205), .Y(n_220) );
INVx1_ASAP7_75t_L g488 ( .A(n_205), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
INVx2_ASAP7_75t_L g292 ( .A(n_208), .Y(n_292) );
AOI21x1_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_211), .Y(n_208) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_209), .A2(n_210), .B(n_211), .Y(n_259) );
INVx1_ASAP7_75t_L g234 ( .A(n_212), .Y(n_234) );
OAI21x1_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_222), .B(n_228), .Y(n_213) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_220), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AO32x1_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_250), .A3(n_265), .B1(n_268), .B2(n_272), .Y(n_230) );
AOI32xp33_ASAP7_75t_L g443 ( .A1(n_231), .A2(n_383), .A3(n_444), .B1(n_445), .B2(n_446), .Y(n_443) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_235), .Y(n_231) );
AND2x2_ASAP7_75t_L g305 ( .A(n_232), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g311 ( .A(n_232), .B(n_252), .Y(n_311) );
AND2x2_ASAP7_75t_L g363 ( .A(n_232), .B(n_343), .Y(n_363) );
AND2x4_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
INVx1_ASAP7_75t_L g298 ( .A(n_233), .Y(n_298) );
INVx1_ASAP7_75t_L g352 ( .A(n_235), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_235), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g411 ( .A(n_235), .B(n_341), .Y(n_411) );
AND2x2_ASAP7_75t_L g472 ( .A(n_235), .B(n_362), .Y(n_472) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g278 ( .A(n_236), .B(n_274), .Y(n_278) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
BUFx3_ASAP7_75t_L g275 ( .A(n_237), .Y(n_275) );
OAI21x1_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_241), .B(n_249), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
BUFx3_ASAP7_75t_L g289 ( .A(n_240), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_247), .B(n_248), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_250), .B(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_251), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_252), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g465 ( .A(n_252), .B(n_395), .Y(n_465) );
AND2x2_ASAP7_75t_L g469 ( .A(n_252), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_263), .Y(n_252) );
INVx2_ASAP7_75t_L g271 ( .A(n_253), .Y(n_271) );
INVx1_ASAP7_75t_L g445 ( .A(n_253), .Y(n_445) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_259), .B(n_260), .Y(n_253) );
NAND2xp33_ASAP7_75t_L g290 ( .A(n_254), .B(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_R g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx2_ASAP7_75t_L g270 ( .A(n_263), .Y(n_270) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVxp67_ASAP7_75t_L g349 ( .A(n_264), .Y(n_349) );
NAND2x1p5_ASAP7_75t_L g430 ( .A(n_265), .B(n_431), .Y(n_430) );
BUFx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_266), .B(n_367), .Y(n_434) );
AND2x2_ASAP7_75t_L g467 ( .A(n_266), .B(n_352), .Y(n_467) );
BUFx2_ASAP7_75t_L g322 ( .A(n_267), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_268), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_269), .B(n_394), .Y(n_393) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx2_ASAP7_75t_L g427 ( .A(n_270), .Y(n_427) );
AND2x2_ASAP7_75t_L g353 ( .A(n_271), .B(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g478 ( .A(n_273), .B(n_329), .Y(n_478) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx3_ASAP7_75t_L g333 ( .A(n_275), .Y(n_333) );
AND2x2_ASAP7_75t_L g388 ( .A(n_275), .B(n_370), .Y(n_388) );
OAI211xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_280), .B(n_284), .C(n_299), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND2x2_ASAP7_75t_L g419 ( .A(n_278), .B(n_322), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_278), .B(n_368), .Y(n_448) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
BUFx2_ASAP7_75t_L g295 ( .A(n_282), .Y(n_295) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_283), .B(n_358), .Y(n_441) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_283), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_295), .B(n_296), .Y(n_284) );
INVx1_ASAP7_75t_L g418 ( .A(n_285), .Y(n_418) );
INVx1_ASAP7_75t_L g477 ( .A(n_286), .Y(n_477) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_293), .Y(n_286) );
OR2x2_ASAP7_75t_L g313 ( .A(n_287), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g350 ( .A(n_287), .Y(n_350) );
INVx1_ASAP7_75t_L g385 ( .A(n_287), .Y(n_385) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g314 ( .A(n_293), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_293), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g439 ( .A(n_293), .Y(n_439) );
BUFx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g337 ( .A(n_294), .Y(n_337) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g342 ( .A(n_298), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g407 ( .A(n_300), .B(n_408), .Y(n_407) );
OAI21xp5_ASAP7_75t_SL g449 ( .A1(n_300), .A2(n_450), .B(n_451), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g451 ( .A1(n_300), .A2(n_452), .B(n_455), .C(n_457), .Y(n_451) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g369 ( .A(n_301), .B(n_370), .Y(n_369) );
NAND4xp25_ASAP7_75t_L g302 ( .A(n_303), .B(n_318), .C(n_326), .D(n_344), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_310), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_305), .A2(n_387), .B1(n_389), .B2(n_392), .Y(n_386) );
AND2x4_ASAP7_75t_L g403 ( .A(n_306), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
AND2x2_ASAP7_75t_L g315 ( .A(n_308), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g457 ( .A(n_308), .B(n_458), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B(n_315), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x4_ASAP7_75t_L g444 ( .A(n_316), .B(n_329), .Y(n_444) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g399 ( .A(n_317), .Y(n_399) );
INVxp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
AOI32xp33_ASAP7_75t_L g344 ( .A1(n_321), .A2(n_345), .A3(n_348), .B1(n_351), .B2(n_353), .Y(n_344) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g461 ( .A(n_324), .B(n_333), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_334), .B1(n_338), .B2(n_342), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_331), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g339 ( .A(n_329), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g376 ( .A(n_330), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g347 ( .A(n_333), .Y(n_347) );
INVx1_ASAP7_75t_L g367 ( .A(n_333), .Y(n_367) );
AND2x2_ASAP7_75t_L g398 ( .A(n_333), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g410 ( .A(n_333), .Y(n_410) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_334), .A2(n_392), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g413 ( .A(n_336), .Y(n_413) );
BUFx3_ASAP7_75t_L g404 ( .A(n_337), .Y(n_404) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g382 ( .A(n_340), .Y(n_382) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g351 ( .A(n_341), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g357 ( .A(n_341), .B(n_358), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_342), .A2(n_444), .B(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g378 ( .A(n_343), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g436 ( .A(n_343), .Y(n_436) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g373 ( .A(n_347), .Y(n_373) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx2_ASAP7_75t_L g384 ( .A(n_349), .Y(n_384) );
INVx2_ASAP7_75t_L g395 ( .A(n_354), .Y(n_395) );
NAND4xp25_ASAP7_75t_L g355 ( .A(n_356), .B(n_364), .C(n_380), .D(n_386), .Y(n_355) );
OAI21xp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_359), .B(n_363), .Y(n_356) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_362), .Y(n_359) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_362), .B(n_373), .Y(n_372) );
OAI31xp33_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_371), .A3(n_374), .B(n_378), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
NOR2xp67_ASAP7_75t_L g423 ( .A(n_367), .B(n_369), .Y(n_423) );
INVx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g387 ( .A(n_377), .B(n_388), .Y(n_387) );
BUFx2_ASAP7_75t_L g431 ( .A(n_377), .Y(n_431) );
INVx1_ASAP7_75t_L g458 ( .A(n_377), .Y(n_458) );
AND2x2_ASAP7_75t_L g453 ( .A(n_379), .B(n_454), .Y(n_453) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
AOI32xp33_ASAP7_75t_L g432 ( .A1(n_384), .A2(n_412), .A3(n_433), .B1(n_435), .B2(n_440), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_384), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g475 ( .A(n_384), .Y(n_475) );
INVx2_ASAP7_75t_L g447 ( .A(n_387), .Y(n_447) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_395), .Y(n_402) );
OAI21xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_400), .B(n_405), .Y(n_396) );
INVxp67_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
OAI21xp33_ASAP7_75t_SL g428 ( .A1(n_403), .A2(n_424), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g464 ( .A(n_404), .Y(n_464) );
INVx2_ASAP7_75t_L g470 ( .A(n_404), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_411), .B(n_412), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NOR3xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_442), .C(n_459), .Y(n_414) );
NAND4xp25_ASAP7_75t_SL g415 ( .A(n_416), .B(n_421), .C(n_428), .D(n_432), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_419), .B2(n_420), .Y(n_416) );
BUFx2_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2xp33_ASAP7_75t_SL g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g476 ( .A(n_439), .Y(n_476) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_449), .Y(n_442) );
INVx1_ASAP7_75t_L g454 ( .A(n_445), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND4xp25_ASAP7_75t_L g459 ( .A(n_460), .B(n_466), .C(n_468), .D(n_471), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2x1p5_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B1(n_477), .B2(n_478), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
CKINVDCx6p67_ASAP7_75t_R g479 ( .A(n_480), .Y(n_479) );
CKINVDCx11_ASAP7_75t_R g480 ( .A(n_481), .Y(n_480) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_487), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AO21x2_ASAP7_75t_L g736 ( .A1(n_487), .A2(n_675), .B(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OAI221xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_494), .B1(n_669), .B2(n_679), .C(n_729), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_494), .A2(n_730), .B1(n_733), .B2(n_734), .Y(n_729) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_550), .C(n_638), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_534), .B(n_540), .Y(n_496) );
INVx2_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_504), .Y(n_499) );
AND2x6_ASAP7_75t_L g510 ( .A(n_500), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x4_ASAP7_75t_L g517 ( .A(n_501), .B(n_518), .Y(n_517) );
OR2x2_ASAP7_75t_L g535 ( .A(n_501), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g588 ( .A(n_502), .B(n_545), .Y(n_588) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx2_ASAP7_75t_L g523 ( .A(n_503), .Y(n_523) );
AND2x4_ASAP7_75t_L g567 ( .A(n_503), .B(n_545), .Y(n_567) );
OR2x2_ASAP7_75t_L g711 ( .A(n_503), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g721 ( .A(n_503), .B(n_712), .Y(n_721) );
INVx2_ASAP7_75t_SL g556 ( .A(n_504), .Y(n_556) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
AND2x4_ASAP7_75t_L g519 ( .A(n_506), .B(n_515), .Y(n_519) );
INVx1_ASAP7_75t_L g533 ( .A(n_506), .Y(n_533) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g574 ( .A(n_507), .B(n_508), .Y(n_574) );
INVx2_ASAP7_75t_L g515 ( .A(n_508), .Y(n_515) );
CKINVDCx14_ASAP7_75t_R g509 ( .A(n_510), .Y(n_509) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx4_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx12f_ASAP7_75t_L g554 ( .A(n_513), .Y(n_554) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_513), .Y(n_571) );
AND2x4_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
AND2x4_ASAP7_75t_L g537 ( .A(n_514), .B(n_525), .Y(n_537) );
INVx1_ASAP7_75t_L g581 ( .A(n_514), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_517), .B(n_520), .Y(n_516) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_518), .Y(n_584) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_519), .Y(n_529) );
INVx2_ASAP7_75t_L g564 ( .A(n_519), .Y(n_564) );
CKINVDCx14_ASAP7_75t_R g521 ( .A(n_522), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
AND2x4_ASAP7_75t_L g531 ( .A(n_523), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g539 ( .A(n_523), .Y(n_539) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_524), .B(n_708), .C(n_710), .Y(n_707) );
AND2x4_ASAP7_75t_L g718 ( .A(n_524), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g580 ( .A(n_525), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx5_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
CKINVDCx8_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
INVx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OR2x2_ASAP7_75t_L g538 ( .A(n_536), .B(n_539), .Y(n_538) );
BUFx2_ASAP7_75t_L g559 ( .A(n_536), .Y(n_559) );
INVx8_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_543), .B(n_547), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g712 ( .A(n_546), .Y(n_712) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g668 ( .A(n_548), .Y(n_668) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g566 ( .A(n_549), .Y(n_566) );
INVx2_ASAP7_75t_L g587 ( .A(n_549), .Y(n_587) );
AND3x2_ASAP7_75t_SL g591 ( .A(n_549), .B(n_592), .C(n_595), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_565), .B1(n_568), .B2(n_586), .C(n_589), .Y(n_550) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B1(n_560), .B2(n_561), .Y(n_557) );
OAI221xp5_ASAP7_75t_L g596 ( .A1(n_558), .A2(n_597), .B1(n_605), .B2(n_610), .C(n_611), .Y(n_596) );
AOI222xp33_ASAP7_75t_L g652 ( .A1(n_560), .A2(n_653), .B1(n_656), .B2(n_657), .C1(n_659), .C2(n_660), .Y(n_652) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx4_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x6_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
BUFx4f_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B1(n_582), .B2(n_585), .Y(n_575) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x6_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
OR2x6_ASAP7_75t_L g621 ( .A(n_587), .B(n_622), .Y(n_621) );
OAI22xp5_ASAP7_75t_SL g589 ( .A1(n_590), .A2(n_596), .B1(n_620), .B2(n_624), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g645 ( .A(n_593), .Y(n_645) );
AND2x4_ASAP7_75t_L g657 ( .A(n_593), .B(n_658), .Y(n_657) );
AND2x4_ASAP7_75t_SL g660 ( .A(n_593), .B(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx4_ASAP7_75t_L g649 ( .A(n_600), .Y(n_649) );
INVx5_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g637 ( .A(n_601), .Y(n_637) );
AND2x4_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx1_ASAP7_75t_L g616 ( .A(n_602), .Y(n_616) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_602), .Y(n_658) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g609 ( .A(n_603), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_603), .B(n_604), .Y(n_628) );
INVx2_ASAP7_75t_L g608 ( .A(n_604), .Y(n_608) );
BUFx4f_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
BUFx3_ASAP7_75t_L g630 ( .A(n_606), .Y(n_630) );
BUFx12f_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2x1p5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
AND2x4_ASAP7_75t_L g655 ( .A(n_608), .B(n_609), .Y(n_655) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx5_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g661 ( .A(n_615), .Y(n_661) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g644 ( .A(n_618), .B(n_645), .Y(n_644) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
BUFx4f_ASAP7_75t_L g634 ( .A(n_619), .Y(n_634) );
BUFx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OAI221xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_629), .B1(n_630), .B2(n_631), .C(n_632), .Y(n_624) );
INVx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx3_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_SL g640 ( .A(n_627), .B(n_641), .Y(n_640) );
OR2x6_ASAP7_75t_L g651 ( .A(n_627), .B(n_645), .Y(n_651) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
BUFx3_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_650), .B(n_664), .Y(n_638) );
INVx3_ASAP7_75t_R g648 ( .A(n_641), .Y(n_648) );
AND2x4_ASAP7_75t_L g663 ( .A(n_641), .B(n_655), .Y(n_663) );
BUFx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
CKINVDCx5p33_ASAP7_75t_R g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x4_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
CKINVDCx8_ASAP7_75t_R g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_670), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_671), .Y(n_670) );
BUFx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
BUFx6f_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_677), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
BUFx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g705 ( .A(n_676), .Y(n_705) );
AND2x2_ASAP7_75t_L g737 ( .A(n_677), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_678), .B(n_705), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_699), .B1(n_722), .B2(n_723), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_680), .A2(n_722), .B1(n_731), .B2(n_732), .Y(n_730) );
XNOR2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_691), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_686), .B1(n_687), .B2(n_690), .Y(n_681) );
INVx1_ASAP7_75t_L g690 ( .A(n_682), .Y(n_690) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
XOR2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B1(n_694), .B2(n_698), .Y(n_691) );
INVx1_ASAP7_75t_L g698 ( .A(n_692), .Y(n_698) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx3_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
BUFx3_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx5_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx3_ASAP7_75t_L g731 ( .A(n_702), .Y(n_731) );
AND2x6_ASAP7_75t_L g702 ( .A(n_703), .B(n_713), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_706), .Y(n_703) );
INVxp67_ASAP7_75t_L g727 ( .A(n_704), .Y(n_727) );
INVx1_ASAP7_75t_L g738 ( .A(n_705), .Y(n_738) );
INVxp67_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_707), .B(n_717), .Y(n_728) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
CKINVDCx11_ASAP7_75t_R g715 ( .A(n_709), .Y(n_715) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_716), .Y(n_713) );
CKINVDCx5p33_ASAP7_75t_R g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
BUFx6f_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
BUFx6f_ASAP7_75t_L g732 ( .A(n_725), .Y(n_732) );
INVx4_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_735), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_736), .Y(n_735) );
endmodule