module real_jpeg_21302_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_0),
.A2(n_66),
.B1(n_67),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_0),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_0),
.A2(n_41),
.B1(n_48),
.B2(n_115),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_115),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_115),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_2),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_2),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_2),
.A2(n_41),
.B1(n_48),
.B2(n_68),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_68),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_68),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_3),
.A2(n_66),
.B1(n_67),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_3),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_3),
.A2(n_41),
.B1(n_48),
.B2(n_74),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_74),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_74),
.Y(n_162)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_4),
.A2(n_41),
.B1(n_48),
.B2(n_70),
.Y(n_72)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_6),
.A2(n_66),
.B1(n_67),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_6),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_6),
.A2(n_41),
.B1(n_48),
.B2(n_93),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_93),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_93),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_7),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_7),
.B(n_72),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_L g179 ( 
.A1(n_7),
.A2(n_16),
.B(n_33),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_133),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_7),
.A2(n_55),
.B1(n_57),
.B2(n_188),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_7),
.B(n_88),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g217 ( 
.A1(n_7),
.A2(n_48),
.B(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_9),
.A2(n_41),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_47),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_47),
.Y(n_147)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_10),
.A2(n_171),
.B1(n_172),
.B2(n_174),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_12),
.A2(n_66),
.B1(n_67),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_12),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_12),
.A2(n_41),
.B1(n_48),
.B2(n_135),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_135),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_135),
.Y(n_188)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_42),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_14),
.A2(n_30),
.A3(n_48),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_15),
.A2(n_41),
.B1(n_48),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_50),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_50),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_16),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_16),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_16),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

BUFx3_ASAP7_75t_SL g30 ( 
.A(n_17),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_117),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_116),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_96),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_22),
.B(n_96),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_76),
.B2(n_95),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_52),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_39),
.B(n_51),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_26),
.B(n_39),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_27),
.A2(n_32),
.B1(n_35),
.B2(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_27),
.A2(n_32),
.B1(n_60),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_27),
.A2(n_32),
.B1(n_83),
.B2(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_27),
.A2(n_32),
.B1(n_108),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_27),
.A2(n_32),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_27),
.A2(n_32),
.B1(n_183),
.B2(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_27),
.A2(n_32),
.B1(n_203),
.B2(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_27),
.A2(n_32),
.B1(n_126),
.B2(n_221),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_29),
.B(n_42),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_30),
.A2(n_31),
.B(n_133),
.C(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_32),
.B(n_133),
.Y(n_186)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_34),
.B(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_44),
.B1(n_45),
.B2(n_49),
.Y(n_39)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_40),
.A2(n_44),
.B1(n_86),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_40),
.A2(n_44),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_40),
.A2(n_44),
.B1(n_111),
.B2(n_130),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_40),
.A2(n_44),
.B1(n_157),
.B2(n_217),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_42),
.Y(n_43)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_41),
.A2(n_71),
.B1(n_132),
.B2(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_41),
.B(n_133),
.Y(n_214)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_48),
.B(n_70),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_61),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_59),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_62),
.B1(n_63),
.B2(n_75),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_54),
.A2(n_59),
.B1(n_75),
.B2(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_57),
.B(n_58),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_58),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_55),
.A2(n_57),
.B1(n_79),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_55),
.A2(n_57),
.B1(n_106),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_55),
.A2(n_56),
.B1(n_147),
.B2(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_55),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_55),
.A2(n_57),
.B1(n_173),
.B2(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_55),
.A2(n_80),
.B1(n_175),
.B2(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_55),
.A2(n_80),
.B1(n_162),
.B2(n_205),
.Y(n_211)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_59),
.Y(n_102)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_70),
.B(n_71),
.C(n_72),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_70),
.Y(n_71)
);

HAxp5_ASAP7_75t_SL g132 ( 
.A(n_67),
.B(n_133),
.CON(n_132),
.SN(n_132)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_69),
.A2(n_72),
.B1(n_132),
.B2(n_134),
.Y(n_131)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_84),
.C(n_89),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_78),
.B(n_82),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_80),
.B(n_133),
.Y(n_191)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_89),
.B1(n_90),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_84),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_87),
.A2(n_88),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_91),
.A2(n_94),
.B1(n_114),
.B2(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.C(n_103),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_101),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_103),
.B(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_109),
.C(n_112),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_104),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_107),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_259),
.B(n_264),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_163),
.B(n_246),
.C(n_258),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_148),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_120),
.B(n_148),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_136),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_122),
.B(n_123),
.C(n_136),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.C(n_131),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_131),
.B(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_134),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_143),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_138),
.B(n_142),
.C(n_143),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_141),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_146),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_153),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_149),
.B(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.C(n_160),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_155),
.B(n_231),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_159),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_245),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_240),
.B(n_244),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_226),
.B(n_239),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_207),
.B(n_225),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_195),
.B(n_206),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_184),
.B(n_194),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_176),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_176),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_180),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_189),
.B(n_193),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_187),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_197),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_204),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_202),
.C(n_204),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_209),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_215),
.B1(n_223),
.B2(n_224),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_210),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_212),
.Y(n_235)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_219),
.B1(n_220),
.B2(n_222),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_216),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_222),
.C(n_223),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_227),
.B(n_228),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_233),
.B2(n_234),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_236),
.C(n_237),
.Y(n_241)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_235),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_236),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_241),
.B(n_242),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_247),
.B(n_248),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_257),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_249),
.Y(n_257)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_255),
.C(n_257),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_260),
.B(n_261),
.Y(n_264)
);


endmodule