module fake_jpeg_4566_n_206 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_17),
.B1(n_24),
.B2(n_16),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_19),
.B(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_6),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_35),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_17),
.B1(n_13),
.B2(n_22),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_49),
.B1(n_24),
.B2(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_30),
.A2(n_17),
.B1(n_24),
.B2(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_16),
.B1(n_24),
.B2(n_33),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_28),
.A2(n_17),
.B1(n_13),
.B2(n_22),
.Y(n_49)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_59),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_47),
.B1(n_41),
.B2(n_37),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_63),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_62),
.B(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_65),
.B(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_27),
.B(n_33),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_34),
.B(n_63),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_37),
.B(n_18),
.C(n_35),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_49),
.B1(n_26),
.B2(n_42),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_26),
.B1(n_30),
.B2(n_38),
.Y(n_93)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_78),
.Y(n_91)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_34),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_81),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_54),
.B(n_37),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_51),
.Y(n_82)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_53),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_83),
.A2(n_65),
.B1(n_56),
.B2(n_62),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_70),
.C(n_68),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_96),
.B(n_77),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_94),
.B1(n_98),
.B2(n_99),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_69),
.A2(n_26),
.B1(n_42),
.B2(n_30),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_73),
.Y(n_109)
);

AO21x1_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_53),
.B(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_97),
.B(n_81),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_71),
.A2(n_36),
.B1(n_40),
.B2(n_38),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_74),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_106),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_100),
.B(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_85),
.B(n_76),
.Y(n_111)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_72),
.C(n_93),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_80),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_86),
.C(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_114),
.B(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_82),
.Y(n_115)
);

FAx1_ASAP7_75t_SL g120 ( 
.A(n_116),
.B(n_117),
.CI(n_91),
.CON(n_120),
.SN(n_120)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_84),
.Y(n_117)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_113),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_108),
.B(n_116),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_125),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_90),
.C(n_91),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_123),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_128),
.B1(n_112),
.B2(n_135),
.Y(n_137)
);

AOI211xp5_ASAP7_75t_SL g128 ( 
.A1(n_104),
.A2(n_99),
.B(n_96),
.C(n_67),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_96),
.B(n_32),
.C(n_19),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_131),
.A2(n_134),
.B1(n_106),
.B2(n_19),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_50),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_107),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_36),
.B1(n_40),
.B2(n_51),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_137),
.B(n_134),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_144),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_127),
.C(n_130),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_140),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_126),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_142),
.B(n_146),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_107),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_135),
.A2(n_60),
.B1(n_23),
.B2(n_39),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_132),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_128),
.A2(n_23),
.B1(n_78),
.B2(n_32),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_102),
.B1(n_23),
.B2(n_29),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_131),
.A2(n_102),
.B1(n_21),
.B2(n_15),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_150),
.B1(n_121),
.B2(n_45),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_20),
.B1(n_14),
.B2(n_45),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_82),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_152),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_25),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_119),
.C(n_129),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_155),
.C(n_157),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_129),
.C(n_127),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_120),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_159),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_21),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_141),
.B(n_144),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_162),
.B(n_165),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_152),
.B(n_15),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_151),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_45),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_166),
.A2(n_173),
.B1(n_163),
.B2(n_156),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_148),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_167),
.A2(n_170),
.B(n_172),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_159),
.B(n_139),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_169),
.B(n_174),
.Y(n_184)
);

NOR2xp67_ASAP7_75t_SL g170 ( 
.A(n_161),
.B(n_14),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_21),
.B1(n_20),
.B2(n_14),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_9),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_157),
.A2(n_9),
.B1(n_12),
.B2(n_11),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_161),
.B(n_25),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_177),
.B(n_25),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_158),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_185),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_176),
.Y(n_179)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_175),
.A2(n_8),
.B1(n_11),
.B2(n_10),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_8),
.C(n_11),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_183),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_171),
.B(n_25),
.Y(n_183)
);

OAI221xp5_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_21),
.B1(n_14),
.B2(n_20),
.C(n_3),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_186),
.B(n_5),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_184),
.A2(n_7),
.B(n_10),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_188),
.B(n_190),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_181),
.A2(n_7),
.B(n_10),
.Y(n_190)
);

AOI21x1_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_0),
.B(n_1),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_184),
.C(n_9),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_197),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_198),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_191),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_0),
.Y(n_198)
);

NAND3xp33_ASAP7_75t_SL g199 ( 
.A(n_194),
.B(n_3),
.C(n_4),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_199),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_201),
.A2(n_14),
.B(n_20),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_203),
.A2(n_21),
.B(n_25),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_200),
.C(n_20),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_205),
.Y(n_206)
);


endmodule