module fake_jpeg_25609_n_81 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_81);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_81;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_7),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx9p33_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx5_ASAP7_75t_SL g34 ( 
.A(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_1),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_24),
.Y(n_30)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_24),
.B(n_9),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_13),
.Y(n_37)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_28),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_23),
.B(n_30),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_44),
.C(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_17),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_29),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_34),
.B1(n_18),
.B2(n_16),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_39),
.B1(n_45),
.B2(n_44),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_34),
.B1(n_17),
.B2(n_15),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

A2O1A1O1Ixp25_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_17),
.B(n_15),
.C(n_29),
.D(n_1),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_2),
.B(n_3),
.Y(n_61)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_56),
.B(n_57),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_55),
.A2(n_45),
.B1(n_29),
.B2(n_43),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_60),
.B(n_47),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_43),
.B1(n_6),
.B2(n_4),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_61),
.A2(n_48),
.B(n_2),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_61),
.B(n_53),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_50),
.B(n_51),
.Y(n_66)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

FAx1_ASAP7_75t_SL g68 ( 
.A(n_67),
.B(n_59),
.CI(n_2),
.CON(n_68),
.SN(n_68)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_4),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_63),
.B1(n_62),
.B2(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_71),
.B(n_73),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_72),
.C(n_69),
.Y(n_76)
);

AOI21x1_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_77),
.B(n_69),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_68),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_5),
.Y(n_79)
);

AO21x1_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_7),
.B(n_8),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_80),
.B(n_54),
.Y(n_81)
);


endmodule