module fake_ariane_240_n_1695 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1695);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1695;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_146;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_145;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1429;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_147;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx2_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_35),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_52),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_59),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_73),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_16),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_61),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_25),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_66),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_92),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_121),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_89),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_136),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_34),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_50),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_90),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_70),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_49),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_108),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_56),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_7),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_44),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_20),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_93),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_8),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_3),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_47),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_47),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_54),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_23),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_94),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_6),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_75),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_31),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_38),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_5),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_40),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_81),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_129),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_85),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_124),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_1),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_104),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_7),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_122),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_33),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_82),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_38),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_87),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_14),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_1),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_21),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_130),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_115),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_46),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_34),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_48),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_16),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_9),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_60),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_120),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_96),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_98),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_67),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_20),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_51),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_55),
.Y(n_223)
);

BUFx2_ASAP7_75t_R g224 ( 
.A(n_37),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_3),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_77),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_86),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_80),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_144),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_101),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_76),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_68),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_52),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_135),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_25),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_26),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_84),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_53),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_21),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_111),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_43),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_14),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_27),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_64),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_50),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_9),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_123),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_107),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_40),
.Y(n_249)
);

BUFx8_ASAP7_75t_SL g250 ( 
.A(n_51),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_57),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_5),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_131),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_53),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_91),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_39),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_69),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_31),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_43),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_27),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_36),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_134),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_72),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_22),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_128),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_99),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g267 ( 
.A(n_126),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_6),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_110),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_114),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_18),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_39),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_32),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_102),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_32),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_26),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_105),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_24),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_141),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_8),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_78),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_37),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_103),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_137),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_71),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_65),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_15),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_127),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_4),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_46),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_133),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_83),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_18),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_30),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_13),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_109),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_178),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_222),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_250),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_160),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_219),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_222),
.Y(n_302)
);

INVxp33_ASAP7_75t_SL g303 ( 
.A(n_147),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_222),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_277),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_222),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_261),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_283),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_147),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_222),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_149),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_149),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_170),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_146),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_152),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_152),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_163),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_146),
.Y(n_318)
);

INVxp33_ASAP7_75t_SL g319 ( 
.A(n_166),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_190),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_181),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_163),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_180),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_180),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_226),
.Y(n_325)
);

INVxp33_ASAP7_75t_SL g326 ( 
.A(n_166),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_233),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_226),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_193),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_272),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_229),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_229),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_230),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_230),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_150),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_154),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_235),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_156),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_191),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_272),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_191),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g342 ( 
.A(n_167),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_182),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_185),
.Y(n_344)
);

INVxp33_ASAP7_75t_SL g345 ( 
.A(n_173),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_187),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_192),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_218),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_281),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_206),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_218),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_208),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_249),
.Y(n_353)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_173),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_214),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_221),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_198),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_225),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_200),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g360 ( 
.A(n_239),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_242),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_259),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_246),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_194),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_202),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_232),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_254),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_258),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_204),
.Y(n_369)
);

INVxp33_ASAP7_75t_SL g370 ( 
.A(n_175),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_260),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_268),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_364),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_313),
.A2(n_224),
.B1(n_295),
.B2(n_256),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_364),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_300),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_298),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_298),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_302),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_302),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_304),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_304),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_301),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_306),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_306),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_323),
.B(n_145),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_310),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_330),
.B(n_189),
.Y(n_389)
);

AND2x6_ASAP7_75t_L g390 ( 
.A(n_314),
.B(n_183),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_310),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_311),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_311),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_312),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_312),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_315),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_305),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_297),
.A2(n_273),
.B1(n_264),
.B2(n_238),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_330),
.Y(n_400)
);

BUFx8_ASAP7_75t_L g401 ( 
.A(n_314),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_366),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_316),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_316),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_340),
.B(n_269),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_317),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_317),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_322),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_325),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_325),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_366),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_328),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_309),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_328),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_331),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_331),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_308),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_332),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_323),
.B(n_148),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_320),
.Y(n_421)
);

OA21x2_ASAP7_75t_L g422 ( 
.A1(n_332),
.A2(n_157),
.B(n_155),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_333),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_340),
.B(n_251),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_297),
.A2(n_360),
.B1(n_342),
.B2(n_349),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_314),
.B(n_255),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_333),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_321),
.Y(n_428)
);

OA21x2_ASAP7_75t_L g429 ( 
.A1(n_334),
.A2(n_161),
.B(n_158),
.Y(n_429)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_323),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_334),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_323),
.B(n_251),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_318),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_335),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_335),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_336),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_318),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_318),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_339),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_339),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_336),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_339),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_341),
.B(n_255),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_373),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_421),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_373),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_377),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_376),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_373),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_377),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_375),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_433),
.B(n_341),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_324),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_433),
.B(n_349),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_389),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_341),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_375),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_401),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_430),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_438),
.Y(n_460)
);

AOI21x1_ASAP7_75t_L g461 ( 
.A1(n_375),
.A2(n_420),
.B(n_422),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_421),
.B(n_329),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_400),
.B(n_307),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_389),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_437),
.B(n_348),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_405),
.B(n_357),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_378),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_379),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_405),
.B(n_359),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_378),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_380),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_430),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_376),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_379),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_424),
.B(n_363),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_379),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_379),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_425),
.A2(n_363),
.B1(n_241),
.B2(n_175),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_430),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_405),
.B(n_365),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_425),
.A2(n_176),
.B1(n_271),
.B2(n_236),
.Y(n_481)
);

NAND2xp33_ASAP7_75t_L g482 ( 
.A(n_402),
.B(n_369),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_379),
.Y(n_483)
);

OR2x6_ASAP7_75t_L g484 ( 
.A(n_424),
.B(n_338),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_380),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_389),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_422),
.A2(n_319),
.B1(n_354),
.B2(n_370),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_426),
.B(n_348),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_430),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_437),
.B(n_348),
.Y(n_490)
);

NOR2x1p5_ASAP7_75t_L g491 ( 
.A(n_402),
.B(n_299),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_381),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_430),
.Y(n_493)
);

AND2x2_ASAP7_75t_SL g494 ( 
.A(n_422),
.B(n_183),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_381),
.Y(n_495)
);

BUFx6f_ASAP7_75t_SL g496 ( 
.A(n_426),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_383),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_385),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_383),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_384),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_400),
.B(n_303),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_414),
.B(n_338),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_412),
.B(n_326),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_383),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_385),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_383),
.Y(n_506)
);

BUFx4f_ASAP7_75t_L g507 ( 
.A(n_390),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_387),
.B(n_345),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_383),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_437),
.B(n_351),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_376),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_376),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_386),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_401),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_386),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_437),
.B(n_351),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_401),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_376),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_434),
.B(n_343),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_376),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_376),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_388),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_397),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_388),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_426),
.B(n_443),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_412),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_376),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g528 ( 
.A(n_432),
.B(n_266),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_391),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_391),
.Y(n_530)
);

AO22x2_ASAP7_75t_L g531 ( 
.A1(n_426),
.A2(n_284),
.B1(n_282),
.B2(n_280),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_422),
.A2(n_351),
.B1(n_294),
.B2(n_243),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_394),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_394),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_414),
.B(n_344),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_394),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_394),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_394),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_387),
.B(n_151),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_394),
.Y(n_540)
);

NOR2x1p5_ASAP7_75t_L g541 ( 
.A(n_418),
.B(n_176),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_394),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_435),
.B(n_344),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_394),
.Y(n_544)
);

CKINVDCx6p67_ASAP7_75t_R g545 ( 
.A(n_428),
.Y(n_545)
);

AND3x2_ASAP7_75t_L g546 ( 
.A(n_426),
.B(n_347),
.C(n_346),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_395),
.Y(n_547)
);

NOR3xp33_ASAP7_75t_L g548 ( 
.A(n_374),
.B(n_241),
.C(n_236),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_395),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_395),
.Y(n_550)
);

NAND3xp33_ASAP7_75t_L g551 ( 
.A(n_420),
.B(n_172),
.C(n_169),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_390),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_443),
.B(n_346),
.Y(n_553)
);

AND3x2_ASAP7_75t_L g554 ( 
.A(n_443),
.B(n_350),
.C(n_347),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_438),
.B(n_439),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_395),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_395),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_395),
.Y(n_558)
);

INVx11_ASAP7_75t_L g559 ( 
.A(n_401),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_L g560 ( 
.A(n_422),
.B(n_429),
.C(n_435),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_436),
.B(n_350),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_436),
.B(n_352),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_395),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_429),
.A2(n_243),
.B1(n_371),
.B2(n_368),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_395),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_401),
.Y(n_566)
);

CKINVDCx6p67_ASAP7_75t_R g567 ( 
.A(n_428),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_438),
.B(n_352),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_411),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_411),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_443),
.B(n_441),
.Y(n_571)
);

CKINVDCx6p67_ASAP7_75t_R g572 ( 
.A(n_390),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_411),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_411),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_411),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_443),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_441),
.B(n_151),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_411),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_399),
.B(n_153),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_432),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_439),
.B(n_355),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_411),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_393),
.B(n_355),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_399),
.B(n_153),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_411),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_439),
.B(n_356),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_418),
.Y(n_587)
);

OR2x6_ASAP7_75t_L g588 ( 
.A(n_374),
.B(n_356),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_419),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_419),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_419),
.Y(n_591)
);

BUFx10_ASAP7_75t_L g592 ( 
.A(n_390),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_L g593 ( 
.A(n_390),
.B(n_440),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_508),
.A2(n_432),
.B1(n_442),
.B2(n_440),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_475),
.B(n_440),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_478),
.A2(n_429),
.B1(n_442),
.B2(n_406),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_475),
.B(n_442),
.Y(n_597)
);

OAI22xp33_ASAP7_75t_L g598 ( 
.A1(n_481),
.A2(n_295),
.B1(n_245),
.B2(n_293),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_467),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_475),
.B(n_393),
.Y(n_600)
);

OAI221xp5_ASAP7_75t_L g601 ( 
.A1(n_478),
.A2(n_290),
.B1(n_293),
.B2(n_245),
.C(n_289),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_470),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_475),
.B(n_393),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_449),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_453),
.B(n_580),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_500),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_453),
.B(n_393),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_484),
.B(n_392),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_500),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_445),
.B(n_393),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_523),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_445),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_470),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_455),
.B(n_398),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_459),
.B(n_398),
.Y(n_615)
);

NAND3xp33_ASAP7_75t_L g616 ( 
.A(n_501),
.B(n_256),
.C(n_252),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_449),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_464),
.B(n_327),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_580),
.B(n_398),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_464),
.B(n_337),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_455),
.Y(n_621)
);

A2O1A1Ixp33_ASAP7_75t_L g622 ( 
.A1(n_576),
.A2(n_398),
.B(n_416),
.C(n_392),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_583),
.B(n_398),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_583),
.B(n_416),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_459),
.B(n_416),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_484),
.B(n_396),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_486),
.B(n_353),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_481),
.A2(n_429),
.B1(n_410),
.B2(n_396),
.Y(n_628)
);

NOR2xp67_ASAP7_75t_L g629 ( 
.A(n_523),
.B(n_416),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_484),
.B(n_416),
.Y(n_630)
);

O2A1O1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_553),
.A2(n_571),
.B(n_539),
.C(n_525),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_471),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_459),
.B(n_419),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_451),
.Y(n_634)
);

AND2x4_ASAP7_75t_SL g635 ( 
.A(n_484),
.B(n_362),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_526),
.B(n_358),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_502),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_485),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_466),
.B(n_469),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_451),
.Y(n_640)
);

OAI221xp5_ASAP7_75t_L g641 ( 
.A1(n_487),
.A2(n_271),
.B1(n_252),
.B2(n_287),
.C(n_289),
.Y(n_641)
);

AND2x6_ASAP7_75t_L g642 ( 
.A(n_559),
.B(n_403),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_472),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_480),
.B(n_403),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_472),
.B(n_479),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_447),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_587),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_526),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_460),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_484),
.B(n_404),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_502),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_485),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_576),
.B(n_404),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_519),
.B(n_406),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_519),
.B(n_407),
.Y(n_655)
);

INVx8_ASAP7_75t_L g656 ( 
.A(n_496),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_564),
.A2(n_429),
.B1(n_408),
.B2(n_409),
.Y(n_657)
);

INVxp67_ASAP7_75t_SL g658 ( 
.A(n_472),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_479),
.B(n_419),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_460),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_460),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_492),
.Y(n_662)
);

AOI221xp5_ASAP7_75t_L g663 ( 
.A1(n_579),
.A2(n_290),
.B1(n_287),
.B2(n_368),
.C(n_358),
.Y(n_663)
);

O2A1O1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_495),
.A2(n_409),
.B(n_410),
.C(n_413),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_496),
.A2(n_415),
.B1(n_413),
.B2(n_284),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_496),
.A2(n_415),
.B1(n_159),
.B2(n_168),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_495),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_531),
.A2(n_423),
.B1(n_419),
.B2(n_431),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_479),
.B(n_419),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_543),
.B(n_417),
.Y(n_670)
);

INVxp67_ASAP7_75t_SL g671 ( 
.A(n_489),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_444),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_454),
.B(n_431),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_488),
.B(n_361),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_498),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_452),
.B(n_431),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_498),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_543),
.B(n_417),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_489),
.B(n_419),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_561),
.B(n_417),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_561),
.B(n_427),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_562),
.B(n_427),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_562),
.B(n_427),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_577),
.B(n_207),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_447),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_488),
.B(n_423),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_488),
.B(n_489),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_535),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_462),
.B(n_211),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_493),
.B(n_423),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_444),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_488),
.B(n_423),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_505),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_446),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_493),
.B(n_212),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_446),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_505),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_457),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_531),
.A2(n_423),
.B1(n_243),
.B2(n_266),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_513),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_493),
.B(n_423),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_545),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_448),
.B(n_423),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_457),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_448),
.B(n_423),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_468),
.Y(n_706)
);

AND2x4_ASAP7_75t_SL g707 ( 
.A(n_545),
.B(n_367),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_513),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_568),
.B(n_165),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_531),
.A2(n_532),
.B1(n_584),
.B2(n_588),
.Y(n_710)
);

AND2x4_ASAP7_75t_SL g711 ( 
.A(n_567),
.B(n_367),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_535),
.B(n_213),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_463),
.B(n_215),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_528),
.B(n_162),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_528),
.B(n_162),
.Y(n_715)
);

BUFx5_ASAP7_75t_L g716 ( 
.A(n_592),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_515),
.B(n_275),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_528),
.B(n_164),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_468),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_450),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_482),
.B(n_371),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_567),
.B(n_372),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_515),
.B(n_276),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_546),
.B(n_168),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_474),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_503),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_SL g727 ( 
.A(n_458),
.B(n_278),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_541),
.B(n_588),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_448),
.B(n_171),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_522),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_522),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_491),
.B(n_171),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_560),
.A2(n_228),
.B(n_205),
.C(n_244),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_507),
.Y(n_734)
);

A2O1A1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_560),
.A2(n_179),
.B(n_177),
.C(n_196),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_524),
.Y(n_736)
);

OAI21xp5_ASAP7_75t_L g737 ( 
.A1(n_494),
.A2(n_174),
.B(n_270),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_474),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_448),
.B(n_209),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_524),
.A2(n_237),
.B1(n_292),
.B2(n_231),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_448),
.B(n_210),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_588),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_473),
.B(n_210),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_476),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_529),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_476),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_477),
.Y(n_747)
);

NAND2x1p5_ASAP7_75t_L g748 ( 
.A(n_514),
.B(n_285),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_554),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_477),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_483),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_541),
.B(n_223),
.Y(n_752)
);

AO22x1_ASAP7_75t_L g753 ( 
.A1(n_685),
.A2(n_548),
.B1(n_566),
.B2(n_517),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_599),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_604),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_608),
.B(n_473),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_602),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_639),
.B(n_588),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_608),
.B(n_517),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_604),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_613),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_673),
.B(n_614),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_SL g763 ( 
.A1(n_742),
.A2(n_588),
.B1(n_531),
.B2(n_566),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_673),
.B(n_530),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_632),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_612),
.B(n_494),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_608),
.B(n_483),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_617),
.Y(n_768)
);

BUFx12f_ASAP7_75t_L g769 ( 
.A(n_611),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_605),
.B(n_581),
.Y(n_770)
);

O2A1O1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_598),
.A2(n_509),
.B(n_497),
.C(n_506),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_713),
.A2(n_551),
.B1(n_494),
.B2(n_509),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_638),
.Y(n_773)
);

A2O1A1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_737),
.A2(n_551),
.B(n_504),
.C(n_499),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_626),
.B(n_674),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_707),
.Y(n_776)
);

OR2x6_ASAP7_75t_L g777 ( 
.A(n_656),
.B(n_552),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_646),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_652),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_713),
.A2(n_506),
.B1(n_504),
.B2(n_499),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_626),
.B(n_687),
.Y(n_781)
);

INVx5_ASAP7_75t_L g782 ( 
.A(n_656),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_721),
.B(n_586),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_707),
.Y(n_784)
);

BUFx4f_ASAP7_75t_L g785 ( 
.A(n_656),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_607),
.B(n_497),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_626),
.Y(n_787)
);

INVx5_ASAP7_75t_L g788 ( 
.A(n_642),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_637),
.B(n_461),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_651),
.B(n_461),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_662),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_606),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_712),
.B(n_555),
.Y(n_793)
);

INVx1_ASAP7_75t_SL g794 ( 
.A(n_618),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_639),
.A2(n_542),
.B1(n_590),
.B2(n_537),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_620),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_734),
.Y(n_797)
);

NAND3xp33_ASAP7_75t_SL g798 ( 
.A(n_601),
.B(n_237),
.C(n_231),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_667),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_630),
.B(n_473),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_675),
.Y(n_801)
);

XOR2xp5_ASAP7_75t_L g802 ( 
.A(n_606),
.B(n_456),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_617),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_634),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_629),
.B(n_473),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_711),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_712),
.B(n_465),
.Y(n_807)
);

OR2x4_ASAP7_75t_L g808 ( 
.A(n_717),
.B(n_547),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_677),
.B(n_473),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_693),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_711),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_717),
.B(n_490),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_723),
.B(n_510),
.Y(n_813)
);

AND2x6_ASAP7_75t_L g814 ( 
.A(n_734),
.B(n_697),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_700),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_723),
.B(n_516),
.Y(n_816)
);

INVx6_ASAP7_75t_L g817 ( 
.A(n_674),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_634),
.Y(n_818)
);

NAND3xp33_ASAP7_75t_SL g819 ( 
.A(n_689),
.B(n_247),
.C(n_248),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_708),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_636),
.B(n_542),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_647),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_710),
.A2(n_572),
.B1(n_552),
.B2(n_390),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_688),
.B(n_590),
.Y(n_824)
);

INVx5_ASAP7_75t_L g825 ( 
.A(n_642),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_641),
.A2(n_572),
.B1(n_552),
.B2(n_390),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_730),
.B(n_520),
.Y(n_827)
);

INVxp67_ASAP7_75t_SL g828 ( 
.A(n_595),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_SL g829 ( 
.A1(n_635),
.A2(n_285),
.B1(n_296),
.B2(n_253),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_645),
.A2(n_518),
.B(n_521),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_645),
.A2(n_518),
.B(n_521),
.Y(n_831)
);

AO21x1_ASAP7_75t_L g832 ( 
.A1(n_729),
.A2(n_538),
.B(n_537),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_731),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_609),
.Y(n_834)
);

OR2x6_ASAP7_75t_L g835 ( 
.A(n_609),
.B(n_552),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_736),
.B(n_520),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_640),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_644),
.B(n_511),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_600),
.B(n_511),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_627),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_603),
.B(n_512),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_603),
.B(n_512),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_621),
.B(n_527),
.Y(n_843)
);

AND2x6_ASAP7_75t_L g844 ( 
.A(n_745),
.B(n_533),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_642),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_597),
.A2(n_390),
.B1(n_533),
.B2(n_591),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_640),
.Y(n_847)
);

OAI21xp5_ASAP7_75t_L g848 ( 
.A1(n_622),
.A2(n_527),
.B(n_534),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_642),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_701),
.A2(n_520),
.B(n_534),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_635),
.B(n_536),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_709),
.B(n_536),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_670),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_672),
.Y(n_854)
);

INVx4_ASAP7_75t_L g855 ( 
.A(n_642),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_726),
.B(n_520),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_691),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_678),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_654),
.B(n_540),
.Y(n_859)
);

INVx5_ASAP7_75t_L g860 ( 
.A(n_649),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_749),
.B(n_540),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_680),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_722),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_720),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_610),
.B(n_538),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_681),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_623),
.A2(n_558),
.B(n_549),
.C(n_557),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_655),
.B(n_544),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_727),
.A2(n_570),
.B1(n_549),
.B2(n_557),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_694),
.B(n_696),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_694),
.B(n_547),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_682),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_686),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_648),
.Y(n_874)
);

OAI22xp33_ASAP7_75t_L g875 ( 
.A1(n_650),
.A2(n_247),
.B1(n_286),
.B2(n_288),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_698),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_702),
.B(n_752),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_628),
.A2(n_390),
.B1(n_575),
.B2(n_591),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_683),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_699),
.A2(n_550),
.B1(n_565),
.B2(n_589),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_748),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_698),
.Y(n_882)
);

CKINVDCx14_ASAP7_75t_R g883 ( 
.A(n_728),
.Y(n_883)
);

NAND2x1p5_ASAP7_75t_L g884 ( 
.A(n_649),
.B(n_507),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_610),
.B(n_616),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_668),
.A2(n_574),
.B1(n_565),
.B2(n_589),
.Y(n_886)
);

OAI221xp5_ASAP7_75t_L g887 ( 
.A1(n_663),
.A2(n_563),
.B1(n_570),
.B2(n_573),
.C(n_558),
.Y(n_887)
);

NAND2x1p5_ASAP7_75t_L g888 ( 
.A(n_660),
.B(n_507),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_732),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_692),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_695),
.B(n_624),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_643),
.B(n_556),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_689),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_660),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_661),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_704),
.Y(n_896)
);

AND2x6_ASAP7_75t_SL g897 ( 
.A(n_684),
.B(n_199),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_658),
.B(n_569),
.Y(n_898)
);

AOI21xp33_ASAP7_75t_L g899 ( 
.A1(n_684),
.A2(n_573),
.B(n_563),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_704),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_706),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_661),
.Y(n_902)
);

NOR2x2_ASAP7_75t_L g903 ( 
.A(n_706),
.B(n_569),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_748),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_751),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_724),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_719),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_716),
.B(n_547),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_725),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_666),
.B(n_574),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_716),
.B(n_547),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_671),
.B(n_575),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_725),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_738),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_738),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_744),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_746),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_746),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_716),
.B(n_547),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_665),
.B(n_578),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_740),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_653),
.B(n_578),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_594),
.A2(n_582),
.B1(n_585),
.B2(n_593),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_747),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_676),
.B(n_582),
.Y(n_925)
);

O2A1O1Ixp5_ASAP7_75t_SL g926 ( 
.A1(n_899),
.A2(n_729),
.B(n_743),
.C(n_741),
.Y(n_926)
);

INVx8_ASAP7_75t_L g927 ( 
.A(n_782),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_762),
.A2(n_619),
.B1(n_596),
.B2(n_631),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_893),
.B(n_714),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_921),
.A2(n_664),
.B(n_741),
.C(n_743),
.Y(n_930)
);

BUFx4f_ASAP7_75t_L g931 ( 
.A(n_769),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_764),
.A2(n_690),
.B(n_679),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_758),
.B(n_750),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_754),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_758),
.B(n_739),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_757),
.Y(n_936)
);

OR2x6_ASAP7_75t_SL g937 ( 
.A(n_778),
.B(n_248),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_885),
.A2(n_735),
.B(n_733),
.C(n_718),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_909),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_793),
.B(n_750),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_775),
.B(n_751),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_774),
.A2(n_615),
.B(n_625),
.Y(n_942)
);

O2A1O1Ixp5_ASAP7_75t_L g943 ( 
.A1(n_832),
.A2(n_739),
.B(n_703),
.C(n_705),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_925),
.A2(n_633),
.B(n_659),
.Y(n_944)
);

AO32x1_ASAP7_75t_L g945 ( 
.A1(n_789),
.A2(n_585),
.A3(n_227),
.B1(n_234),
.B2(n_240),
.Y(n_945)
);

OR2x6_ASAP7_75t_L g946 ( 
.A(n_775),
.B(n_715),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_782),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_863),
.B(n_615),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_822),
.Y(n_949)
);

O2A1O1Ixp5_ASAP7_75t_L g950 ( 
.A1(n_807),
.A2(n_703),
.B(n_705),
.C(n_669),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_853),
.A2(n_657),
.B1(n_625),
.B2(n_659),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_908),
.A2(n_716),
.B(n_220),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_858),
.A2(n_262),
.B1(n_257),
.B2(n_286),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_761),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_834),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_R g956 ( 
.A(n_834),
.B(n_257),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_911),
.A2(n_216),
.B(n_184),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_SL g958 ( 
.A(n_855),
.B(n_592),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_772),
.A2(n_296),
.B(n_263),
.C(n_292),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_782),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_819),
.A2(n_265),
.B(n_291),
.C(n_288),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_765),
.Y(n_962)
);

OAI21xp33_ASAP7_75t_SL g963 ( 
.A1(n_781),
.A2(n_0),
.B(n_2),
.Y(n_963)
);

OAI21x1_ASAP7_75t_L g964 ( 
.A1(n_848),
.A2(n_592),
.B(n_267),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_SL g965 ( 
.A1(n_864),
.A2(n_291),
.B1(n_265),
.B2(n_263),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_782),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_798),
.A2(n_382),
.B(n_279),
.C(n_274),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_785),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_798),
.A2(n_382),
.B(n_195),
.C(n_217),
.Y(n_969)
);

OAI21x1_ASAP7_75t_L g970 ( 
.A1(n_830),
.A2(n_267),
.B(n_194),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_909),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_919),
.A2(n_201),
.B(n_197),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_787),
.B(n_382),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_915),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_796),
.Y(n_975)
);

BUFx12f_ASAP7_75t_L g976 ( 
.A(n_792),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_773),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_779),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_915),
.Y(n_979)
);

AOI21x1_ASAP7_75t_L g980 ( 
.A1(n_805),
.A2(n_382),
.B(n_267),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_862),
.A2(n_382),
.B(n_188),
.C(n_186),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_866),
.B(n_872),
.Y(n_982)
);

INVxp67_ASAP7_75t_SL g983 ( 
.A(n_787),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_785),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_812),
.A2(n_0),
.B(n_2),
.C(n_4),
.Y(n_985)
);

O2A1O1Ixp5_ASAP7_75t_L g986 ( 
.A1(n_805),
.A2(n_382),
.B(n_11),
.C(n_12),
.Y(n_986)
);

AO22x1_ASAP7_75t_L g987 ( 
.A1(n_889),
.A2(n_203),
.B1(n_183),
.B2(n_382),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_879),
.A2(n_382),
.B1(n_203),
.B2(n_183),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_874),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_863),
.B(n_817),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_864),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_856),
.A2(n_203),
.B(n_183),
.C(n_194),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_783),
.B(n_10),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_835),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_797),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_759),
.B(n_267),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_854),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_817),
.B(n_10),
.Y(n_998)
);

BUFx2_ASAP7_75t_SL g999 ( 
.A(n_792),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_770),
.B(n_194),
.Y(n_1000)
);

OR2x2_ASAP7_75t_SL g1001 ( 
.A(n_897),
.B(n_203),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_856),
.A2(n_203),
.B(n_267),
.C(n_194),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_776),
.B(n_784),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_791),
.A2(n_13),
.B1(n_15),
.B2(n_17),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_813),
.A2(n_17),
.B(n_19),
.C(n_22),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_SL g1006 ( 
.A(n_855),
.B(n_267),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_903),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_SL g1008 ( 
.A(n_788),
.B(n_267),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_794),
.B(n_19),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_799),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_801),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_840),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_781),
.A2(n_194),
.B1(n_267),
.B2(n_28),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_806),
.B(n_194),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_810),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_817),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_816),
.A2(n_194),
.B(n_24),
.C(n_28),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_859),
.A2(n_63),
.B(n_140),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_815),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_883),
.B(n_29),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_883),
.B(n_29),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_774),
.A2(n_831),
.B(n_865),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_820),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_833),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_828),
.B(n_766),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_877),
.B(n_30),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_857),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_868),
.A2(n_74),
.B(n_139),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_802),
.B(n_33),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_875),
.A2(n_35),
.B(n_36),
.C(n_41),
.Y(n_1030)
);

NOR2xp67_ASAP7_75t_SL g1031 ( 
.A(n_788),
.B(n_41),
.Y(n_1031)
);

OR2x2_ASAP7_75t_L g1032 ( 
.A(n_811),
.B(n_42),
.Y(n_1032)
);

NOR2x1_ASAP7_75t_L g1033 ( 
.A(n_881),
.B(n_95),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_906),
.Y(n_1034)
);

NOR3xp33_ASAP7_75t_L g1035 ( 
.A(n_753),
.B(n_42),
.C(n_44),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_R g1036 ( 
.A(n_845),
.B(n_849),
.Y(n_1036)
);

OR2x6_ASAP7_75t_L g1037 ( 
.A(n_777),
.B(n_45),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_821),
.B(n_48),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_797),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_808),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_829),
.B(n_49),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_L g1042 ( 
.A(n_875),
.B(n_58),
.C(n_62),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_896),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_865),
.A2(n_117),
.B(n_125),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_851),
.Y(n_1045)
);

INVx6_ASAP7_75t_L g1046 ( 
.A(n_881),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_771),
.A2(n_142),
.B(n_867),
.C(n_843),
.Y(n_1047)
);

AOI21xp33_ASAP7_75t_L g1048 ( 
.A1(n_763),
.A2(n_790),
.B(n_852),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_809),
.A2(n_827),
.B(n_836),
.C(n_824),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_922),
.A2(n_850),
.B(n_898),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_861),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_835),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_900),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_892),
.A2(n_912),
.B(n_871),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_808),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_SL g1056 ( 
.A1(n_942),
.A2(n_869),
.B(n_842),
.Y(n_1056)
);

AOI221xp5_ASAP7_75t_SL g1057 ( 
.A1(n_1030),
.A2(n_887),
.B1(n_786),
.B2(n_836),
.C(n_827),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_931),
.Y(n_1058)
);

OAI21xp33_ASAP7_75t_L g1059 ( 
.A1(n_935),
.A2(n_829),
.B(n_763),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_970),
.A2(n_871),
.B(n_809),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_1017),
.A2(n_756),
.B(n_800),
.C(n_835),
.Y(n_1061)
);

AO32x2_ASAP7_75t_L g1062 ( 
.A1(n_928),
.A2(n_903),
.A3(n_870),
.B1(n_800),
.B2(n_902),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_1037),
.A2(n_756),
.B1(n_878),
.B2(n_780),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_948),
.B(n_797),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1025),
.B(n_902),
.Y(n_1065)
);

AO31x2_ASAP7_75t_L g1066 ( 
.A1(n_1050),
.A2(n_938),
.A3(n_1047),
.B(n_1002),
.Y(n_1066)
);

INVx4_ASAP7_75t_L g1067 ( 
.A(n_968),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_934),
.Y(n_1068)
);

BUFx12f_ASAP7_75t_L g1069 ( 
.A(n_976),
.Y(n_1069)
);

INVx5_ASAP7_75t_L g1070 ( 
.A(n_1037),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_1022),
.A2(n_882),
.B(n_876),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_928),
.A2(n_838),
.B(n_923),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_936),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_933),
.B(n_873),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_982),
.B(n_873),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_1022),
.A2(n_964),
.B(n_1054),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_949),
.B(n_861),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_940),
.B(n_890),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_926),
.A2(n_795),
.B(n_839),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_950),
.A2(n_841),
.B(n_886),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_943),
.A2(n_924),
.B(n_918),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_989),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_944),
.A2(n_907),
.B(n_913),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_1012),
.Y(n_1084)
);

NAND2x1_ASAP7_75t_L g1085 ( 
.A(n_994),
.B(n_814),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_1007),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_931),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_955),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1037),
.A2(n_878),
.B1(n_823),
.B2(n_825),
.Y(n_1089)
);

AO22x2_ASAP7_75t_L g1090 ( 
.A1(n_1007),
.A2(n_910),
.B1(n_917),
.B2(n_847),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_961),
.A2(n_890),
.B(n_920),
.C(n_845),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1020),
.B(n_904),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_991),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_983),
.B(n_941),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_954),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_997),
.Y(n_1096)
);

AO21x2_ASAP7_75t_L g1097 ( 
.A1(n_1048),
.A2(n_901),
.B(n_914),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1021),
.B(n_904),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_975),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_968),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1027),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_956),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_962),
.B(n_767),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_977),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_965),
.B(n_895),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_932),
.A2(n_886),
.B(n_880),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1029),
.B(n_895),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1044),
.A2(n_952),
.B(n_951),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_968),
.Y(n_1109)
);

NOR2x1_ASAP7_75t_R g1110 ( 
.A(n_984),
.B(n_797),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_951),
.A2(n_860),
.B(n_849),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_SL g1112 ( 
.A1(n_967),
.A2(n_969),
.B(n_1038),
.C(n_959),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_978),
.B(n_767),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_930),
.A2(n_860),
.B(n_880),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1010),
.B(n_767),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1013),
.A2(n_823),
.B(n_826),
.C(n_894),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1049),
.A2(n_916),
.B(n_888),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1018),
.A2(n_884),
.B(n_760),
.Y(n_1118)
);

CKINVDCx11_ASAP7_75t_R g1119 ( 
.A(n_937),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1006),
.A2(n_860),
.B(n_895),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_958),
.A2(n_895),
.B(n_905),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_1026),
.Y(n_1122)
);

O2A1O1Ixp5_ASAP7_75t_SL g1123 ( 
.A1(n_929),
.A2(n_844),
.B(n_905),
.C(n_768),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1028),
.A2(n_755),
.B(n_837),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_1034),
.Y(n_1125)
);

AO21x2_ASAP7_75t_L g1126 ( 
.A1(n_1048),
.A2(n_818),
.B(n_804),
.Y(n_1126)
);

OA21x2_ASAP7_75t_L g1127 ( 
.A1(n_992),
.A2(n_803),
.B(n_846),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_958),
.A2(n_777),
.B(n_846),
.Y(n_1128)
);

OA21x2_ASAP7_75t_L g1129 ( 
.A1(n_1000),
.A2(n_826),
.B(n_844),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_993),
.A2(n_814),
.B(n_767),
.C(n_844),
.Y(n_1130)
);

OA21x2_ASAP7_75t_L g1131 ( 
.A1(n_1000),
.A2(n_844),
.B(n_814),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_1016),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_984),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_984),
.Y(n_1134)
);

NAND3x1_ASAP7_75t_L g1135 ( 
.A(n_1041),
.B(n_1035),
.C(n_998),
.Y(n_1135)
);

INVx1_ASAP7_75t_SL g1136 ( 
.A(n_1051),
.Y(n_1136)
);

AOI221x1_ASAP7_75t_L g1137 ( 
.A1(n_1042),
.A2(n_1004),
.B1(n_988),
.B2(n_981),
.C(n_953),
.Y(n_1137)
);

O2A1O1Ixp5_ASAP7_75t_SL g1138 ( 
.A1(n_1004),
.A2(n_1014),
.B(n_1043),
.C(n_1053),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_SL g1139 ( 
.A1(n_1052),
.A2(n_985),
.B(n_1005),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1008),
.A2(n_988),
.B(n_987),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1009),
.A2(n_953),
.B1(n_1055),
.B2(n_1045),
.Y(n_1141)
);

AO31x2_ASAP7_75t_L g1142 ( 
.A1(n_939),
.A2(n_974),
.A3(n_971),
.B(n_979),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_947),
.B(n_960),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1011),
.B(n_1015),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_945),
.A2(n_1019),
.B(n_1024),
.Y(n_1145)
);

NOR2xp67_ASAP7_75t_SL g1146 ( 
.A(n_999),
.B(n_966),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1033),
.A2(n_986),
.B(n_996),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1023),
.A2(n_972),
.B(n_957),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1052),
.B(n_946),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_990),
.A2(n_1040),
.B1(n_946),
.B2(n_1003),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_946),
.B(n_973),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1032),
.B(n_1046),
.Y(n_1152)
);

OAI22x1_ASAP7_75t_L g1153 ( 
.A1(n_1001),
.A2(n_963),
.B1(n_945),
.B2(n_1031),
.Y(n_1153)
);

AOI221x1_ASAP7_75t_L g1154 ( 
.A1(n_995),
.A2(n_1039),
.B1(n_947),
.B2(n_960),
.C(n_966),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_947),
.B(n_960),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_995),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_927),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_1039),
.B(n_1046),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_927),
.B(n_1036),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_935),
.A2(n_758),
.B(n_713),
.C(n_793),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_938),
.A2(n_928),
.B(n_1022),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_968),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_935),
.B(n_762),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1020),
.B(n_464),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_935),
.B(n_762),
.Y(n_1165)
);

AO31x2_ASAP7_75t_L g1166 ( 
.A1(n_1050),
.A2(n_832),
.A3(n_938),
.B(n_1047),
.Y(n_1166)
);

AO32x2_ASAP7_75t_L g1167 ( 
.A1(n_928),
.A2(n_1004),
.A3(n_951),
.B1(n_988),
.B2(n_953),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_935),
.B(n_762),
.Y(n_1168)
);

INVx2_ASAP7_75t_SL g1169 ( 
.A(n_931),
.Y(n_1169)
);

NOR2xp67_ASAP7_75t_L g1170 ( 
.A(n_976),
.B(n_612),
.Y(n_1170)
);

AO32x2_ASAP7_75t_L g1171 ( 
.A1(n_928),
.A2(n_1004),
.A3(n_951),
.B1(n_988),
.B2(n_953),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_935),
.A2(n_893),
.B1(n_445),
.B2(n_758),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_927),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_968),
.B(n_775),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1050),
.A2(n_762),
.B(n_891),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_989),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_935),
.B(n_762),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_935),
.A2(n_762),
.B1(n_758),
.B2(n_764),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_935),
.B(n_762),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_970),
.A2(n_1050),
.B(n_980),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_927),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1020),
.B(n_464),
.Y(n_1182)
);

NOR2x1_ASAP7_75t_SL g1183 ( 
.A(n_1037),
.B(n_1052),
.Y(n_1183)
);

AO21x1_ASAP7_75t_L g1184 ( 
.A1(n_935),
.A2(n_1044),
.B(n_758),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_949),
.B(n_464),
.Y(n_1185)
);

NAND2x1p5_ASAP7_75t_L g1186 ( 
.A(n_1070),
.B(n_1085),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1108),
.A2(n_1160),
.B(n_1178),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1060),
.A2(n_1175),
.B(n_1083),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_1099),
.B(n_1185),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1178),
.A2(n_1122),
.B(n_1172),
.Y(n_1190)
);

INVx2_ASAP7_75t_R g1191 ( 
.A(n_1070),
.Y(n_1191)
);

INVx8_ASAP7_75t_L g1192 ( 
.A(n_1070),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1176),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1059),
.A2(n_1184),
.B1(n_1161),
.B2(n_1182),
.Y(n_1194)
);

NAND2x1p5_ASAP7_75t_L g1195 ( 
.A(n_1070),
.B(n_1146),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1144),
.Y(n_1196)
);

AOI221xp5_ASAP7_75t_L g1197 ( 
.A1(n_1161),
.A2(n_1168),
.B1(n_1163),
.B2(n_1165),
.C(n_1177),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1168),
.A2(n_1179),
.B(n_1177),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1071),
.A2(n_1111),
.B(n_1081),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1131),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1144),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1157),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1124),
.A2(n_1118),
.B(n_1123),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1145),
.A2(n_1137),
.A3(n_1114),
.B(n_1153),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1142),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1068),
.Y(n_1206)
);

OA21x2_ASAP7_75t_L g1207 ( 
.A1(n_1072),
.A2(n_1079),
.B(n_1080),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1073),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1167),
.B(n_1171),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1142),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1142),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1164),
.A2(n_1179),
.B1(n_1089),
.B2(n_1141),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1135),
.A2(n_1084),
.B1(n_1099),
.B2(n_1089),
.Y(n_1213)
);

BUFx8_ASAP7_75t_L g1214 ( 
.A(n_1069),
.Y(n_1214)
);

INVxp67_ASAP7_75t_SL g1215 ( 
.A(n_1065),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1082),
.B(n_1077),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1082),
.Y(n_1217)
);

CKINVDCx6p67_ASAP7_75t_R g1218 ( 
.A(n_1087),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1167),
.B(n_1171),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1105),
.A2(n_1063),
.B1(n_1088),
.B2(n_1093),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_SL g1221 ( 
.A1(n_1183),
.A2(n_1139),
.B(n_1056),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1109),
.Y(n_1222)
);

AO21x1_ASAP7_75t_L g1223 ( 
.A1(n_1063),
.A2(n_1061),
.B(n_1091),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_SL g1224 ( 
.A1(n_1090),
.A2(n_1086),
.B1(n_1107),
.B2(n_1106),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1095),
.Y(n_1225)
);

AOI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1074),
.A2(n_1078),
.B(n_1064),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_SL g1227 ( 
.A1(n_1103),
.A2(n_1113),
.B(n_1115),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1075),
.B(n_1065),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1149),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1117),
.A2(n_1148),
.B(n_1138),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1167),
.B(n_1171),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1128),
.A2(n_1147),
.B(n_1131),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1116),
.A2(n_1086),
.B1(n_1075),
.B2(n_1150),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1129),
.A2(n_1120),
.B(n_1121),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1129),
.A2(n_1074),
.B(n_1078),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1096),
.Y(n_1236)
);

AO21x2_ASAP7_75t_L g1237 ( 
.A1(n_1097),
.A2(n_1126),
.B(n_1130),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1058),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1151),
.B(n_1154),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_SL g1240 ( 
.A1(n_1169),
.A2(n_1094),
.B(n_1104),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1101),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_1132),
.Y(n_1242)
);

AO21x2_ASAP7_75t_L g1243 ( 
.A1(n_1097),
.A2(n_1126),
.B(n_1112),
.Y(n_1243)
);

NAND3xp33_ASAP7_75t_SL g1244 ( 
.A(n_1102),
.B(n_1125),
.C(n_1134),
.Y(n_1244)
);

NOR2xp67_ASAP7_75t_L g1245 ( 
.A(n_1067),
.B(n_1100),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1119),
.A2(n_1092),
.B1(n_1098),
.B2(n_1136),
.Y(n_1246)
);

AO21x2_ASAP7_75t_L g1247 ( 
.A1(n_1143),
.A2(n_1155),
.B(n_1062),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1127),
.A2(n_1173),
.B(n_1181),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1136),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1173),
.A2(n_1181),
.B(n_1166),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1166),
.A2(n_1066),
.B(n_1152),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1166),
.A2(n_1066),
.B(n_1062),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1156),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1066),
.A2(n_1062),
.B(n_1057),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1158),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1170),
.A2(n_1159),
.B(n_1158),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1133),
.Y(n_1257)
);

NAND2x1p5_ASAP7_75t_L g1258 ( 
.A(n_1133),
.B(n_1162),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1067),
.A2(n_1174),
.B(n_1110),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1133),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1162),
.Y(n_1261)
);

AO21x2_ASAP7_75t_L g1262 ( 
.A1(n_1162),
.A2(n_1108),
.B(n_1140),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1180),
.A2(n_1076),
.B(n_970),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1142),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1144),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1144),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1059),
.A2(n_758),
.B1(n_1041),
.B2(n_588),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1058),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1160),
.A2(n_1172),
.B1(n_893),
.B2(n_1178),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1176),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1144),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1180),
.A2(n_1076),
.B(n_970),
.Y(n_1272)
);

NAND2x1p5_ASAP7_75t_L g1273 ( 
.A(n_1070),
.B(n_1085),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1180),
.A2(n_1076),
.B(n_970),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1144),
.Y(n_1275)
);

O2A1O1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1160),
.A2(n_1178),
.B(n_1122),
.C(n_713),
.Y(n_1276)
);

NAND3xp33_ASAP7_75t_L g1277 ( 
.A(n_1172),
.B(n_893),
.C(n_1160),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1160),
.A2(n_1178),
.B(n_713),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1144),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1059),
.A2(n_758),
.B1(n_1041),
.B2(n_588),
.Y(n_1280)
);

NAND2x1p5_ASAP7_75t_L g1281 ( 
.A(n_1070),
.B(n_1085),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1160),
.A2(n_1172),
.B1(n_893),
.B2(n_1178),
.Y(n_1282)
);

OAI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1172),
.A2(n_1163),
.B1(n_1168),
.B2(n_1165),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1180),
.A2(n_1076),
.B(n_970),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1144),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1070),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1176),
.Y(n_1287)
);

OAI222xp33_ASAP7_75t_L g1288 ( 
.A1(n_1172),
.A2(n_588),
.B1(n_763),
.B2(n_478),
.C1(n_481),
.C2(n_710),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1160),
.A2(n_1172),
.B1(n_893),
.B2(n_1178),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1172),
.A2(n_1163),
.B1(n_1168),
.B2(n_1165),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1142),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1160),
.A2(n_1172),
.B1(n_893),
.B2(n_1178),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1160),
.A2(n_1178),
.B(n_1122),
.C(n_713),
.Y(n_1293)
);

AOI221xp5_ASAP7_75t_L g1294 ( 
.A1(n_1122),
.A2(n_598),
.B1(n_601),
.B2(n_713),
.C(n_641),
.Y(n_1294)
);

NOR2xp67_ASAP7_75t_L g1295 ( 
.A(n_1169),
.B(n_792),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1070),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1180),
.A2(n_1076),
.B(n_970),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1157),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1144),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1108),
.A2(n_1160),
.B(n_1178),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1144),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1084),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1144),
.Y(n_1303)
);

AOI222xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1122),
.A2(n_374),
.B1(n_345),
.B2(n_319),
.C1(n_354),
.C2(n_326),
.Y(n_1304)
);

AO21x1_ASAP7_75t_L g1305 ( 
.A1(n_1108),
.A2(n_1161),
.B(n_1178),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1144),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1144),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_1215),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1228),
.B(n_1197),
.Y(n_1309)
);

AOI221x1_ASAP7_75t_SL g1310 ( 
.A1(n_1283),
.A2(n_1290),
.B1(n_1292),
.B2(n_1282),
.C(n_1289),
.Y(n_1310)
);

OA21x2_ASAP7_75t_L g1311 ( 
.A1(n_1230),
.A2(n_1300),
.B(n_1187),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1305),
.A2(n_1293),
.B(n_1276),
.Y(n_1312)
);

O2A1O1Ixp5_ASAP7_75t_L g1313 ( 
.A1(n_1305),
.A2(n_1269),
.B(n_1223),
.C(n_1290),
.Y(n_1313)
);

OA21x2_ASAP7_75t_L g1314 ( 
.A1(n_1230),
.A2(n_1254),
.B(n_1252),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1283),
.A2(n_1190),
.B(n_1277),
.C(n_1294),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1288),
.A2(n_1220),
.B(n_1213),
.C(n_1198),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1302),
.A2(n_1267),
.B(n_1280),
.C(n_1240),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1216),
.B(n_1242),
.Y(n_1318)
);

OA21x2_ASAP7_75t_L g1319 ( 
.A1(n_1254),
.A2(n_1252),
.B(n_1203),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1203),
.A2(n_1188),
.B(n_1232),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1189),
.B(n_1249),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1196),
.B(n_1201),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1253),
.B(n_1246),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_SL g1324 ( 
.A1(n_1195),
.A2(n_1233),
.B(n_1256),
.Y(n_1324)
);

O2A1O1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1267),
.A2(n_1280),
.B(n_1194),
.C(n_1221),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1194),
.A2(n_1212),
.B1(n_1246),
.B2(n_1224),
.Y(n_1326)
);

NAND2xp33_ASAP7_75t_SL g1327 ( 
.A(n_1238),
.B(n_1268),
.Y(n_1327)
);

O2A1O1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1212),
.A2(n_1227),
.B(n_1244),
.C(n_1225),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1209),
.B(n_1219),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1193),
.A2(n_1270),
.B1(n_1287),
.B2(n_1218),
.Y(n_1330)
);

OA22x2_ASAP7_75t_L g1331 ( 
.A1(n_1209),
.A2(n_1219),
.B1(n_1231),
.B2(n_1255),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1231),
.B(n_1265),
.Y(n_1332)
);

INVx3_ASAP7_75t_SL g1333 ( 
.A(n_1238),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1266),
.B(n_1271),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1206),
.B(n_1208),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1275),
.B(n_1279),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1218),
.A2(n_1202),
.B1(n_1298),
.B2(n_1207),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1202),
.A2(n_1298),
.B1(n_1306),
.B2(n_1303),
.Y(n_1338)
);

O2A1O1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1304),
.A2(n_1262),
.B(n_1257),
.C(n_1261),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1285),
.Y(n_1340)
);

AOI21x1_ASAP7_75t_SL g1341 ( 
.A1(n_1239),
.A2(n_1214),
.B(n_1268),
.Y(n_1341)
);

AOI211xp5_ASAP7_75t_L g1342 ( 
.A1(n_1295),
.A2(n_1307),
.B(n_1301),
.C(n_1299),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_1222),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1260),
.B(n_1229),
.Y(n_1344)
);

AOI221xp5_ASAP7_75t_L g1345 ( 
.A1(n_1262),
.A2(n_1229),
.B1(n_1247),
.B2(n_1192),
.C(n_1259),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1186),
.A2(n_1281),
.B1(n_1273),
.B2(n_1245),
.Y(n_1346)
);

OA22x2_ASAP7_75t_L g1347 ( 
.A1(n_1286),
.A2(n_1296),
.B1(n_1251),
.B2(n_1235),
.Y(n_1347)
);

O2A1O1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1258),
.A2(n_1286),
.B(n_1200),
.C(n_1247),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1258),
.A2(n_1191),
.B(n_1243),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1226),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1214),
.Y(n_1351)
);

O2A1O1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1200),
.A2(n_1243),
.B(n_1236),
.C(n_1241),
.Y(n_1352)
);

NOR2x1_ASAP7_75t_SL g1353 ( 
.A(n_1191),
.B(n_1237),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1204),
.B(n_1250),
.Y(n_1354)
);

O2A1O1Ixp5_ASAP7_75t_L g1355 ( 
.A1(n_1205),
.A2(n_1264),
.B(n_1210),
.C(n_1211),
.Y(n_1355)
);

A2O1A1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1232),
.A2(n_1234),
.B(n_1248),
.C(n_1210),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1248),
.B(n_1234),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1199),
.A2(n_1272),
.B(n_1284),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1264),
.A2(n_1291),
.B(n_1199),
.C(n_1272),
.Y(n_1359)
);

O2A1O1Ixp5_ASAP7_75t_L g1360 ( 
.A1(n_1291),
.A2(n_1263),
.B(n_1274),
.C(n_1284),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1297),
.A2(n_1277),
.B1(n_1160),
.B2(n_1172),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1242),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1216),
.B(n_1217),
.Y(n_1363)
);

O2A1O1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1278),
.A2(n_1269),
.B(n_1289),
.C(n_1282),
.Y(n_1364)
);

AND2x6_ASAP7_75t_L g1365 ( 
.A(n_1239),
.B(n_1209),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1216),
.B(n_1217),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1216),
.B(n_1217),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1216),
.B(n_1217),
.Y(n_1368)
);

CKINVDCx16_ASAP7_75t_R g1369 ( 
.A(n_1202),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1215),
.B(n_1228),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1189),
.B(n_1249),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1216),
.B(n_1217),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1230),
.A2(n_1300),
.B(n_1187),
.Y(n_1373)
);

OA21x2_ASAP7_75t_L g1374 ( 
.A1(n_1230),
.A2(n_1300),
.B(n_1187),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1242),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1242),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1230),
.A2(n_1300),
.B(n_1187),
.Y(n_1377)
);

NOR2x1_ASAP7_75t_SL g1378 ( 
.A(n_1213),
.B(n_1070),
.Y(n_1378)
);

OA21x2_ASAP7_75t_L g1379 ( 
.A1(n_1230),
.A2(n_1300),
.B(n_1187),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1216),
.B(n_1217),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1278),
.A2(n_1160),
.B(n_1178),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1242),
.Y(n_1382)
);

O2A1O1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1278),
.A2(n_1269),
.B(n_1289),
.C(n_1282),
.Y(n_1383)
);

OA21x2_ASAP7_75t_L g1384 ( 
.A1(n_1230),
.A2(n_1300),
.B(n_1187),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1329),
.B(n_1331),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1334),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1329),
.B(n_1332),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1334),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1308),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1335),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1331),
.B(n_1314),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1340),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1313),
.A2(n_1315),
.B(n_1381),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1357),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1365),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1332),
.B(n_1370),
.Y(n_1396)
);

AOI221xp5_ASAP7_75t_L g1397 ( 
.A1(n_1310),
.A2(n_1309),
.B1(n_1383),
.B2(n_1364),
.C(n_1326),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1370),
.B(n_1321),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1319),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1322),
.Y(n_1400)
);

NAND2xp33_ASAP7_75t_SL g1401 ( 
.A(n_1333),
.B(n_1351),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1336),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_1343),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1309),
.B(n_1312),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1350),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1314),
.B(n_1319),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1357),
.B(n_1365),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1371),
.B(n_1362),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1365),
.Y(n_1409)
);

INVxp67_ASAP7_75t_L g1410 ( 
.A(n_1375),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_SL g1411 ( 
.A1(n_1316),
.A2(n_1346),
.B(n_1378),
.Y(n_1411)
);

INVx2_ASAP7_75t_SL g1412 ( 
.A(n_1347),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1376),
.B(n_1382),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1355),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1320),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1318),
.B(n_1363),
.Y(n_1416)
);

OR2x6_ASAP7_75t_L g1417 ( 
.A(n_1349),
.B(n_1348),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1320),
.Y(n_1418)
);

AO21x2_ASAP7_75t_L g1419 ( 
.A1(n_1352),
.A2(n_1354),
.B(n_1312),
.Y(n_1419)
);

AO21x2_ASAP7_75t_L g1420 ( 
.A1(n_1352),
.A2(n_1356),
.B(n_1359),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1347),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1358),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1311),
.B(n_1384),
.Y(n_1423)
);

INVx2_ASAP7_75t_SL g1424 ( 
.A(n_1344),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1365),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1365),
.Y(n_1426)
);

OA21x2_ASAP7_75t_L g1427 ( 
.A1(n_1360),
.A2(n_1345),
.B(n_1361),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1407),
.B(n_1353),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1405),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1404),
.B(n_1384),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1399),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1386),
.B(n_1373),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1386),
.B(n_1373),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1393),
.B(n_1337),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1391),
.B(n_1379),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1399),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1422),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1391),
.B(n_1379),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1391),
.B(n_1385),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1385),
.B(n_1377),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1403),
.Y(n_1441)
);

OR2x2_ASAP7_75t_SL g1442 ( 
.A(n_1427),
.B(n_1369),
.Y(n_1442)
);

AOI21xp33_ASAP7_75t_SL g1443 ( 
.A1(n_1393),
.A2(n_1330),
.B(n_1338),
.Y(n_1443)
);

BUFx3_ASAP7_75t_L g1444 ( 
.A(n_1395),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1385),
.B(n_1377),
.Y(n_1445)
);

NAND2x1p5_ASAP7_75t_L g1446 ( 
.A(n_1427),
.B(n_1374),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1397),
.B(n_1342),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1407),
.B(n_1374),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1407),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1407),
.B(n_1372),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1387),
.B(n_1366),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1405),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1407),
.B(n_1367),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1406),
.Y(n_1454)
);

INVxp67_ASAP7_75t_L g1455 ( 
.A(n_1421),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1406),
.B(n_1368),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1439),
.B(n_1409),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1431),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1447),
.A2(n_1397),
.B(n_1411),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1431),
.Y(n_1460)
);

AO21x2_ASAP7_75t_L g1461 ( 
.A1(n_1430),
.A2(n_1420),
.B(n_1414),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1434),
.A2(n_1412),
.B1(n_1421),
.B2(n_1427),
.Y(n_1462)
);

OAI33xp33_ASAP7_75t_L g1463 ( 
.A1(n_1447),
.A2(n_1410),
.A3(n_1413),
.B1(n_1408),
.B2(n_1400),
.B3(n_1396),
.Y(n_1463)
);

NOR4xp25_ASAP7_75t_SL g1464 ( 
.A(n_1443),
.B(n_1409),
.C(n_1389),
.D(n_1327),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1429),
.Y(n_1465)
);

NAND2xp33_ASAP7_75t_R g1466 ( 
.A(n_1434),
.B(n_1389),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1429),
.Y(n_1467)
);

AOI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1443),
.A2(n_1412),
.B1(n_1317),
.B2(n_1325),
.C(n_1388),
.Y(n_1468)
);

AOI322xp5_ASAP7_75t_L g1469 ( 
.A1(n_1439),
.A2(n_1412),
.A3(n_1323),
.B1(n_1426),
.B2(n_1425),
.C1(n_1345),
.C2(n_1380),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1441),
.B(n_1396),
.Y(n_1470)
);

OAI221xp5_ASAP7_75t_L g1471 ( 
.A1(n_1443),
.A2(n_1427),
.B1(n_1417),
.B2(n_1328),
.C(n_1339),
.Y(n_1471)
);

NAND3xp33_ASAP7_75t_L g1472 ( 
.A(n_1430),
.B(n_1427),
.C(n_1410),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1452),
.Y(n_1473)
);

AOI221xp5_ASAP7_75t_L g1474 ( 
.A1(n_1439),
.A2(n_1388),
.B1(n_1406),
.B2(n_1419),
.C(n_1400),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_R g1475 ( 
.A(n_1441),
.B(n_1401),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1456),
.B(n_1392),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1449),
.B(n_1450),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1451),
.B(n_1403),
.Y(n_1478)
);

NAND3xp33_ASAP7_75t_SL g1479 ( 
.A(n_1446),
.B(n_1413),
.C(n_1392),
.Y(n_1479)
);

AO21x2_ASAP7_75t_L g1480 ( 
.A1(n_1432),
.A2(n_1420),
.B(n_1414),
.Y(n_1480)
);

AOI21xp33_ASAP7_75t_L g1481 ( 
.A1(n_1432),
.A2(n_1417),
.B(n_1419),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1452),
.Y(n_1482)
);

AND2x2_ASAP7_75t_SL g1483 ( 
.A(n_1449),
.B(n_1426),
.Y(n_1483)
);

OAI33xp33_ASAP7_75t_L g1484 ( 
.A1(n_1454),
.A2(n_1408),
.A3(n_1398),
.B1(n_1390),
.B2(n_1416),
.B3(n_1402),
.Y(n_1484)
);

A2O1A1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1440),
.A2(n_1425),
.B(n_1414),
.C(n_1387),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1449),
.B(n_1424),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1446),
.A2(n_1417),
.B(n_1324),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1444),
.B(n_1424),
.Y(n_1488)
);

AOI33xp33_ASAP7_75t_L g1489 ( 
.A1(n_1435),
.A2(n_1390),
.A3(n_1402),
.B1(n_1423),
.B2(n_1424),
.B3(n_1418),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1451),
.B(n_1416),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1428),
.B(n_1394),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1458),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1459),
.B(n_1451),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1483),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1458),
.Y(n_1495)
);

INVx1_ASAP7_75t_SL g1496 ( 
.A(n_1480),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1460),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1477),
.B(n_1440),
.Y(n_1498)
);

BUFx12f_ASAP7_75t_L g1499 ( 
.A(n_1483),
.Y(n_1499)
);

OA21x2_ASAP7_75t_L g1500 ( 
.A1(n_1472),
.A2(n_1415),
.B(n_1418),
.Y(n_1500)
);

INVxp67_ASAP7_75t_L g1501 ( 
.A(n_1472),
.Y(n_1501)
);

OAI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1471),
.A2(n_1446),
.B(n_1455),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1477),
.B(n_1440),
.Y(n_1503)
);

INVxp67_ASAP7_75t_L g1504 ( 
.A(n_1461),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1483),
.B(n_1444),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1465),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1467),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1491),
.B(n_1428),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1467),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1468),
.A2(n_1446),
.B(n_1417),
.Y(n_1510)
);

OA21x2_ASAP7_75t_L g1511 ( 
.A1(n_1481),
.A2(n_1437),
.B(n_1436),
.Y(n_1511)
);

AND2x4_ASAP7_75t_SL g1512 ( 
.A(n_1457),
.B(n_1428),
.Y(n_1512)
);

OA21x2_ASAP7_75t_L g1513 ( 
.A1(n_1474),
.A2(n_1437),
.B(n_1436),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1473),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1473),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1482),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1482),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1501),
.B(n_1490),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1507),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1512),
.B(n_1457),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1500),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1493),
.B(n_1489),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1507),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1509),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1499),
.B(n_1475),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_R g1526 ( 
.A(n_1499),
.B(n_1466),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1512),
.B(n_1464),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1494),
.B(n_1487),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1512),
.B(n_1464),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1501),
.B(n_1490),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1509),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1512),
.B(n_1486),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1512),
.B(n_1486),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1493),
.B(n_1478),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1494),
.B(n_1491),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1501),
.B(n_1445),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1494),
.B(n_1491),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1517),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1517),
.Y(n_1539)
);

OAI33xp33_ASAP7_75t_L g1540 ( 
.A1(n_1504),
.A2(n_1470),
.A3(n_1454),
.B1(n_1476),
.B2(n_1433),
.B3(n_1488),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1506),
.B(n_1485),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1506),
.B(n_1435),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1494),
.B(n_1491),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1499),
.B(n_1450),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1510),
.B(n_1435),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1514),
.B(n_1454),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1510),
.B(n_1438),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1514),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1510),
.B(n_1513),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1499),
.B(n_1450),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1514),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1499),
.A2(n_1442),
.B1(n_1462),
.B2(n_1444),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1515),
.Y(n_1553)
);

NAND4xp25_ASAP7_75t_L g1554 ( 
.A(n_1502),
.B(n_1479),
.C(n_1448),
.D(n_1469),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1505),
.B(n_1453),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1515),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1515),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1505),
.B(n_1453),
.Y(n_1558)
);

INVx6_ASAP7_75t_L g1559 ( 
.A(n_1508),
.Y(n_1559)
);

INVx4_ASAP7_75t_L g1560 ( 
.A(n_1508),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1521),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1534),
.B(n_1498),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1557),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1518),
.B(n_1516),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1518),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1548),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1548),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1551),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1522),
.B(n_1530),
.Y(n_1569)
);

BUFx12f_ASAP7_75t_L g1570 ( 
.A(n_1528),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1544),
.B(n_1550),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1525),
.B(n_1463),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1551),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1521),
.Y(n_1574)
);

AND2x2_ASAP7_75t_SL g1575 ( 
.A(n_1541),
.B(n_1527),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1530),
.B(n_1498),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1519),
.B(n_1498),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1553),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1540),
.B(n_1484),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1553),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1536),
.B(n_1516),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1526),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1544),
.B(n_1498),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1550),
.B(n_1503),
.Y(n_1584)
);

NAND3xp33_ASAP7_75t_L g1585 ( 
.A(n_1554),
.B(n_1502),
.C(n_1513),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1520),
.B(n_1503),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1546),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1556),
.Y(n_1588)
);

INVxp67_ASAP7_75t_SL g1589 ( 
.A(n_1549),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1556),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1519),
.B(n_1503),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1523),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1546),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1552),
.A2(n_1442),
.B1(n_1502),
.B2(n_1513),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1523),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1520),
.B(n_1560),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1571),
.B(n_1565),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1565),
.B(n_1524),
.Y(n_1598)
);

NAND2x1_ASAP7_75t_L g1599 ( 
.A(n_1596),
.B(n_1559),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1571),
.B(n_1527),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1585),
.A2(n_1513),
.B1(n_1547),
.B2(n_1545),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1566),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1582),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1583),
.B(n_1529),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1566),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1583),
.B(n_1584),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1567),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1570),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1579),
.B(n_1524),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1575),
.B(n_1531),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1567),
.Y(n_1611)
);

CKINVDCx16_ASAP7_75t_R g1612 ( 
.A(n_1570),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1568),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1576),
.B(n_1531),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1575),
.A2(n_1513),
.B1(n_1528),
.B2(n_1461),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1589),
.A2(n_1513),
.B1(n_1528),
.B2(n_1461),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1561),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1564),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1564),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1568),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1573),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1597),
.Y(n_1622)
);

NOR2x1p5_ASAP7_75t_L g1623 ( 
.A(n_1599),
.B(n_1569),
.Y(n_1623)
);

AOI32xp33_ASAP7_75t_L g1624 ( 
.A1(n_1601),
.A2(n_1572),
.A3(n_1594),
.B1(n_1528),
.B2(n_1529),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1597),
.B(n_1603),
.Y(n_1625)
);

OAI22xp33_ASAP7_75t_SL g1626 ( 
.A1(n_1609),
.A2(n_1504),
.B1(n_1496),
.B2(n_1559),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1606),
.B(n_1562),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1615),
.A2(n_1513),
.B1(n_1561),
.B2(n_1574),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1600),
.A2(n_1574),
.B1(n_1500),
.B2(n_1480),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1606),
.B(n_1563),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1612),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1616),
.A2(n_1500),
.B1(n_1496),
.B2(n_1504),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1612),
.B(n_1596),
.Y(n_1633)
);

A2O1A1Ixp33_ASAP7_75t_L g1634 ( 
.A1(n_1610),
.A2(n_1469),
.B(n_1496),
.C(n_1581),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1618),
.B(n_1563),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1619),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1600),
.A2(n_1500),
.B1(n_1480),
.B2(n_1584),
.Y(n_1637)
);

AOI32xp33_ASAP7_75t_L g1638 ( 
.A1(n_1604),
.A2(n_1595),
.A3(n_1592),
.B1(n_1593),
.B2(n_1587),
.Y(n_1638)
);

OAI222xp33_ASAP7_75t_L g1639 ( 
.A1(n_1617),
.A2(n_1595),
.B1(n_1592),
.B2(n_1581),
.C1(n_1573),
.C2(n_1590),
.Y(n_1639)
);

AOI322xp5_ASAP7_75t_L g1640 ( 
.A1(n_1608),
.A2(n_1577),
.A3(n_1591),
.B1(n_1593),
.B2(n_1587),
.C1(n_1586),
.C2(n_1542),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1631),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1623),
.B(n_1604),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1625),
.B(n_1598),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1622),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1627),
.B(n_1614),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1630),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1635),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1636),
.Y(n_1648)
);

BUFx2_ASAP7_75t_L g1649 ( 
.A(n_1633),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1628),
.A2(n_1617),
.B1(n_1500),
.B2(n_1511),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1639),
.B(n_1599),
.Y(n_1651)
);

NOR3x1_ASAP7_75t_L g1652 ( 
.A(n_1649),
.B(n_1614),
.C(n_1605),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1649),
.B(n_1639),
.Y(n_1653)
);

OAI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1650),
.A2(n_1624),
.B1(n_1634),
.B2(n_1632),
.C(n_1637),
.Y(n_1654)
);

OAI221xp5_ASAP7_75t_SL g1655 ( 
.A1(n_1651),
.A2(n_1638),
.B1(n_1640),
.B2(n_1629),
.C(n_1617),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1641),
.Y(n_1656)
);

NAND3xp33_ASAP7_75t_SL g1657 ( 
.A(n_1644),
.B(n_1642),
.C(n_1643),
.Y(n_1657)
);

OAI32xp33_ASAP7_75t_L g1658 ( 
.A1(n_1645),
.A2(n_1611),
.A3(n_1621),
.B1(n_1620),
.B2(n_1613),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1648),
.Y(n_1659)
);

AOI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1642),
.A2(n_1626),
.B(n_1621),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1645),
.B(n_1596),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1661),
.B(n_1648),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_SL g1663 ( 
.A(n_1656),
.B(n_1647),
.Y(n_1663)
);

NOR3xp33_ASAP7_75t_L g1664 ( 
.A(n_1657),
.B(n_1647),
.C(n_1648),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1659),
.Y(n_1665)
);

BUFx2_ASAP7_75t_L g1666 ( 
.A(n_1653),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1655),
.A2(n_1646),
.B(n_1620),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1667),
.A2(n_1660),
.B(n_1658),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1662),
.Y(n_1669)
);

NAND3xp33_ASAP7_75t_L g1670 ( 
.A(n_1664),
.B(n_1654),
.C(n_1613),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1663),
.B(n_1602),
.Y(n_1671)
);

AOI221xp5_ASAP7_75t_L g1672 ( 
.A1(n_1666),
.A2(n_1611),
.B1(n_1607),
.B2(n_1605),
.C(n_1602),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1665),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_R g1674 ( 
.A(n_1669),
.B(n_1652),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1668),
.A2(n_1607),
.B(n_1538),
.Y(n_1675)
);

AOI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1670),
.A2(n_1590),
.B1(n_1588),
.B2(n_1578),
.C(n_1580),
.Y(n_1676)
);

OAI21xp33_ASAP7_75t_SL g1677 ( 
.A1(n_1671),
.A2(n_1560),
.B(n_1580),
.Y(n_1677)
);

OAI211xp5_ASAP7_75t_L g1678 ( 
.A1(n_1673),
.A2(n_1560),
.B(n_1588),
.C(n_1578),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1674),
.B(n_1672),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1678),
.Y(n_1680)
);

NAND4xp75_ASAP7_75t_L g1681 ( 
.A(n_1675),
.B(n_1586),
.C(n_1539),
.D(n_1538),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1680),
.B(n_1677),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1682),
.B(n_1681),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1683),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1683),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_SL g1686 ( 
.A1(n_1684),
.A2(n_1679),
.B1(n_1676),
.B2(n_1559),
.Y(n_1686)
);

OAI31xp33_ASAP7_75t_SL g1687 ( 
.A1(n_1685),
.A2(n_1679),
.A3(n_1539),
.B(n_1543),
.Y(n_1687)
);

AOI22x1_ASAP7_75t_L g1688 ( 
.A1(n_1687),
.A2(n_1686),
.B1(n_1535),
.B2(n_1537),
.Y(n_1688)
);

OAI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1687),
.A2(n_1535),
.B(n_1537),
.Y(n_1689)
);

XOR2xp5_ASAP7_75t_L g1690 ( 
.A(n_1688),
.B(n_1341),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_SL g1691 ( 
.A1(n_1690),
.A2(n_1689),
.B1(n_1559),
.B2(n_1500),
.Y(n_1691)
);

AOI322xp5_ASAP7_75t_L g1692 ( 
.A1(n_1691),
.A2(n_1543),
.A3(n_1558),
.B1(n_1555),
.B2(n_1497),
.C1(n_1495),
.C2(n_1492),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_SL g1693 ( 
.A1(n_1692),
.A2(n_1558),
.B1(n_1555),
.B2(n_1532),
.Y(n_1693)
);

AOI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1693),
.A2(n_1533),
.B1(n_1532),
.B2(n_1503),
.Y(n_1694)
);

AOI211xp5_ASAP7_75t_L g1695 ( 
.A1(n_1694),
.A2(n_1516),
.B(n_1533),
.C(n_1495),
.Y(n_1695)
);


endmodule