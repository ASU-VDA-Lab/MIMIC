module fake_aes_10661_n_1197 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_323, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1197);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1197;
wire n_1173;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_667;
wire n_496;
wire n_801;
wire n_988;
wire n_1059;
wire n_1158;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_1196;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_1122;
wire n_779;
wire n_993;
wire n_528;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_1175;
wire n_853;
wire n_1161;
wire n_987;
wire n_1030;
wire n_765;
wire n_1177;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_545;
wire n_896;
wire n_1185;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_1163;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_617;
wire n_384;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_1090;
wire n_1191;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_1194;
wire n_694;
wire n_1179;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_1174;
wire n_1005;
wire n_951;
wire n_702;
wire n_1024;
wire n_1016;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_1097;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_1169;
wire n_652;
wire n_968;
wire n_975;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_955;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_1188;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1011;
wire n_880;
wire n_1101;
wire n_1155;
wire n_630;
wire n_511;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_1180;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_624;
wire n_426;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_1160;
wire n_1184;
wire n_1018;
wire n_1195;
wire n_738;
wire n_979;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_1138;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_399;
wire n_892;
wire n_1171;
wire n_665;
wire n_571;
wire n_1154;
wire n_459;
wire n_863;
wire n_907;
wire n_708;
wire n_1062;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_950;
wire n_1046;
wire n_460;
wire n_1183;
wire n_478;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_1167;
wire n_864;
wire n_1186;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_1157;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_990;
wire n_751;
wire n_800;
wire n_626;
wire n_941;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_1178;
wire n_931;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_1041;
wire n_578;
wire n_926;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_601;
wire n_439;
wire n_996;
wire n_1176;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_1181;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_806;
wire n_881;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_935;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_654;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_1170;
wire n_419;
wire n_1193;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_1125;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_1060;
wire n_1133;
wire n_908;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_1159;
wire n_553;
wire n_440;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_912;
wire n_947;
wire n_1043;
wire n_924;
wire n_378;
wire n_582;
wire n_1141;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_1189;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_1172;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_1165;
wire n_930;
wire n_994;
wire n_1182;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_1168;
wire n_377;
wire n_510;
wire n_343;
wire n_1112;
wire n_1075;
wire n_675;
wire n_967;
wire n_504;
wire n_581;
wire n_458;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_1084;
wire n_722;
wire n_855;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_1164;
wire n_1038;
wire n_341;
wire n_1162;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_695;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_1104;
wire n_1187;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_1190;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1146;
wire n_1108;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_1192;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_1166;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_819;
wire n_772;
wire n_405;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
wire n_1127;
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_217), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_287), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_312), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_276), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_170), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_93), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_12), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_31), .Y(n_331) );
INVx1_ASAP7_75t_SL g332 ( .A(n_199), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_76), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_224), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_120), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_315), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_250), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_252), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_4), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_207), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_271), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_210), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_197), .Y(n_343) );
CKINVDCx16_ASAP7_75t_R g344 ( .A(n_239), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_189), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_184), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_63), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_111), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_221), .Y(n_349) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_151), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_169), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_99), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_24), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_28), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_139), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_3), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_62), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g358 ( .A(n_82), .Y(n_358) );
INVxp67_ASAP7_75t_L g359 ( .A(n_268), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_302), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_43), .Y(n_361) );
CKINVDCx14_ASAP7_75t_R g362 ( .A(n_55), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_172), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_108), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_57), .Y(n_365) );
INVx2_ASAP7_75t_SL g366 ( .A(n_35), .Y(n_366) );
BUFx3_ASAP7_75t_L g367 ( .A(n_218), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_19), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_237), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_232), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_164), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_192), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_103), .Y(n_373) );
CKINVDCx14_ASAP7_75t_R g374 ( .A(n_292), .Y(n_374) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_149), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_262), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_1), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_34), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_49), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_242), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_240), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_307), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_1), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_129), .Y(n_384) );
BUFx10_ASAP7_75t_L g385 ( .A(n_201), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_215), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_125), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_267), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_320), .Y(n_389) );
INVx1_ASAP7_75t_SL g390 ( .A(n_304), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_40), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_233), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_167), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_305), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_114), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_92), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_38), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_162), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_37), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_275), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_191), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_195), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_182), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_15), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_288), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_264), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_256), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_298), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_16), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_41), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_126), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_319), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_244), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_253), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_0), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_72), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_67), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_112), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_249), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_209), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_251), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_246), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_281), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_318), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_91), .Y(n_425) );
CKINVDCx16_ASAP7_75t_R g426 ( .A(n_80), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_285), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_22), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_277), .Y(n_429) );
CKINVDCx14_ASAP7_75t_R g430 ( .A(n_113), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_30), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_133), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_20), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_15), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_241), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_140), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_158), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_238), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_86), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_212), .Y(n_440) );
INVx2_ASAP7_75t_SL g441 ( .A(n_127), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_21), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_142), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_282), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_200), .Y(n_445) );
BUFx3_ASAP7_75t_L g446 ( .A(n_299), .Y(n_446) );
INVxp33_ASAP7_75t_L g447 ( .A(n_118), .Y(n_447) );
BUFx5_ASAP7_75t_L g448 ( .A(n_110), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_313), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_115), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_309), .Y(n_451) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_296), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_10), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_42), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_10), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_2), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_81), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_5), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_20), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_109), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_31), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_243), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_168), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_254), .Y(n_464) );
NOR2xp67_ASAP7_75t_L g465 ( .A(n_79), .B(n_32), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_136), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_202), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_248), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_51), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_216), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_117), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_266), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_152), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_247), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_124), .Y(n_475) );
INVx1_ASAP7_75t_SL g476 ( .A(n_231), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_303), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_190), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_301), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_132), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_179), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_321), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_150), .Y(n_483) );
CKINVDCx16_ASAP7_75t_R g484 ( .A(n_116), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_211), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_188), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_235), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_213), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_270), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_47), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_121), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_73), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_185), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_348), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_370), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_344), .A2(n_3), .B1(n_0), .B2(n_2), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_438), .B(n_4), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_348), .Y(n_498) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_330), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_366), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_433), .B(n_5), .Y(n_501) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_360), .Y(n_502) );
AND2x6_ASAP7_75t_L g503 ( .A(n_363), .B(n_44), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_436), .B(n_6), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_350), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_448), .Y(n_506) );
OA21x2_ASAP7_75t_L g507 ( .A1(n_333), .A2(n_46), .B(n_45), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_339), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_441), .B(n_6), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_358), .A2(n_9), .B1(n_7), .B2(n_8), .Y(n_510) );
INVx4_ASAP7_75t_L g511 ( .A(n_324), .Y(n_511) );
INVx2_ASAP7_75t_SL g512 ( .A(n_385), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_426), .A2(n_484), .B1(n_368), .B2(n_397), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_448), .Y(n_514) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_360), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_391), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_399), .B(n_7), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_364), .A2(n_11), .B1(n_8), .B2(n_9), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_410), .B(n_11), .Y(n_519) );
INVx5_ASAP7_75t_L g520 ( .A(n_385), .Y(n_520) );
BUFx2_ASAP7_75t_L g521 ( .A(n_331), .Y(n_521) );
INVx5_ASAP7_75t_L g522 ( .A(n_360), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_415), .Y(n_523) );
BUFx12f_ASAP7_75t_L g524 ( .A(n_353), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_431), .Y(n_525) );
INVx1_ASAP7_75t_SL g526 ( .A(n_521), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_499), .B(n_434), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_506), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_514), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_515), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_515), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_501), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_501), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_511), .B(n_447), .Y(n_534) );
NAND2xp33_ASAP7_75t_L g535 ( .A(n_503), .B(n_448), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_495), .B(n_447), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_499), .B(n_362), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_500), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_494), .Y(n_539) );
BUFx2_ASAP7_75t_L g540 ( .A(n_524), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_515), .Y(n_541) );
INVx3_ASAP7_75t_L g542 ( .A(n_498), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_504), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_504), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_509), .B(n_448), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_509), .B(n_448), .Y(n_546) );
AOI21x1_ASAP7_75t_L g547 ( .A1(n_507), .A2(n_336), .B(n_334), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_508), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_511), .B(n_359), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_515), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_516), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_523), .Y(n_552) );
O2A1O1Ixp5_ASAP7_75t_L g553 ( .A1(n_545), .A2(n_497), .B(n_452), .C(n_517), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_543), .B(n_520), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_526), .B(n_505), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_544), .B(n_513), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_528), .B(n_337), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_534), .B(n_520), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_528), .B(n_340), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_536), .B(n_520), .Y(n_560) );
INVxp67_ASAP7_75t_L g561 ( .A(n_537), .Y(n_561) );
BUFx3_ASAP7_75t_L g562 ( .A(n_529), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_536), .B(n_520), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_542), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_538), .Y(n_565) );
CKINVDCx11_ASAP7_75t_R g566 ( .A(n_540), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_542), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_548), .B(n_512), .Y(n_568) );
INVxp67_ASAP7_75t_L g569 ( .A(n_549), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_549), .B(n_525), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_529), .B(n_341), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_551), .B(n_345), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_532), .A2(n_510), .B1(n_518), .B2(n_496), .Y(n_573) );
NOR2xp67_ASAP7_75t_L g574 ( .A(n_527), .B(n_510), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_539), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_552), .B(n_347), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_533), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_535), .A2(n_503), .B1(n_519), .B2(n_517), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_545), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_546), .B(n_355), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_546), .Y(n_581) );
BUFx3_ASAP7_75t_L g582 ( .A(n_530), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_535), .A2(n_503), .B1(n_519), .B2(n_454), .Y(n_583) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_547), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_531), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_531), .B(n_503), .Y(n_586) );
INVx3_ASAP7_75t_L g587 ( .A(n_541), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_541), .B(n_518), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_550), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_550), .Y(n_590) );
CKINVDCx6p67_ASAP7_75t_R g591 ( .A(n_540), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_543), .A2(n_445), .B1(n_475), .B2(n_395), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_543), .B(n_357), .Y(n_593) );
NOR2xp67_ASAP7_75t_L g594 ( .A(n_555), .B(n_12), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_578), .A2(n_507), .B(n_452), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_570), .B(n_354), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_562), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_574), .A2(n_374), .B1(n_430), .B2(n_453), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_578), .A2(n_369), .B(n_365), .Y(n_599) );
AND2x2_ASAP7_75t_SL g600 ( .A(n_592), .B(n_455), .Y(n_600) );
OR2x6_ASAP7_75t_L g601 ( .A(n_561), .B(n_456), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_570), .B(n_356), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_569), .B(n_325), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_556), .B(n_377), .Y(n_604) );
A2O1A1Ixp33_ASAP7_75t_L g605 ( .A1(n_553), .A2(n_459), .B(n_465), .C(n_386), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_577), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_573), .A2(n_430), .B1(n_374), .B2(n_383), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_583), .A2(n_404), .B1(n_409), .B2(n_378), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_593), .B(n_428), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_586), .A2(n_387), .B(n_382), .Y(n_610) );
A2O1A1Ixp33_ASAP7_75t_L g611 ( .A1(n_581), .A2(n_393), .B(n_394), .C(n_392), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_583), .B(n_326), .Y(n_612) );
INVxp67_ASAP7_75t_L g613 ( .A(n_554), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_580), .A2(n_401), .B(n_398), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_565), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_588), .A2(n_458), .B1(n_461), .B2(n_442), .Y(n_616) );
INVx3_ASAP7_75t_L g617 ( .A(n_591), .Y(n_617) );
AO21x1_ASAP7_75t_L g618 ( .A1(n_580), .A2(n_417), .B(n_412), .Y(n_618) );
INVxp67_ASAP7_75t_SL g619 ( .A(n_575), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_560), .A2(n_420), .B(n_419), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_563), .B(n_328), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_579), .A2(n_427), .B(n_421), .Y(n_622) );
AO21x1_ASAP7_75t_L g623 ( .A1(n_557), .A2(n_435), .B(n_429), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_558), .A2(n_444), .B(n_443), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g625 ( .A1(n_572), .A2(n_451), .B(n_450), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_568), .B(n_329), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_584), .A2(n_473), .B(n_471), .Y(n_627) );
INVx3_ASAP7_75t_L g628 ( .A(n_564), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_572), .A2(n_480), .B1(n_481), .B2(n_478), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_584), .A2(n_576), .B(n_559), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_567), .B(n_335), .Y(n_631) );
O2A1O1Ixp33_ASAP7_75t_L g632 ( .A1(n_576), .A2(n_489), .B(n_491), .C(n_482), .Y(n_632) );
INVx2_ASAP7_75t_SL g633 ( .A(n_557), .Y(n_633) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_584), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_L g635 ( .A1(n_559), .A2(n_332), .B(n_472), .C(n_390), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_571), .B(n_338), .Y(n_636) );
INVx3_ASAP7_75t_L g637 ( .A(n_582), .Y(n_637) );
AO32x1_ASAP7_75t_L g638 ( .A1(n_584), .A2(n_414), .A3(n_423), .B1(n_372), .B2(n_327), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_585), .A2(n_432), .B(n_425), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_615), .B(n_566), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_619), .A2(n_476), .B1(n_343), .B2(n_346), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_630), .A2(n_590), .B(n_589), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_596), .B(n_342), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_604), .B(n_582), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_606), .Y(n_645) );
NOR2x1_ASAP7_75t_SL g646 ( .A(n_601), .B(n_363), .Y(n_646) );
NAND2xp33_ASAP7_75t_L g647 ( .A(n_634), .B(n_448), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_595), .A2(n_587), .B(n_449), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_602), .A2(n_351), .B1(n_352), .B2(n_349), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_633), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_617), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_597), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_613), .B(n_361), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_600), .B(n_13), .Y(n_654) );
NOR2x1_ASAP7_75t_SL g655 ( .A(n_598), .B(n_367), .Y(n_655) );
OAI21x1_ASAP7_75t_L g656 ( .A1(n_627), .A2(n_375), .B(n_360), .Y(n_656) );
AO31x2_ASAP7_75t_L g657 ( .A1(n_618), .A2(n_502), .A3(n_375), .B(n_522), .Y(n_657) );
A2O1A1Ixp33_ASAP7_75t_L g658 ( .A1(n_599), .A2(n_446), .B(n_367), .C(n_375), .Y(n_658) );
NOR2xp33_ASAP7_75t_SL g659 ( .A(n_634), .B(n_371), .Y(n_659) );
OAI21xp5_ASAP7_75t_L g660 ( .A1(n_605), .A2(n_446), .B(n_376), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_628), .Y(n_661) );
NOR2x1_ASAP7_75t_L g662 ( .A(n_594), .B(n_502), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_616), .B(n_373), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_628), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_626), .B(n_13), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_609), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_622), .B(n_379), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_611), .B(n_380), .Y(n_668) );
AOI21x1_ASAP7_75t_SL g669 ( .A1(n_621), .A2(n_522), .B(n_384), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_612), .A2(n_388), .B(n_381), .Y(n_670) );
AOI21x1_ASAP7_75t_SL g671 ( .A1(n_636), .A2(n_522), .B(n_396), .Y(n_671) );
OAI21x1_ASAP7_75t_SL g672 ( .A1(n_623), .A2(n_14), .B(n_16), .Y(n_672) );
CKINVDCx8_ASAP7_75t_R g673 ( .A(n_634), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_625), .B(n_607), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_608), .B(n_14), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_610), .A2(n_400), .B(n_389), .Y(n_676) );
AOI31xp67_ASAP7_75t_L g677 ( .A1(n_638), .A2(n_502), .A3(n_522), .B(n_50), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_629), .B(n_603), .Y(n_678) );
OAI22x1_ASAP7_75t_L g679 ( .A1(n_631), .A2(n_403), .B1(n_405), .B2(n_402), .Y(n_679) );
OAI21x1_ASAP7_75t_L g680 ( .A1(n_637), .A2(n_52), .B(n_48), .Y(n_680) );
OAI21xp33_ASAP7_75t_L g681 ( .A1(n_620), .A2(n_407), .B(n_406), .Y(n_681) );
AO21x2_ASAP7_75t_L g682 ( .A1(n_638), .A2(n_54), .B(n_53), .Y(n_682) );
AO21x1_ASAP7_75t_L g683 ( .A1(n_624), .A2(n_639), .B(n_635), .Y(n_683) );
INVx5_ASAP7_75t_L g684 ( .A(n_632), .Y(n_684) );
BUFx2_ASAP7_75t_L g685 ( .A(n_614), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_594), .B(n_408), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_615), .B(n_411), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_615), .B(n_413), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_604), .B(n_493), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_615), .Y(n_690) );
AND2x4_ASAP7_75t_L g691 ( .A(n_690), .B(n_17), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_640), .B(n_416), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_666), .B(n_17), .Y(n_693) );
OAI21xp5_ASAP7_75t_L g694 ( .A1(n_674), .A2(n_422), .B(n_418), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_645), .Y(n_695) );
OA21x2_ASAP7_75t_L g696 ( .A1(n_648), .A2(n_437), .B(n_424), .Y(n_696) );
OAI21x1_ASAP7_75t_L g697 ( .A1(n_671), .A2(n_58), .B(n_56), .Y(n_697) );
OR2x2_ASAP7_75t_L g698 ( .A(n_654), .B(n_18), .Y(n_698) );
OA21x2_ASAP7_75t_L g699 ( .A1(n_680), .A2(n_440), .B(n_439), .Y(n_699) );
AO21x2_ASAP7_75t_L g700 ( .A1(n_682), .A2(n_60), .B(n_59), .Y(n_700) );
CKINVDCx8_ASAP7_75t_R g701 ( .A(n_684), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_652), .Y(n_702) );
OA21x2_ASAP7_75t_L g703 ( .A1(n_658), .A2(n_460), .B(n_457), .Y(n_703) );
OAI21x1_ASAP7_75t_L g704 ( .A1(n_669), .A2(n_64), .B(n_61), .Y(n_704) );
AO21x2_ASAP7_75t_L g705 ( .A1(n_682), .A2(n_66), .B(n_65), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g706 ( .A(n_660), .B(n_463), .C(n_462), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_685), .Y(n_707) );
OAI21x1_ASAP7_75t_L g708 ( .A1(n_656), .A2(n_69), .B(n_68), .Y(n_708) );
OAI21xp5_ASAP7_75t_L g709 ( .A1(n_678), .A2(n_466), .B(n_464), .Y(n_709) );
OAI21x1_ASAP7_75t_L g710 ( .A1(n_642), .A2(n_71), .B(n_70), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_675), .A2(n_468), .B1(n_469), .B2(n_467), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_661), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_664), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_689), .B(n_470), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_663), .B(n_474), .Y(n_715) );
AO21x2_ASAP7_75t_L g716 ( .A1(n_655), .A2(n_75), .B(n_74), .Y(n_716) );
INVx4_ASAP7_75t_L g717 ( .A(n_684), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_650), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_672), .Y(n_719) );
OAI21x1_ASAP7_75t_L g720 ( .A1(n_662), .A2(n_78), .B(n_77), .Y(n_720) );
BUFx2_ASAP7_75t_L g721 ( .A(n_651), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_665), .B(n_21), .Y(n_722) );
BUFx2_ASAP7_75t_L g723 ( .A(n_679), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g724 ( .A1(n_644), .A2(n_479), .B(n_477), .Y(n_724) );
OAI21xp5_ASAP7_75t_L g725 ( .A1(n_667), .A2(n_485), .B(n_483), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_684), .A2(n_492), .B1(n_490), .B2(n_488), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_657), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_653), .B(n_23), .Y(n_728) );
AOI21x1_ASAP7_75t_L g729 ( .A1(n_686), .A2(n_487), .B(n_486), .Y(n_729) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_659), .A2(n_23), .B1(n_24), .B2(n_25), .Y(n_730) );
AO21x2_ASAP7_75t_L g731 ( .A1(n_683), .A2(n_84), .B(n_83), .Y(n_731) );
O2A1O1Ixp33_ASAP7_75t_L g732 ( .A1(n_643), .A2(n_25), .B(n_26), .C(n_27), .Y(n_732) );
CKINVDCx5p33_ASAP7_75t_R g733 ( .A(n_641), .Y(n_733) );
OR2x2_ASAP7_75t_L g734 ( .A(n_687), .B(n_26), .Y(n_734) );
OR2x2_ASAP7_75t_L g735 ( .A(n_688), .B(n_27), .Y(n_735) );
INVx5_ASAP7_75t_L g736 ( .A(n_673), .Y(n_736) );
AO222x2_ASAP7_75t_L g737 ( .A1(n_649), .A2(n_28), .B1(n_29), .B2(n_30), .C1(n_32), .C2(n_33), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_657), .Y(n_738) );
BUFx10_ASAP7_75t_L g739 ( .A(n_659), .Y(n_739) );
AO21x2_ASAP7_75t_L g740 ( .A1(n_647), .A2(n_87), .B(n_85), .Y(n_740) );
AND2x4_ASAP7_75t_L g741 ( .A(n_668), .B(n_29), .Y(n_741) );
OA21x2_ASAP7_75t_L g742 ( .A1(n_677), .A2(n_89), .B(n_88), .Y(n_742) );
NAND2x1p5_ASAP7_75t_L g743 ( .A(n_676), .B(n_33), .Y(n_743) );
NOR2x1_ASAP7_75t_SL g744 ( .A(n_681), .B(n_90), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_670), .Y(n_745) );
OAI21x1_ASAP7_75t_SL g746 ( .A1(n_646), .A2(n_35), .B(n_36), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_690), .Y(n_747) );
OR2x2_ASAP7_75t_L g748 ( .A(n_640), .B(n_36), .Y(n_748) );
A2O1A1Ixp33_ASAP7_75t_L g749 ( .A1(n_674), .A2(n_37), .B(n_38), .C(n_39), .Y(n_749) );
NAND3xp33_ASAP7_75t_L g750 ( .A(n_658), .B(n_39), .C(n_40), .Y(n_750) );
AND2x4_ASAP7_75t_L g751 ( .A(n_690), .B(n_41), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_695), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_695), .Y(n_753) );
INVx3_ASAP7_75t_L g754 ( .A(n_736), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_698), .B(n_691), .Y(n_755) );
INVx1_ASAP7_75t_SL g756 ( .A(n_739), .Y(n_756) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_707), .Y(n_757) );
INVx5_ASAP7_75t_L g758 ( .A(n_736), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_702), .Y(n_759) );
INVx4_ASAP7_75t_L g760 ( .A(n_736), .Y(n_760) );
INVx3_ASAP7_75t_L g761 ( .A(n_701), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_691), .B(n_42), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_751), .B(n_94), .Y(n_763) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_707), .Y(n_764) );
AND2x4_ASAP7_75t_L g765 ( .A(n_751), .B(n_95), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g766 ( .A(n_721), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_712), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_713), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_713), .Y(n_769) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_738), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_718), .Y(n_771) );
OAI21x1_ASAP7_75t_L g772 ( .A1(n_697), .A2(n_96), .B(n_97), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_693), .Y(n_773) );
BUFx3_ASAP7_75t_L g774 ( .A(n_739), .Y(n_774) );
AND2x2_ASAP7_75t_L g775 ( .A(n_733), .B(n_98), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_748), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_734), .Y(n_777) );
INVx3_ASAP7_75t_L g778 ( .A(n_717), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_735), .Y(n_779) );
OAI21x1_ASAP7_75t_L g780 ( .A1(n_704), .A2(n_100), .B(n_101), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_728), .B(n_102), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_741), .B(n_104), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_741), .B(n_105), .Y(n_783) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_727), .Y(n_784) );
OA21x2_ASAP7_75t_L g785 ( .A1(n_719), .A2(n_106), .B(n_107), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_711), .B(n_119), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_723), .A2(n_122), .B1(n_123), .B2(n_128), .Y(n_787) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_717), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_746), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_722), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_719), .Y(n_791) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_699), .Y(n_792) );
BUFx3_ASAP7_75t_L g793 ( .A(n_743), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_749), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_732), .Y(n_795) );
BUFx2_ASAP7_75t_SL g796 ( .A(n_737), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_745), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_692), .B(n_130), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_745), .Y(n_799) );
AND2x2_ASAP7_75t_L g800 ( .A(n_730), .B(n_131), .Y(n_800) );
INVx3_ASAP7_75t_L g801 ( .A(n_716), .Y(n_801) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_699), .Y(n_802) );
INVx1_ASAP7_75t_SL g803 ( .A(n_703), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_729), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_720), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_715), .B(n_134), .Y(n_806) );
INVx5_ASAP7_75t_L g807 ( .A(n_744), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_724), .B(n_135), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_694), .B(n_137), .Y(n_809) );
AOI21x1_ASAP7_75t_L g810 ( .A1(n_742), .A2(n_323), .B(n_141), .Y(n_810) );
AO21x2_ASAP7_75t_L g811 ( .A1(n_744), .A2(n_138), .B(n_143), .Y(n_811) );
A2O1A1Ixp33_ASAP7_75t_L g812 ( .A1(n_750), .A2(n_144), .B(n_145), .C(n_146), .Y(n_812) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_731), .Y(n_813) );
INVx3_ASAP7_75t_L g814 ( .A(n_740), .Y(n_814) );
O2A1O1Ixp33_ASAP7_75t_L g815 ( .A1(n_709), .A2(n_147), .B(n_148), .C(n_153), .Y(n_815) );
OA21x2_ASAP7_75t_L g816 ( .A1(n_710), .A2(n_154), .B(n_155), .Y(n_816) );
INVx2_ASAP7_75t_SL g817 ( .A(n_696), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_706), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_714), .B(n_156), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_708), .Y(n_820) );
BUFx3_ASAP7_75t_L g821 ( .A(n_726), .Y(n_821) );
INVx2_ASAP7_75t_L g822 ( .A(n_700), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_700), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_725), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_705), .Y(n_825) );
OR2x2_ASAP7_75t_L g826 ( .A(n_742), .B(n_322), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_747), .Y(n_827) );
OAI21x1_ASAP7_75t_L g828 ( .A1(n_697), .A2(n_157), .B(n_159), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_737), .B(n_160), .Y(n_829) );
NAND2xp33_ASAP7_75t_R g830 ( .A(n_699), .B(n_161), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_695), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_695), .Y(n_832) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_707), .Y(n_833) );
INVx2_ASAP7_75t_L g834 ( .A(n_695), .Y(n_834) );
NAND2xp33_ASAP7_75t_R g835 ( .A(n_699), .B(n_163), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_695), .Y(n_836) );
INVx3_ASAP7_75t_L g837 ( .A(n_736), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_695), .Y(n_838) );
NOR2x1p5_ASAP7_75t_L g839 ( .A(n_760), .B(n_165), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_755), .B(n_166), .Y(n_840) );
BUFx2_ASAP7_75t_L g841 ( .A(n_788), .Y(n_841) );
HB1xp67_ASAP7_75t_L g842 ( .A(n_784), .Y(n_842) );
AND2x2_ASAP7_75t_L g843 ( .A(n_762), .B(n_171), .Y(n_843) );
AND2x2_ASAP7_75t_L g844 ( .A(n_776), .B(n_173), .Y(n_844) );
AND2x2_ASAP7_75t_L g845 ( .A(n_777), .B(n_174), .Y(n_845) );
INVx5_ASAP7_75t_L g846 ( .A(n_758), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_759), .Y(n_847) );
INVx2_ASAP7_75t_L g848 ( .A(n_827), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_752), .Y(n_849) );
BUFx2_ASAP7_75t_L g850 ( .A(n_778), .Y(n_850) );
AND2x2_ASAP7_75t_L g851 ( .A(n_779), .B(n_175), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_753), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_838), .Y(n_853) );
BUFx2_ASAP7_75t_L g854 ( .A(n_778), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_771), .B(n_176), .Y(n_855) );
INVx3_ASAP7_75t_L g856 ( .A(n_758), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_829), .B(n_177), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_834), .B(n_178), .Y(n_858) );
INVx2_ASAP7_75t_L g859 ( .A(n_797), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_831), .Y(n_860) );
INVx2_ASAP7_75t_L g861 ( .A(n_799), .Y(n_861) );
INVx2_ASAP7_75t_L g862 ( .A(n_791), .Y(n_862) );
INVx2_ASAP7_75t_L g863 ( .A(n_770), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_832), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_836), .Y(n_865) );
AND2x4_ASAP7_75t_L g866 ( .A(n_765), .B(n_180), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_829), .B(n_181), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_767), .Y(n_868) );
AND2x4_ASAP7_75t_SL g869 ( .A(n_765), .B(n_183), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_770), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_775), .B(n_186), .Y(n_871) );
INVx5_ASAP7_75t_L g872 ( .A(n_758), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_768), .Y(n_873) );
NOR2xp33_ASAP7_75t_L g874 ( .A(n_796), .B(n_187), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_769), .Y(n_875) );
AND2x4_ASAP7_75t_L g876 ( .A(n_757), .B(n_193), .Y(n_876) );
HB1xp67_ASAP7_75t_L g877 ( .A(n_784), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_790), .B(n_194), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_757), .Y(n_879) );
NOR2xp33_ASAP7_75t_L g880 ( .A(n_824), .B(n_196), .Y(n_880) );
INVxp67_ASAP7_75t_SL g881 ( .A(n_764), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_764), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_763), .B(n_782), .Y(n_883) );
OR2x2_ASAP7_75t_L g884 ( .A(n_833), .B(n_198), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_820), .Y(n_885) );
INVx2_ASAP7_75t_L g886 ( .A(n_833), .Y(n_886) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_792), .Y(n_887) );
OR2x2_ASAP7_75t_L g888 ( .A(n_756), .B(n_203), .Y(n_888) );
INVx2_ASAP7_75t_L g889 ( .A(n_773), .Y(n_889) );
HB1xp67_ASAP7_75t_L g890 ( .A(n_792), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_774), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_783), .B(n_204), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_774), .Y(n_893) );
INVx3_ASAP7_75t_L g894 ( .A(n_758), .Y(n_894) );
AND2x2_ASAP7_75t_L g895 ( .A(n_756), .B(n_781), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_761), .B(n_205), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_794), .B(n_206), .Y(n_897) );
BUFx6f_ASAP7_75t_L g898 ( .A(n_793), .Y(n_898) );
BUFx2_ASAP7_75t_L g899 ( .A(n_760), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_793), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_789), .Y(n_901) );
INVx3_ASAP7_75t_L g902 ( .A(n_754), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_804), .Y(n_903) );
BUFx2_ASAP7_75t_L g904 ( .A(n_754), .Y(n_904) );
NOR2xp67_ASAP7_75t_L g905 ( .A(n_837), .B(n_208), .Y(n_905) );
INVx2_ASAP7_75t_L g906 ( .A(n_823), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_821), .B(n_214), .Y(n_907) );
NAND2x1p5_ASAP7_75t_L g908 ( .A(n_837), .B(n_219), .Y(n_908) );
INVxp67_ASAP7_75t_SL g909 ( .A(n_802), .Y(n_909) );
INVxp67_ASAP7_75t_SL g910 ( .A(n_802), .Y(n_910) );
BUFx2_ASAP7_75t_L g911 ( .A(n_766), .Y(n_911) );
INVx4_ASAP7_75t_L g912 ( .A(n_766), .Y(n_912) );
INVx2_ASAP7_75t_L g913 ( .A(n_822), .Y(n_913) );
AND2x2_ASAP7_75t_L g914 ( .A(n_821), .B(n_220), .Y(n_914) );
AND2x4_ASAP7_75t_L g915 ( .A(n_807), .B(n_222), .Y(n_915) );
INVx2_ASAP7_75t_L g916 ( .A(n_825), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_795), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_818), .B(n_223), .Y(n_918) );
INVx2_ASAP7_75t_L g919 ( .A(n_805), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_808), .B(n_225), .Y(n_920) );
INVxp67_ASAP7_75t_L g921 ( .A(n_817), .Y(n_921) );
AND2x4_ASAP7_75t_L g922 ( .A(n_807), .B(n_226), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_798), .B(n_227), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_824), .A2(n_228), .B1(n_229), .B2(n_230), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_800), .B(n_234), .Y(n_925) );
AND2x2_ASAP7_75t_L g926 ( .A(n_786), .B(n_236), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_801), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_806), .B(n_245), .Y(n_928) );
INVx3_ASAP7_75t_L g929 ( .A(n_807), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_809), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_809), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_803), .Y(n_932) );
INVxp67_ASAP7_75t_L g933 ( .A(n_830), .Y(n_933) );
INVx2_ASAP7_75t_L g934 ( .A(n_807), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_806), .B(n_255), .Y(n_935) );
OR2x2_ASAP7_75t_L g936 ( .A(n_819), .B(n_257), .Y(n_936) );
AND2x2_ASAP7_75t_L g937 ( .A(n_819), .B(n_258), .Y(n_937) );
INVx2_ASAP7_75t_L g938 ( .A(n_814), .Y(n_938) );
HB1xp67_ASAP7_75t_L g939 ( .A(n_830), .Y(n_939) );
INVxp67_ASAP7_75t_SL g940 ( .A(n_835), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_787), .B(n_259), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_903), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_889), .B(n_787), .Y(n_943) );
INVxp67_ASAP7_75t_SL g944 ( .A(n_842), .Y(n_944) );
NOR2xp67_ASAP7_75t_L g945 ( .A(n_846), .B(n_872), .Y(n_945) );
OR2x2_ASAP7_75t_L g946 ( .A(n_841), .B(n_879), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_895), .B(n_813), .Y(n_947) );
INVxp67_ASAP7_75t_SL g948 ( .A(n_842), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_875), .B(n_814), .Y(n_949) );
BUFx2_ASAP7_75t_L g950 ( .A(n_899), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_849), .B(n_785), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_850), .B(n_854), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_883), .B(n_811), .Y(n_953) );
OR2x2_ASAP7_75t_L g954 ( .A(n_886), .B(n_826), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_852), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_853), .B(n_812), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_848), .B(n_811), .Y(n_957) );
AND2x4_ASAP7_75t_L g958 ( .A(n_881), .B(n_812), .Y(n_958) );
OR2x2_ASAP7_75t_L g959 ( .A(n_886), .B(n_816), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_881), .B(n_816), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_860), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_864), .Y(n_962) );
BUFx2_ASAP7_75t_L g963 ( .A(n_898), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_865), .B(n_815), .Y(n_964) );
OR2x2_ASAP7_75t_L g965 ( .A(n_882), .B(n_828), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_868), .B(n_815), .Y(n_966) );
OR2x2_ASAP7_75t_L g967 ( .A(n_877), .B(n_780), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_873), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_847), .Y(n_969) );
OR2x2_ASAP7_75t_L g970 ( .A(n_877), .B(n_772), .Y(n_970) );
AND2x2_ASAP7_75t_L g971 ( .A(n_891), .B(n_810), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_917), .B(n_835), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_893), .B(n_260), .Y(n_973) );
AOI21xp5_ASAP7_75t_SL g974 ( .A1(n_866), .A2(n_261), .B(n_263), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_862), .Y(n_975) );
AND2x4_ASAP7_75t_SL g976 ( .A(n_912), .B(n_265), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_862), .Y(n_977) );
INVxp67_ASAP7_75t_SL g978 ( .A(n_921), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_930), .B(n_269), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_863), .Y(n_980) );
INVxp67_ASAP7_75t_L g981 ( .A(n_911), .Y(n_981) );
NAND2xp33_ASAP7_75t_SL g982 ( .A(n_839), .B(n_272), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_863), .Y(n_983) );
HB1xp67_ASAP7_75t_L g984 ( .A(n_904), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_870), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_900), .B(n_273), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_870), .Y(n_987) );
AOI221xp5_ASAP7_75t_L g988 ( .A1(n_874), .A2(n_274), .B1(n_278), .B2(n_279), .C(n_280), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_840), .B(n_283), .Y(n_989) );
INVx3_ASAP7_75t_L g990 ( .A(n_929), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_931), .B(n_284), .Y(n_991) );
HB1xp67_ASAP7_75t_L g992 ( .A(n_876), .Y(n_992) );
NOR2xp33_ASAP7_75t_L g993 ( .A(n_912), .B(n_286), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_907), .B(n_289), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_914), .B(n_290), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_859), .B(n_291), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_861), .B(n_293), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_861), .B(n_294), .Y(n_998) );
CKINVDCx20_ASAP7_75t_R g999 ( .A(n_874), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_901), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_857), .B(n_295), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_867), .B(n_297), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_884), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_876), .B(n_300), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_902), .B(n_306), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_887), .Y(n_1006) );
INVx3_ASAP7_75t_L g1007 ( .A(n_929), .Y(n_1007) );
OR2x2_ASAP7_75t_L g1008 ( .A(n_887), .B(n_308), .Y(n_1008) );
AND2x4_ASAP7_75t_L g1009 ( .A(n_846), .B(n_310), .Y(n_1009) );
BUFx6f_ASAP7_75t_L g1010 ( .A(n_846), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_843), .B(n_311), .Y(n_1011) );
HB1xp67_ASAP7_75t_L g1012 ( .A(n_921), .Y(n_1012) );
AND2x4_ASAP7_75t_L g1013 ( .A(n_872), .B(n_314), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_890), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_844), .B(n_316), .Y(n_1015) );
OR2x2_ASAP7_75t_L g1016 ( .A(n_890), .B(n_317), .Y(n_1016) );
OR2x2_ASAP7_75t_L g1017 ( .A(n_909), .B(n_910), .Y(n_1017) );
AND2x4_ASAP7_75t_L g1018 ( .A(n_872), .B(n_934), .Y(n_1018) );
AND2x4_ASAP7_75t_L g1019 ( .A(n_872), .B(n_934), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_906), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_885), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_845), .B(n_851), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_939), .B(n_878), .Y(n_1023) );
BUFx2_ASAP7_75t_R g1024 ( .A(n_856), .Y(n_1024) );
AND2x4_ASAP7_75t_L g1025 ( .A(n_940), .B(n_894), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_880), .B(n_933), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_952), .B(n_939), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_947), .B(n_940), .Y(n_1028) );
NOR2xp33_ASAP7_75t_L g1029 ( .A(n_1012), .B(n_933), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_950), .B(n_910), .Y(n_1030) );
INVx2_ASAP7_75t_SL g1031 ( .A(n_1018), .Y(n_1031) );
NAND2xp5_ASAP7_75t_L g1032 ( .A(n_942), .B(n_909), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_984), .B(n_932), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_1006), .B(n_919), .Y(n_1034) );
INVx3_ASAP7_75t_L g1035 ( .A(n_1018), .Y(n_1035) );
OR2x2_ASAP7_75t_L g1036 ( .A(n_946), .B(n_913), .Y(n_1036) );
AND2x4_ASAP7_75t_L g1037 ( .A(n_1025), .B(n_938), .Y(n_1037) );
OR2x2_ASAP7_75t_L g1038 ( .A(n_978), .B(n_913), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_955), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_1023), .B(n_938), .Y(n_1040) );
INVxp33_ASAP7_75t_L g1041 ( .A(n_945), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_953), .B(n_927), .Y(n_1042) );
INVxp67_ASAP7_75t_L g1043 ( .A(n_1017), .Y(n_1043) );
INVx2_ASAP7_75t_L g1044 ( .A(n_977), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_992), .B(n_927), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_981), .B(n_869), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_961), .B(n_869), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_962), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_968), .Y(n_1049) );
OR2x2_ASAP7_75t_L g1050 ( .A(n_944), .B(n_916), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_948), .B(n_918), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1000), .Y(n_1052) );
NOR2xp33_ASAP7_75t_L g1053 ( .A(n_1026), .B(n_880), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_1025), .B(n_888), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_969), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1014), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_980), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_983), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_963), .B(n_866), .Y(n_1059) );
OR2x2_ASAP7_75t_L g1060 ( .A(n_985), .B(n_916), .Y(n_1060) );
INVx2_ASAP7_75t_L g1061 ( .A(n_977), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_987), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1020), .Y(n_1063) );
INVx2_ASAP7_75t_SL g1064 ( .A(n_1019), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_975), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1021), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_1003), .B(n_896), .Y(n_1067) );
AND2x4_ASAP7_75t_L g1068 ( .A(n_990), .B(n_915), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_1022), .B(n_871), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_949), .Y(n_1070) );
INVx2_ASAP7_75t_L g1071 ( .A(n_959), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_965), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_990), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1007), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1007), .B(n_925), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_972), .B(n_858), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1040), .B(n_960), .Y(n_1077) );
INVxp67_ASAP7_75t_SL g1078 ( .A(n_1038), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_1043), .B(n_964), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1042), .B(n_957), .Y(n_1080) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1071), .Y(n_1081) );
NOR2x1p5_ASAP7_75t_L g1082 ( .A(n_1035), .B(n_1010), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_1028), .B(n_971), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1039), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_1043), .B(n_966), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_1027), .B(n_958), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_1071), .B(n_958), .Y(n_1087) );
HB1xp67_ASAP7_75t_L g1088 ( .A(n_1030), .Y(n_1088) );
INVx2_ASAP7_75t_L g1089 ( .A(n_1044), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_1070), .B(n_956), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1048), .Y(n_1091) );
INVx2_ASAP7_75t_SL g1092 ( .A(n_1035), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1054), .B(n_954), .Y(n_1093) );
OR2x2_ASAP7_75t_L g1094 ( .A(n_1036), .B(n_967), .Y(n_1094) );
BUFx2_ASAP7_75t_L g1095 ( .A(n_1031), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_1033), .B(n_970), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1049), .Y(n_1097) );
INVx1_ASAP7_75t_SL g1098 ( .A(n_1064), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1072), .B(n_951), .Y(n_1099) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1052), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1055), .Y(n_1101) );
INVxp67_ASAP7_75t_L g1102 ( .A(n_1029), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1045), .B(n_1024), .Y(n_1103) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_1032), .B(n_1016), .Y(n_1104) );
OR2x2_ASAP7_75t_L g1105 ( .A(n_1032), .B(n_1050), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1056), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1057), .Y(n_1107) );
OR2x2_ASAP7_75t_L g1108 ( .A(n_1060), .B(n_1008), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1058), .Y(n_1109) );
INVx2_ASAP7_75t_L g1110 ( .A(n_1061), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1062), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_1029), .B(n_943), .Y(n_1112) );
OR2x2_ASAP7_75t_L g1113 ( .A(n_1034), .B(n_1010), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1063), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1105), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1078), .B(n_1076), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1078), .B(n_1076), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1088), .B(n_1037), .Y(n_1118) );
OAI21xp33_ASAP7_75t_SL g1119 ( .A1(n_1082), .A2(n_1041), .B(n_1046), .Y(n_1119) );
HB1xp67_ASAP7_75t_L g1120 ( .A(n_1088), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1084), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1091), .Y(n_1122) );
NOR2xp67_ASAP7_75t_R g1123 ( .A(n_1095), .B(n_1010), .Y(n_1123) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_1098), .A2(n_1041), .B1(n_999), .B2(n_1068), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_1079), .B(n_1066), .Y(n_1125) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1097), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1086), .B(n_1037), .Y(n_1127) );
INVx2_ASAP7_75t_L g1128 ( .A(n_1089), .Y(n_1128) );
NAND3xp33_ASAP7_75t_L g1129 ( .A(n_1085), .B(n_1053), .C(n_1074), .Y(n_1129) );
AOI32xp33_ASAP7_75t_L g1130 ( .A1(n_1103), .A2(n_982), .A3(n_976), .B1(n_1069), .B2(n_924), .Y(n_1130) );
AND2x4_ASAP7_75t_L g1131 ( .A(n_1092), .B(n_1073), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1100), .Y(n_1132) );
OR2x2_ASAP7_75t_L g1133 ( .A(n_1094), .B(n_1034), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1107), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1099), .B(n_1065), .Y(n_1135) );
INVxp67_ASAP7_75t_L g1136 ( .A(n_1090), .Y(n_1136) );
AOI22xp5_ASAP7_75t_L g1137 ( .A1(n_1102), .A2(n_1053), .B1(n_1047), .B2(n_1067), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1109), .Y(n_1138) );
AOI222xp33_ASAP7_75t_L g1139 ( .A1(n_1119), .A2(n_1102), .B1(n_1112), .B2(n_1087), .C1(n_1099), .C2(n_1101), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_1136), .B(n_1083), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1141 ( .A(n_1116), .B(n_1083), .Y(n_1141) );
NOR2xp67_ASAP7_75t_L g1142 ( .A(n_1119), .B(n_1120), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1133), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1117), .B(n_1087), .Y(n_1144) );
OR2x2_ASAP7_75t_L g1145 ( .A(n_1135), .B(n_1081), .Y(n_1145) );
INVxp67_ASAP7_75t_L g1146 ( .A(n_1124), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1118), .B(n_1086), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1121), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1122), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1126), .Y(n_1150) );
AND2x4_ASAP7_75t_L g1151 ( .A(n_1129), .B(n_1092), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1132), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1134), .Y(n_1153) );
OAI21xp33_ASAP7_75t_L g1154 ( .A1(n_1130), .A2(n_1096), .B(n_1093), .Y(n_1154) );
AOI22xp5_ASAP7_75t_L g1155 ( .A1(n_1146), .A2(n_1137), .B1(n_1115), .B2(n_1125), .Y(n_1155) );
OAI221xp5_ASAP7_75t_SL g1156 ( .A1(n_1154), .A2(n_1104), .B1(n_1108), .B2(n_1113), .C(n_1075), .Y(n_1156) );
NAND4xp25_ASAP7_75t_L g1157 ( .A(n_1139), .B(n_993), .C(n_988), .D(n_924), .Y(n_1157) );
O2A1O1Ixp5_ASAP7_75t_L g1158 ( .A1(n_1151), .A2(n_1138), .B(n_1131), .C(n_1106), .Y(n_1158) );
OAI21xp5_ASAP7_75t_L g1159 ( .A1(n_1142), .A2(n_1131), .B(n_974), .Y(n_1159) );
INVxp67_ASAP7_75t_L g1160 ( .A(n_1148), .Y(n_1160) );
OAI222xp33_ASAP7_75t_L g1161 ( .A1(n_1151), .A2(n_1127), .B1(n_1077), .B2(n_1123), .C1(n_1059), .C2(n_1111), .Y(n_1161) );
OAI21xp5_ASAP7_75t_L g1162 ( .A1(n_1149), .A2(n_1004), .B(n_1068), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1143), .B(n_1114), .Y(n_1163) );
AOI322xp5_ASAP7_75t_L g1164 ( .A1(n_1140), .A2(n_1077), .A3(n_1080), .B1(n_1081), .B2(n_1128), .C1(n_1051), .C2(n_1068), .Y(n_1164) );
OAI211xp5_ASAP7_75t_L g1165 ( .A1(n_1141), .A2(n_1001), .B(n_1002), .C(n_1011), .Y(n_1165) );
AOI22xp5_ASAP7_75t_L g1166 ( .A1(n_1165), .A2(n_1153), .B1(n_1152), .B2(n_1150), .Y(n_1166) );
NAND3xp33_ASAP7_75t_L g1167 ( .A(n_1156), .B(n_1144), .C(n_1145), .Y(n_1167) );
NAND3xp33_ASAP7_75t_SL g1168 ( .A(n_1158), .B(n_908), .C(n_936), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1155), .B(n_1147), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1160), .B(n_1080), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_1164), .B(n_1089), .Y(n_1171) );
NAND3xp33_ASAP7_75t_SL g1172 ( .A(n_1159), .B(n_908), .C(n_989), .Y(n_1172) );
NOR3xp33_ASAP7_75t_L g1173 ( .A(n_1157), .B(n_1005), .C(n_991), .Y(n_1173) );
AOI22xp5_ASAP7_75t_L g1174 ( .A1(n_1168), .A2(n_1163), .B1(n_1162), .B2(n_1161), .Y(n_1174) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1170), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1167), .Y(n_1176) );
NAND3xp33_ASAP7_75t_L g1177 ( .A(n_1171), .B(n_979), .C(n_973), .Y(n_1177) );
NOR2x1_ASAP7_75t_L g1178 ( .A(n_1172), .B(n_1013), .Y(n_1178) );
NAND3xp33_ASAP7_75t_L g1179 ( .A(n_1173), .B(n_986), .C(n_897), .Y(n_1179) );
NAND4xp75_ASAP7_75t_L g1180 ( .A(n_1176), .B(n_1169), .C(n_1166), .D(n_905), .Y(n_1180) );
NOR2xp67_ASAP7_75t_L g1181 ( .A(n_1175), .B(n_1177), .Y(n_1181) );
NAND2x1_ASAP7_75t_SL g1182 ( .A(n_1178), .B(n_1009), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1179), .Y(n_1183) );
NOR2xp33_ASAP7_75t_L g1184 ( .A(n_1183), .B(n_1174), .Y(n_1184) );
XNOR2x1_ASAP7_75t_L g1185 ( .A(n_1180), .B(n_1009), .Y(n_1185) );
XNOR2xp5_ASAP7_75t_L g1186 ( .A(n_1181), .B(n_1013), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1182), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1184), .B(n_1110), .Y(n_1188) );
INVx2_ASAP7_75t_L g1189 ( .A(n_1187), .Y(n_1189) );
AOI32xp33_ASAP7_75t_L g1190 ( .A1(n_1185), .A2(n_941), .A3(n_892), .B1(n_928), .B2(n_935), .Y(n_1190) );
OAI22xp5_ASAP7_75t_L g1191 ( .A1(n_1189), .A2(n_1186), .B1(n_1188), .B2(n_1190), .Y(n_1191) );
AO22x2_ASAP7_75t_SL g1192 ( .A1(n_1191), .A2(n_923), .B1(n_937), .B2(n_920), .Y(n_1192) );
XNOR2xp5_ASAP7_75t_L g1193 ( .A(n_1192), .B(n_1015), .Y(n_1193) );
AOI22xp5_ASAP7_75t_L g1194 ( .A1(n_1193), .A2(n_994), .B1(n_995), .B2(n_926), .Y(n_1194) );
OAI21xp5_ASAP7_75t_SL g1195 ( .A1(n_1194), .A2(n_922), .B(n_855), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_1195), .B(n_998), .Y(n_1196) );
AOI21xp5_ASAP7_75t_L g1197 ( .A1(n_1196), .A2(n_996), .B(n_997), .Y(n_1197) );
endmodule