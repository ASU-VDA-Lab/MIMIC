module real_jpeg_10691_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_283, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_283;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_1),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_1),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

AOI21xp33_ASAP7_75t_L g199 ( 
.A1(n_1),
.A2(n_16),
.B(n_32),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_2),
.A2(n_26),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_2),
.A2(n_35),
.B1(n_57),
.B2(n_58),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_2),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_3),
.A2(n_57),
.B1(n_58),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_3),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_116),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_116),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_3),
.A2(n_26),
.B1(n_34),
.B2(n_116),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_4),
.A2(n_49),
.B1(n_57),
.B2(n_58),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_5),
.A2(n_26),
.B1(n_34),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_5),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_5),
.A2(n_57),
.B1(n_58),
.B2(n_99),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_99),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_99),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_SL g54 ( 
.A1(n_8),
.A2(n_45),
.B(n_55),
.C(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_8),
.B(n_45),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx6f_ASAP7_75t_SL g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_11),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_11),
.A2(n_57),
.B1(n_58),
.B2(n_125),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_125),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_11),
.A2(n_26),
.B1(n_34),
.B2(n_125),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_12),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_12),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_51),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_13),
.A2(n_51),
.B1(n_57),
.B2(n_58),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_15),
.A2(n_26),
.B1(n_34),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_15),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_15),
.A2(n_57),
.B1(n_58),
.B2(n_82),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_15),
.A2(n_45),
.B1(n_46),
.B2(n_82),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_82),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_16),
.A2(n_45),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_16),
.B(n_45),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_16),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_16),
.A2(n_72),
.B1(n_75),
.B2(n_134),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_16),
.A2(n_31),
.B(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_16),
.B(n_31),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_16),
.B(n_180),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_16),
.A2(n_26),
.B1(n_34),
.B2(n_136),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_17),
.A2(n_26),
.B1(n_34),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_17),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_17),
.A2(n_37),
.B1(n_45),
.B2(n_46),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_17),
.A2(n_37),
.B1(n_57),
.B2(n_58),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_105),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_83),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_21),
.B(n_83),
.Y(n_104)
);

BUFx24_ASAP7_75t_SL g282 ( 
.A(n_21),
.Y(n_282)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_63),
.CI(n_68),
.CON(n_21),
.SN(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_38),
.B2(n_39),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_25),
.A2(n_30),
.B1(n_33),
.B2(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_25),
.A2(n_30),
.B1(n_81),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_25),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_25),
.A2(n_30),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_25),
.A2(n_30),
.B1(n_98),
.B2(n_233),
.Y(n_250)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_28),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_26),
.A2(n_28),
.B(n_136),
.C(n_199),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_30),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_42),
.Y(n_43)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_52),
.B1(n_53),
.B2(n_62),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_44),
.B1(n_48),
.B2(n_50),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_44),
.B1(n_48),
.B2(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_41),
.A2(n_44),
.B1(n_65),
.B2(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_41),
.A2(n_44),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_41),
.A2(n_44),
.B1(n_160),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_41),
.A2(n_44),
.B1(n_176),
.B2(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_41),
.A2(n_44),
.B1(n_217),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_41),
.A2(n_44),
.B1(n_102),
.B2(n_229),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_43),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_44),
.B(n_136),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_45),
.B(n_47),
.Y(n_164)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_46),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_56),
.B(n_60),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_56),
.B1(n_60),
.B2(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_56),
.B1(n_67),
.B2(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_54),
.A2(n_56),
.B1(n_78),
.B2(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_54),
.A2(n_56),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_54),
.A2(n_56),
.B1(n_124),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_54),
.A2(n_56),
.B1(n_149),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_54),
.A2(n_56),
.B1(n_156),
.B2(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_54),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_54),
.A2(n_56),
.B1(n_95),
.B2(n_239),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_56),
.B(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_56),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_57),
.B(n_59),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_57),
.B(n_140),
.Y(n_139)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_58),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_64),
.B(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_79),
.B(n_80),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_70),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_77),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_71),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_79),
.B1(n_80),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_71),
.A2(n_77),
.B1(n_79),
.B2(n_264),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B(n_76),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_75),
.B1(n_76),
.B2(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_72),
.A2(n_75),
.B1(n_115),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_72),
.A2(n_75),
.B1(n_118),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_72),
.A2(n_75),
.B1(n_151),
.B2(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_72),
.A2(n_75),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_72),
.A2(n_75),
.B1(n_93),
.B2(n_203),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_73),
.A2(n_74),
.B1(n_114),
.B2(n_117),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_73),
.A2(n_74),
.B1(n_168),
.B2(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_74),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_75),
.B(n_136),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_77),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_80),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.C(n_89),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_84),
.B(n_88),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_89),
.A2(n_90),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.C(n_100),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_91),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_92),
.B(n_94),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI321xp33_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_258),
.A3(n_269),
.B1(n_275),
.B2(n_280),
.C(n_283),
.Y(n_105)
);

NOR3xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_223),
.C(n_254),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_192),
.B(n_222),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_170),
.B(n_191),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_153),
.B(n_169),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_143),
.B(n_152),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_131),
.B(n_142),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_119),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_119),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_126),
.B2(n_130),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_130),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_123),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_126),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_137),
.B(n_141),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_135),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_144),
.B(n_145),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_146),
.B(n_154),
.Y(n_169)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_148),
.CI(n_150),
.CON(n_146),
.SN(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_154),
.Y(n_171)
);

FAx1_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_157),
.CI(n_161),
.CON(n_154),
.SN(n_154)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_159),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_166),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_172),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_184),
.B2(n_185),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_187),
.C(n_189),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_177),
.B1(n_178),
.B2(n_183),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_175),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_181),
.C(n_183),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_180),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_182),
.Y(n_202)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_186),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_187),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_188),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_193),
.B(n_194),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_207),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_196),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_196),
.B(n_206),
.C(n_207),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_201),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_204),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_218),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_215),
.B2(n_216),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_215),
.C(n_218),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_213),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_221),
.Y(n_232)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI21xp33_ASAP7_75t_L g276 ( 
.A1(n_224),
.A2(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_241),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_225),
.B(n_241),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_236),
.C(n_240),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_235),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_230),
.B1(n_231),
.B2(n_234),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_228),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_SL g252 ( 
.A(n_230),
.B(n_234),
.C(n_235),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_240),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_238),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_252),
.B2(n_253),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_245),
.C(n_253),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_249),
.C(n_251),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_248),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_252),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_256),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_266),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_259),
.B(n_266),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.C(n_265),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_274),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_263),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_270),
.A2(n_276),
.B(n_279),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_271),
.B(n_272),
.Y(n_279)
);


endmodule