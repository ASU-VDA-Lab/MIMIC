module fake_jpeg_7117_n_142 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_22),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_21),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_32),
.Y(n_53)
);

NOR2xp67_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_21),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_16),
.B(n_25),
.C(n_15),
.Y(n_54)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_35),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_30),
.B(n_28),
.C(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_51),
.B(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_17),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_63),
.Y(n_69)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_57),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_30),
.B1(n_16),
.B2(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_65),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_26),
.B1(n_20),
.B2(n_24),
.Y(n_57)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_45),
.B(n_35),
.C(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_17),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_20),
.B1(n_26),
.B2(n_13),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_23),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_18),
.B1(n_24),
.B2(n_23),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_34),
.B1(n_41),
.B2(n_39),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_74),
.B1(n_82),
.B2(n_75),
.Y(n_88)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_80),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_74),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_17),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_91),
.B1(n_94),
.B2(n_96),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_93),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_61),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_61),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_51),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_86),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_72),
.C(n_70),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_106),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_97),
.A2(n_67),
.B1(n_68),
.B2(n_78),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_108),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_89),
.A2(n_67),
.B1(n_70),
.B2(n_51),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_70),
.B1(n_19),
.B2(n_13),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_41),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_111),
.B(n_112),
.Y(n_120)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_113),
.B(n_118),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_106),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_115),
.B(n_116),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_84),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_114),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_122),
.Y(n_128)
);

OAI31xp33_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_101),
.A3(n_90),
.B(n_105),
.Y(n_121)
);

AOI31xp67_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_18),
.A3(n_2),
.B(n_0),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_101),
.C(n_39),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_117),
.C(n_19),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_122),
.B(n_14),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_120),
.B(n_125),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_124),
.A2(n_76),
.B1(n_2),
.B2(n_6),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_130),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_132),
.B(n_133),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_10),
.B(n_4),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_131),
.B(n_126),
.Y(n_136)
);

AOI21x1_ASAP7_75t_SL g139 ( 
.A1(n_136),
.A2(n_137),
.B(n_9),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_8),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_135),
.A2(n_76),
.B1(n_9),
.B2(n_11),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_139),
.B(n_11),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_12),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_2),
.Y(n_142)
);


endmodule