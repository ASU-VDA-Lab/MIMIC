module fake_netlist_5_537_n_664 (n_137, n_91, n_82, n_122, n_10, n_140, n_24, n_124, n_86, n_136, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_664);

input n_137;
input n_91;
input n_82;
input n_122;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_664;

wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_418;
wire n_248;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_619;
wire n_408;
wire n_376;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_483;
wire n_544;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_501;
wire n_245;
wire n_280;
wire n_590;
wire n_629;
wire n_378;
wire n_551;
wire n_581;
wire n_382;
wire n_554;
wire n_254;
wire n_583;
wire n_302;
wire n_265;
wire n_526;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_455;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_507;
wire n_497;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_506;
wire n_610;
wire n_509;
wire n_568;
wire n_373;
wire n_147;
wire n_307;
wire n_633;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_546;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_264;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_243;
wire n_183;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_415;
wire n_141;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_584;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_638;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_332;
wire n_170;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_627;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_572;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_269;
wire n_529;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_262;
wire n_238;
wire n_639;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_256;
wire n_305;
wire n_533;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_56),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_29),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_89),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_43),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_37),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_121),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

BUFx10_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_33),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_11),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_79),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_57),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_74),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_19),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_108),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_66),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_50),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_72),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_51),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_35),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_67),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_133),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_49),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_122),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_126),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_10),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_47),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_26),
.Y(n_176)
);

BUFx10_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_130),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_97),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_86),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_124),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_20),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_132),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_83),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_3),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_118),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_27),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_96),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_128),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_103),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_14),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_12),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_81),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_127),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_140),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_6),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_109),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_25),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_18),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_1),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_34),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_9),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_87),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_16),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_12),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_15),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_111),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_208),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_206),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_0),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_173),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_151),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_159),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_153),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_171),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_145),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_144),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_145),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_155),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_170),
.B(n_0),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_192),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_L g226 ( 
.A(n_152),
.B(n_1),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_196),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_193),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_146),
.Y(n_230)
);

NOR2xp67_ASAP7_75t_L g231 ( 
.A(n_152),
.B(n_2),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_204),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_141),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_207),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_178),
.B(n_2),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_142),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_143),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_147),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_148),
.Y(n_239)
);

NOR2xp67_ASAP7_75t_L g240 ( 
.A(n_162),
.B(n_3),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_150),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g242 ( 
.A(n_149),
.Y(n_242)
);

NOR2xp67_ASAP7_75t_L g243 ( 
.A(n_162),
.B(n_4),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_164),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_154),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_176),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_165),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_156),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_168),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_185),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_174),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_179),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_184),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_180),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_157),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_189),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_236),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_219),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_210),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_220),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_221),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

OA21x2_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_176),
.B(n_197),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_254),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_236),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_R g267 ( 
.A(n_225),
.B(n_227),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_237),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_237),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_245),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_216),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_222),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_210),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_225),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_215),
.B(n_190),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_245),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_201),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_214),
.B(n_153),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_197),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_212),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_246),
.Y(n_283)
);

NAND2xp33_ASAP7_75t_R g284 ( 
.A(n_227),
.B(n_4),
.Y(n_284)
);

OA21x2_ASAP7_75t_L g285 ( 
.A1(n_246),
.A2(n_209),
.B(n_205),
.Y(n_285)
);

NOR2xp67_ASAP7_75t_L g286 ( 
.A(n_232),
.B(n_195),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_242),
.B(n_199),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_233),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_218),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_212),
.B(n_202),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_224),
.B(n_153),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_249),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_239),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_251),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_252),
.B(n_203),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_211),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_256),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_253),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_241),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_217),
.B(n_158),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_255),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_223),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_235),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_226),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_232),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_229),
.B(n_217),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_213),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_234),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_234),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_288),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_160),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_161),
.Y(n_312)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_274),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_260),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_163),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_261),
.Y(n_318)
);

OR2x6_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_250),
.Y(n_319)
);

NAND3xp33_ASAP7_75t_L g320 ( 
.A(n_279),
.B(n_243),
.C(n_240),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_228),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_263),
.Y(n_322)
);

AND3x2_ASAP7_75t_L g323 ( 
.A(n_276),
.B(n_177),
.C(n_231),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_307),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_267),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_306),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_307),
.A2(n_290),
.B1(n_291),
.B2(n_280),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_166),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_269),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_271),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_298),
.B(n_177),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_265),
.Y(n_332)
);

INVx5_ASAP7_75t_L g333 ( 
.A(n_275),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_275),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_292),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_302),
.B(n_167),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_265),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_265),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_286),
.B(n_177),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_281),
.B(n_198),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_308),
.B(n_169),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_308),
.B(n_267),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_300),
.B(n_194),
.Y(n_344)
);

OR2x6_ASAP7_75t_L g345 ( 
.A(n_298),
.B(n_180),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_296),
.Y(n_346)
);

BUFx4f_ASAP7_75t_L g347 ( 
.A(n_275),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_285),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_302),
.B(n_172),
.Y(n_349)
);

NAND2xp33_ASAP7_75t_L g350 ( 
.A(n_277),
.B(n_287),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_275),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_304),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_273),
.Y(n_353)
);

NAND2xp33_ASAP7_75t_L g354 ( 
.A(n_295),
.B(n_180),
.Y(n_354)
);

INVx5_ASAP7_75t_L g355 ( 
.A(n_259),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_293),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_294),
.Y(n_357)
);

BUFx4f_ASAP7_75t_L g358 ( 
.A(n_285),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_297),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_257),
.B(n_266),
.Y(n_360)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_285),
.Y(n_361)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_264),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_273),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_297),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_258),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_299),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_258),
.Y(n_367)
);

NAND2x1p5_ASAP7_75t_L g368 ( 
.A(n_259),
.B(n_180),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_283),
.B(n_175),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_283),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_264),
.Y(n_371)
);

BUFx10_ASAP7_75t_L g372 ( 
.A(n_268),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_264),
.Y(n_373)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_270),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_272),
.B(n_181),
.Y(n_375)
);

AND3x4_ASAP7_75t_L g376 ( 
.A(n_284),
.B(n_5),
.C(n_6),
.Y(n_376)
);

OR2x6_ASAP7_75t_L g377 ( 
.A(n_284),
.B(n_5),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g378 ( 
.A1(n_348),
.A2(n_309),
.B1(n_305),
.B2(n_278),
.Y(n_378)
);

A2O1A1Ixp33_ASAP7_75t_L g379 ( 
.A1(n_358),
.A2(n_188),
.B(n_183),
.C(n_186),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_338),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_371),
.B(n_373),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_327),
.B(n_282),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_331),
.B(n_282),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_348),
.A2(n_282),
.B1(n_187),
.B2(n_182),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_315),
.B(n_301),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_21),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_324),
.A2(n_350),
.B1(n_328),
.B2(n_341),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_311),
.A2(n_289),
.B1(n_262),
.B2(n_70),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_364),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_325),
.B(n_289),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_370),
.Y(n_392)
);

AND2x2_ASAP7_75t_SL g393 ( 
.A(n_374),
.B(n_360),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

BUFx8_ASAP7_75t_L g395 ( 
.A(n_375),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_312),
.A2(n_262),
.B1(n_69),
.B2(n_71),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_371),
.B(n_22),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_317),
.B(n_7),
.Y(n_398)
);

A2O1A1Ixp33_ASAP7_75t_SL g399 ( 
.A1(n_344),
.A2(n_68),
.B(n_137),
.C(n_136),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_316),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_318),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_313),
.B(n_7),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_359),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_351),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_363),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_343),
.B(n_8),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_313),
.B(n_23),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_313),
.B(n_362),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_346),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_336),
.B(n_349),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_362),
.B(n_24),
.Y(n_411)
);

O2A1O1Ixp5_ASAP7_75t_L g412 ( 
.A1(n_361),
.A2(n_73),
.B(n_131),
.C(n_125),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_322),
.B(n_28),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_352),
.B(n_8),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g415 ( 
.A1(n_361),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_329),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_320),
.B(n_13),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_375),
.B(n_13),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_330),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_335),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_357),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_321),
.B(n_14),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_369),
.B(n_15),
.Y(n_423)
);

INVx5_ASAP7_75t_L g424 ( 
.A(n_332),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_369),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_310),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_314),
.B(n_77),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_351),
.Y(n_428)
);

AND2x4_ASAP7_75t_SL g429 ( 
.A(n_372),
.B(n_78),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_R g430 ( 
.A(n_356),
.B(n_76),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_337),
.B(n_80),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_365),
.B(n_16),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_334),
.B(n_82),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_351),
.B(n_75),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_342),
.B(n_17),
.Y(n_435)
);

NAND2xp33_ASAP7_75t_L g436 ( 
.A(n_332),
.B(n_84),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_332),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_319),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_345),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_339),
.B(n_65),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_354),
.A2(n_85),
.B1(n_30),
.B2(n_31),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_339),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_377),
.Y(n_443)
);

INVx5_ASAP7_75t_L g444 ( 
.A(n_339),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_410),
.B(n_374),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_394),
.Y(n_446)
);

INVx5_ASAP7_75t_L g447 ( 
.A(n_404),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_381),
.B(n_340),
.Y(n_448)
);

NOR3xp33_ASAP7_75t_SL g449 ( 
.A(n_418),
.B(n_367),
.C(n_366),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_405),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_443),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_426),
.Y(n_452)
);

INVx5_ASAP7_75t_L g453 ( 
.A(n_404),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_416),
.B(n_319),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_380),
.Y(n_455)
);

A2O1A1Ixp33_ASAP7_75t_L g456 ( 
.A1(n_406),
.A2(n_376),
.B(n_377),
.C(n_347),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_388),
.B(n_372),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_381),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_392),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_428),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_395),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_400),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_437),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_403),
.Y(n_464)
);

BUFx4f_ASAP7_75t_L g465 ( 
.A(n_432),
.Y(n_465)
);

INVx5_ASAP7_75t_L g466 ( 
.A(n_404),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_391),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_384),
.B(n_345),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_382),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_419),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_401),
.B(n_355),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_420),
.B(n_355),
.Y(n_472)
);

CKINVDCx6p67_ASAP7_75t_R g473 ( 
.A(n_393),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_421),
.B(n_355),
.Y(n_474)
);

OR2x6_ASAP7_75t_L g475 ( 
.A(n_438),
.B(n_368),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_398),
.B(n_425),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_395),
.Y(n_477)
);

NOR3xp33_ASAP7_75t_SL g478 ( 
.A(n_383),
.B(n_323),
.C(n_17),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_409),
.B(n_333),
.Y(n_479)
);

NOR3xp33_ASAP7_75t_SL g480 ( 
.A(n_423),
.B(n_32),
.C(n_36),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_442),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_390),
.B(n_333),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_430),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_411),
.B(n_387),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_435),
.B(n_333),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_415),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_442),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_434),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_484),
.A2(n_397),
.B(n_387),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_484),
.A2(n_397),
.B(n_411),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_488),
.A2(n_408),
.B(n_444),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_462),
.Y(n_492)
);

OAI22x1_ASAP7_75t_L g493 ( 
.A1(n_467),
.A2(n_389),
.B1(n_422),
.B2(n_386),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_465),
.Y(n_494)
);

NAND2x1p5_ASAP7_75t_L g495 ( 
.A(n_447),
.B(n_444),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_465),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_448),
.A2(n_408),
.B(n_424),
.Y(n_497)
);

OR2x6_ASAP7_75t_L g498 ( 
.A(n_461),
.B(n_417),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_470),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_469),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_458),
.B(n_378),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_452),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_458),
.B(n_414),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_468),
.B(n_483),
.Y(n_504)
);

OAI21x1_ASAP7_75t_L g505 ( 
.A1(n_481),
.A2(n_431),
.B(n_427),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_481),
.A2(n_431),
.B(n_427),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_445),
.B(n_385),
.Y(n_507)
);

AND2x2_ASAP7_75t_SL g508 ( 
.A(n_486),
.B(n_396),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_460),
.A2(n_433),
.B(n_440),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_460),
.A2(n_433),
.B(n_440),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_476),
.A2(n_379),
.B(n_412),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_463),
.A2(n_434),
.B(n_407),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_446),
.B(n_439),
.Y(n_513)
);

AOI211x1_ASAP7_75t_L g514 ( 
.A1(n_457),
.A2(n_402),
.B(n_413),
.C(n_407),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_486),
.B(n_444),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_459),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_470),
.A2(n_441),
.B(n_399),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_463),
.A2(n_444),
.B(n_424),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_464),
.B(n_429),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_508),
.A2(n_457),
.B(n_456),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_503),
.B(n_456),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_516),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_516),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_512),
.A2(n_482),
.B(n_464),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_509),
.A2(n_459),
.B(n_471),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_510),
.A2(n_487),
.B(n_479),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_505),
.A2(n_479),
.B(n_436),
.Y(n_527)
);

OAI21x1_ASAP7_75t_L g528 ( 
.A1(n_505),
.A2(n_447),
.B(n_453),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_506),
.A2(n_447),
.B(n_453),
.Y(n_529)
);

OA21x2_ASAP7_75t_L g530 ( 
.A1(n_490),
.A2(n_511),
.B(n_489),
.Y(n_530)
);

OAI21x1_ASAP7_75t_SL g531 ( 
.A1(n_490),
.A2(n_480),
.B(n_473),
.Y(n_531)
);

OAI22xp33_ASAP7_75t_L g532 ( 
.A1(n_494),
.A2(n_473),
.B1(n_452),
.B2(n_461),
.Y(n_532)
);

AOI221xp5_ASAP7_75t_SL g533 ( 
.A1(n_493),
.A2(n_451),
.B1(n_450),
.B2(n_478),
.C(n_449),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_508),
.A2(n_466),
.B1(n_447),
.B2(n_453),
.Y(n_534)
);

AO21x1_ASAP7_75t_L g535 ( 
.A1(n_515),
.A2(n_485),
.B(n_454),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g536 ( 
.A1(n_506),
.A2(n_466),
.B(n_453),
.Y(n_536)
);

OA21x2_ASAP7_75t_L g537 ( 
.A1(n_489),
.A2(n_485),
.B(n_474),
.Y(n_537)
);

AO21x2_ASAP7_75t_L g538 ( 
.A1(n_517),
.A2(n_485),
.B(n_474),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_499),
.B(n_474),
.Y(n_539)
);

NAND2x1p5_ASAP7_75t_L g540 ( 
.A(n_515),
.B(n_466),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_492),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_501),
.B(n_472),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_514),
.Y(n_543)
);

O2A1O1Ixp33_ASAP7_75t_SL g544 ( 
.A1(n_507),
.A2(n_519),
.B(n_491),
.C(n_497),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_518),
.Y(n_545)
);

OA21x2_ASAP7_75t_L g546 ( 
.A1(n_497),
.A2(n_472),
.B(n_454),
.Y(n_546)
);

AOI21xp33_ASAP7_75t_L g547 ( 
.A1(n_520),
.A2(n_498),
.B(n_496),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_539),
.B(n_504),
.Y(n_548)
);

OR2x6_ASAP7_75t_L g549 ( 
.A(n_535),
.B(n_500),
.Y(n_549)
);

OAI21x1_ASAP7_75t_L g550 ( 
.A1(n_525),
.A2(n_491),
.B(n_495),
.Y(n_550)
);

OR2x6_ASAP7_75t_L g551 ( 
.A(n_535),
.B(n_455),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_539),
.B(n_498),
.Y(n_552)
);

NAND3x1_ASAP7_75t_L g553 ( 
.A(n_521),
.B(n_542),
.C(n_533),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_541),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_540),
.A2(n_498),
.B1(n_502),
.B2(n_513),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_541),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_522),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_522),
.B(n_502),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_523),
.B(n_454),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_544),
.A2(n_466),
.B(n_424),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_531),
.A2(n_475),
.B1(n_472),
.B2(n_455),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_523),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_543),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_543),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_534),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_538),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_538),
.B(n_475),
.Y(n_567)
);

NAND2xp33_ASAP7_75t_SL g568 ( 
.A(n_538),
.B(n_477),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_R g569 ( 
.A1(n_532),
.A2(n_477),
.B(n_475),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_531),
.B(n_495),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_546),
.Y(n_571)
);

OR2x6_ASAP7_75t_L g572 ( 
.A(n_540),
.B(n_41),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_540),
.A2(n_424),
.B1(n_44),
.B2(n_45),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_545),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_546),
.A2(n_42),
.B1(n_46),
.B2(n_48),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_546),
.B(n_52),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_524),
.B(n_53),
.Y(n_577)
);

AOI221xp5_ASAP7_75t_SL g578 ( 
.A1(n_545),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.C(n_59),
.Y(n_578)
);

OAI211xp5_ASAP7_75t_SL g579 ( 
.A1(n_547),
.A2(n_546),
.B(n_537),
.C(n_526),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_556),
.Y(n_580)
);

OAI211xp5_ASAP7_75t_SL g581 ( 
.A1(n_561),
.A2(n_537),
.B(n_526),
.C(n_530),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_563),
.Y(n_582)
);

OAI211xp5_ASAP7_75t_L g583 ( 
.A1(n_575),
.A2(n_530),
.B(n_537),
.C(n_527),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_563),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_564),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_552),
.A2(n_537),
.B1(n_530),
.B2(n_527),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_554),
.Y(n_587)
);

INVx8_ASAP7_75t_L g588 ( 
.A(n_572),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_557),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_548),
.B(n_60),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_552),
.A2(n_530),
.B1(n_525),
.B2(n_524),
.Y(n_591)
);

AOI211xp5_ASAP7_75t_L g592 ( 
.A1(n_555),
.A2(n_536),
.B(n_529),
.C(n_528),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_562),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_574),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_567),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_548),
.B(n_536),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_549),
.A2(n_529),
.B1(n_528),
.B2(n_63),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_558),
.B(n_61),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_549),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_569),
.A2(n_62),
.B1(n_88),
.B2(n_90),
.Y(n_600)
);

AND3x1_ASAP7_75t_L g601 ( 
.A(n_559),
.B(n_92),
.C(n_94),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_580),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_595),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_582),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_585),
.B(n_566),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_599),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_584),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_591),
.B(n_571),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_589),
.Y(n_609)
);

INVxp67_ASAP7_75t_SL g610 ( 
.A(n_592),
.Y(n_610)
);

OAI22xp33_ASAP7_75t_L g611 ( 
.A1(n_588),
.A2(n_572),
.B1(n_565),
.B2(n_551),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_586),
.B(n_571),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_596),
.B(n_576),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_587),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_594),
.B(n_551),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_593),
.Y(n_616)
);

AO21x2_ASAP7_75t_L g617 ( 
.A1(n_610),
.A2(n_579),
.B(n_583),
.Y(n_617)
);

OAI21x1_ASAP7_75t_L g618 ( 
.A1(n_608),
.A2(n_550),
.B(n_560),
.Y(n_618)
);

OAI31xp33_ASAP7_75t_L g619 ( 
.A1(n_611),
.A2(n_600),
.A3(n_568),
.B(n_590),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_607),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_607),
.Y(n_621)
);

BUFx10_ASAP7_75t_L g622 ( 
.A(n_616),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_603),
.B(n_553),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_613),
.B(n_577),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_620),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_620),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_624),
.B(n_606),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_621),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_621),
.B(n_608),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_622),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_R g631 ( 
.A(n_623),
.B(n_612),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_627),
.B(n_624),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_625),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_629),
.B(n_613),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_630),
.B(n_622),
.Y(n_635)
);

OAI21xp33_ASAP7_75t_L g636 ( 
.A1(n_631),
.A2(n_615),
.B(n_600),
.Y(n_636)
);

NOR3xp33_ASAP7_75t_SL g637 ( 
.A(n_636),
.B(n_619),
.C(n_581),
.Y(n_637)
);

OAI221xp5_ASAP7_75t_L g638 ( 
.A1(n_636),
.A2(n_602),
.B1(n_606),
.B2(n_615),
.C(n_601),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_L g639 ( 
.A(n_635),
.B(n_588),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_634),
.B(n_617),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_632),
.B(n_602),
.Y(n_641)
);

NAND2x1_ASAP7_75t_L g642 ( 
.A(n_641),
.B(n_633),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_638),
.A2(n_617),
.B(n_588),
.Y(n_643)
);

OAI21xp33_ASAP7_75t_L g644 ( 
.A1(n_637),
.A2(n_612),
.B(n_628),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_642),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_643),
.A2(n_639),
.B(n_640),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_645),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_647),
.B(n_644),
.Y(n_648)
);

XNOR2x1_ASAP7_75t_L g649 ( 
.A(n_648),
.B(n_598),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_649),
.B(n_646),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_650),
.Y(n_651)
);

AOI222xp33_ASAP7_75t_L g652 ( 
.A1(n_651),
.A2(n_622),
.B1(n_573),
.B2(n_625),
.C1(n_577),
.C2(n_597),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_652),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_653),
.B(n_617),
.Y(n_654)
);

OAI21xp33_ASAP7_75t_SL g655 ( 
.A1(n_654),
.A2(n_626),
.B(n_604),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_655),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_656),
.A2(n_578),
.B(n_626),
.Y(n_657)
);

AOI21xp33_ASAP7_75t_L g658 ( 
.A1(n_656),
.A2(n_95),
.B(n_98),
.Y(n_658)
);

AOI222xp33_ASAP7_75t_L g659 ( 
.A1(n_657),
.A2(n_622),
.B1(n_609),
.B2(n_614),
.C1(n_583),
.C2(n_605),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_SL g660 ( 
.A1(n_658),
.A2(n_609),
.B1(n_614),
.B2(n_605),
.Y(n_660)
);

AOI222xp33_ASAP7_75t_L g661 ( 
.A1(n_660),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.C1(n_104),
.C2(n_105),
.Y(n_661)
);

AOI222xp33_ASAP7_75t_L g662 ( 
.A1(n_659),
.A2(n_106),
.B1(n_107),
.B2(n_110),
.C1(n_112),
.C2(n_113),
.Y(n_662)
);

OAI221xp5_ASAP7_75t_L g663 ( 
.A1(n_661),
.A2(n_662),
.B1(n_570),
.B2(n_115),
.C(n_116),
.Y(n_663)
);

AOI211xp5_ASAP7_75t_L g664 ( 
.A1(n_663),
.A2(n_138),
.B(n_618),
.C(n_570),
.Y(n_664)
);


endmodule