module fake_jpeg_9550_n_284 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_284);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_14;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_20),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_17),
.Y(n_32)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_29),
.B(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_52),
.Y(n_63)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_30),
.B(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_54),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_17),
.B(n_15),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_16),
.B1(n_18),
.B2(n_25),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_58),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_61),
.Y(n_87)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_47),
.B1(n_53),
.B2(n_54),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_62),
.A2(n_64),
.B1(n_68),
.B2(n_70),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_20),
.B1(n_27),
.B2(n_35),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_67),
.Y(n_96)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_19),
.B1(n_36),
.B2(n_33),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_38),
.A2(n_20),
.B1(n_19),
.B2(n_24),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_75),
.B1(n_27),
.B2(n_44),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_52),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_20),
.B1(n_27),
.B2(n_22),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_19),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_80),
.A2(n_60),
.B(n_19),
.C(n_68),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_63),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_84),
.Y(n_118)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_71),
.B(n_57),
.Y(n_99)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_86),
.A2(n_90),
.B1(n_44),
.B2(n_27),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_98),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_91),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_64),
.A2(n_73),
.B1(n_59),
.B2(n_65),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_92),
.A2(n_95),
.B1(n_60),
.B2(n_56),
.Y(n_110)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_44),
.B1(n_43),
.B2(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_100),
.B(n_106),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_57),
.B(n_40),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_19),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_105),
.C(n_108),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_16),
.B(n_18),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_19),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_40),
.B(n_48),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_68),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_56),
.Y(n_109)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_120),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_68),
.Y(n_112)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_66),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_41),
.Y(n_121)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_121),
.A2(n_98),
.B1(n_90),
.B2(n_85),
.Y(n_125)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_87),
.Y(n_126)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_102),
.A2(n_106),
.B1(n_100),
.B2(n_110),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_127),
.A2(n_132),
.B(n_137),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_105),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_131),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_120),
.B(n_22),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_140),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_103),
.A2(n_93),
.B1(n_78),
.B2(n_86),
.Y(n_130)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_41),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_37),
.C(n_36),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_37),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_141),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_16),
.B(n_18),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_111),
.Y(n_139)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_13),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_99),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

OA21x2_ASAP7_75t_L g147 ( 
.A1(n_136),
.A2(n_123),
.B(n_127),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_147),
.A2(n_165),
.B(n_21),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_148),
.B(n_158),
.Y(n_184)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_153),
.Y(n_181)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_112),
.B(n_118),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_136),
.B(n_138),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_103),
.B1(n_84),
.B2(n_93),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_161),
.Y(n_171)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_135),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_133),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_168),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_0),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_140),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_166),
.Y(n_188)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_169),
.A2(n_170),
.B(n_178),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_142),
.B(n_135),
.Y(n_170)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_142),
.B(n_104),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_172),
.A2(n_46),
.B(n_21),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_128),
.C(n_141),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_186),
.C(n_145),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_149),
.A2(n_111),
.B1(n_114),
.B2(n_117),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_174),
.A2(n_189),
.B1(n_24),
.B2(n_26),
.Y(n_210)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_149),
.A2(n_104),
.B1(n_117),
.B2(n_115),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_187),
.B1(n_190),
.B2(n_163),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_23),
.B(n_22),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_94),
.B1(n_91),
.B2(n_79),
.Y(n_183)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_46),
.C(n_77),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_156),
.A2(n_79),
.B1(n_77),
.B2(n_25),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_25),
.B1(n_15),
.B2(n_21),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_147),
.A2(n_77),
.B1(n_89),
.B2(n_15),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_157),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_176),
.Y(n_192)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_203),
.C(n_186),
.Y(n_213)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_151),
.C(n_152),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_195),
.B(n_201),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_165),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_206),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_175),
.B(n_157),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_202),
.B(n_205),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_145),
.C(n_153),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_147),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_191),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_89),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_207),
.A2(n_210),
.B1(n_190),
.B2(n_177),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_171),
.B(n_12),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_189),
.Y(n_215)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_214),
.C(n_216),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_182),
.C(n_180),
.Y(n_214)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_182),
.C(n_169),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_205),
.A2(n_179),
.B1(n_188),
.B2(n_184),
.Y(n_217)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_184),
.C(n_188),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_26),
.C(n_24),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_174),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_222),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_200),
.A2(n_179),
.B1(n_172),
.B2(n_187),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_223),
.A2(n_224),
.B1(n_194),
.B2(n_196),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_172),
.B1(n_183),
.B2(n_178),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_226),
.B(n_207),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_234),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_233),
.A2(n_240),
.B1(n_13),
.B2(n_2),
.Y(n_251)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_225),
.A2(n_199),
.B1(n_172),
.B2(n_209),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_241),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_198),
.B1(n_202),
.B2(n_197),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_236),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_254)
);

FAx1_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_198),
.CI(n_1),
.CON(n_238),
.SN(n_238)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_0),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_221),
.C(n_26),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_211),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_13),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_242),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_245)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_239),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_244),
.Y(n_257)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_248),
.C(n_249),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_24),
.B1(n_10),
.B2(n_9),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_10),
.B1(n_26),
.B2(n_2),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_1),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_251),
.B(n_13),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_14),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_238),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_254),
.A2(n_242),
.B1(n_3),
.B2(n_4),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_250),
.A2(n_234),
.B1(n_238),
.B2(n_231),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_264),
.B1(n_245),
.B2(n_246),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_261),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_252),
.A2(n_228),
.B1(n_14),
.B2(n_4),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_SL g265 ( 
.A1(n_262),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_14),
.B(n_4),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_6),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_268),
.C(n_269),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_253),
.C(n_246),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_273),
.A2(n_274),
.B(n_275),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_260),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_263),
.B(n_271),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_256),
.B(n_258),
.Y(n_278)
);

AOI21x1_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_276),
.B(n_265),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g280 ( 
.A1(n_279),
.A2(n_6),
.B(n_7),
.Y(n_280)
);

NAND3xp33_ASAP7_75t_SL g281 ( 
.A(n_280),
.B(n_6),
.C(n_7),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_281),
.A2(n_7),
.B1(n_8),
.B2(n_14),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_14),
.B(n_270),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_14),
.Y(n_284)
);


endmodule