module fake_jpeg_13187_n_142 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_142);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_20),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_23),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_67),
.B(n_52),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_50),
.B1(n_53),
.B2(n_56),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_76),
.B1(n_79),
.B2(n_42),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_58),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_55),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_59),
.A2(n_52),
.B1(n_57),
.B2(n_46),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_47),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_45),
.C(n_49),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_81),
.A2(n_42),
.B(n_2),
.Y(n_91)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_88),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_92),
.Y(n_110)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_44),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_86),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_69),
.B(n_0),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_87),
.B(n_89),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_76),
.B(n_1),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_91),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_1),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_96),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_3),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_16),
.B1(n_40),
.B2(n_39),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_18),
.B1(n_37),
.B2(n_36),
.Y(n_107)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_15),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_107),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_95),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_113),
.B1(n_10),
.B2(n_11),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_83),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_111),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_84),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_10),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_5),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_93),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_19),
.B(n_35),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_115),
.A2(n_106),
.B1(n_110),
.B2(n_114),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_110),
.A2(n_22),
.B1(n_31),
.B2(n_12),
.Y(n_117)
);

OAI22x1_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_120),
.B1(n_107),
.B2(n_113),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_27),
.C(n_29),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_125),
.C(n_102),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_122),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_11),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_123),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_103),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_130),
.B1(n_117),
.B2(n_116),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_132),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_119),
.B1(n_120),
.B2(n_124),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_133),
.A2(n_119),
.B(n_126),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_118),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_135),
.B(n_126),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_104),
.B(n_14),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_13),
.CI(n_28),
.CON(n_140),
.SN(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_41),
.C(n_112),
.Y(n_141)
);

BUFx24_ASAP7_75t_SL g142 ( 
.A(n_141),
.Y(n_142)
);


endmodule