module fake_jpeg_25072_n_161 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_161);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_13),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_9),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_0),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_71),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_64),
.B(n_0),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_46),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_48),
.B1(n_44),
.B2(n_52),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_84),
.B1(n_60),
.B2(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_55),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_44),
.B1(n_43),
.B2(n_56),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_65),
.B1(n_47),
.B2(n_49),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_99),
.B1(n_74),
.B2(n_51),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_91),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_59),
.B1(n_42),
.B2(n_63),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_92),
.A2(n_98),
.B1(n_91),
.B2(n_79),
.Y(n_109)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_1),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_97),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_96),
.Y(n_105)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_63),
.B1(n_70),
.B2(n_66),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_62),
.B1(n_57),
.B2(n_61),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_1),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_95),
.A2(n_86),
.B1(n_87),
.B2(n_89),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_104),
.A2(n_108),
.B(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_5),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_99),
.A2(n_57),
.B1(n_22),
.B2(n_41),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_18),
.B(n_40),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_3),
.B(n_4),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_2),
.Y(n_118)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_112),
.B(n_114),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_107),
.B1(n_101),
.B2(n_106),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_119),
.B1(n_120),
.B2(n_5),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_103),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_116),
.Y(n_121)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_79),
.C(n_98),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_31),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_23),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_126),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_28),
.B(n_37),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_32),
.B(n_12),
.Y(n_141)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_129),
.Y(n_144)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_130),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_21),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_118),
.B(n_6),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_125),
.B1(n_129),
.B2(n_121),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_7),
.C(n_8),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_145),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_146),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_124),
.B(n_14),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_128),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_137),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_150),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_149),
.B(n_138),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_142),
.B1(n_139),
.B2(n_151),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_144),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_140),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_143),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_148),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_135),
.C(n_15),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_36),
.Y(n_161)
);


endmodule