module fake_jpeg_3186_n_150 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_150);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_4),
.B(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_38),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_21),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_29),
.Y(n_46)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_23),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_47),
.B1(n_49),
.B2(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_27),
.B1(n_26),
.B2(n_22),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_32),
.A2(n_21),
.B1(n_29),
.B2(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_52),
.B(n_22),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_25),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_14),
.B1(n_28),
.B2(n_25),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_54),
.A2(n_61),
.B1(n_42),
.B2(n_40),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_55),
.B(n_56),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_51),
.A2(n_39),
.B1(n_38),
.B2(n_18),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_41),
.B(n_52),
.Y(n_59)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_50),
.Y(n_81)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_15),
.B1(n_30),
.B2(n_3),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_15),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_7),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_74),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_47),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_64),
.B1(n_63),
.B2(n_61),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_81),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_40),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_43),
.B(n_33),
.C(n_42),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_42),
.B(n_60),
.C(n_33),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_73),
.C(n_81),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_95),
.C(n_2),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_86),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_94),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_98),
.B1(n_83),
.B2(n_79),
.Y(n_105)
);

AO22x1_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_64),
.B1(n_57),
.B2(n_55),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_SL g95 ( 
.A(n_72),
.B(n_43),
.C(n_70),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_97),
.B(n_101),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_69),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_91),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_77),
.B1(n_71),
.B2(n_3),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_103),
.B(n_0),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_102),
.A2(n_76),
.B1(n_85),
.B2(n_82),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_90),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_68),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_109),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_77),
.Y(n_109)
);

OAI21x1_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_112),
.B(n_106),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_110),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_0),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_116),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_117),
.B(n_119),
.Y(n_129)
);

OAI21x1_ASAP7_75t_L g118 ( 
.A1(n_116),
.A2(n_100),
.B(n_95),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_118),
.A2(n_8),
.B(n_10),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_115),
.B(n_90),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_122),
.B1(n_126),
.B2(n_100),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_103),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_111),
.A2(n_100),
.B1(n_4),
.B2(n_6),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_2),
.B1(n_4),
.B2(n_8),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_110),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_130),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_132),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_7),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_120),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_126),
.B(n_124),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_138),
.Y(n_140)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_127),
.C(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_141),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_130),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_142),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_145),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_136),
.C(n_122),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_140),
.Y(n_147)
);

NAND3xp33_ASAP7_75t_SL g148 ( 
.A(n_147),
.B(n_145),
.C(n_119),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_148),
.A2(n_146),
.B(n_11),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_2),
.Y(n_150)
);


endmodule