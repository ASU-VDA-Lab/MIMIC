module fake_netlist_6_2676_n_1553 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_334, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_332, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1553);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_332;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1553;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_1094;
wire n_953;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_811;
wire n_683;
wire n_1207;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_380;
wire n_1535;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1240;

INVx1_ASAP7_75t_L g336 ( 
.A(n_334),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_291),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_106),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_63),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_155),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_272),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_74),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_93),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_304),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_68),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_24),
.Y(n_346)
);

BUFx5_ASAP7_75t_L g347 ( 
.A(n_323),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_207),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_151),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_205),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_54),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_257),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_76),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_53),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_275),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_137),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_171),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_265),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_42),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_222),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_16),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_11),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_12),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_201),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_326),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_69),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_231),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_133),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_177),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_210),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_7),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_211),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_79),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_206),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_92),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_109),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_85),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_101),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_281),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_236),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_288),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_125),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_64),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_232),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_327),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_264),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_227),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_97),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_25),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_224),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_188),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_258),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_278),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_105),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_285),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_176),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_111),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_189),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_263),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_282),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_245),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_62),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_305),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_301),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_219),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_251),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_294),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_297),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_139),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_131),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_252),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_98),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_115),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_128),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_306),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_283),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_107),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_42),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_299),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_333),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_141),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_150),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_311),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_123),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_279),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_136),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_114),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_108),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_269),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_203),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_198),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_35),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_72),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_287),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_130),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_78),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_331),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_238),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_273),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_72),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_310),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_164),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_132),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_175),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_179),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_170),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_173),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_254),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_248),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_244),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_325),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_335),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_81),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_262),
.Y(n_454)
);

BUFx10_ASAP7_75t_L g455 ( 
.A(n_329),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_33),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_7),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_32),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_324),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_148),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_160),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_104),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_75),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_199),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_22),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_307),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_14),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_11),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_161),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_193),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_314),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_68),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_169),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_289),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_40),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_62),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_81),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_28),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_67),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_330),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_292),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_16),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_276),
.Y(n_483)
);

INVxp33_ASAP7_75t_L g484 ( 
.A(n_180),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_65),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_75),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_18),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_0),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_135),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_121),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_235),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_144),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_204),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_44),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_73),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_39),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_53),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_242),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_143),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_58),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_250),
.Y(n_501)
);

BUFx5_ASAP7_75t_L g502 ( 
.A(n_134),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_240),
.Y(n_503)
);

INVxp67_ASAP7_75t_SL g504 ( 
.A(n_23),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_96),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_268),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_218),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_290),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_223),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_116),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_315),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_22),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_284),
.Y(n_513)
);

BUFx10_ASAP7_75t_L g514 ( 
.A(n_159),
.Y(n_514)
);

INVx4_ASAP7_75t_R g515 ( 
.A(n_37),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_214),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_256),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_267),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_302),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_67),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_74),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_127),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_309),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_166),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_5),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_80),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_229),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_99),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_255),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_145),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_226),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_124),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_32),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_216),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_57),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_138),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_88),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_178),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_243),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_212),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_308),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g542 ( 
.A(n_41),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_35),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_185),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_126),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_163),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_220),
.Y(n_547)
);

BUFx5_ASAP7_75t_L g548 ( 
.A(n_293),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_48),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_300),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_64),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_20),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_286),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_316),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_234),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_57),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_0),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_61),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_91),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_41),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_246),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_52),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_475),
.B(n_1),
.Y(n_563)
);

BUFx12f_ASAP7_75t_L g564 ( 
.A(n_542),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_341),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_389),
.B(n_1),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_341),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_457),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_341),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_389),
.B(n_2),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_443),
.B(n_2),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_484),
.B(n_3),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_479),
.B(n_3),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_457),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_487),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_443),
.B(n_4),
.Y(n_576)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_349),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_338),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_468),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_369),
.B(n_448),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_442),
.B(n_4),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_455),
.Y(n_582)
);

INVx5_ASAP7_75t_L g583 ( 
.A(n_349),
.Y(n_583)
);

BUFx8_ASAP7_75t_SL g584 ( 
.A(n_440),
.Y(n_584)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_349),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_487),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_398),
.B(n_5),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_407),
.Y(n_588)
);

INVx5_ASAP7_75t_L g589 ( 
.A(n_407),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_369),
.B(n_6),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_484),
.B(n_6),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_462),
.B(n_8),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_361),
.Y(n_593)
);

CKINVDCx6p67_ASAP7_75t_R g594 ( 
.A(n_542),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_407),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_407),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_490),
.Y(n_597)
);

BUFx8_ASAP7_75t_SL g598 ( 
.A(n_494),
.Y(n_598)
);

BUFx12f_ASAP7_75t_L g599 ( 
.A(n_455),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_448),
.B(n_8),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_490),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_490),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_468),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_468),
.B(n_9),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_490),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_339),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_468),
.B(n_9),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_558),
.B(n_10),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_503),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_558),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_342),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_558),
.B(n_10),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_538),
.B(n_12),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_558),
.B(n_13),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_526),
.Y(n_615)
);

BUFx12f_ASAP7_75t_L g616 ( 
.A(n_514),
.Y(n_616)
);

INVx5_ASAP7_75t_L g617 ( 
.A(n_503),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_538),
.B(n_13),
.Y(n_618)
);

BUFx8_ASAP7_75t_SL g619 ( 
.A(n_549),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_346),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_514),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_343),
.B(n_14),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_418),
.B(n_15),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_453),
.B(n_15),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_561),
.B(n_17),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_503),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_353),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_379),
.B(n_17),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_393),
.B(n_18),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_362),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_503),
.Y(n_631)
);

BUFx8_ASAP7_75t_SL g632 ( 
.A(n_552),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_488),
.B(n_19),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_412),
.B(n_19),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_344),
.Y(n_635)
);

BUFx8_ASAP7_75t_SL g636 ( 
.A(n_560),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_347),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_347),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_473),
.B(n_20),
.Y(n_639)
);

INVxp33_ASAP7_75t_SL g640 ( 
.A(n_345),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_348),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_351),
.Y(n_642)
);

CKINVDCx16_ASAP7_75t_R g643 ( 
.A(n_372),
.Y(n_643)
);

BUFx8_ASAP7_75t_L g644 ( 
.A(n_383),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_456),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_474),
.B(n_21),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_391),
.B(n_21),
.Y(n_647)
);

BUFx12f_ASAP7_75t_L g648 ( 
.A(n_562),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_357),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_358),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_516),
.B(n_23),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_510),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_510),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_336),
.B(n_24),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_404),
.B(n_25),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_481),
.B(n_26),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_458),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_354),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_347),
.Y(n_659)
);

BUFx12f_ASAP7_75t_L g660 ( 
.A(n_359),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_532),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_489),
.B(n_26),
.Y(n_662)
);

CKINVDCx16_ASAP7_75t_R g663 ( 
.A(n_529),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_476),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_478),
.B(n_27),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_340),
.B(n_27),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_360),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_347),
.Y(n_668)
);

BUFx12f_ASAP7_75t_L g669 ( 
.A(n_363),
.Y(n_669)
);

INVx5_ASAP7_75t_L g670 ( 
.A(n_532),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_482),
.B(n_28),
.Y(n_671)
);

XNOR2xp5_ASAP7_75t_L g672 ( 
.A(n_366),
.B(n_29),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_521),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_531),
.B(n_29),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_502),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_502),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_557),
.B(n_30),
.Y(n_677)
);

BUFx8_ASAP7_75t_L g678 ( 
.A(n_543),
.Y(n_678)
);

BUFx12f_ASAP7_75t_L g679 ( 
.A(n_371),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_504),
.B(n_30),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_350),
.B(n_31),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_352),
.B(n_31),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_355),
.B(n_33),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_356),
.B(n_34),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_364),
.B(n_34),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_373),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_402),
.B(n_36),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_432),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_365),
.B(n_36),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_370),
.B(n_37),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_376),
.B(n_38),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_532),
.Y(n_692)
);

INVx5_ASAP7_75t_L g693 ( 
.A(n_532),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_433),
.B(n_38),
.Y(n_694)
);

BUFx2_ASAP7_75t_L g695 ( 
.A(n_436),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_546),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_380),
.B(n_39),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_546),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_546),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_546),
.Y(n_700)
);

INVx5_ASAP7_75t_L g701 ( 
.A(n_502),
.Y(n_701)
);

BUFx8_ASAP7_75t_SL g702 ( 
.A(n_337),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_381),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_367),
.Y(n_704)
);

AND2x6_ASAP7_75t_L g705 ( 
.A(n_384),
.B(n_86),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_385),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_386),
.B(n_40),
.Y(n_707)
);

INVx5_ASAP7_75t_L g708 ( 
.A(n_502),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_463),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_388),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_392),
.Y(n_711)
);

INVx5_ASAP7_75t_L g712 ( 
.A(n_502),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_397),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_579),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_647),
.A2(n_406),
.B1(n_420),
.B2(n_400),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_662),
.A2(n_480),
.B1(n_491),
.B2(n_441),
.Y(n_716)
);

AO22x2_ASAP7_75t_L g717 ( 
.A1(n_622),
.A2(n_403),
.B1(n_408),
.B2(n_399),
.Y(n_717)
);

AO22x2_ASAP7_75t_L g718 ( 
.A1(n_622),
.A2(n_590),
.B1(n_618),
.B2(n_613),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_603),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_702),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_674),
.A2(n_513),
.B1(n_537),
.B2(n_493),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_643),
.A2(n_467),
.B1(n_472),
.B2(n_465),
.Y(n_722)
);

OAI22xp33_ASAP7_75t_SL g723 ( 
.A1(n_566),
.A2(n_485),
.B1(n_486),
.B2(n_477),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_SL g724 ( 
.A1(n_672),
.A2(n_495),
.B1(n_497),
.B2(n_496),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_603),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_610),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_703),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_686),
.B(n_492),
.Y(n_728)
);

OAI22xp33_ASAP7_75t_L g729 ( 
.A1(n_566),
.A2(n_512),
.B1(n_520),
.B2(n_500),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_663),
.A2(n_533),
.B1(n_535),
.B2(n_525),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_SL g731 ( 
.A1(n_570),
.A2(n_556),
.B1(n_551),
.B2(n_524),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_565),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_565),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_565),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_587),
.A2(n_541),
.B1(n_523),
.B2(n_374),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_686),
.B(n_368),
.Y(n_736)
);

NAND2xp33_ASAP7_75t_SL g737 ( 
.A(n_563),
.B(n_375),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_710),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_582),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_569),
.Y(n_740)
);

AOI22x1_ASAP7_75t_L g741 ( 
.A1(n_590),
.A2(n_411),
.B1(n_413),
.B2(n_410),
.Y(n_741)
);

OA22x2_ASAP7_75t_L g742 ( 
.A1(n_575),
.A2(n_415),
.B1(n_421),
.B2(n_414),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_592),
.A2(n_378),
.B1(n_382),
.B2(n_377),
.Y(n_743)
);

AO22x2_ASAP7_75t_L g744 ( 
.A1(n_613),
.A2(n_423),
.B1(n_424),
.B2(n_422),
.Y(n_744)
);

OAI22xp33_ASAP7_75t_L g745 ( 
.A1(n_570),
.A2(n_427),
.B1(n_428),
.B2(n_426),
.Y(n_745)
);

OAI22xp33_ASAP7_75t_L g746 ( 
.A1(n_621),
.A2(n_593),
.B1(n_581),
.B2(n_623),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_578),
.Y(n_747)
);

OAI22xp33_ASAP7_75t_L g748 ( 
.A1(n_621),
.A2(n_438),
.B1(n_445),
.B2(n_434),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_709),
.B(n_387),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_649),
.B(n_447),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_709),
.B(n_390),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_569),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_572),
.A2(n_395),
.B1(n_396),
.B2(n_394),
.Y(n_753)
);

AO22x2_ASAP7_75t_L g754 ( 
.A1(n_618),
.A2(n_460),
.B1(n_461),
.B2(n_459),
.Y(n_754)
);

OR2x6_ASAP7_75t_L g755 ( 
.A(n_648),
.B(n_466),
.Y(n_755)
);

OAI22xp33_ASAP7_75t_L g756 ( 
.A1(n_581),
.A2(n_498),
.B1(n_501),
.B2(n_471),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_569),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_564),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_658),
.B(n_695),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_667),
.B(n_704),
.Y(n_760)
);

BUFx6f_ASAP7_75t_SL g761 ( 
.A(n_580),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_SL g762 ( 
.A1(n_591),
.A2(n_517),
.B1(n_522),
.B2(n_508),
.Y(n_762)
);

OAI22xp33_ASAP7_75t_L g763 ( 
.A1(n_623),
.A2(n_540),
.B1(n_530),
.B2(n_405),
.Y(n_763)
);

AO22x2_ASAP7_75t_L g764 ( 
.A1(n_573),
.A2(n_515),
.B1(n_45),
.B2(n_43),
.Y(n_764)
);

BUFx6f_ASAP7_75t_SL g765 ( 
.A(n_580),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_591),
.A2(n_409),
.B1(n_416),
.B2(n_401),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_642),
.B(n_417),
.Y(n_767)
);

OA22x2_ASAP7_75t_L g768 ( 
.A1(n_568),
.A2(n_425),
.B1(n_429),
.B2(n_419),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_604),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_640),
.B(n_430),
.Y(n_770)
);

OR2x6_ASAP7_75t_L g771 ( 
.A(n_660),
.B(n_43),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_688),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_588),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_635),
.B(n_431),
.Y(n_774)
);

OAI22xp33_ASAP7_75t_SL g775 ( 
.A1(n_571),
.A2(n_559),
.B1(n_555),
.B2(n_554),
.Y(n_775)
);

XNOR2xp5_ASAP7_75t_L g776 ( 
.A(n_677),
.B(n_44),
.Y(n_776)
);

OAI22xp33_ASAP7_75t_SL g777 ( 
.A1(n_576),
.A2(n_553),
.B1(n_550),
.B2(n_435),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_588),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_588),
.Y(n_779)
);

OAI22xp33_ASAP7_75t_R g780 ( 
.A1(n_628),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_641),
.B(n_437),
.Y(n_781)
);

OAI22xp33_ASAP7_75t_L g782 ( 
.A1(n_633),
.A2(n_439),
.B1(n_444),
.B2(n_446),
.Y(n_782)
);

OAI22xp33_ASAP7_75t_L g783 ( 
.A1(n_633),
.A2(n_449),
.B1(n_450),
.B2(n_451),
.Y(n_783)
);

OAI22xp33_ASAP7_75t_R g784 ( 
.A1(n_628),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_650),
.B(n_452),
.Y(n_785)
);

OAI22xp33_ASAP7_75t_L g786 ( 
.A1(n_681),
.A2(n_454),
.B1(n_464),
.B2(n_469),
.Y(n_786)
);

AO22x2_ASAP7_75t_L g787 ( 
.A1(n_600),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_SL g788 ( 
.A1(n_629),
.A2(n_470),
.B1(n_483),
.B2(n_499),
.Y(n_788)
);

BUFx10_ASAP7_75t_L g789 ( 
.A(n_629),
.Y(n_789)
);

BUFx10_ASAP7_75t_L g790 ( 
.A(n_655),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_595),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_655),
.A2(n_527),
.B1(n_547),
.B2(n_545),
.Y(n_792)
);

OAI22xp33_ASAP7_75t_L g793 ( 
.A1(n_681),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_656),
.A2(n_528),
.B1(n_544),
.B2(n_539),
.Y(n_794)
);

OAI22xp33_ASAP7_75t_L g795 ( 
.A1(n_684),
.A2(n_509),
.B1(n_511),
.B2(n_518),
.Y(n_795)
);

AND2x2_ASAP7_75t_SL g796 ( 
.A(n_656),
.B(n_49),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_595),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_669),
.A2(n_536),
.B1(n_534),
.B2(n_519),
.Y(n_798)
);

OAI22xp33_ASAP7_75t_SL g799 ( 
.A1(n_576),
.A2(n_548),
.B1(n_502),
.B2(n_52),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_604),
.Y(n_800)
);

OAI22xp33_ASAP7_75t_L g801 ( 
.A1(n_684),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_679),
.A2(n_548),
.B1(n_56),
.B2(n_58),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_599),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_680),
.A2(n_625),
.B1(n_694),
.B2(n_687),
.Y(n_804)
);

OAI22xp33_ASAP7_75t_L g805 ( 
.A1(n_691),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_624),
.B(n_87),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_595),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_596),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_607),
.Y(n_809)
);

OAI22xp33_ASAP7_75t_L g810 ( 
.A1(n_691),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_810)
);

OAI22xp33_ASAP7_75t_SL g811 ( 
.A1(n_707),
.A2(n_548),
.B1(n_61),
.B2(n_63),
.Y(n_811)
);

OAI22xp33_ASAP7_75t_SL g812 ( 
.A1(n_707),
.A2(n_548),
.B1(n_65),
.B2(n_66),
.Y(n_812)
);

INVxp33_ASAP7_75t_L g813 ( 
.A(n_584),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_574),
.Y(n_814)
);

XNOR2xp5_ASAP7_75t_L g815 ( 
.A(n_715),
.B(n_598),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_727),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_738),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_757),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_757),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_778),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_714),
.Y(n_821)
);

XNOR2x2_ASAP7_75t_L g822 ( 
.A(n_787),
.B(n_665),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_778),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_750),
.B(n_625),
.Y(n_824)
);

AND2x2_ASAP7_75t_SL g825 ( 
.A(n_796),
.B(n_654),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_728),
.B(n_594),
.Y(n_826)
);

XNOR2xp5_ASAP7_75t_L g827 ( 
.A(n_716),
.B(n_619),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_759),
.B(n_586),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_726),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_797),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_719),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_769),
.B(n_706),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_800),
.B(n_577),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_797),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_814),
.Y(n_835)
);

XNOR2xp5_ASAP7_75t_L g836 ( 
.A(n_721),
.B(n_632),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_809),
.B(n_706),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_732),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_747),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_733),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_734),
.Y(n_841)
);

INVxp33_ASAP7_75t_L g842 ( 
.A(n_724),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_806),
.B(n_654),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_740),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_772),
.B(n_606),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_752),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_735),
.B(n_606),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_773),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_736),
.B(n_611),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_749),
.B(n_577),
.Y(n_850)
);

CKINVDCx20_ASAP7_75t_R g851 ( 
.A(n_731),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_781),
.A2(n_661),
.B(n_567),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_751),
.B(n_611),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_779),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_791),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_718),
.Y(n_856)
);

AND2x2_ASAP7_75t_SL g857 ( 
.A(n_806),
.B(n_666),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_807),
.Y(n_858)
);

XOR2xp5_ASAP7_75t_L g859 ( 
.A(n_813),
.B(n_636),
.Y(n_859)
);

XOR2xp5_ASAP7_75t_L g860 ( 
.A(n_720),
.B(n_627),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_808),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_725),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_718),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_774),
.A2(n_661),
.B(n_567),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_785),
.B(n_804),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_742),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_741),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_767),
.B(n_577),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_786),
.B(n_583),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_739),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_741),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_746),
.B(n_706),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_771),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_793),
.B(n_666),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_761),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_795),
.B(n_682),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_761),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_760),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_765),
.Y(n_879)
);

XOR2xp5_ASAP7_75t_L g880 ( 
.A(n_798),
.B(n_627),
.Y(n_880)
);

XNOR2x2_ASAP7_75t_L g881 ( 
.A(n_787),
.B(n_665),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_717),
.B(n_630),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_744),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_789),
.B(n_615),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_744),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_765),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_782),
.B(n_583),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_717),
.B(n_630),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_768),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_754),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_754),
.Y(n_891)
);

XOR2xp5_ASAP7_75t_L g892 ( 
.A(n_776),
.B(n_722),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_762),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_783),
.B(n_583),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_789),
.B(n_615),
.Y(n_895)
);

INVxp33_ASAP7_75t_SL g896 ( 
.A(n_788),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_799),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_790),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_790),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_748),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_802),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_811),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_771),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_812),
.Y(n_904)
);

XOR2xp5_ASAP7_75t_L g905 ( 
.A(n_730),
.B(n_89),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_821),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_821),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_849),
.B(n_853),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_831),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_884),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_857),
.B(n_764),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_857),
.B(n_753),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_895),
.Y(n_913)
);

OR2x2_ASAP7_75t_L g914 ( 
.A(n_847),
.B(n_729),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_831),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_878),
.B(n_770),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_829),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_845),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_824),
.B(n_764),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_829),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_863),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_843),
.B(n_766),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_843),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_824),
.B(n_682),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_843),
.B(n_828),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_882),
.B(n_683),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_882),
.B(n_683),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_878),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_888),
.B(n_685),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_862),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_888),
.B(n_685),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_856),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_832),
.B(n_792),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_865),
.B(n_689),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_832),
.B(n_689),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_816),
.Y(n_936)
);

INVx8_ASAP7_75t_L g937 ( 
.A(n_873),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_817),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_837),
.B(n_690),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_825),
.A2(n_780),
.B1(n_784),
.B2(n_745),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_838),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_837),
.B(n_690),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_840),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_856),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_883),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_866),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_867),
.B(n_794),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_835),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_825),
.B(n_697),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_841),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_844),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_872),
.B(n_697),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_846),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_848),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_871),
.B(n_743),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_854),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_897),
.B(n_639),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_874),
.B(n_737),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_855),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_902),
.B(n_646),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_874),
.B(n_705),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_858),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_904),
.B(n_646),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_889),
.B(n_651),
.Y(n_964)
);

BUFx12f_ASAP7_75t_SL g965 ( 
.A(n_826),
.Y(n_965)
);

OAI21x1_ASAP7_75t_L g966 ( 
.A1(n_864),
.A2(n_608),
.B(n_607),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_883),
.B(n_885),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_876),
.B(n_705),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_870),
.B(n_651),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_870),
.B(n_664),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_861),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_818),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_876),
.A2(n_705),
.B(n_763),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_893),
.B(n_664),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_850),
.B(n_705),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_893),
.B(n_885),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_868),
.B(n_775),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_833),
.B(n_777),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_839),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_900),
.B(n_756),
.Y(n_980)
);

BUFx8_ASAP7_75t_L g981 ( 
.A(n_873),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_819),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_820),
.Y(n_983)
);

AND2x6_ASAP7_75t_L g984 ( 
.A(n_890),
.B(n_612),
.Y(n_984)
);

BUFx5_ASAP7_75t_L g985 ( 
.A(n_891),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_869),
.B(n_723),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_901),
.B(n_755),
.Y(n_987)
);

INVxp67_ASAP7_75t_SL g988 ( 
.A(n_823),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_839),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_830),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_898),
.B(n_673),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_899),
.B(n_673),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_834),
.B(n_620),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_887),
.B(n_711),
.Y(n_994)
);

INVxp67_ASAP7_75t_SL g995 ( 
.A(n_894),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_875),
.B(n_877),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_822),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_842),
.B(n_645),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_852),
.B(n_711),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_822),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_842),
.B(n_657),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_918),
.B(n_892),
.Y(n_1002)
);

INVx5_ASAP7_75t_L g1003 ( 
.A(n_945),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_924),
.B(n_896),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_945),
.Y(n_1005)
);

AND2x6_ASAP7_75t_L g1006 ( 
.A(n_949),
.B(n_873),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_923),
.B(n_879),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_907),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_SL g1009 ( 
.A(n_928),
.B(n_896),
.Y(n_1009)
);

BUFx12f_ASAP7_75t_L g1010 ( 
.A(n_981),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_945),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_918),
.B(n_881),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_923),
.B(n_886),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_908),
.B(n_880),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_907),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_937),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_908),
.B(n_873),
.Y(n_1017)
);

OR2x6_ASAP7_75t_L g1018 ( 
.A(n_937),
.B(n_903),
.Y(n_1018)
);

AOI21x1_ASAP7_75t_L g1019 ( 
.A1(n_975),
.A2(n_638),
.B(n_637),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_924),
.B(n_801),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_948),
.B(n_903),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_952),
.B(n_805),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_948),
.B(n_903),
.Y(n_1023)
);

BUFx4f_ASAP7_75t_L g1024 ( 
.A(n_937),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_914),
.B(n_881),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_952),
.B(n_810),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_909),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_945),
.Y(n_1028)
);

BUFx4f_ASAP7_75t_L g1029 ( 
.A(n_937),
.Y(n_1029)
);

CKINVDCx8_ASAP7_75t_R g1030 ( 
.A(n_937),
.Y(n_1030)
);

NAND2x1p5_ASAP7_75t_L g1031 ( 
.A(n_928),
.B(n_903),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_948),
.B(n_755),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_945),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_SL g1034 ( 
.A(n_928),
.B(n_851),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_920),
.Y(n_1035)
);

BUFx12f_ASAP7_75t_L g1036 ( 
.A(n_981),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_920),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_981),
.Y(n_1038)
);

BUFx12f_ASAP7_75t_L g1039 ( 
.A(n_981),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_967),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_909),
.Y(n_1041)
);

AND2x2_ASAP7_75t_SL g1042 ( 
.A(n_997),
.B(n_612),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_906),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_934),
.B(n_659),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_914),
.B(n_851),
.Y(n_1045)
);

BUFx8_ASAP7_75t_SL g1046 ( 
.A(n_989),
.Y(n_1046)
);

AND2x2_ASAP7_75t_SL g1047 ( 
.A(n_997),
.B(n_614),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_920),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_920),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_991),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_998),
.B(n_803),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_967),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_934),
.B(n_668),
.Y(n_1053)
);

INVx4_ASAP7_75t_L g1054 ( 
.A(n_967),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_998),
.B(n_758),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1001),
.B(n_815),
.Y(n_1056)
);

BUFx4f_ASAP7_75t_L g1057 ( 
.A(n_987),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_915),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_947),
.B(n_675),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1001),
.B(n_827),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_965),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_967),
.B(n_671),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_921),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_925),
.B(n_671),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_906),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_932),
.B(n_860),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_944),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_925),
.B(n_608),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_983),
.Y(n_1069)
);

OR2x6_ASAP7_75t_L g1070 ( 
.A(n_911),
.B(n_616),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_921),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_983),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_946),
.B(n_90),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_965),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_915),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_936),
.B(n_94),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_979),
.B(n_836),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_926),
.B(n_676),
.Y(n_1078)
);

NAND2xp33_ASAP7_75t_L g1079 ( 
.A(n_985),
.B(n_958),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_926),
.B(n_614),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_979),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_910),
.B(n_905),
.Y(n_1082)
);

NAND2x1p5_ASAP7_75t_L g1083 ( 
.A(n_1024),
.B(n_983),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1043),
.Y(n_1084)
);

INVx3_ASAP7_75t_SL g1085 ( 
.A(n_1081),
.Y(n_1085)
);

BUFx2_ASAP7_75t_SL g1086 ( 
.A(n_1038),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_1017),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1043),
.Y(n_1088)
);

BUFx2_ASAP7_75t_SL g1089 ( 
.A(n_1038),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1065),
.Y(n_1090)
);

AND2x6_ASAP7_75t_L g1091 ( 
.A(n_1040),
.B(n_911),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1055),
.B(n_913),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_1067),
.Y(n_1093)
);

BUFx5_ASAP7_75t_L g1094 ( 
.A(n_1011),
.Y(n_1094)
);

BUFx12f_ASAP7_75t_L g1095 ( 
.A(n_1010),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1075),
.Y(n_1096)
);

BUFx8_ASAP7_75t_L g1097 ( 
.A(n_1061),
.Y(n_1097)
);

BUFx4f_ASAP7_75t_SL g1098 ( 
.A(n_1036),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1075),
.Y(n_1099)
);

BUFx5_ASAP7_75t_L g1100 ( 
.A(n_1033),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1059),
.B(n_919),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_1016),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_1046),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_1018),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_1074),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1059),
.B(n_919),
.Y(n_1106)
);

BUFx2_ASAP7_75t_SL g1107 ( 
.A(n_1030),
.Y(n_1107)
);

CKINVDCx14_ASAP7_75t_R g1108 ( 
.A(n_1056),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1058),
.Y(n_1109)
);

INVx5_ASAP7_75t_L g1110 ( 
.A(n_1018),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1021),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_1067),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_1068),
.Y(n_1113)
);

BUFx4f_ASAP7_75t_SL g1114 ( 
.A(n_1039),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_1012),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_1040),
.Y(n_1116)
);

NAND2x1p5_ASAP7_75t_L g1117 ( 
.A(n_1024),
.B(n_983),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1051),
.B(n_1064),
.Y(n_1118)
);

INVxp67_ASAP7_75t_SL g1119 ( 
.A(n_1040),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_1046),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1008),
.Y(n_1121)
);

INVxp67_ASAP7_75t_SL g1122 ( 
.A(n_1040),
.Y(n_1122)
);

INVxp67_ASAP7_75t_SL g1123 ( 
.A(n_1069),
.Y(n_1123)
);

INVx5_ASAP7_75t_SL g1124 ( 
.A(n_1018),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1080),
.B(n_985),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1008),
.Y(n_1126)
);

INVx5_ASAP7_75t_L g1127 ( 
.A(n_1006),
.Y(n_1127)
);

NAND2x1p5_ASAP7_75t_L g1128 ( 
.A(n_1029),
.B(n_917),
.Y(n_1128)
);

BUFx10_ASAP7_75t_L g1129 ( 
.A(n_1032),
.Y(n_1129)
);

INVx8_ASAP7_75t_L g1130 ( 
.A(n_1003),
.Y(n_1130)
);

BUFx12f_ASAP7_75t_L g1131 ( 
.A(n_1032),
.Y(n_1131)
);

NOR2x1_ASAP7_75t_L g1132 ( 
.A(n_1016),
.B(n_916),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1080),
.B(n_985),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_1002),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_1021),
.Y(n_1135)
);

BUFx4f_ASAP7_75t_L g1136 ( 
.A(n_1006),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1015),
.Y(n_1137)
);

INVx4_ASAP7_75t_L g1138 ( 
.A(n_1003),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1027),
.Y(n_1139)
);

INVx1_ASAP7_75t_SL g1140 ( 
.A(n_1004),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_1004),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1052),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1027),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_1023),
.B(n_921),
.Y(n_1144)
);

INVx8_ASAP7_75t_L g1145 ( 
.A(n_1003),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_1052),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_1057),
.Y(n_1147)
);

BUFx12f_ASAP7_75t_L g1148 ( 
.A(n_1070),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1045),
.B(n_969),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1050),
.B(n_1007),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1041),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1041),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1109),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1084),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1088),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1126),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_SL g1157 ( 
.A1(n_1140),
.A2(n_1034),
.B1(n_1045),
.B2(n_1000),
.Y(n_1157)
);

NAND2x1p5_ASAP7_75t_L g1158 ( 
.A(n_1127),
.B(n_1029),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1149),
.A2(n_1025),
.B1(n_940),
.B2(n_1000),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1101),
.B(n_1022),
.Y(n_1160)
);

BUFx12f_ASAP7_75t_L g1161 ( 
.A(n_1097),
.Y(n_1161)
);

CKINVDCx6p67_ASAP7_75t_R g1162 ( 
.A(n_1085),
.Y(n_1162)
);

CKINVDCx11_ASAP7_75t_R g1163 ( 
.A(n_1095),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1104),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_SL g1165 ( 
.A1(n_1141),
.A2(n_1009),
.B1(n_1060),
.B2(n_1047),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1090),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1137),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_1093),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_1093),
.Y(n_1169)
);

BUFx10_ASAP7_75t_L g1170 ( 
.A(n_1103),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1143),
.Y(n_1171)
);

OAI22xp33_ASAP7_75t_R g1172 ( 
.A1(n_1134),
.A2(n_784),
.B1(n_780),
.B2(n_1066),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1096),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_SL g1174 ( 
.A1(n_1141),
.A2(n_1009),
.B1(n_1047),
.B2(n_1042),
.Y(n_1174)
);

BUFx4f_ASAP7_75t_SL g1175 ( 
.A(n_1131),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1134),
.A2(n_1014),
.B1(n_1082),
.B2(n_912),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_1097),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1127),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1118),
.A2(n_1042),
.B1(n_1057),
.B2(n_1073),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1099),
.Y(n_1180)
);

INVx6_ASAP7_75t_L g1181 ( 
.A(n_1129),
.Y(n_1181)
);

OAI22xp33_ASAP7_75t_SL g1182 ( 
.A1(n_1101),
.A2(n_1020),
.B1(n_1026),
.B2(n_1022),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1121),
.Y(n_1183)
);

OAI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1115),
.A2(n_987),
.B1(n_1077),
.B2(n_1020),
.Y(n_1184)
);

INVx6_ASAP7_75t_L g1185 ( 
.A(n_1129),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1113),
.A2(n_1073),
.B1(n_984),
.B2(n_933),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_SL g1187 ( 
.A1(n_1108),
.A2(n_1115),
.B1(n_1070),
.B2(n_1148),
.Y(n_1187)
);

CKINVDCx11_ASAP7_75t_R g1188 ( 
.A(n_1120),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1127),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_1112),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_SL g1191 ( 
.A1(n_1123),
.A2(n_1076),
.B(n_968),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1105),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1139),
.Y(n_1193)
);

INVxp67_ASAP7_75t_L g1194 ( 
.A(n_1112),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1151),
.Y(n_1195)
);

NAND2x1p5_ASAP7_75t_L g1196 ( 
.A(n_1110),
.B(n_1063),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_1111),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_SL g1198 ( 
.A1(n_1091),
.A2(n_973),
.B1(n_1026),
.B2(n_1006),
.Y(n_1198)
);

CKINVDCx11_ASAP7_75t_R g1199 ( 
.A(n_1104),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1092),
.B(n_1062),
.Y(n_1200)
);

BUFx4f_ASAP7_75t_L g1201 ( 
.A(n_1104),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1087),
.A2(n_984),
.B1(n_1006),
.B2(n_986),
.Y(n_1202)
);

BUFx4f_ASAP7_75t_SL g1203 ( 
.A(n_1147),
.Y(n_1203)
);

INVx6_ASAP7_75t_L g1204 ( 
.A(n_1110),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1152),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_1135),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1106),
.A2(n_955),
.B1(n_1071),
.B2(n_1063),
.Y(n_1207)
);

NAND2x1p5_ASAP7_75t_L g1208 ( 
.A(n_1110),
.B(n_1063),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1091),
.A2(n_984),
.B1(n_922),
.B2(n_995),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_1098),
.Y(n_1210)
);

INVx6_ASAP7_75t_L g1211 ( 
.A(n_1150),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1116),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1094),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1094),
.Y(n_1214)
);

INVx6_ASAP7_75t_L g1215 ( 
.A(n_1144),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1114),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1091),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1144),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1130),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1119),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1119),
.Y(n_1221)
);

INVx5_ASAP7_75t_L g1222 ( 
.A(n_1204),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1178),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_SL g1224 ( 
.A1(n_1157),
.A2(n_1091),
.B1(n_1136),
.B2(n_980),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_SL g1225 ( 
.A1(n_1157),
.A2(n_1086),
.B1(n_1089),
.B2(n_1123),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1153),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1165),
.A2(n_984),
.B1(n_939),
.B2(n_942),
.Y(n_1227)
);

OR2x2_ASAP7_75t_SL g1228 ( 
.A(n_1211),
.B(n_977),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1165),
.A2(n_1133),
.B1(n_1125),
.B2(n_1063),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_1210),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1188),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1174),
.A2(n_984),
.B1(n_978),
.B2(n_938),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1200),
.B(n_970),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_1162),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1174),
.A2(n_984),
.B1(n_938),
.B2(n_936),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_SL g1236 ( 
.A1(n_1187),
.A2(n_1124),
.B1(n_1107),
.B2(n_1079),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1159),
.B(n_970),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1184),
.A2(n_992),
.B1(n_991),
.B2(n_1007),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1172),
.A2(n_939),
.B1(n_942),
.B2(n_935),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1194),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1176),
.A2(n_992),
.B1(n_1013),
.B2(n_935),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1179),
.A2(n_859),
.B1(n_1070),
.B2(n_1013),
.Y(n_1242)
);

BUFx4f_ASAP7_75t_SL g1243 ( 
.A(n_1161),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_SL g1244 ( 
.A1(n_1182),
.A2(n_1124),
.B1(n_1079),
.B2(n_678),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1186),
.A2(n_1122),
.B1(n_1031),
.B2(n_1124),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_SL g1246 ( 
.A1(n_1217),
.A2(n_678),
.B1(n_644),
.B2(n_974),
.Y(n_1246)
);

CKINVDCx6p67_ASAP7_75t_R g1247 ( 
.A(n_1163),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_1177),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1198),
.A2(n_1044),
.B1(n_1053),
.B2(n_1132),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1218),
.B(n_1168),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1192),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1160),
.A2(n_644),
.B1(n_974),
.B2(n_961),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1154),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_1216),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1193),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1198),
.A2(n_1122),
.B1(n_1031),
.B2(n_1072),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1178),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_SL g1258 ( 
.A1(n_1160),
.A2(n_1169),
.B1(n_1190),
.B2(n_1168),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1170),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1169),
.B(n_976),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1190),
.B(n_969),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1206),
.B(n_994),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1206),
.B(n_976),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1155),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1209),
.A2(n_1202),
.B1(n_1197),
.B2(n_1207),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1199),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1194),
.A2(n_1069),
.B1(n_1072),
.B2(n_1128),
.Y(n_1267)
);

OAI21xp33_ASAP7_75t_L g1268 ( 
.A1(n_1191),
.A2(n_993),
.B(n_963),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1166),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1211),
.A2(n_1128),
.B1(n_1054),
.B2(n_1117),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1173),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_1175),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_SL g1273 ( 
.A1(n_1212),
.A2(n_996),
.B1(n_634),
.B2(n_963),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1201),
.A2(n_1054),
.B1(n_1117),
.B2(n_1083),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1180),
.Y(n_1275)
);

BUFx12f_ASAP7_75t_L g1276 ( 
.A(n_1170),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1215),
.A2(n_996),
.B1(n_960),
.B2(n_957),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1205),
.A2(n_930),
.B1(n_1078),
.B2(n_953),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1183),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1203),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1156),
.B(n_957),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1201),
.A2(n_1083),
.B1(n_1146),
.B2(n_1142),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1220),
.A2(n_1146),
.B1(n_1142),
.B2(n_1028),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1195),
.A2(n_943),
.B1(n_962),
.B2(n_953),
.Y(n_1284)
);

OAI21xp33_ASAP7_75t_L g1285 ( 
.A1(n_1221),
.A2(n_993),
.B(n_960),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1239),
.A2(n_1228),
.B1(n_1236),
.B2(n_1224),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1239),
.A2(n_1242),
.B1(n_1237),
.B2(n_1252),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1273),
.A2(n_1204),
.B1(n_1164),
.B2(n_1185),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1252),
.A2(n_996),
.B1(n_941),
.B2(n_951),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_SL g1290 ( 
.A1(n_1246),
.A2(n_996),
.B(n_1158),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1250),
.B(n_1167),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1240),
.B(n_1171),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_SL g1293 ( 
.A1(n_1268),
.A2(n_1158),
.B(n_1196),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1227),
.A2(n_950),
.B1(n_956),
.B2(n_951),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1227),
.A2(n_950),
.B1(n_959),
.B2(n_956),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1226),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1236),
.A2(n_1285),
.B1(n_1232),
.B2(n_1244),
.Y(n_1297)
);

AOI221xp5_ASAP7_75t_L g1298 ( 
.A1(n_1263),
.A2(n_959),
.B1(n_964),
.B2(n_990),
.C(n_972),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1245),
.A2(n_1164),
.B1(n_1181),
.B2(n_1189),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_SL g1300 ( 
.A1(n_1229),
.A2(n_1189),
.B1(n_1208),
.B2(n_1196),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1256),
.A2(n_1208),
.B1(n_1100),
.B2(n_1094),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1244),
.A2(n_971),
.B1(n_982),
.B2(n_990),
.Y(n_1302)
);

OAI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1261),
.A2(n_1214),
.B1(n_1213),
.B2(n_1219),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1233),
.A2(n_971),
.B1(n_982),
.B2(n_972),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1265),
.A2(n_971),
.B1(n_954),
.B2(n_548),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1225),
.A2(n_954),
.B1(n_1094),
.B2(n_1100),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1260),
.B(n_1094),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1243),
.A2(n_1266),
.B1(n_1276),
.B2(n_1222),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1225),
.A2(n_1238),
.B1(n_1241),
.B2(n_1246),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1281),
.A2(n_711),
.B1(n_713),
.B2(n_931),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1235),
.A2(n_954),
.B1(n_1100),
.B2(n_988),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1222),
.A2(n_1145),
.B1(n_1219),
.B2(n_1102),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1258),
.B(n_966),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1258),
.A2(n_954),
.B1(n_1028),
.B2(n_1005),
.Y(n_1314)
);

NAND3xp33_ASAP7_75t_L g1315 ( 
.A(n_1277),
.B(n_713),
.C(n_999),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_SL g1316 ( 
.A1(n_1222),
.A2(n_1102),
.B1(n_985),
.B2(n_964),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1262),
.A2(n_929),
.B1(n_927),
.B2(n_1048),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1253),
.Y(n_1318)
);

INVx6_ASAP7_75t_L g1319 ( 
.A(n_1251),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1255),
.B(n_966),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1249),
.A2(n_1037),
.B1(n_1049),
.B2(n_1035),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1234),
.A2(n_1259),
.B1(n_1272),
.B2(n_1230),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1264),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1284),
.A2(n_1138),
.B1(n_1019),
.B2(n_985),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1223),
.B(n_1257),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1274),
.A2(n_985),
.B1(n_708),
.B2(n_712),
.Y(n_1326)
);

AOI222xp33_ASAP7_75t_L g1327 ( 
.A1(n_1269),
.A2(n_708),
.B1(n_701),
.B2(n_712),
.C1(n_70),
.C2(n_71),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1248),
.A2(n_1270),
.B1(n_1247),
.B2(n_1282),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1267),
.A2(n_701),
.B1(n_700),
.B2(n_699),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1223),
.A2(n_1257),
.B1(n_1275),
.B2(n_1279),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_SL g1331 ( 
.A1(n_1231),
.A2(n_60),
.B1(n_66),
.B2(n_69),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1278),
.A2(n_585),
.B1(n_589),
.B2(n_605),
.Y(n_1332)
);

NOR3xp33_ASAP7_75t_L g1333 ( 
.A(n_1283),
.B(n_70),
.C(n_73),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1271),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1280),
.B(n_95),
.Y(n_1335)
);

OAI222xp33_ASAP7_75t_L g1336 ( 
.A1(n_1254),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.C1(n_79),
.C2(n_80),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1239),
.A2(n_585),
.B1(n_589),
.B2(n_605),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1273),
.A2(n_652),
.B1(n_699),
.B2(n_698),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_SL g1339 ( 
.A1(n_1273),
.A2(n_631),
.B1(n_698),
.B2(n_696),
.Y(n_1339)
);

AOI221xp5_ASAP7_75t_L g1340 ( 
.A1(n_1239),
.A2(n_700),
.B1(n_696),
.B2(n_692),
.C(n_653),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1224),
.A2(n_696),
.B1(n_626),
.B2(n_692),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1250),
.B(n_82),
.Y(n_1342)
);

INVx4_ASAP7_75t_L g1343 ( 
.A(n_1222),
.Y(n_1343)
);

OAI211xp5_ASAP7_75t_SL g1344 ( 
.A1(n_1252),
.A2(n_82),
.B(n_83),
.C(n_84),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1296),
.B(n_83),
.Y(n_1345)
);

NAND3xp33_ASAP7_75t_L g1346 ( 
.A(n_1327),
.B(n_597),
.C(n_601),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1286),
.B(n_84),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1318),
.B(n_100),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1291),
.B(n_597),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_SL g1350 ( 
.A1(n_1287),
.A2(n_653),
.B(n_652),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1344),
.A2(n_693),
.B(n_670),
.Y(n_1351)
);

NAND3xp33_ASAP7_75t_L g1352 ( 
.A(n_1333),
.B(n_631),
.C(n_601),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1309),
.A2(n_631),
.B1(n_601),
.B2(n_602),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1292),
.B(n_602),
.Y(n_1354)
);

NOR3xp33_ASAP7_75t_L g1355 ( 
.A(n_1336),
.B(n_102),
.C(n_103),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1334),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1290),
.A2(n_652),
.B1(n_602),
.B2(n_609),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1288),
.B(n_1303),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1307),
.B(n_1323),
.Y(n_1359)
);

OAI221xp5_ASAP7_75t_L g1360 ( 
.A1(n_1289),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.C(n_117),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1342),
.B(n_118),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1325),
.B(n_119),
.Y(n_1362)
);

OAI21xp33_ASAP7_75t_L g1363 ( 
.A1(n_1297),
.A2(n_120),
.B(n_122),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1330),
.B(n_129),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1320),
.B(n_1299),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1328),
.B(n_140),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1303),
.B(n_142),
.Y(n_1367)
);

OAI221xp5_ASAP7_75t_SL g1368 ( 
.A1(n_1302),
.A2(n_146),
.B1(n_147),
.B2(n_149),
.C(n_152),
.Y(n_1368)
);

NAND3xp33_ASAP7_75t_L g1369 ( 
.A(n_1331),
.B(n_617),
.C(n_661),
.Y(n_1369)
);

OAI221xp5_ASAP7_75t_L g1370 ( 
.A1(n_1338),
.A2(n_153),
.B1(n_154),
.B2(n_156),
.C(n_157),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1300),
.B(n_158),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1313),
.B(n_162),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_SL g1373 ( 
.A1(n_1337),
.A2(n_165),
.B(n_167),
.Y(n_1373)
);

OAI21xp33_ASAP7_75t_L g1374 ( 
.A1(n_1339),
.A2(n_168),
.B(n_172),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1319),
.B(n_1306),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1319),
.B(n_174),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1298),
.B(n_617),
.C(n_567),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1319),
.B(n_1301),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_SL g1379 ( 
.A(n_1343),
.B(n_181),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1341),
.A2(n_1308),
.B1(n_1294),
.B2(n_1295),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1312),
.B(n_182),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1305),
.B(n_183),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1317),
.B(n_184),
.Y(n_1383)
);

NAND4xp25_ASAP7_75t_L g1384 ( 
.A(n_1340),
.B(n_186),
.C(n_187),
.D(n_190),
.Y(n_1384)
);

NOR3xp33_ASAP7_75t_L g1385 ( 
.A(n_1315),
.B(n_191),
.C(n_192),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1304),
.B(n_194),
.Y(n_1386)
);

NAND3xp33_ASAP7_75t_L g1387 ( 
.A(n_1310),
.B(n_195),
.C(n_196),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1343),
.B(n_197),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1310),
.B(n_1314),
.Y(n_1389)
);

NAND3xp33_ASAP7_75t_L g1390 ( 
.A(n_1293),
.B(n_200),
.C(n_202),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1322),
.B(n_1311),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1321),
.B(n_208),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1335),
.B(n_209),
.Y(n_1393)
);

NAND3xp33_ASAP7_75t_L g1394 ( 
.A(n_1347),
.B(n_1316),
.C(n_1329),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1358),
.B(n_1326),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1356),
.B(n_1324),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1359),
.B(n_1332),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1378),
.B(n_213),
.Y(n_1398)
);

NOR3xp33_ASAP7_75t_L g1399 ( 
.A(n_1346),
.B(n_215),
.C(n_217),
.Y(n_1399)
);

NAND3xp33_ASAP7_75t_L g1400 ( 
.A(n_1355),
.B(n_221),
.C(n_225),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1363),
.A2(n_228),
.B1(n_230),
.B2(n_233),
.Y(n_1401)
);

NAND3xp33_ASAP7_75t_L g1402 ( 
.A(n_1358),
.B(n_237),
.C(n_239),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1375),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_L g1404 ( 
.A(n_1369),
.B(n_241),
.C(n_247),
.Y(n_1404)
);

AOI221xp5_ASAP7_75t_L g1405 ( 
.A1(n_1350),
.A2(n_1353),
.B1(n_1368),
.B2(n_1365),
.C(n_1352),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1345),
.B(n_249),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1354),
.B(n_253),
.Y(n_1407)
);

AO21x2_ASAP7_75t_L g1408 ( 
.A1(n_1372),
.A2(n_259),
.B(n_260),
.Y(n_1408)
);

NOR3xp33_ASAP7_75t_L g1409 ( 
.A(n_1390),
.B(n_261),
.C(n_266),
.Y(n_1409)
);

NAND4xp75_ASAP7_75t_L g1410 ( 
.A(n_1366),
.B(n_270),
.C(n_271),
.D(n_274),
.Y(n_1410)
);

AO21x2_ASAP7_75t_L g1411 ( 
.A1(n_1385),
.A2(n_277),
.B(n_280),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1349),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1379),
.B(n_295),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1391),
.B(n_296),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1361),
.B(n_298),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1348),
.B(n_303),
.Y(n_1416)
);

NAND4xp75_ASAP7_75t_L g1417 ( 
.A(n_1381),
.B(n_312),
.C(n_313),
.D(n_317),
.Y(n_1417)
);

AO21x2_ASAP7_75t_L g1418 ( 
.A1(n_1385),
.A2(n_318),
.B(n_319),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1367),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1362),
.B(n_320),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1357),
.B(n_321),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1376),
.B(n_322),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1412),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1395),
.A2(n_1380),
.B1(n_1384),
.B2(n_1374),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1396),
.Y(n_1425)
);

NAND3xp33_ASAP7_75t_SL g1426 ( 
.A(n_1395),
.B(n_1405),
.C(n_1400),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1396),
.Y(n_1427)
);

INVxp67_ASAP7_75t_L g1428 ( 
.A(n_1403),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1419),
.B(n_1371),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1398),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1419),
.B(n_1364),
.Y(n_1431)
);

XNOR2xp5_ASAP7_75t_L g1432 ( 
.A(n_1398),
.B(n_1393),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1397),
.B(n_1389),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1411),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1408),
.B(n_1388),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1408),
.B(n_1377),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1408),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1411),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1411),
.B(n_1383),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1418),
.B(n_1373),
.Y(n_1440)
);

NAND4xp75_ASAP7_75t_L g1441 ( 
.A(n_1413),
.B(n_1351),
.C(n_1386),
.D(n_1392),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1418),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1418),
.B(n_1387),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1414),
.B(n_1382),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1415),
.B(n_1360),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1407),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1406),
.B(n_328),
.Y(n_1447)
);

INVx2_ASAP7_75t_SL g1448 ( 
.A(n_1422),
.Y(n_1448)
);

XOR2x2_ASAP7_75t_L g1449 ( 
.A(n_1410),
.B(n_1370),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1422),
.B(n_332),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1423),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1425),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1425),
.Y(n_1453)
);

INVxp67_ASAP7_75t_L g1454 ( 
.A(n_1433),
.Y(n_1454)
);

XNOR2xp5_ASAP7_75t_L g1455 ( 
.A(n_1426),
.B(n_1420),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1427),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1427),
.Y(n_1457)
);

XNOR2xp5_ASAP7_75t_L g1458 ( 
.A(n_1432),
.B(n_1449),
.Y(n_1458)
);

INVx1_ASAP7_75t_SL g1459 ( 
.A(n_1430),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1437),
.Y(n_1460)
);

XOR2x2_ASAP7_75t_L g1461 ( 
.A(n_1424),
.B(n_1394),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1433),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1437),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1432),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1446),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1448),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1434),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1428),
.B(n_1420),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1448),
.Y(n_1469)
);

INVx1_ASAP7_75t_SL g1470 ( 
.A(n_1429),
.Y(n_1470)
);

XNOR2x2_ASAP7_75t_L g1471 ( 
.A(n_1449),
.B(n_1402),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1445),
.A2(n_1409),
.B1(n_1399),
.B2(n_1417),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1463),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1467),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1467),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1467),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1452),
.Y(n_1477)
);

AOI22x1_ASAP7_75t_L g1478 ( 
.A1(n_1458),
.A2(n_1434),
.B1(n_1440),
.B2(n_1443),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1452),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1451),
.Y(n_1480)
);

XOR2x2_ASAP7_75t_L g1481 ( 
.A(n_1458),
.B(n_1424),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1464),
.A2(n_1443),
.B1(n_1434),
.B2(n_1439),
.Y(n_1482)
);

AOI22x1_ASAP7_75t_L g1483 ( 
.A1(n_1455),
.A2(n_1440),
.B1(n_1443),
.B2(n_1439),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1453),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1453),
.Y(n_1485)
);

INVx5_ASAP7_75t_L g1486 ( 
.A(n_1461),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1468),
.Y(n_1487)
);

OA22x2_ASAP7_75t_L g1488 ( 
.A1(n_1455),
.A2(n_1442),
.B1(n_1435),
.B2(n_1438),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1472),
.A2(n_1442),
.B1(n_1438),
.B2(n_1436),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1454),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1457),
.Y(n_1491)
);

XNOR2x1_ASAP7_75t_L g1492 ( 
.A(n_1461),
.B(n_1441),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1459),
.A2(n_1441),
.B1(n_1435),
.B2(n_1444),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1480),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1490),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1490),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1477),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1487),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1486),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1479),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1485),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1491),
.Y(n_1502)
);

INVx2_ASAP7_75t_SL g1503 ( 
.A(n_1487),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1473),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1499),
.A2(n_1486),
.B1(n_1492),
.B2(n_1481),
.Y(n_1505)
);

AOI22x1_ASAP7_75t_L g1506 ( 
.A1(n_1498),
.A2(n_1486),
.B1(n_1503),
.B2(n_1496),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1495),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1494),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1497),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1500),
.Y(n_1510)
);

INVx8_ASAP7_75t_L g1511 ( 
.A(n_1499),
.Y(n_1511)
);

INVxp67_ASAP7_75t_L g1512 ( 
.A(n_1503),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1501),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1505),
.B(n_1486),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1512),
.B(n_1502),
.Y(n_1515)
);

AOI221x1_ASAP7_75t_SL g1516 ( 
.A1(n_1507),
.A2(n_1493),
.B1(n_1482),
.B2(n_1489),
.C(n_1504),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1509),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1508),
.Y(n_1518)
);

OAI31xp33_ASAP7_75t_L g1519 ( 
.A1(n_1506),
.A2(n_1493),
.A3(n_1482),
.B(n_1489),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1511),
.A2(n_1483),
.B1(n_1478),
.B2(n_1488),
.Y(n_1520)
);

OAI22x1_ASAP7_75t_L g1521 ( 
.A1(n_1510),
.A2(n_1469),
.B1(n_1471),
.B2(n_1476),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1518),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1514),
.A2(n_1488),
.B1(n_1511),
.B2(n_1513),
.Y(n_1523)
);

AO22x2_ASAP7_75t_L g1524 ( 
.A1(n_1517),
.A2(n_1475),
.B1(n_1474),
.B2(n_1473),
.Y(n_1524)
);

AOI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1520),
.A2(n_1462),
.B1(n_1466),
.B2(n_1446),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1518),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1515),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1521),
.Y(n_1528)
);

INVxp67_ASAP7_75t_SL g1529 ( 
.A(n_1522),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1526),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1524),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1527),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1529),
.Y(n_1533)
);

AO22x2_ASAP7_75t_L g1534 ( 
.A1(n_1530),
.A2(n_1528),
.B1(n_1516),
.B2(n_1519),
.Y(n_1534)
);

AOI221xp5_ASAP7_75t_SL g1535 ( 
.A1(n_1531),
.A2(n_1523),
.B1(n_1525),
.B2(n_1471),
.C(n_1460),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1530),
.A2(n_1484),
.B(n_1465),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1533),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1534),
.A2(n_1532),
.B1(n_1469),
.B2(n_1468),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1536),
.Y(n_1539)
);

INVxp67_ASAP7_75t_SL g1540 ( 
.A(n_1538),
.Y(n_1540)
);

OAI22x1_ASAP7_75t_L g1541 ( 
.A1(n_1537),
.A2(n_1534),
.B1(n_1535),
.B2(n_1532),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_SL g1542 ( 
.A1(n_1539),
.A2(n_1447),
.B1(n_1450),
.B2(n_1484),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1541),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1542),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1540),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1545),
.A2(n_1447),
.B1(n_1450),
.B2(n_1415),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1543),
.A2(n_1457),
.B1(n_1470),
.B2(n_1456),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1546),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1547),
.Y(n_1549)
);

OAI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1549),
.A2(n_1544),
.B1(n_1404),
.B2(n_1401),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1550),
.Y(n_1551)
);

AO22x2_ASAP7_75t_L g1552 ( 
.A1(n_1551),
.A2(n_1548),
.B1(n_1421),
.B2(n_1416),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1552),
.A2(n_1416),
.B1(n_1429),
.B2(n_1431),
.Y(n_1553)
);


endmodule