module fake_jpeg_25699_n_162 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_25),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_22),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_33),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_10),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_66),
.Y(n_79)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_0),
.C(n_1),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_0),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_54),
.B1(n_46),
.B2(n_49),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_74),
.A2(n_78),
.B1(n_56),
.B2(n_50),
.Y(n_99)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

CKINVDCx6p67_ASAP7_75t_R g102 ( 
.A(n_77),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_54),
.B1(n_46),
.B2(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_86),
.Y(n_87)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_88),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_57),
.B1(n_44),
.B2(n_60),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_94),
.B1(n_96),
.B2(n_98),
.Y(n_109)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_91),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_77),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_79),
.A2(n_47),
.B1(n_53),
.B2(n_81),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_64),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_3),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_82),
.A2(n_57),
.B1(n_59),
.B2(n_58),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_52),
.B1(n_45),
.B2(n_61),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_100),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_61),
.B1(n_56),
.B2(n_50),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_2),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_48),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_111),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_2),
.B(n_3),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_4),
.B(n_6),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_102),
.B1(n_7),
.B2(n_8),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_113),
.B(n_4),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_106),
.A2(n_89),
.B1(n_95),
.B2(n_90),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_101),
.B1(n_10),
.B2(n_11),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_102),
.C(n_109),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_31),
.C(n_42),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_118),
.B(n_119),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_12),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_6),
.B(n_7),
.C(n_9),
.Y(n_121)
);

HAxp5_ASAP7_75t_SL g125 ( 
.A(n_121),
.B(n_110),
.CON(n_125),
.SN(n_125)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_130),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_114),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_126),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_135),
.Y(n_143)
);

NAND2x1_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_9),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_134),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_121),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_131),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_119),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_135)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_137),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_17),
.B1(n_19),
.B2(n_23),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_147),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_132),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_128),
.C(n_134),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_129),
.C(n_141),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_139),
.B1(n_133),
.B2(n_124),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_153),
.A2(n_130),
.B(n_148),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_149),
.Y(n_156)
);

NOR2xp67_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_145),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_142),
.B(n_144),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_146),
.A3(n_125),
.B1(n_143),
.B2(n_151),
.C1(n_35),
.C2(n_38),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_160),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_30),
.Y(n_162)
);


endmodule