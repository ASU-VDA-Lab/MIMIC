module real_aes_7447_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_1), .A2(n_104), .B1(n_115), .B2(n_751), .Y(n_103) );
INVx1_ASAP7_75t_L g514 ( .A(n_2), .Y(n_514) );
INVx1_ASAP7_75t_L g155 ( .A(n_3), .Y(n_155) );
OAI22xp5_ASAP7_75t_SL g738 ( .A1(n_4), .A2(n_739), .B1(n_742), .B2(n_743), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_4), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g125 ( .A1(n_5), .A2(n_126), .B1(n_127), .B2(n_450), .Y(n_125) );
INVx1_ASAP7_75t_L g450 ( .A(n_5), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_6), .A2(n_41), .B1(n_180), .B2(n_470), .Y(n_499) );
AOI21xp33_ASAP7_75t_L g199 ( .A1(n_7), .A2(n_171), .B(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_8), .B(n_169), .Y(n_525) );
AND2x6_ASAP7_75t_L g148 ( .A(n_9), .B(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_10), .A2(n_253), .B(n_254), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_11), .B(n_42), .Y(n_114) );
INVx1_ASAP7_75t_L g205 ( .A(n_12), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_13), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g140 ( .A(n_14), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_15), .B(n_161), .Y(n_478) );
INVx1_ASAP7_75t_L g259 ( .A(n_16), .Y(n_259) );
INVx1_ASAP7_75t_L g508 ( .A(n_17), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_18), .B(n_136), .Y(n_530) );
AO32x2_ASAP7_75t_L g497 ( .A1(n_19), .A2(n_135), .A3(n_169), .B1(n_472), .B2(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_20), .B(n_180), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_21), .B(n_176), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_22), .B(n_136), .Y(n_516) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_23), .A2(n_34), .B1(n_447), .B2(n_448), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_23), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_24), .A2(n_53), .B1(n_180), .B2(n_470), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_25), .B(n_171), .Y(n_216) );
AOI22xp33_ASAP7_75t_SL g471 ( .A1(n_26), .A2(n_79), .B1(n_161), .B2(n_180), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_27), .B(n_180), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_28), .B(n_183), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_29), .A2(n_257), .B(n_258), .C(n_260), .Y(n_256) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_30), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_31), .B(n_166), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_32), .B(n_159), .Y(n_158) );
AOI222xp33_ASAP7_75t_L g455 ( .A1(n_33), .A2(n_456), .B1(n_738), .B2(n_744), .C1(n_747), .C2(n_748), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_34), .Y(n_448) );
INVx1_ASAP7_75t_L g194 ( .A(n_35), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_36), .B(n_166), .Y(n_495) );
INVx2_ASAP7_75t_L g146 ( .A(n_37), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_38), .B(n_180), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_39), .B(n_166), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_40), .A2(n_148), .B(n_151), .C(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g192 ( .A(n_43), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_44), .B(n_159), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_45), .B(n_180), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_46), .B(n_452), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_47), .A2(n_89), .B1(n_223), .B2(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_48), .B(n_180), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_49), .B(n_180), .Y(n_509) );
CKINVDCx16_ASAP7_75t_R g195 ( .A(n_50), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_51), .B(n_513), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_52), .B(n_171), .Y(n_236) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_54), .A2(n_63), .B1(n_161), .B2(n_180), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_55), .A2(n_151), .B1(n_161), .B2(n_190), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_56), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_57), .B(n_180), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g142 ( .A(n_58), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_59), .B(n_180), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_60), .A2(n_179), .B(n_203), .C(n_204), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_61), .Y(n_250) );
INVx1_ASAP7_75t_L g201 ( .A(n_62), .Y(n_201) );
INVx1_ASAP7_75t_L g149 ( .A(n_64), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_65), .B(n_180), .Y(n_515) );
INVx1_ASAP7_75t_L g139 ( .A(n_66), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_67), .Y(n_120) );
AO32x2_ASAP7_75t_L g467 ( .A1(n_68), .A2(n_169), .A3(n_228), .B1(n_468), .B2(n_472), .Y(n_467) );
INVx1_ASAP7_75t_L g547 ( .A(n_69), .Y(n_547) );
INVx1_ASAP7_75t_L g490 ( .A(n_70), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_71), .A2(n_78), .B1(n_740), .B2(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_71), .Y(n_741) );
A2O1A1Ixp33_ASAP7_75t_SL g175 ( .A1(n_72), .A2(n_176), .B(n_177), .C(n_179), .Y(n_175) );
INVxp67_ASAP7_75t_L g178 ( .A(n_73), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_74), .B(n_161), .Y(n_491) );
INVx1_ASAP7_75t_L g108 ( .A(n_75), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_76), .Y(n_197) );
INVx1_ASAP7_75t_L g243 ( .A(n_77), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_78), .Y(n_740) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_80), .A2(n_148), .B(n_151), .C(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_81), .B(n_470), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_82), .B(n_161), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_83), .B(n_156), .Y(n_219) );
INVx2_ASAP7_75t_L g137 ( .A(n_84), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_85), .B(n_176), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_86), .B(n_161), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_87), .A2(n_148), .B(n_151), .C(n_154), .Y(n_150) );
OR2x2_ASAP7_75t_L g110 ( .A(n_88), .B(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g459 ( .A(n_88), .B(n_112), .Y(n_459) );
INVx2_ASAP7_75t_L g737 ( .A(n_88), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_90), .A2(n_102), .B1(n_161), .B2(n_162), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_91), .B(n_166), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_92), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_93), .A2(n_148), .B(n_151), .C(n_231), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_94), .Y(n_238) );
INVx1_ASAP7_75t_L g174 ( .A(n_95), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_96), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_97), .B(n_156), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_98), .B(n_161), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_99), .B(n_169), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_100), .B(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_101), .A2(n_171), .B(n_172), .Y(n_170) );
CKINVDCx6p67_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g752 ( .A(n_105), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_SL g124 ( .A(n_110), .Y(n_124) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_110), .Y(n_453) );
NOR2x2_ASAP7_75t_L g750 ( .A(n_111), .B(n_737), .Y(n_750) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g736 ( .A(n_112), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_454), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
NAND3xp33_ASAP7_75t_L g454 ( .A(n_117), .B(n_451), .C(n_455), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_125), .B(n_451), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_445), .B1(n_446), .B2(n_449), .Y(n_127) );
INVx2_ASAP7_75t_L g449 ( .A(n_128), .Y(n_449) );
OAI22xp5_ASAP7_75t_SL g456 ( .A1(n_128), .A2(n_457), .B1(n_460), .B2(n_734), .Y(n_456) );
OR4x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_334), .C(n_394), .D(n_421), .Y(n_128) );
NAND4xp25_ASAP7_75t_SL g129 ( .A(n_130), .B(n_282), .C(n_313), .D(n_330), .Y(n_129) );
O2A1O1Ixp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_207), .B(n_209), .C(n_262), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_185), .Y(n_131) );
INVx1_ASAP7_75t_L g324 ( .A(n_132), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_132), .A2(n_365), .B1(n_413), .B2(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_167), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_133), .B(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g275 ( .A(n_133), .B(n_187), .Y(n_275) );
AND2x2_ASAP7_75t_L g317 ( .A(n_133), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_133), .B(n_208), .Y(n_329) );
INVx1_ASAP7_75t_L g369 ( .A(n_133), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_133), .B(n_423), .Y(n_422) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g297 ( .A(n_134), .B(n_187), .Y(n_297) );
INVx3_ASAP7_75t_L g301 ( .A(n_134), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_134), .B(n_359), .Y(n_358) );
AO21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_141), .B(n_163), .Y(n_134) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_135), .A2(n_188), .B(n_196), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_135), .B(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g224 ( .A(n_135), .Y(n_224) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_136), .Y(n_169) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_137), .B(n_138), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
OAI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_150), .Y(n_141) );
OAI22xp33_ASAP7_75t_L g188 ( .A1(n_143), .A2(n_181), .B1(n_189), .B2(n_195), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g242 ( .A1(n_143), .A2(n_243), .B(n_244), .Y(n_242) );
NAND2x1p5_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
AND2x4_ASAP7_75t_L g171 ( .A(n_144), .B(n_148), .Y(n_171) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx1_ASAP7_75t_L g513 ( .A(n_145), .Y(n_513) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g152 ( .A(n_146), .Y(n_152) );
INVx1_ASAP7_75t_L g162 ( .A(n_146), .Y(n_162) );
INVx1_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx3_ASAP7_75t_L g157 ( .A(n_147), .Y(n_157) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_147), .Y(n_159) );
INVx1_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_147), .Y(n_191) );
INVx4_ASAP7_75t_SL g181 ( .A(n_148), .Y(n_181) );
BUFx3_ASAP7_75t_L g472 ( .A(n_148), .Y(n_472) );
OAI21xp5_ASAP7_75t_L g475 ( .A1(n_148), .A2(n_476), .B(n_480), .Y(n_475) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_148), .A2(n_489), .B(n_492), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_148), .A2(n_507), .B(n_511), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_148), .A2(n_519), .B(n_522), .Y(n_518) );
INVx5_ASAP7_75t_L g173 ( .A(n_151), .Y(n_173) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
BUFx3_ASAP7_75t_L g223 ( .A(n_152), .Y(n_223) );
INVx1_ASAP7_75t_L g470 ( .A(n_152), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_158), .C(n_160), .Y(n_154) );
O2A1O1Ixp5_ASAP7_75t_SL g489 ( .A1(n_156), .A2(n_179), .B(n_490), .C(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g500 ( .A(n_156), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_156), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_156), .A2(n_544), .B(n_545), .Y(n_543) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_157), .B(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_157), .B(n_205), .Y(n_204) );
OAI22xp5_ASAP7_75t_SL g468 ( .A1(n_157), .A2(n_159), .B1(n_469), .B2(n_471), .Y(n_468) );
INVx2_ASAP7_75t_L g203 ( .A(n_159), .Y(n_203) );
INVx4_ASAP7_75t_L g234 ( .A(n_159), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_159), .A2(n_499), .B1(n_500), .B2(n_501), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_159), .A2(n_500), .B1(n_533), .B2(n_534), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_160), .A2(n_508), .B(n_509), .C(n_510), .Y(n_507) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_165), .B(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_165), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g228 ( .A(n_166), .Y(n_228) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_166), .A2(n_252), .B(n_261), .Y(n_251) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_166), .A2(n_475), .B(n_483), .Y(n_474) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_166), .A2(n_488), .B(n_495), .Y(n_487) );
AND2x2_ASAP7_75t_L g388 ( .A(n_167), .B(n_198), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_167), .B(n_301), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_167), .B(n_416), .Y(n_415) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g208 ( .A(n_168), .B(n_187), .Y(n_208) );
INVx1_ASAP7_75t_L g270 ( .A(n_168), .Y(n_270) );
BUFx2_ASAP7_75t_L g274 ( .A(n_168), .Y(n_274) );
AND2x2_ASAP7_75t_L g318 ( .A(n_168), .B(n_186), .Y(n_318) );
OR2x2_ASAP7_75t_L g357 ( .A(n_168), .B(n_186), .Y(n_357) );
AND2x2_ASAP7_75t_L g382 ( .A(n_168), .B(n_198), .Y(n_382) );
AND2x2_ASAP7_75t_L g441 ( .A(n_168), .B(n_271), .Y(n_441) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_182), .Y(n_168) );
INVx4_ASAP7_75t_L g184 ( .A(n_169), .Y(n_184) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_169), .A2(n_518), .B(n_525), .Y(n_517) );
BUFx2_ASAP7_75t_L g253 ( .A(n_171), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_175), .C(n_181), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_173), .A2(n_181), .B(n_201), .C(n_202), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_173), .A2(n_181), .B(n_255), .C(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g479 ( .A(n_176), .Y(n_479) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_180), .Y(n_235) );
OA21x2_ASAP7_75t_L g198 ( .A1(n_183), .A2(n_199), .B(n_206), .Y(n_198) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_SL g225 ( .A(n_184), .B(n_226), .Y(n_225) );
NAND3xp33_ASAP7_75t_L g531 ( .A(n_184), .B(n_472), .C(n_532), .Y(n_531) );
AO21x1_ASAP7_75t_L g578 ( .A1(n_184), .A2(n_532), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g416 ( .A(n_185), .Y(n_416) );
OR2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_198), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_186), .B(n_198), .Y(n_302) );
AND2x2_ASAP7_75t_L g312 ( .A(n_186), .B(n_301), .Y(n_312) );
BUFx2_ASAP7_75t_L g323 ( .A(n_186), .Y(n_323) );
INVx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g345 ( .A(n_187), .B(n_198), .Y(n_345) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_187), .Y(n_400) );
OAI22xp5_ASAP7_75t_SL g190 ( .A1(n_191), .A2(n_192), .B1(n_193), .B2(n_194), .Y(n_190) );
INVx2_ASAP7_75t_L g193 ( .A(n_191), .Y(n_193) );
INVx4_ASAP7_75t_L g257 ( .A(n_191), .Y(n_257) );
AND2x2_ASAP7_75t_SL g207 ( .A(n_198), .B(n_208), .Y(n_207) );
INVx1_ASAP7_75t_SL g271 ( .A(n_198), .Y(n_271) );
BUFx2_ASAP7_75t_L g296 ( .A(n_198), .Y(n_296) );
INVx2_ASAP7_75t_L g315 ( .A(n_198), .Y(n_315) );
AND2x2_ASAP7_75t_L g377 ( .A(n_198), .B(n_301), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_203), .A2(n_481), .B(n_482), .Y(n_480) );
O2A1O1Ixp5_ASAP7_75t_L g546 ( .A1(n_203), .A2(n_512), .B(n_547), .C(n_548), .Y(n_546) );
AOI321xp33_ASAP7_75t_L g396 ( .A1(n_207), .A2(n_397), .A3(n_398), .B1(n_399), .B2(n_401), .C(n_402), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_208), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_208), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g390 ( .A(n_208), .B(n_369), .Y(n_390) );
AND2x2_ASAP7_75t_L g423 ( .A(n_208), .B(n_315), .Y(n_423) );
INVx1_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_239), .Y(n_210) );
OR2x2_ASAP7_75t_L g325 ( .A(n_211), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_227), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx3_ASAP7_75t_L g277 ( .A(n_214), .Y(n_277) );
AND2x2_ASAP7_75t_L g287 ( .A(n_214), .B(n_241), .Y(n_287) );
AND2x2_ASAP7_75t_L g292 ( .A(n_214), .B(n_267), .Y(n_292) );
INVx1_ASAP7_75t_L g309 ( .A(n_214), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_214), .B(n_290), .Y(n_328) );
AND2x2_ASAP7_75t_L g333 ( .A(n_214), .B(n_266), .Y(n_333) );
OR2x2_ASAP7_75t_L g365 ( .A(n_214), .B(n_354), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_214), .B(n_278), .Y(n_404) );
AND2x2_ASAP7_75t_L g438 ( .A(n_214), .B(n_264), .Y(n_438) );
OR2x6_ASAP7_75t_L g214 ( .A(n_215), .B(n_225), .Y(n_214) );
AOI21xp5_ASAP7_75t_SL g215 ( .A1(n_216), .A2(n_217), .B(n_224), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_221), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_221), .A2(n_246), .B(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g260 ( .A(n_223), .Y(n_260) );
INVx1_ASAP7_75t_L g248 ( .A(n_224), .Y(n_248) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_224), .A2(n_506), .B(n_516), .Y(n_505) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_224), .A2(n_542), .B(n_549), .Y(n_541) );
INVx1_ASAP7_75t_L g265 ( .A(n_227), .Y(n_265) );
INVx2_ASAP7_75t_L g280 ( .A(n_227), .Y(n_280) );
AND2x2_ASAP7_75t_L g320 ( .A(n_227), .B(n_291), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_227), .B(n_267), .Y(n_342) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_237), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_236), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_235), .Y(n_231) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g426 ( .A(n_240), .B(n_277), .Y(n_426) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_251), .Y(n_240) );
INVx2_ASAP7_75t_L g267 ( .A(n_241), .Y(n_267) );
AND2x2_ASAP7_75t_L g420 ( .A(n_241), .B(n_280), .Y(n_420) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_248), .B(n_249), .Y(n_241) );
AND2x2_ASAP7_75t_L g266 ( .A(n_251), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g281 ( .A(n_251), .Y(n_281) );
INVx1_ASAP7_75t_L g291 ( .A(n_251), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_257), .B(n_259), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_257), .A2(n_493), .B(n_494), .Y(n_492) );
INVx1_ASAP7_75t_L g510 ( .A(n_257), .Y(n_510) );
OAI22xp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_268), .B1(n_272), .B2(n_276), .Y(n_262) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_263), .A2(n_381), .B1(n_418), .B2(n_419), .Y(n_417) );
INVx1_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_L g332 ( .A(n_265), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_266), .B(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g327 ( .A(n_267), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_267), .B(n_280), .Y(n_354) );
INVx1_ASAP7_75t_L g370 ( .A(n_267), .Y(n_370) );
AND2x2_ASAP7_75t_L g311 ( .A(n_269), .B(n_312), .Y(n_311) );
INVx3_ASAP7_75t_SL g350 ( .A(n_269), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_269), .B(n_275), .Y(n_427) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx1_ASAP7_75t_L g436 ( .A(n_272), .Y(n_436) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_273), .B(n_369), .Y(n_411) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx3_ASAP7_75t_SL g316 ( .A(n_275), .Y(n_316) );
NAND2x1_ASAP7_75t_SL g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x2_ASAP7_75t_L g337 ( .A(n_277), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g344 ( .A(n_277), .B(n_281), .Y(n_344) );
AND2x2_ASAP7_75t_L g349 ( .A(n_277), .B(n_290), .Y(n_349) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_277), .Y(n_398) );
OAI311xp33_ASAP7_75t_L g421 ( .A1(n_278), .A2(n_422), .A3(n_424), .B1(n_425), .C1(n_435), .Y(n_421) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g434 ( .A(n_279), .B(n_307), .Y(n_434) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
AND2x2_ASAP7_75t_L g290 ( .A(n_280), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g338 ( .A(n_280), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g393 ( .A(n_280), .Y(n_393) );
INVx1_ASAP7_75t_L g286 ( .A(n_281), .Y(n_286) );
INVx1_ASAP7_75t_L g306 ( .A(n_281), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_281), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g339 ( .A(n_281), .Y(n_339) );
AOI221xp5_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_285), .B1(n_293), .B2(n_298), .C(n_303), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_288), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx4_ASAP7_75t_L g307 ( .A(n_287), .Y(n_307) );
AND2x2_ASAP7_75t_L g401 ( .A(n_287), .B(n_320), .Y(n_401) );
AND2x2_ASAP7_75t_L g408 ( .A(n_287), .B(n_290), .Y(n_408) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_290), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g319 ( .A(n_292), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_295), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g444 ( .A(n_297), .B(n_388), .Y(n_444) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g429 ( .A(n_301), .B(n_357), .Y(n_429) );
OAI211xp5_ASAP7_75t_L g394 ( .A1(n_302), .A2(n_395), .B(n_396), .C(n_409), .Y(n_394) );
AOI21xp33_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_308), .B(n_310), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NOR2xp67_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g373 ( .A(n_307), .Y(n_373) );
OAI221xp5_ASAP7_75t_L g402 ( .A1(n_308), .A2(n_403), .B1(n_404), .B2(n_405), .C(n_406), .Y(n_402) );
AND2x2_ASAP7_75t_L g379 ( .A(n_309), .B(n_320), .Y(n_379) );
AND2x2_ASAP7_75t_L g432 ( .A(n_309), .B(n_327), .Y(n_432) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_312), .B(n_350), .Y(n_374) );
O2A1O1Ixp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_317), .B(n_319), .C(n_321), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AND2x2_ASAP7_75t_L g360 ( .A(n_315), .B(n_318), .Y(n_360) );
OR2x2_ASAP7_75t_L g403 ( .A(n_315), .B(n_357), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_316), .B(n_382), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_316), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_SL g347 ( .A(n_317), .Y(n_347) );
INVx1_ASAP7_75t_L g413 ( .A(n_320), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_325), .B1(n_328), .B2(n_329), .Y(n_321) );
INVx1_ASAP7_75t_L g336 ( .A(n_322), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_323), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g399 ( .A(n_324), .B(n_400), .Y(n_399) );
INVxp67_ASAP7_75t_L g385 ( .A(n_326), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_327), .B(n_413), .Y(n_412) );
OAI22xp33_ASAP7_75t_L g386 ( .A1(n_328), .A2(n_387), .B1(n_389), .B2(n_391), .Y(n_386) );
INVx1_ASAP7_75t_L g395 ( .A(n_331), .Y(n_395) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
AND2x2_ASAP7_75t_L g437 ( .A(n_332), .B(n_432), .Y(n_437) );
AOI222xp33_ASAP7_75t_L g366 ( .A1(n_333), .A2(n_367), .B1(n_370), .B2(n_371), .C1(n_374), .C2(n_375), .Y(n_366) );
NAND4xp25_ASAP7_75t_SL g334 ( .A(n_335), .B(n_355), .C(n_366), .D(n_378), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B1(n_340), .B2(n_345), .C(n_346), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_338), .B(n_373), .Y(n_372) );
INVxp67_ASAP7_75t_L g364 ( .A(n_339), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_340), .A2(n_410), .B1(n_412), .B2(n_414), .C(n_417), .Y(n_409) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g352 ( .A(n_344), .B(n_353), .Y(n_352) );
OAI21xp33_ASAP7_75t_L g406 ( .A1(n_345), .A2(n_407), .B(n_408), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B1(n_350), .B2(n_351), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_358), .B(n_361), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g397 ( .A(n_368), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_369), .B(n_388), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_369), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_373), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g405 ( .A(n_377), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_383), .B2(n_385), .C(n_386), .Y(n_378) );
INVxp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI222xp33_ASAP7_75t_L g425 ( .A1(n_388), .A2(n_426), .B1(n_427), .B2(n_428), .C1(n_430), .C2(n_433), .Y(n_425) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_392), .B(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g424 ( .A(n_398), .Y(n_424) );
INVxp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVxp33_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_437), .B1(n_438), .B2(n_439), .C(n_442), .Y(n_435) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_449), .A2(n_457), .B1(n_745), .B2(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g746 ( .A(n_460), .Y(n_746) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND3x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_654), .C(n_702), .Y(n_461) );
NOR4xp25_ASAP7_75t_L g462 ( .A(n_463), .B(n_582), .C(n_627), .D(n_641), .Y(n_462) );
OAI311xp33_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_502), .A3(n_526), .B1(n_535), .C1(n_550), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_473), .Y(n_464) );
OAI21xp33_ASAP7_75t_L g535 ( .A1(n_465), .A2(n_536), .B(n_538), .Y(n_535) );
AND2x2_ASAP7_75t_L g643 ( .A(n_465), .B(n_570), .Y(n_643) );
AND2x2_ASAP7_75t_L g700 ( .A(n_465), .B(n_586), .Y(n_700) );
BUFx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g593 ( .A(n_466), .B(n_496), .Y(n_593) );
AND2x2_ASAP7_75t_L g650 ( .A(n_466), .B(n_598), .Y(n_650) );
INVx1_ASAP7_75t_L g691 ( .A(n_466), .Y(n_691) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_467), .Y(n_559) );
AND2x2_ASAP7_75t_L g600 ( .A(n_467), .B(n_496), .Y(n_600) );
AND2x2_ASAP7_75t_L g604 ( .A(n_467), .B(n_497), .Y(n_604) );
INVx1_ASAP7_75t_L g616 ( .A(n_467), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_472), .A2(n_543), .B(n_546), .Y(n_542) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_484), .Y(n_473) );
AND2x2_ASAP7_75t_L g537 ( .A(n_474), .B(n_496), .Y(n_537) );
INVx2_ASAP7_75t_L g571 ( .A(n_474), .Y(n_571) );
AND2x2_ASAP7_75t_L g586 ( .A(n_474), .B(n_497), .Y(n_586) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_474), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_474), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g606 ( .A(n_474), .B(n_569), .Y(n_606) );
INVx1_ASAP7_75t_L g618 ( .A(n_474), .Y(n_618) );
INVx1_ASAP7_75t_L g659 ( .A(n_474), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_474), .B(n_559), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B(n_479), .Y(n_476) );
NOR2xp67_ASAP7_75t_L g484 ( .A(n_485), .B(n_496), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g536 ( .A(n_486), .B(n_537), .Y(n_536) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_486), .Y(n_564) );
AND2x2_ASAP7_75t_SL g617 ( .A(n_486), .B(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g621 ( .A(n_486), .B(n_496), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_486), .B(n_616), .Y(n_679) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g569 ( .A(n_487), .Y(n_569) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_487), .Y(n_585) );
OR2x2_ASAP7_75t_L g658 ( .A(n_487), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g565 ( .A(n_497), .Y(n_565) );
AND2x2_ASAP7_75t_L g570 ( .A(n_497), .B(n_571), .Y(n_570) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_500), .A2(n_512), .B(n_514), .C(n_515), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_500), .A2(n_523), .B(n_524), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_502), .B(n_553), .Y(n_716) );
INVx1_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g686 ( .A(n_503), .B(n_528), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_517), .Y(n_503) );
AND2x2_ASAP7_75t_L g562 ( .A(n_504), .B(n_553), .Y(n_562) );
INVx2_ASAP7_75t_L g574 ( .A(n_504), .Y(n_574) );
AND2x2_ASAP7_75t_L g608 ( .A(n_504), .B(n_556), .Y(n_608) );
AND2x2_ASAP7_75t_L g675 ( .A(n_504), .B(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_505), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g555 ( .A(n_505), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g595 ( .A(n_505), .B(n_517), .Y(n_595) );
AND2x2_ASAP7_75t_L g612 ( .A(n_505), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g538 ( .A(n_517), .B(n_539), .Y(n_538) );
INVx3_ASAP7_75t_L g556 ( .A(n_517), .Y(n_556) );
AND2x2_ASAP7_75t_L g561 ( .A(n_517), .B(n_541), .Y(n_561) );
AND2x2_ASAP7_75t_L g634 ( .A(n_517), .B(n_613), .Y(n_634) );
AND2x2_ASAP7_75t_L g699 ( .A(n_517), .B(n_689), .Y(n_699) );
OAI311xp33_ASAP7_75t_L g582 ( .A1(n_526), .A2(n_583), .A3(n_587), .B1(n_589), .C1(n_609), .Y(n_582) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g594 ( .A(n_527), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g653 ( .A(n_527), .B(n_561), .Y(n_653) );
AND2x2_ASAP7_75t_L g727 ( .A(n_527), .B(n_608), .Y(n_727) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_528), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g662 ( .A(n_528), .Y(n_662) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx3_ASAP7_75t_L g553 ( .A(n_529), .Y(n_553) );
NOR2x1_ASAP7_75t_L g625 ( .A(n_529), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g682 ( .A(n_529), .B(n_556), .Y(n_682) );
AND2x4_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g579 ( .A(n_530), .Y(n_579) );
AND2x2_ASAP7_75t_L g557 ( .A(n_537), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g610 ( .A(n_537), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g690 ( .A(n_537), .B(n_691), .Y(n_690) );
AOI221xp5_ASAP7_75t_L g589 ( .A1(n_538), .A2(n_570), .B1(n_590), .B2(n_594), .C(n_596), .Y(n_589) );
INVx1_ASAP7_75t_L g714 ( .A(n_539), .Y(n_714) );
OR2x2_ASAP7_75t_L g680 ( .A(n_540), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g575 ( .A(n_541), .B(n_556), .Y(n_575) );
OR2x2_ASAP7_75t_L g577 ( .A(n_541), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g602 ( .A(n_541), .Y(n_602) );
INVx2_ASAP7_75t_L g613 ( .A(n_541), .Y(n_613) );
AND2x2_ASAP7_75t_L g640 ( .A(n_541), .B(n_578), .Y(n_640) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_541), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_557), .B1(n_560), .B2(n_563), .C(n_566), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
AND2x2_ASAP7_75t_L g651 ( .A(n_553), .B(n_561), .Y(n_651) );
AND2x2_ASAP7_75t_L g701 ( .A(n_553), .B(n_555), .Y(n_701) );
INVx2_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g588 ( .A(n_555), .B(n_559), .Y(n_588) );
AND2x2_ASAP7_75t_L g667 ( .A(n_555), .B(n_640), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_556), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g626 ( .A(n_556), .Y(n_626) );
OAI21xp33_ASAP7_75t_L g636 ( .A1(n_557), .A2(n_637), .B(n_639), .Y(n_636) );
OR2x2_ASAP7_75t_L g580 ( .A(n_558), .B(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g646 ( .A(n_558), .B(n_606), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_558), .B(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g623 ( .A(n_559), .B(n_592), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_559), .B(n_706), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_560), .B(n_586), .Y(n_696) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
AND2x2_ASAP7_75t_L g619 ( .A(n_561), .B(n_574), .Y(n_619) );
INVx1_ASAP7_75t_L g635 ( .A(n_562), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_572), .B1(n_576), .B2(n_580), .Y(n_566) );
INVx2_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx2_ASAP7_75t_L g598 ( .A(n_569), .Y(n_598) );
INVx1_ASAP7_75t_L g611 ( .A(n_569), .Y(n_611) );
INVx1_ASAP7_75t_L g581 ( .A(n_570), .Y(n_581) );
AND2x2_ASAP7_75t_L g652 ( .A(n_570), .B(n_598), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_570), .B(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
OR2x2_ASAP7_75t_L g576 ( .A(n_573), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_573), .B(n_689), .Y(n_688) );
NOR2xp67_ASAP7_75t_L g720 ( .A(n_573), .B(n_721), .Y(n_720) );
INVx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g723 ( .A(n_575), .B(n_675), .Y(n_723) );
INVx1_ASAP7_75t_SL g689 ( .A(n_577), .Y(n_689) );
AND2x2_ASAP7_75t_L g629 ( .A(n_578), .B(n_613), .Y(n_629) );
INVx1_ASAP7_75t_L g676 ( .A(n_578), .Y(n_676) );
OAI222xp33_ASAP7_75t_L g717 ( .A1(n_583), .A2(n_673), .B1(n_718), .B2(n_719), .C1(n_722), .C2(n_724), .Y(n_717) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx1_ASAP7_75t_L g638 ( .A(n_585), .Y(n_638) );
AND2x2_ASAP7_75t_L g649 ( .A(n_586), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g718 ( .A(n_586), .B(n_691), .Y(n_718) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_588), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g693 ( .A(n_590), .Y(n_693) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_SL g631 ( .A(n_593), .Y(n_631) );
AND2x2_ASAP7_75t_L g710 ( .A(n_593), .B(n_671), .Y(n_710) );
AND2x2_ASAP7_75t_L g733 ( .A(n_593), .B(n_617), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_595), .B(n_629), .Y(n_628) );
OAI32xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_599), .A3(n_601), .B1(n_603), .B2(n_607), .Y(n_596) );
BUFx2_ASAP7_75t_L g671 ( .A(n_598), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_599), .B(n_617), .Y(n_698) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g637 ( .A(n_600), .B(n_638), .Y(n_637) );
AND2x4_ASAP7_75t_L g705 ( .A(n_600), .B(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g694 ( .A(n_601), .B(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
AND2x2_ASAP7_75t_L g665 ( .A(n_604), .B(n_638), .Y(n_665) );
INVx2_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
OAI221xp5_ASAP7_75t_SL g627 ( .A1(n_606), .A2(n_628), .B1(n_630), .B2(n_632), .C(n_636), .Y(n_627) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g639 ( .A(n_608), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g645 ( .A(n_608), .B(n_629), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_612), .B1(n_614), .B2(n_619), .C(n_620), .Y(n_609) );
INVx1_ASAP7_75t_L g728 ( .A(n_610), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_611), .B(n_705), .Y(n_704) );
NAND2x1p5_ASAP7_75t_L g624 ( .A(n_612), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_617), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g683 ( .A(n_617), .Y(n_683) );
BUFx3_ASAP7_75t_L g706 ( .A(n_618), .Y(n_706) );
INVx1_ASAP7_75t_SL g647 ( .A(n_619), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_619), .B(n_661), .Y(n_660) );
AOI21xp33_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_622), .B(n_624), .Y(n_620) );
OAI221xp5_ASAP7_75t_L g725 ( .A1(n_621), .A2(n_722), .B1(n_726), .B2(n_728), .C(n_729), .Y(n_725) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g668 ( .A(n_626), .B(n_629), .Y(n_668) );
INVx1_ASAP7_75t_L g732 ( .A(n_626), .Y(n_732) );
INVx2_ASAP7_75t_L g721 ( .A(n_629), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_629), .B(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g674 ( .A(n_634), .B(n_675), .Y(n_674) );
OAI221xp5_ASAP7_75t_SL g641 ( .A1(n_642), .A2(n_644), .B1(n_646), .B2(n_647), .C(n_648), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_651), .B1(n_652), .B2(n_653), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_650), .A2(n_712), .B1(n_713), .B2(n_715), .Y(n_711) );
OAI21xp5_ASAP7_75t_L g729 ( .A1(n_653), .A2(n_730), .B(n_733), .Y(n_729) );
NOR4xp25_ASAP7_75t_SL g654 ( .A(n_655), .B(n_663), .C(n_672), .D(n_692), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_660), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .B1(n_669), .B2(n_670), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g708 ( .A(n_668), .Y(n_708) );
OAI221xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_677), .B1(n_680), .B2(n_683), .C(n_684), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g695 ( .A(n_675), .Y(n_695) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OAI21xp5_ASAP7_75t_SL g684 ( .A1(n_685), .A2(n_687), .B(n_690), .Y(n_684) );
INVx1_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OAI211xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_694), .B(n_696), .C(n_697), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B1(n_700), .B2(n_701), .Y(n_697) );
CKINVDCx14_ASAP7_75t_R g707 ( .A(n_701), .Y(n_707) );
NOR3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_717), .C(n_725), .Y(n_702) );
OAI221xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_707), .B1(n_708), .B2(n_709), .C(n_711), .Y(n_703) );
INVxp67_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
CKINVDCx16_ASAP7_75t_R g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g745 ( .A(n_735), .Y(n_745) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
CKINVDCx16_ASAP7_75t_R g747 ( .A(n_738), .Y(n_747) );
INVx1_ASAP7_75t_L g742 ( .A(n_739), .Y(n_742) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx3_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
endmodule