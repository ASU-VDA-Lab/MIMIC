module fake_jpeg_20323_n_105 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

AND2x4_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_20),
.B1(n_18),
.B2(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_31),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_20),
.B1(n_18),
.B2(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_32),
.B(n_36),
.Y(n_48)
);

NOR2x1_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_35),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_17),
.B(n_16),
.C(n_13),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_41),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_17),
.B(n_16),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_28),
.B(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_12),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_9),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_11),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_22),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_22),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_54),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_22),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_57),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_27),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_38),
.B1(n_37),
.B2(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_65),
.Y(n_73)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_68),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_47),
.B1(n_48),
.B2(n_4),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_50),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_56),
.C(n_57),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_77),
.C(n_81),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_76),
.B(n_79),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_56),
.C(n_53),
.Y(n_77)
);

AO21x1_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_51),
.B(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_49),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_60),
.C(n_55),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_72),
.B1(n_69),
.B2(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_70),
.B1(n_64),
.B2(n_72),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_78),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_66),
.C(n_59),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_63),
.C(n_59),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_91),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_59),
.B(n_80),
.Y(n_92)
);

OA21x2_ASAP7_75t_SL g96 ( 
.A1(n_92),
.A2(n_93),
.B(n_4),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_48),
.C(n_2),
.Y(n_93)
);

AOI322xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_88),
.A3(n_82),
.B1(n_85),
.B2(n_87),
.C1(n_83),
.C2(n_1),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_95),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_2),
.C(n_4),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_97),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_99),
.A2(n_100),
.B(n_101),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_97),
.B(n_5),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_5),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_5),
.C(n_6),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_98),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_102),
.Y(n_105)
);


endmodule