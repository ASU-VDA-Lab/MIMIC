module fake_jpeg_14936_n_68 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_68);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_68;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

BUFx5_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_5),
.B(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_3),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_22),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_16),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_20),
.A2(n_24),
.B1(n_16),
.B2(n_5),
.Y(n_33)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_15),
.A2(n_10),
.B(n_14),
.C(n_13),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_14),
.B(n_10),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_16),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

NAND2xp33_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_11),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_13),
.B(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_8),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_4),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_5),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_11),
.C(n_17),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_30),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_31),
.B(n_32),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_37),
.B1(n_18),
.B2(n_19),
.Y(n_43)
);

NOR3xp33_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_30),
.C(n_39),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_39),
.B(n_17),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_20),
.A2(n_17),
.B1(n_8),
.B2(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_9),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_9),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_45),
.B(n_46),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_48),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_33),
.B1(n_37),
.B2(n_29),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_26),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_9),
.B1(n_18),
.B2(n_40),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_34),
.B(n_45),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_56),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_49),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_55),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

XOR2x1_ASAP7_75t_SL g57 ( 
.A(n_55),
.B(n_44),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_58),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_60),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_47),
.C(n_57),
.Y(n_64)
);

NAND4xp25_ASAP7_75t_SL g66 ( 
.A(n_64),
.B(n_48),
.C(n_61),
.D(n_59),
.Y(n_66)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

OAI221xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_66),
.B1(n_63),
.B2(n_50),
.C(n_35),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_64),
.C(n_41),
.Y(n_68)
);


endmodule