module fake_jpeg_3242_n_112 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_9),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_45),
.Y(n_47)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_33),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_42),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_29),
.B1(n_35),
.B2(n_38),
.Y(n_52)
);

AO22x1_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_55),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_34),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_59),
.Y(n_71)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_30),
.B1(n_32),
.B2(n_36),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_60),
.A2(n_42),
.B1(n_38),
.B2(n_31),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_32),
.C(n_30),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_65),
.B(n_17),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_54),
.B1(n_31),
.B2(n_3),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_63),
.A2(n_55),
.B1(n_52),
.B2(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_68),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_70),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_61),
.B1(n_58),
.B2(n_56),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_70),
.B1(n_66),
.B2(n_71),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_12),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_79),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_74),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_75),
.B(n_4),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_84),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_16),
.C(n_27),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_88),
.C(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_90),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_28),
.B(n_24),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_19),
.B(n_21),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_23),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_96),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_100),
.B(n_102),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_101),
.B(n_98),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_97),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_94),
.B1(n_91),
.B2(n_103),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_93),
.C(n_100),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_92),
.Y(n_108)
);

MAJx2_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_90),
.C(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_99),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_20),
.C(n_22),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_8),
.C(n_9),
.Y(n_112)
);


endmodule