module real_jpeg_9084_n_12 (n_5, n_4, n_8, n_0, n_278, n_1, n_11, n_2, n_6, n_277, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_278;
input n_1;
input n_11;
input n_2;
input n_6;
input n_277;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_262;
wire n_19;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_205;
wire n_110;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_130;
wire n_144;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_167;
wire n_244;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_1),
.A2(n_29),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_1),
.A2(n_29),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_1),
.A2(n_11),
.B1(n_29),
.B2(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_2),
.A2(n_87),
.B1(n_88),
.B2(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_2),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_2),
.A2(n_10),
.B(n_87),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_3),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_174),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_3),
.A2(n_87),
.B1(n_88),
.B2(n_174),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_6),
.A2(n_40),
.B(n_45),
.C(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_6),
.B(n_40),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_6),
.A2(n_10),
.B(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_SL g74 ( 
.A(n_7),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_9),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_9),
.A2(n_40),
.B1(n_41),
.B2(n_156),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_9),
.A2(n_87),
.B1(n_88),
.B2(n_156),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_9),
.A2(n_11),
.B1(n_134),
.B2(n_156),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_10),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_10),
.B(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_10),
.A2(n_35),
.B1(n_87),
.B2(n_88),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_10),
.A2(n_74),
.B(n_88),
.C(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_10),
.B(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_10),
.A2(n_11),
.B1(n_35),
.B2(n_134),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_11),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_11),
.A2(n_114),
.B(n_115),
.C(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_11),
.B(n_115),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_11),
.A2(n_35),
.B(n_115),
.C(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_263),
.Y(n_12)
);

OAI321xp33_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_231),
.A3(n_256),
.B1(n_261),
.B2(n_262),
.C(n_277),
.Y(n_13)
);

AOI321xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_185),
.A3(n_205),
.B1(n_225),
.B2(n_230),
.C(n_278),
.Y(n_14)
);

NOR3xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_148),
.C(n_182),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_121),
.B(n_147),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_102),
.B(n_120),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_80),
.B(n_101),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_65),
.B(n_79),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_55),
.B(n_64),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.Y(n_21)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_22),
.B(n_36),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_22),
.A2(n_57),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_22),
.B(n_106),
.C(n_112),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_30),
.B(n_31),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_24),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_25),
.B(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_30),
.B(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_30),
.A2(n_99),
.B1(n_155),
.B2(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_31),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_32),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_35),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_33),
.A2(n_154),
.B(n_157),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_34),
.B(n_98),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_41),
.B(n_46),
.C(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_35),
.B(n_45),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_35),
.A2(n_40),
.B(n_75),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_37),
.B(n_52),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_37),
.A2(n_54),
.B1(n_85),
.B2(n_93),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_37),
.B(n_85),
.C(n_100),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_37),
.A2(n_54),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_44),
.B(n_47),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_39),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_40),
.A2(n_41),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_45),
.B(n_49),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_45),
.A2(n_201),
.B(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_45),
.A2(n_49),
.B1(n_201),
.B2(n_212),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_47),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_48),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_54),
.B(n_153),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_60),
.B(n_63),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_61),
.B(n_62),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_68),
.B1(n_69),
.B2(n_78),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_70),
.C(n_77),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_62),
.A2(n_78),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_62),
.B(n_141),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_67),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_86),
.B(n_89),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_86),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_72),
.B(n_107),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_72),
.A2(n_107),
.B1(n_238),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_74),
.B(n_88),
.C(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_73),
.A2(n_237),
.B(n_239),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_74),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_88),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_76),
.A2(n_77),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_76),
.A2(n_77),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_76),
.B(n_171),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_105),
.C(n_119),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_82),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_94),
.B2(n_100),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_85),
.A2(n_93),
.B1(n_127),
.B2(n_130),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_85),
.B(n_127),
.C(n_132),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_85),
.A2(n_93),
.B1(n_161),
.B2(n_162),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_85),
.B(n_161),
.C(n_195),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_87),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_89),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_90),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_94),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_97),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_98),
.B(n_173),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_104),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_117),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_116),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_106),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_106),
.A2(n_116),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_106),
.B(n_161),
.C(n_164),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_133),
.B(n_135),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_114),
.A2(n_136),
.B1(n_137),
.B2(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_114),
.B(n_137),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_114),
.A2(n_270),
.B(n_271),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_116),
.A2(n_211),
.B(n_213),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_116),
.B(n_211),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_118),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_122),
.B(n_123),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_139),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_124),
.B(n_140),
.C(n_146),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_131),
.B2(n_132),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_127),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_129),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_131),
.A2(n_132),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_131),
.A2(n_132),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_131),
.A2(n_132),
.B1(n_248),
.B2(n_254),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_131),
.B(n_240),
.C(n_243),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_131),
.B(n_254),
.C(n_255),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_132),
.B(n_176),
.C(n_178),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_133),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_135),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_136),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_140),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_144),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g226 ( 
.A1(n_149),
.A2(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_165),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_150),
.B(n_165),
.Y(n_228)
);

FAx1_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_158),
.CI(n_159),
.CON(n_150),
.SN(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_161),
.A2(n_162),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_161),
.B(n_241),
.C(n_252),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_181),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_175),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_175),
.C(n_181),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_180),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_184),
.Y(n_227)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_186),
.A2(n_226),
.B(n_229),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_187),
.B(n_188),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_204),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_196),
.B2(n_197),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_197),
.C(n_204),
.Y(n_206)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_192),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_203),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_199),
.B1(n_217),
.B2(n_220),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_200),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_199),
.A2(n_215),
.B(n_217),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_200),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_207),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_223),
.B2(n_224),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_214),
.B1(n_221),
.B2(n_222),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_210),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_222),
.C(n_224),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_212),
.B(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_233),
.C(n_244),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_213),
.B(n_233),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_214),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_217),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_223),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_246),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_246),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_240),
.B1(n_241),
.B2(n_243),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_236),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_240),
.A2(n_241),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_244),
.A2(n_245),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_255),
.Y(n_246)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_248),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_257),
.B(n_258),
.Y(n_261)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_259),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_274),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_273),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_273),
.Y(n_274)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_266),
.Y(n_275)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_269),
.CI(n_272),
.CON(n_266),
.SN(n_266)
);


endmodule