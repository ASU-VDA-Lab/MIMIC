module fake_jpeg_21838_n_349 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_50),
.A2(n_35),
.B1(n_17),
.B2(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_69),
.B1(n_28),
.B2(n_22),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_34),
.B1(n_17),
.B2(n_25),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_55),
.A2(n_49),
.B1(n_20),
.B2(n_21),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_34),
.B1(n_17),
.B2(n_25),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_64),
.B1(n_18),
.B2(n_49),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_31),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_63),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_31),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_18),
.B1(n_31),
.B2(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_41),
.A2(n_37),
.B1(n_28),
.B2(n_27),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx2_ASAP7_75t_SL g105 ( 
.A(n_70),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_42),
.B(n_33),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_71),
.B(n_26),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_33),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_74),
.B(n_99),
.Y(n_107)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_86),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_50),
.B1(n_46),
.B2(n_39),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_78),
.A2(n_106),
.B1(n_99),
.B2(n_81),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_81),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_80),
.A2(n_100),
.B1(n_72),
.B2(n_52),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_85),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_83),
.A2(n_95),
.B1(n_103),
.B2(n_29),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_62),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_46),
.B1(n_39),
.B2(n_47),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_88),
.A2(n_72),
.B1(n_61),
.B2(n_29),
.Y(n_132)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_27),
.B(n_26),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_69),
.Y(n_109)
);

BUFx8_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_56),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_93),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_45),
.Y(n_94)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_55),
.A2(n_49),
.B1(n_20),
.B2(n_30),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_45),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_66),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_63),
.Y(n_99)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_60),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_101),
.B(n_21),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_63),
.B(n_38),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_58),
.C(n_67),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_51),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_51),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_112),
.B(n_121),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_69),
.B(n_66),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_113),
.A2(n_24),
.B(n_36),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_SL g143 ( 
.A1(n_114),
.A2(n_131),
.B(n_105),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_69),
.B(n_47),
.C(n_51),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_134),
.B(n_132),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_69),
.B1(n_67),
.B2(n_61),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_123),
.A2(n_135),
.B1(n_89),
.B2(n_85),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_130),
.B1(n_132),
.B2(n_136),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_79),
.A2(n_58),
.B1(n_38),
.B2(n_72),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_75),
.A2(n_47),
.B1(n_36),
.B2(n_32),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_80),
.A2(n_30),
.B1(n_43),
.B2(n_40),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_111),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

AOI32xp33_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_104),
.A3(n_102),
.B1(n_80),
.B2(n_88),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_24),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_80),
.B1(n_104),
.B2(n_102),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

INVxp67_ASAP7_75t_SL g168 ( 
.A(n_140),
.Y(n_168)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_141),
.B(n_148),
.Y(n_193)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_144),
.B1(n_160),
.B2(n_110),
.Y(n_176)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_118),
.B1(n_117),
.B2(n_122),
.Y(n_184)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_116),
.A2(n_75),
.B1(n_74),
.B2(n_93),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_150),
.B1(n_157),
.B2(n_159),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_116),
.A2(n_92),
.B1(n_97),
.B2(n_96),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_135),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_152),
.B(n_154),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_113),
.A2(n_77),
.B(n_87),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_153),
.A2(n_156),
.B(n_165),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_91),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g155 ( 
.A1(n_109),
.A2(n_87),
.B(n_82),
.C(n_44),
.D(n_43),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_134),
.C(n_109),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_100),
.B1(n_87),
.B2(n_76),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_91),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_163),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_131),
.B1(n_123),
.B2(n_130),
.Y(n_159)
);

AO22x1_ASAP7_75t_SL g160 ( 
.A1(n_114),
.A2(n_100),
.B1(n_32),
.B2(n_36),
.Y(n_160)
);

XNOR2x1_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_40),
.Y(n_161)
);

XNOR2x1_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_0),
.Y(n_199)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_121),
.B(n_13),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_164),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_128),
.A2(n_44),
.B(n_43),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_126),
.A2(n_44),
.B1(n_84),
.B2(n_36),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_166),
.A2(n_118),
.B1(n_108),
.B2(n_125),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_167),
.A2(n_73),
.B(n_1),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_169),
.B(n_198),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_127),
.B(n_107),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_172),
.A2(n_199),
.B(n_160),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_137),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_191),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_176),
.A2(n_180),
.B1(n_184),
.B2(n_157),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_167),
.A2(n_107),
.B(n_120),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_190),
.B(n_163),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_120),
.B1(n_111),
.B2(n_124),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_179),
.A2(n_182),
.B1(n_187),
.B2(n_188),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_124),
.B1(n_125),
.B2(n_122),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_195),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_117),
.C(n_108),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_186),
.C(n_197),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_91),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_147),
.A2(n_119),
.B1(n_32),
.B2(n_24),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_147),
.A2(n_73),
.B1(n_1),
.B2(n_2),
.Y(n_188)
);

FAx1_ASAP7_75t_SL g191 ( 
.A(n_158),
.B(n_0),
.CI(n_2),
.CON(n_191),
.SN(n_191)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_140),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_142),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_16),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_141),
.B(n_0),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_200),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_16),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_15),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_148),
.B(n_0),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_162),
.Y(n_202)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_202),
.Y(n_249)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_203),
.B(n_206),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_228),
.B(n_200),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_170),
.Y(n_207)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_211),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_187),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_180),
.Y(n_210)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_210),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_213),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_174),
.A2(n_166),
.B1(n_138),
.B2(n_155),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_214),
.A2(n_225),
.B1(n_192),
.B2(n_7),
.Y(n_252)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_216),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_219),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_144),
.C(n_151),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_227),
.C(n_230),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_172),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_174),
.A2(n_146),
.B1(n_15),
.B2(n_14),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_223),
.A2(n_224),
.B1(n_229),
.B2(n_231),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_199),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_177),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_3),
.C(n_4),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_3),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_176),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_4),
.C(n_5),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_188),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_211),
.A2(n_190),
.B(n_178),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_235),
.A2(n_227),
.B(n_220),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_252),
.Y(n_261)
);

XNOR2x2_ASAP7_75t_SL g238 ( 
.A(n_209),
.B(n_181),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_238),
.B(n_218),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_214),
.B(n_169),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_246),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_191),
.B(n_197),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_247),
.B(n_248),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_195),
.C(n_175),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_212),
.C(n_226),
.Y(n_259)
);

OA21x2_ASAP7_75t_L g247 ( 
.A1(n_229),
.A2(n_191),
.B(n_175),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_205),
.A2(n_171),
.B(n_192),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_12),
.C(n_10),
.Y(n_253)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_206),
.A2(n_10),
.B1(n_12),
.B2(n_9),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_254),
.A2(n_224),
.B1(n_223),
.B2(n_225),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_226),
.B(n_232),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_232),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_218),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_258)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_258),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_260),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_221),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_236),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_269),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_265),
.B(n_266),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_257),
.C(n_239),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_267),
.B(n_270),
.Y(n_297)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_242),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_273),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_240),
.A2(n_204),
.B1(n_207),
.B2(n_230),
.Y(n_274)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_238),
.B(n_216),
.Y(n_275)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_276),
.A2(n_278),
.B(n_264),
.Y(n_288)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_233),
.Y(n_277)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_277),
.Y(n_287)
);

INVxp33_ASAP7_75t_L g279 ( 
.A(n_250),
.Y(n_279)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_233),
.Y(n_280)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_276),
.A2(n_251),
.B1(n_234),
.B2(n_235),
.Y(n_281)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_234),
.B1(n_256),
.B2(n_249),
.Y(n_282)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_269),
.A2(n_246),
.B1(n_243),
.B2(n_256),
.Y(n_286)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_288),
.A2(n_291),
.B(n_268),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_264),
.A2(n_252),
.B(n_247),
.Y(n_291)
);

INVx13_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_254),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_R g293 ( 
.A(n_271),
.B(n_244),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_293),
.A2(n_243),
.B(n_275),
.Y(n_310)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_247),
.Y(n_299)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_299),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_303),
.A2(n_307),
.B(n_310),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_263),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_304),
.B(n_305),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_241),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_266),
.C(n_259),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_311),
.C(n_272),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_288),
.A2(n_268),
.B(n_237),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_260),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_309),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_273),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_272),
.C(n_220),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_290),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_298),
.B(n_262),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_313),
.B(n_286),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_283),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_316),
.C(n_306),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_300),
.A2(n_285),
.B1(n_295),
.B2(n_290),
.Y(n_318)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_318),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_321),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_311),
.B(n_297),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_324),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_301),
.A2(n_291),
.B1(n_289),
.B2(n_296),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_307),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_299),
.A2(n_285),
.B(n_293),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_308),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_327),
.B(n_330),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_287),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_318),
.B(n_303),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_294),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_314),
.C(n_315),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_333),
.A2(n_294),
.B1(n_258),
.B2(n_8),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g334 ( 
.A(n_314),
.B(n_302),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_320),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_335),
.B(n_337),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_338),
.C(n_340),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_329),
.A2(n_325),
.B1(n_324),
.B2(n_310),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_328),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_332),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_342),
.B(n_327),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_336),
.B1(n_339),
.B2(n_344),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_346),
.A2(n_343),
.B(n_342),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_347),
.A2(n_326),
.B1(n_335),
.B2(n_8),
.Y(n_348)
);

XNOR2x2_ASAP7_75t_SL g349 ( 
.A(n_348),
.B(n_8),
.Y(n_349)
);


endmodule