module fake_jpeg_15370_n_126 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_126);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_60),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_0),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_58),
.A2(n_42),
.B1(n_45),
.B2(n_48),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_59),
.A2(n_42),
.B1(n_45),
.B2(n_51),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_40),
.B1(n_39),
.B2(n_44),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_54),
.B1(n_44),
.B2(n_46),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_54),
.B1(n_52),
.B2(n_43),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_70),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_72),
.B(n_3),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_41),
.B1(n_1),
.B2(n_2),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_73),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_79)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_19),
.B1(n_36),
.B2(n_34),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_6),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_22),
.C(n_33),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_85),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_84),
.B1(n_89),
.B2(n_77),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_12),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_63),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_69),
.B1(n_12),
.B2(n_68),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_38),
.Y(n_91)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_94),
.B(n_89),
.Y(n_104)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_103),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_106),
.B(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_105),
.B(n_107),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_94),
.B(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_92),
.B(n_82),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_106),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_112),
.C(n_109),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_114),
.B(n_97),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_96),
.B1(n_76),
.B2(n_81),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_108),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_116),
.B(n_117),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_100),
.B1(n_113),
.B2(n_99),
.Y(n_119)
);

OAI221xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_98),
.B1(n_88),
.B2(n_95),
.C(n_68),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_13),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_14),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_16),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_17),
.C(n_18),
.Y(n_124)
);

AOI321xp33_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_20),
.A3(n_23),
.B1(n_24),
.B2(n_25),
.C(n_26),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_29),
.Y(n_126)
);


endmodule