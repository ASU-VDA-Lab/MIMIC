module fake_jpeg_22123_n_165 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_9),
.B(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_31),
.Y(n_46)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_32),
.A2(n_26),
.B1(n_25),
.B2(n_17),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_33),
.B(n_34),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_38),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_2),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_2),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_43),
.B(n_12),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_23),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_2),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_27),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_21),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_58),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_54),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_33),
.B(n_22),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_70),
.C(n_10),
.Y(n_89)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_60),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_19),
.B(n_23),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_15),
.B(n_29),
.C(n_16),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_63),
.B1(n_37),
.B2(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_66),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_26),
.B1(n_28),
.B2(n_22),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_36),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_65),
.B(n_3),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_36),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_29),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_69),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_18),
.C(n_15),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_31),
.B(n_18),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_11),
.Y(n_90)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_79),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_SL g111 ( 
.A(n_75),
.B(n_85),
.C(n_89),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_78),
.Y(n_104)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_16),
.B1(n_37),
.B2(n_3),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_3),
.B(n_5),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_93),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_52),
.A2(n_65),
.B1(n_64),
.B2(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_76),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_100),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_72),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_50),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_90),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_113),
.B(n_118),
.Y(n_132)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_81),
.B(n_86),
.Y(n_114)
);

AO21x1_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_111),
.B(n_103),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_88),
.C(n_72),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_123),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_82),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_120),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_74),
.C(n_89),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_73),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_124),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_79),
.C(n_73),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_73),
.C(n_80),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_102),
.B1(n_111),
.B2(n_101),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_128),
.A2(n_134),
.B1(n_120),
.B2(n_112),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_130),
.B(n_59),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_106),
.B(n_102),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_75),
.B1(n_112),
.B2(n_93),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_136),
.B(n_115),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_121),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_142),
.B(n_143),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_137),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_133),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_141),
.A2(n_144),
.B1(n_133),
.B2(n_110),
.Y(n_152)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_SL g143 ( 
.A1(n_129),
.A2(n_93),
.B(n_53),
.C(n_126),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_51),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_146),
.C(n_147),
.Y(n_149)
);

A2O1A1O1Ixp25_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_93),
.B(n_59),
.C(n_118),
.D(n_110),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_135),
.C(n_132),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_152),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_131),
.B(n_134),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_151),
.A2(n_143),
.B1(n_139),
.B2(n_96),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_157),
.B(n_149),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_97),
.B1(n_52),
.B2(n_46),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_158),
.C(n_46),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_161),
.B(n_156),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_160),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_157),
.A2(n_153),
.B(n_49),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_156),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_163),
.C(n_53),
.Y(n_165)
);


endmodule