module fake_aes_6640_n_567 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_567);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_567;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_409;
wire n_363;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g74 ( .A(n_15), .Y(n_74) );
CKINVDCx16_ASAP7_75t_R g75 ( .A(n_48), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_18), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_54), .Y(n_77) );
INVxp33_ASAP7_75t_SL g78 ( .A(n_56), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_26), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_45), .Y(n_80) );
BUFx3_ASAP7_75t_L g81 ( .A(n_30), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_29), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_59), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_19), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_6), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_32), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_38), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_34), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_16), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_16), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_44), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_3), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_11), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_43), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_55), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_28), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_1), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_20), .Y(n_98) );
BUFx2_ASAP7_75t_L g99 ( .A(n_66), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_21), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_36), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_60), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_72), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_8), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_33), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_19), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_63), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_27), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_62), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_35), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_67), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_8), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_46), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_73), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_40), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_47), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_53), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_22), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_41), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_58), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_13), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_69), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_99), .B(n_0), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_122), .Y(n_124) );
INVxp67_ASAP7_75t_L g125 ( .A(n_99), .Y(n_125) );
OAI21x1_ASAP7_75t_L g126 ( .A1(n_122), .A2(n_23), .B(n_70), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_122), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_77), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_74), .B(n_0), .Y(n_129) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_89), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_75), .B(n_1), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_110), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_77), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_89), .B(n_2), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_79), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_110), .Y(n_136) );
NOR2xp67_ASAP7_75t_L g137 ( .A(n_104), .B(n_2), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_74), .B(n_3), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_76), .B(n_4), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_86), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_79), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_78), .Y(n_142) );
OAI21x1_ASAP7_75t_L g143 ( .A1(n_80), .A2(n_25), .B(n_68), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_96), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_80), .Y(n_145) );
CKINVDCx16_ASAP7_75t_R g146 ( .A(n_81), .Y(n_146) );
OAI21x1_ASAP7_75t_L g147 ( .A1(n_82), .A2(n_24), .B(n_65), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_76), .B(n_84), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_100), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_82), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_84), .B(n_4), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_101), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_118), .Y(n_153) );
INVxp67_ASAP7_75t_L g154 ( .A(n_90), .Y(n_154) );
CKINVDCx16_ASAP7_75t_R g155 ( .A(n_81), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_90), .B(n_5), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_83), .B(n_5), .Y(n_157) );
INVxp33_ASAP7_75t_SL g158 ( .A(n_92), .Y(n_158) );
BUFx10_ASAP7_75t_L g159 ( .A(n_83), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_87), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_87), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_88), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_88), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_94), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_125), .B(n_107), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_125), .B(n_121), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_139), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_139), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_153), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_139), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_124), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_127), .B(n_121), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_146), .B(n_108), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_159), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_139), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_127), .B(n_112), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_139), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_124), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_146), .B(n_105), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_124), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_127), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_127), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_127), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_153), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_130), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_130), .Y(n_186) );
INVxp67_ASAP7_75t_L g187 ( .A(n_131), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_134), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_159), .B(n_120), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_124), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_124), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_134), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_134), .B(n_112), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_134), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_124), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_134), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_124), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_140), .Y(n_198) );
OAI22xp33_ASAP7_75t_L g199 ( .A1(n_123), .A2(n_92), .B1(n_93), .B2(n_97), .Y(n_199) );
OR2x2_ASAP7_75t_SL g200 ( .A(n_155), .B(n_97), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_138), .Y(n_201) );
AOI22x1_ASAP7_75t_L g202 ( .A1(n_163), .A2(n_120), .B1(n_119), .B2(n_117), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_138), .Y(n_203) );
AND2x6_ASAP7_75t_L g204 ( .A(n_138), .B(n_119), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_126), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_155), .B(n_102), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_154), .B(n_117), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_154), .B(n_93), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_156), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_156), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_156), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_163), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_128), .B(n_98), .Y(n_213) );
NAND2x1p5_ASAP7_75t_L g214 ( .A(n_131), .B(n_98), .Y(n_214) );
AOI22xp33_ASAP7_75t_SL g215 ( .A1(n_131), .A2(n_106), .B1(n_85), .B2(n_114), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_164), .B(n_116), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_132), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_163), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_163), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_159), .B(n_116), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_158), .B(n_109), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_128), .B(n_115), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_133), .B(n_109), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_133), .B(n_114), .Y(n_224) );
NAND3xp33_ASAP7_75t_L g225 ( .A(n_123), .B(n_113), .C(n_111), .Y(n_225) );
OR2x2_ASAP7_75t_L g226 ( .A(n_148), .B(n_115), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_158), .B(n_113), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_163), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_145), .Y(n_229) );
BUFx2_ASAP7_75t_L g230 ( .A(n_204), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_218), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_226), .B(n_159), .Y(n_232) );
NOR2x1p5_ASAP7_75t_SL g233 ( .A(n_212), .B(n_150), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_218), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_218), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_219), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_219), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_199), .B(n_144), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_219), .Y(n_239) );
INVx2_ASAP7_75t_SL g240 ( .A(n_226), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_208), .B(n_159), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_208), .B(n_152), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_221), .B(n_149), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_181), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_201), .B(n_137), .Y(n_245) );
INVx4_ASAP7_75t_L g246 ( .A(n_204), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_180), .Y(n_247) );
INVx4_ASAP7_75t_L g248 ( .A(n_204), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_203), .B(n_209), .Y(n_249) );
BUFx3_ASAP7_75t_L g250 ( .A(n_204), .Y(n_250) );
NOR3xp33_ASAP7_75t_SL g251 ( .A(n_198), .B(n_140), .C(n_142), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_193), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_191), .Y(n_253) );
NOR3xp33_ASAP7_75t_SL g254 ( .A(n_198), .B(n_142), .C(n_157), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_193), .Y(n_255) );
NOR3xp33_ASAP7_75t_SL g256 ( .A(n_169), .B(n_157), .C(n_129), .Y(n_256) );
INVx3_ASAP7_75t_SL g257 ( .A(n_169), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_228), .A2(n_126), .B(n_143), .Y(n_258) );
INVx4_ASAP7_75t_L g259 ( .A(n_204), .Y(n_259) );
INVx4_ASAP7_75t_L g260 ( .A(n_204), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_182), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_205), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_221), .B(n_164), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_183), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_191), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_229), .Y(n_266) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_205), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_185), .B(n_148), .Y(n_268) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_187), .A2(n_137), .B1(n_162), .B2(n_141), .Y(n_269) );
INVx2_ASAP7_75t_SL g270 ( .A(n_172), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_210), .B(n_129), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_191), .Y(n_272) );
INVx2_ASAP7_75t_SL g273 ( .A(n_172), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_214), .Y(n_274) );
CKINVDCx14_ASAP7_75t_R g275 ( .A(n_184), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_193), .Y(n_276) );
INVx3_ASAP7_75t_L g277 ( .A(n_172), .Y(n_277) );
INVx1_ASAP7_75t_SL g278 ( .A(n_184), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_205), .Y(n_279) );
INVx3_ASAP7_75t_L g280 ( .A(n_176), .Y(n_280) );
INVxp67_ASAP7_75t_SL g281 ( .A(n_214), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_186), .B(n_151), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_176), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_205), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_227), .A2(n_162), .B1(n_161), .B2(n_141), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_167), .Y(n_286) );
INVx1_ASAP7_75t_SL g287 ( .A(n_166), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_168), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_166), .Y(n_289) );
NOR2x1_ASAP7_75t_L g290 ( .A(n_225), .B(n_151), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_170), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_222), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_195), .Y(n_293) );
INVx4_ASAP7_75t_L g294 ( .A(n_176), .Y(n_294) );
NAND2xp33_ASAP7_75t_R g295 ( .A(n_173), .B(n_179), .Y(n_295) );
NAND2xp33_ASAP7_75t_SL g296 ( .A(n_175), .B(n_161), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_246), .Y(n_297) );
NAND3xp33_ASAP7_75t_L g298 ( .A(n_256), .B(n_227), .C(n_215), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_240), .B(n_211), .Y(n_299) );
INVxp67_ASAP7_75t_L g300 ( .A(n_281), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_244), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_250), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_246), .B(n_213), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_257), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_244), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_232), .A2(n_174), .B(n_189), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_235), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_261), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_235), .Y(n_309) );
AND2x2_ASAP7_75t_SL g310 ( .A(n_246), .B(n_216), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_257), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_248), .Y(n_312) );
AOI222xp33_ASAP7_75t_L g313 ( .A1(n_287), .A2(n_165), .B1(n_213), .B2(n_207), .C1(n_206), .C2(n_135), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_240), .B(n_213), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_250), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_239), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_248), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_261), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_292), .B(n_224), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g320 ( .A1(n_259), .A2(n_177), .B1(n_200), .B2(n_196), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_264), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_239), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_259), .B(n_260), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_262), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_252), .A2(n_224), .B1(n_223), .B2(n_216), .Y(n_325) );
BUFx8_ASAP7_75t_L g326 ( .A(n_230), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_259), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_260), .B(n_224), .Y(n_328) );
BUFx8_ASAP7_75t_L g329 ( .A(n_274), .Y(n_329) );
BUFx4f_ASAP7_75t_SL g330 ( .A(n_278), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_243), .B(n_200), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_295), .A2(n_223), .B1(n_216), .B2(n_220), .Y(n_332) );
INVx2_ASAP7_75t_SL g333 ( .A(n_260), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_262), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_274), .B(n_223), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_264), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g337 ( .A1(n_289), .A2(n_189), .B1(n_188), .B2(n_194), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_252), .A2(n_192), .B1(n_202), .B2(n_222), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_230), .B(n_135), .Y(n_339) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_262), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_266), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_268), .A2(n_217), .B1(n_145), .B2(n_150), .Y(n_342) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_262), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_294), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_266), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_271), .B(n_217), .Y(n_346) );
NAND2x1_ASAP7_75t_L g347 ( .A(n_252), .B(n_197), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_301), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_332), .A2(n_291), .B1(n_288), .B2(n_286), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_340), .Y(n_350) );
INVx4_ASAP7_75t_L g351 ( .A(n_310), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_323), .B(n_233), .Y(n_352) );
INVx4_ASAP7_75t_SL g353 ( .A(n_323), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_331), .A2(n_275), .B1(n_276), .B2(n_255), .Y(n_354) );
AO31x2_ASAP7_75t_L g355 ( .A1(n_341), .A2(n_160), .A3(n_150), .B(n_145), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_298), .A2(n_276), .B1(n_255), .B2(n_271), .Y(n_356) );
OAI21x1_ASAP7_75t_L g357 ( .A1(n_324), .A2(n_334), .B(n_258), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_346), .B(n_271), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_313), .A2(n_296), .B1(n_285), .B2(n_263), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_310), .A2(n_276), .B1(n_255), .B2(n_242), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_346), .B(n_282), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_340), .Y(n_362) );
OA21x2_ASAP7_75t_L g363 ( .A1(n_324), .A2(n_126), .B(n_147), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_340), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g365 ( .A1(n_306), .A2(n_296), .B(n_279), .Y(n_365) );
INVx4_ASAP7_75t_L g366 ( .A(n_310), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g367 ( .A1(n_330), .A2(n_311), .B1(n_304), .B2(n_329), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_304), .Y(n_368) );
NAND2xp33_ASAP7_75t_R g369 ( .A(n_335), .B(n_251), .Y(n_369) );
INVx4_ASAP7_75t_L g370 ( .A(n_323), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_341), .A2(n_291), .B1(n_288), .B2(n_286), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_335), .A2(n_277), .B1(n_280), .B2(n_273), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_345), .A2(n_270), .B1(n_273), .B2(n_160), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_335), .A2(n_280), .B1(n_277), .B2(n_294), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_301), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_335), .A2(n_280), .B1(n_277), .B2(n_294), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_305), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_351), .A2(n_299), .B1(n_314), .B2(n_320), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_359), .A2(n_325), .B1(n_345), .B2(n_319), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_351), .A2(n_299), .B1(n_314), .B2(n_245), .Y(n_380) );
OAI21x1_ASAP7_75t_L g381 ( .A1(n_357), .A2(n_334), .B(n_305), .Y(n_381) );
INVx4_ASAP7_75t_L g382 ( .A(n_353), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_361), .B(n_282), .Y(n_383) );
OAI221xp5_ASAP7_75t_L g384 ( .A1(n_354), .A2(n_269), .B1(n_254), .B2(n_238), .C(n_249), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_348), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g386 ( .A1(n_351), .A2(n_300), .B1(n_308), .B2(n_318), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_361), .B(n_329), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_348), .B(n_308), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_375), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_375), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_351), .A2(n_245), .B1(n_303), .B2(n_290), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_377), .B(n_318), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_377), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_366), .A2(n_245), .B1(n_303), .B2(n_328), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_366), .B(n_321), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_355), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_358), .B(n_321), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_358), .B(n_336), .Y(n_398) );
OAI21xp33_ASAP7_75t_L g399 ( .A1(n_359), .A2(n_349), .B(n_356), .Y(n_399) );
AO21x2_ASAP7_75t_L g400 ( .A1(n_365), .A2(n_336), .B(n_147), .Y(n_400) );
INVx5_ASAP7_75t_L g401 ( .A(n_366), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_355), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_349), .A2(n_283), .B1(n_339), .B2(n_241), .C(n_160), .Y(n_403) );
INVx2_ASAP7_75t_SL g404 ( .A(n_353), .Y(n_404) );
AOI22xp33_ASAP7_75t_SL g405 ( .A1(n_366), .A2(n_326), .B1(n_303), .B2(n_328), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_385), .B(n_371), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_385), .B(n_371), .Y(n_407) );
NAND3xp33_ASAP7_75t_L g408 ( .A(n_399), .B(n_352), .C(n_369), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_389), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_389), .Y(n_410) );
OA21x2_ASAP7_75t_L g411 ( .A1(n_381), .A2(n_357), .B(n_147), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_401), .B(n_367), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_379), .A2(n_352), .B1(n_370), .B2(n_360), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_401), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_401), .B(n_353), .Y(n_415) );
INVx2_ASAP7_75t_SL g416 ( .A(n_401), .Y(n_416) );
AND2x6_ASAP7_75t_SL g417 ( .A(n_387), .B(n_368), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_389), .Y(n_418) );
AOI222xp33_ASAP7_75t_L g419 ( .A1(n_383), .A2(n_353), .B1(n_373), .B2(n_326), .C1(n_372), .C2(n_376), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_401), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_381), .Y(n_421) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_380), .A2(n_374), .B1(n_373), .B2(n_342), .C(n_338), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_378), .A2(n_337), .B1(n_370), .B2(n_132), .C(n_136), .Y(n_423) );
INVxp67_ASAP7_75t_L g424 ( .A(n_395), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_393), .Y(n_425) );
AOI22xp33_ASAP7_75t_SL g426 ( .A1(n_382), .A2(n_326), .B1(n_370), .B2(n_303), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_379), .A2(n_326), .B1(n_339), .B2(n_328), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_405), .A2(n_339), .B1(n_328), .B2(n_353), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_390), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_390), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_397), .B(n_355), .Y(n_431) );
AOI221xp5_ASAP7_75t_L g432 ( .A1(n_384), .A2(n_136), .B1(n_132), .B2(n_339), .C(n_95), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_397), .B(n_344), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_396), .B(n_355), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_396), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_394), .A2(n_344), .B1(n_317), .B2(n_302), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_434), .B(n_402), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_420), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_408), .A2(n_432), .B1(n_424), .B2(n_423), .C(n_427), .Y(n_439) );
BUFx3_ASAP7_75t_L g440 ( .A(n_420), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_415), .B(n_404), .Y(n_441) );
OAI22xp5_ASAP7_75t_SL g442 ( .A1(n_426), .A2(n_382), .B1(n_404), .B2(n_391), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_414), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_431), .B(n_388), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_431), .B(n_392), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_419), .A2(n_386), .B1(n_403), .B2(n_382), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_417), .B(n_398), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_417), .B(n_91), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_435), .Y(n_449) );
NOR3xp33_ASAP7_75t_L g450 ( .A(n_412), .B(n_94), .C(n_111), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_409), .B(n_392), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_435), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_429), .B(n_400), .Y(n_453) );
OAI31xp33_ASAP7_75t_L g454 ( .A1(n_408), .A2(n_95), .A3(n_317), .B(n_103), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_414), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_409), .B(n_136), .Y(n_456) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_421), .A2(n_143), .B(n_364), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_410), .B(n_400), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_414), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_430), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_418), .B(n_400), .Y(n_461) );
OAI221xp5_ASAP7_75t_L g462 ( .A1(n_428), .A2(n_344), .B1(n_307), .B2(n_309), .C(n_316), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_418), .B(n_6), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_430), .B(n_233), .Y(n_464) );
OAI31xp33_ASAP7_75t_L g465 ( .A1(n_423), .A2(n_323), .A3(n_322), .B(n_307), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_425), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_425), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g468 ( .A1(n_422), .A2(n_237), .B1(n_234), .B2(n_236), .C(n_231), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_411), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_406), .B(n_7), .Y(n_470) );
OAI31xp33_ASAP7_75t_L g471 ( .A1(n_422), .A2(n_297), .A3(n_312), .B(n_327), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_407), .B(n_364), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_407), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_419), .A2(n_363), .B1(n_315), .B2(n_302), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_411), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_440), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_444), .B(n_413), .Y(n_477) );
NOR3xp33_ASAP7_75t_L g478 ( .A(n_448), .B(n_433), .C(n_416), .Y(n_478) );
NAND3xp33_ASAP7_75t_L g479 ( .A(n_447), .B(n_415), .C(n_436), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_445), .B(n_415), .Y(n_480) );
INVx3_ASAP7_75t_L g481 ( .A(n_459), .Y(n_481) );
AND2x4_ASAP7_75t_SL g482 ( .A(n_459), .B(n_362), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_460), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_460), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_466), .Y(n_485) );
INVx2_ASAP7_75t_SL g486 ( .A(n_440), .Y(n_486) );
BUFx2_ASAP7_75t_L g487 ( .A(n_440), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_437), .B(n_411), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_470), .B(n_7), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_455), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_451), .B(n_9), .Y(n_491) );
NAND3x1_ASAP7_75t_SL g492 ( .A(n_454), .B(n_9), .C(n_10), .Y(n_492) );
NOR4xp25_ASAP7_75t_SL g493 ( .A(n_438), .B(n_10), .C(n_11), .D(n_12), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_467), .B(n_13), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_451), .B(n_470), .Y(n_495) );
NAND2xp33_ASAP7_75t_R g496 ( .A(n_438), .B(n_363), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_473), .B(n_14), .Y(n_497) );
NAND4xp25_ASAP7_75t_L g498 ( .A(n_446), .B(n_17), .C(n_18), .D(n_20), .Y(n_498) );
AO21x1_ASAP7_75t_L g499 ( .A1(n_463), .A2(n_17), .B(n_350), .Y(n_499) );
NAND4xp25_ASAP7_75t_L g500 ( .A(n_474), .B(n_237), .C(n_171), .D(n_190), .Y(n_500) );
INVxp67_ASAP7_75t_L g501 ( .A(n_453), .Y(n_501) );
AND3x1_ASAP7_75t_L g502 ( .A(n_450), .B(n_297), .C(n_312), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_442), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_443), .B(n_31), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_449), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_458), .B(n_37), .Y(n_506) );
OAI21xp33_ASAP7_75t_L g507 ( .A1(n_498), .A2(n_453), .B(n_461), .Y(n_507) );
AOI21xp33_ASAP7_75t_SL g508 ( .A1(n_478), .A2(n_465), .B(n_454), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_490), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_479), .A2(n_439), .B1(n_462), .B2(n_459), .Y(n_510) );
NAND2x1p5_ASAP7_75t_L g511 ( .A(n_502), .B(n_441), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_487), .Y(n_512) );
OAI321xp33_ASAP7_75t_L g513 ( .A1(n_489), .A2(n_468), .A3(n_464), .B1(n_452), .B2(n_475), .C(n_472), .Y(n_513) );
AOI21xp33_ASAP7_75t_SL g514 ( .A1(n_478), .A2(n_471), .B(n_456), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_480), .B(n_456), .Y(n_515) );
NOR2x1_ASAP7_75t_L g516 ( .A(n_494), .B(n_469), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_483), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_476), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_477), .A2(n_457), .B1(n_347), .B2(n_284), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_495), .B(n_457), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_485), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_484), .B(n_39), .Y(n_522) );
AOI21xp33_ASAP7_75t_SL g523 ( .A1(n_496), .A2(n_42), .B(n_49), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_499), .A2(n_347), .B1(n_284), .B2(n_267), .Y(n_524) );
OAI21xp33_ASAP7_75t_L g525 ( .A1(n_501), .A2(n_197), .B(n_178), .Y(n_525) );
AOI21xp33_ASAP7_75t_L g526 ( .A1(n_496), .A2(n_50), .B(n_51), .Y(n_526) );
INVx3_ASAP7_75t_L g527 ( .A(n_481), .Y(n_527) );
OAI22xp33_ASAP7_75t_L g528 ( .A1(n_500), .A2(n_297), .B1(n_327), .B2(n_333), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_488), .B(n_52), .Y(n_529) );
AOI332xp33_ASAP7_75t_L g530 ( .A1(n_491), .A2(n_178), .A3(n_57), .B1(n_61), .B2(n_64), .B3(n_71), .C1(n_253), .C2(n_272), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_512), .B(n_486), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_509), .B(n_497), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_521), .Y(n_533) );
AOI211x1_ASAP7_75t_L g534 ( .A1(n_507), .A2(n_506), .B(n_504), .C(n_505), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_509), .B(n_481), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_512), .B(n_508), .Y(n_536) );
NOR4xp25_ASAP7_75t_SL g537 ( .A(n_523), .B(n_492), .C(n_493), .D(n_482), .Y(n_537) );
INVx2_ASAP7_75t_SL g538 ( .A(n_518), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_517), .Y(n_539) );
INVxp67_ASAP7_75t_L g540 ( .A(n_516), .Y(n_540) );
OAI21xp5_ASAP7_75t_SL g541 ( .A1(n_511), .A2(n_482), .B(n_492), .Y(n_541) );
INVxp67_ASAP7_75t_L g542 ( .A(n_520), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_515), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_533), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_541), .A2(n_510), .B(n_513), .Y(n_545) );
AOI221xp5_ASAP7_75t_L g546 ( .A1(n_534), .A2(n_514), .B1(n_513), .B2(n_526), .C(n_527), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_531), .Y(n_547) );
OAI322xp33_ASAP7_75t_L g548 ( .A1(n_542), .A2(n_519), .A3(n_529), .B1(n_524), .B2(n_522), .C1(n_528), .C2(n_530), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_535), .B(n_525), .Y(n_549) );
AO22x1_ASAP7_75t_L g550 ( .A1(n_538), .A2(n_343), .B1(n_279), .B2(n_267), .Y(n_550) );
XOR2x2_ASAP7_75t_L g551 ( .A(n_532), .B(n_343), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_543), .A2(n_279), .B1(n_267), .B2(n_343), .Y(n_552) );
OAI22xp33_ASAP7_75t_SL g553 ( .A1(n_540), .A2(n_247), .B1(n_253), .B2(n_265), .Y(n_553) );
NOR2xp33_ASAP7_75t_R g554 ( .A(n_547), .B(n_539), .Y(n_554) );
INVx2_ASAP7_75t_SL g555 ( .A(n_551), .Y(n_555) );
NOR2xp33_ASAP7_75t_R g556 ( .A(n_549), .B(n_537), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_548), .A2(n_293), .B1(n_553), .B2(n_544), .Y(n_557) );
AND4x1_ASAP7_75t_L g558 ( .A(n_552), .B(n_545), .C(n_536), .D(n_546), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_550), .A2(n_503), .B1(n_545), .B2(n_536), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_555), .B(n_559), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_556), .Y(n_561) );
NAND3xp33_ASAP7_75t_SL g562 ( .A(n_558), .B(n_554), .C(n_557), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_560), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_563), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_564), .Y(n_565) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_565), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_566), .A2(n_561), .B(n_562), .Y(n_567) );
endmodule