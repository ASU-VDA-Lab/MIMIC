module fake_jpeg_17139_n_112 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_112);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_112;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx6_ASAP7_75t_SL g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_12),
.B(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_2),
.Y(n_25)
);

OR2x2_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_2),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_16),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_25),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_13),
.B1(n_18),
.B2(n_15),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_16),
.B1(n_21),
.B2(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_37),
.B(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_45),
.Y(n_58)
);

OA21x2_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_40),
.B(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_24),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_27),
.C(n_20),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_35),
.B1(n_28),
.B2(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_15),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_46),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_19),
.B(n_24),
.C(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_14),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_23),
.B1(n_14),
.B2(n_20),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_35),
.B1(n_28),
.B2(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_3),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_3),
.Y(n_63)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_45),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_51),
.B(n_54),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_42),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_30),
.B(n_35),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_55),
.B(n_4),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_20),
.B(n_17),
.Y(n_55)
);

OAI211xp5_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_63),
.B(n_4),
.C(n_5),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_27),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_32),
.B(n_17),
.Y(n_71)
);

AO22x1_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_39),
.B1(n_41),
.B2(n_37),
.Y(n_64)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_60),
.C(n_54),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_73),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_58),
.B(n_17),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_53),
.C(n_55),
.Y(n_80)
);

NAND2xp67_ASAP7_75t_SL g81 ( 
.A(n_71),
.B(n_76),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_7),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_75),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_77),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_7),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_86),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_51),
.B1(n_59),
.B2(n_57),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_84),
.B1(n_59),
.B2(n_81),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_60),
.C(n_57),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_71),
.B(n_64),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_94),
.Y(n_96)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_86),
.B(n_68),
.CI(n_63),
.CON(n_90),
.SN(n_90)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_91),
.Y(n_97)
);

NOR2xp67_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_76),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_92),
.A2(n_80),
.B1(n_64),
.B2(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_98),
.Y(n_103)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

BUFx4f_ASAP7_75t_SL g99 ( 
.A(n_89),
.Y(n_99)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_99),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_103),
.Y(n_105)
);

OAI21x1_ASAP7_75t_L g102 ( 
.A1(n_95),
.A2(n_90),
.B(n_88),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_97),
.B(n_99),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_105),
.C(n_107),
.Y(n_108)
);

AOI31xp67_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_83),
.A3(n_69),
.B(n_6),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_6),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_100),
.A2(n_69),
.B(n_67),
.Y(n_107)
);

AOI332xp33_ASAP7_75t_L g109 ( 
.A1(n_106),
.A2(n_100),
.A3(n_8),
.B1(n_9),
.B2(n_6),
.B3(n_74),
.C1(n_61),
.C2(n_32),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_110),
.B(n_61),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_108),
.Y(n_112)
);


endmodule