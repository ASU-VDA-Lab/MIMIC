module real_jpeg_22038_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx13_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_1),
.A2(n_55),
.B1(n_56),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_1),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_84),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_2),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_66),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_3),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_3),
.A2(n_55),
.B1(n_56),
.B2(n_75),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_75),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_4),
.A2(n_41),
.B1(n_49),
.B2(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_4),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_49),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_7),
.A2(n_26),
.B(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_7),
.A2(n_103),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_9),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_58),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_9),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_10),
.B(n_38),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g119 ( 
.A1(n_10),
.A2(n_14),
.B(n_28),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_10),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_10),
.A2(n_30),
.B1(n_127),
.B2(n_128),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_10),
.B(n_143),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g156 ( 
.A1(n_10),
.A2(n_38),
.B(n_99),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_14),
.A2(n_55),
.B(n_79),
.C(n_80),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_14),
.B(n_55),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_81),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_14),
.Y(n_81)
);

INVx11_ASAP7_75t_SL g55 ( 
.A(n_15),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_106),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_105),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_89),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_20),
.B(n_89),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_67),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_45),
.B2(n_46),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_29),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_30),
.B(n_65),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_30),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_30),
.A2(n_113),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_30),
.A2(n_115),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_31),
.B(n_65),
.Y(n_104)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_31),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_31),
.B(n_43),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_40),
.B2(n_44),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_41),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_37),
.A2(n_41),
.B(n_44),
.C(n_61),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_51),
.B(n_53),
.C(n_54),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_51),
.Y(n_53)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI32xp33_ASAP7_75t_L g98 ( 
.A1(n_39),
.A2(n_52),
.A3(n_55),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_61),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

HAxp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_43),
.CON(n_40),
.SN(n_40)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_60),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_43),
.A2(n_56),
.B(n_81),
.C(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_43),
.B(n_80),
.Y(n_130)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_59),
.C(n_62),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_47),
.B(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_54),
.B2(n_57),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_48),
.A2(n_50),
.B1(n_54),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_54),
.B1(n_57),
.B2(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_51),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g100 ( 
.A(n_51),
.B(n_56),
.Y(n_100)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_54),
.Y(n_143)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_62),
.B1(n_63),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_76),
.B1(n_77),
.B2(n_88),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_82),
.B(n_85),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_78),
.A2(n_80),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_78),
.A2(n_80),
.B1(n_123),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_78),
.A2(n_80),
.B1(n_95),
.B2(n_146),
.Y(n_158)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_83),
.B(n_87),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.C(n_97),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_90),
.A2(n_91),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_94),
.B(n_97),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_98),
.B(n_101),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B(n_104),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_129),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_163),
.B(n_168),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_150),
.B(n_162),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_137),
.B(n_149),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_124),
.B(n_136),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_116),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_118),
.B(n_120),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_131),
.B(n_135),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_130),
.Y(n_135)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_138),
.B(n_139),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_147),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_145),
.C(n_147),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_152),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_160),
.B2(n_161),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_153),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_155),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_159),
.C(n_160),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_164),
.B(n_165),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);


endmodule