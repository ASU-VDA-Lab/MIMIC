module fake_jpeg_14174_n_251 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_53),
.Y(n_81)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_16),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_65),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_19),
.B(n_23),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g109 ( 
.A(n_54),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_19),
.B(n_3),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_60),
.Y(n_84)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_3),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_68),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_4),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_15),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_67),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_24),
.B(n_6),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_72),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_70),
.B(n_71),
.Y(n_121)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

CKINVDCx9p33_ASAP7_75t_R g72 ( 
.A(n_36),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_25),
.B(n_6),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_25),
.B(n_6),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_76),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_26),
.B(n_7),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_R g77 ( 
.A(n_39),
.B(n_14),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_70),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_79),
.Y(n_89)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_29),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_32),
.B1(n_30),
.B2(n_21),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_83),
.A2(n_45),
.B1(n_54),
.B2(n_47),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_44),
.A2(n_26),
.B1(n_35),
.B2(n_31),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_85),
.A2(n_114),
.B1(n_90),
.B2(n_119),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_72),
.A2(n_21),
.B1(n_32),
.B2(n_30),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_87),
.B(n_98),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_49),
.A2(n_20),
.B1(n_18),
.B2(n_37),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_95),
.A2(n_103),
.B1(n_111),
.B2(n_113),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_37),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_71),
.A2(n_20),
.B1(n_35),
.B2(n_29),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_75),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_43),
.A2(n_31),
.B1(n_9),
.B2(n_11),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_108),
.A2(n_119),
.B1(n_118),
.B2(n_97),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_63),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_8),
.C(n_11),
.Y(n_112)
);

A2O1A1O1Ixp25_ASAP7_75t_L g146 ( 
.A1(n_112),
.A2(n_121),
.B(n_115),
.C(n_109),
.D(n_106),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_56),
.A2(n_12),
.B1(n_62),
.B2(n_58),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_52),
.A2(n_12),
.B1(n_67),
.B2(n_64),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_120),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_78),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_82),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_75),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_124),
.Y(n_160)
);

AO22x1_ASAP7_75t_SL g125 ( 
.A1(n_116),
.A2(n_69),
.B1(n_96),
.B2(n_100),
.Y(n_125)
);

AO21x2_ASAP7_75t_L g166 ( 
.A1(n_125),
.A2(n_155),
.B(n_140),
.Y(n_166)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_69),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_129),
.B(n_132),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_89),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_144),
.Y(n_170)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_81),
.B(n_86),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_92),
.B(n_88),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_134),
.B(n_136),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_83),
.B(n_93),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_91),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_112),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_96),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_143),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_115),
.B(n_87),
.C(n_101),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_143),
.B(n_135),
.Y(n_165)
);

INVx4_ASAP7_75t_SL g141 ( 
.A(n_105),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_141),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_142),
.A2(n_151),
.B(n_154),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_121),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_94),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_149),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_R g181 ( 
.A(n_146),
.B(n_125),
.Y(n_181)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_150),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_SL g167 ( 
.A(n_148),
.B(n_150),
.C(n_144),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_110),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_97),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_122),
.B1(n_105),
.B2(n_107),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_107),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_155),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_89),
.B(n_83),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_98),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_92),
.B(n_81),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_158),
.Y(n_182)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_171),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_166),
.A2(n_127),
.B1(n_157),
.B2(n_131),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_167),
.A2(n_172),
.B1(n_181),
.B2(n_166),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_126),
.A2(n_159),
.B(n_142),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_139),
.B1(n_130),
.B2(n_137),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_159),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g198 ( 
.A(n_174),
.B(n_186),
.Y(n_198)
);

A2O1A1O1Ixp25_ASAP7_75t_L g179 ( 
.A1(n_125),
.A2(n_126),
.B(n_146),
.C(n_156),
.D(n_134),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_179),
.B(n_141),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_152),
.B(n_158),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_133),
.B(n_147),
.Y(n_186)
);

AOI221xp5_ASAP7_75t_L g216 ( 
.A1(n_187),
.A2(n_195),
.B1(n_196),
.B2(n_204),
.C(n_191),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_188),
.B(n_191),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_128),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_190),
.Y(n_217)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_192),
.B(n_193),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_169),
.B(n_141),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_176),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_201),
.Y(n_214)
);

AOI322xp5_ASAP7_75t_SL g195 ( 
.A1(n_182),
.A2(n_163),
.A3(n_178),
.B1(n_171),
.B2(n_164),
.C1(n_173),
.C2(n_179),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_178),
.C(n_164),
.Y(n_196)
);

AO21x2_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_165),
.B(n_167),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_203),
.B1(n_200),
.B2(n_166),
.Y(n_206)
);

BUFx12_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

NAND2x1_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_201),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_175),
.Y(n_210)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_172),
.A2(n_170),
.B1(n_166),
.B2(n_177),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_174),
.Y(n_204)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_186),
.C(n_180),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_205),
.C(n_198),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_160),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_216),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_210),
.A2(n_212),
.B(n_213),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_197),
.A2(n_184),
.B1(n_183),
.B2(n_175),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_188),
.B(n_197),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_185),
.B(n_183),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_203),
.B1(n_192),
.B2(n_202),
.Y(n_218)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_218),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_218),
.B1(n_211),
.B2(n_206),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_205),
.C(n_198),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_222),
.A2(n_197),
.B1(n_210),
.B2(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_207),
.Y(n_233)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_233),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_209),
.C(n_220),
.Y(n_238)
);

AO21x1_ASAP7_75t_L g231 ( 
.A1(n_223),
.A2(n_207),
.B(n_210),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_231),
.A2(n_223),
.B(n_221),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_228),
.A2(n_215),
.B1(n_212),
.B2(n_194),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_215),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_231),
.B1(n_232),
.B2(n_229),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_228),
.Y(n_237)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_237),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_239),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_236),
.A2(n_221),
.B1(n_219),
.B2(n_230),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_241),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_242),
.A2(n_232),
.B(n_222),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_246),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_224),
.C(n_231),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_245),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_249),
.A2(n_248),
.B(n_243),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_240),
.Y(n_251)
);


endmodule