module fake_jpeg_29117_n_33 (n_3, n_2, n_1, n_0, n_4, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_1),
.B(n_2),
.Y(n_6)
);

BUFx2_ASAP7_75t_R g7 ( 
.A(n_0),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_12),
.B(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_8),
.A2(n_4),
.B1(n_9),
.B2(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_25),
.A2(n_16),
.B1(n_19),
.B2(n_20),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_27),
.B1(n_7),
.B2(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_21),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_29),
.C(n_26),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_23),
.C(n_20),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_29),
.C(n_15),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_31),
.A2(n_24),
.B1(n_17),
.B2(n_13),
.Y(n_32)
);

AOI221xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_12),
.B1(n_24),
.B2(n_8),
.C(n_11),
.Y(n_33)
);


endmodule