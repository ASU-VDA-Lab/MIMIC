module fake_jpeg_5598_n_149 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_149);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_22),
.Y(n_56)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_39),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_2),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_46),
.Y(n_70)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_30),
.Y(n_64)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_55),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_52),
.B(n_71),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_19),
.B1(n_25),
.B2(n_18),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_62),
.B1(n_29),
.B2(n_31),
.Y(n_89)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_60),
.Y(n_94)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_67),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_24),
.B1(n_18),
.B2(n_25),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_68),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_33),
.B(n_22),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_66),
.B(n_65),
.Y(n_98)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_30),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_20),
.B1(n_27),
.B2(n_26),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_76),
.B1(n_67),
.B2(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_33),
.A2(n_21),
.B(n_27),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_74),
.A2(n_75),
.B(n_29),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_33),
.A2(n_26),
.B(n_23),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_23),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_91),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_74),
.A2(n_17),
.B(n_6),
.C(n_7),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_98),
.B(n_51),
.Y(n_102)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_76),
.A2(n_32),
.B1(n_29),
.B2(n_31),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_2),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_8),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_54),
.A2(n_31),
.B1(n_32),
.B2(n_9),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_55),
.B1(n_57),
.B2(n_50),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_58),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_85),
.B(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_104),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_110),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_SL g121 ( 
.A1(n_109),
.A2(n_95),
.B(n_80),
.C(n_79),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_94),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_81),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_32),
.B(n_9),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_117),
.B(n_113),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_106),
.B1(n_103),
.B2(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_90),
.B(n_97),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_93),
.C(n_89),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_116),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_121),
.B1(n_123),
.B2(n_106),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_131),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_111),
.B(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_126),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_138),
.B(n_140),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_134),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_127),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_133),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_144),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_146),
.B1(n_145),
.B2(n_111),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_99),
.Y(n_149)
);


endmodule