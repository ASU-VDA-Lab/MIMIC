module fake_jpeg_3017_n_229 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_229);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_5),
.B(n_9),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_4),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_35),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_44),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_22),
.Y(n_77)
);

BUFx24_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_11),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_58),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_86),
.Y(n_91)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_82),
.A2(n_75),
.B1(n_63),
.B2(n_78),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_74),
.B1(n_59),
.B2(n_54),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_75),
.B1(n_60),
.B2(n_56),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_99),
.B1(n_79),
.B2(n_87),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_84),
.B(n_61),
.Y(n_93)
);

OR2x2_ASAP7_75t_SL g103 ( 
.A(n_93),
.B(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_96),
.B(n_74),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_56),
.B1(n_60),
.B2(n_67),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_72),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_73),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_112),
.Y(n_124)
);

HAxp5_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_78),
.CON(n_102),
.SN(n_102)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_105),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_99),
.A2(n_77),
.B1(n_76),
.B2(n_67),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_115),
.B1(n_119),
.B2(n_90),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_71),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_113),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_54),
.B1(n_62),
.B2(n_70),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_107),
.A2(n_118),
.B1(n_1),
.B2(n_6),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_62),
.B1(n_70),
.B2(n_71),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_95),
.A2(n_57),
.B1(n_68),
.B2(n_59),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_97),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_57),
.B1(n_79),
.B2(n_3),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_119)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_136),
.B1(n_137),
.B2(n_13),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_24),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_131),
.Y(n_149)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_130),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_23),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_121),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_141),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_97),
.B1(n_4),
.B2(n_5),
.Y(n_136)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_28),
.C(n_52),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_30),
.C(n_47),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_110),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_33),
.Y(n_166)
);

AO21x2_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_25),
.B(n_50),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_157),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_6),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_144),
.B(n_146),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_7),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_150),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_140),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_21),
.C(n_49),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_152),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_7),
.B(n_8),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_9),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_155),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_10),
.B(n_12),
.C(n_13),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_29),
.C(n_45),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_161),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_12),
.Y(n_159)
);

NAND2xp33_ASAP7_75t_R g167 ( 
.A(n_159),
.B(n_160),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_121),
.A2(n_14),
.B(n_15),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_137),
.A2(n_36),
.B1(n_42),
.B2(n_40),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_163),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_129),
.C(n_120),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_14),
.Y(n_164)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_145),
.B1(n_143),
.B2(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_171),
.Y(n_188)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_143),
.A2(n_136),
.B1(n_138),
.B2(n_122),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_178),
.B1(n_181),
.B2(n_182),
.Y(n_197)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_143),
.A2(n_145),
.B1(n_148),
.B2(n_159),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_122),
.B1(n_17),
.B2(n_20),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_16),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_176),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_198),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_155),
.C(n_162),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_196),
.C(n_192),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_181),
.A2(n_38),
.B1(n_39),
.B2(n_53),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_194),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_172),
.A2(n_20),
.B1(n_177),
.B2(n_171),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_182),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_173),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_174),
.Y(n_213)
);

BUFx24_ASAP7_75t_SL g201 ( 
.A(n_189),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_204),
.Y(n_212)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_202),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_179),
.C(n_170),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_175),
.C(n_169),
.Y(n_211)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_188),
.A2(n_172),
.B1(n_178),
.B2(n_167),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_207),
.B(n_199),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_168),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_193),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_205),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_214),
.Y(n_217)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_208),
.B(n_186),
.CI(n_206),
.CON(n_215),
.SN(n_215)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_210),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_217),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

XNOR2x1_ASAP7_75t_SL g223 ( 
.A(n_222),
.B(n_220),
.Y(n_223)
);

NOR3xp33_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_211),
.C(n_216),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_224),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_226),
.A2(n_212),
.B(n_213),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_215),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_209),
.Y(n_229)
);


endmodule