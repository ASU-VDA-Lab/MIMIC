module fake_jpeg_16992_n_69 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_69);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_69;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_6),
.B(n_8),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

FAx1_ASAP7_75t_SL g19 ( 
.A(n_14),
.B(n_3),
.CI(n_5),
.CON(n_19),
.SN(n_19)
);

FAx1_ASAP7_75t_SL g42 ( 
.A(n_19),
.B(n_24),
.CI(n_20),
.CON(n_42),
.SN(n_42)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_28),
.Y(n_35)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_10),
.A2(n_1),
.B1(n_7),
.B2(n_8),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_1),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_9),
.A2(n_15),
.B(n_11),
.C(n_13),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_17),
.B(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_36),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_15),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_42),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_39),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_42),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_21),
.A2(n_18),
.B1(n_25),
.B2(n_10),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_33),
.B1(n_38),
.B2(n_30),
.Y(n_50)
);

INVxp67_ASAP7_75t_SL g44 ( 
.A(n_32),
.Y(n_44)
);

HAxp5_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_48),
.CON(n_55),
.SN(n_55)
);

OAI21xp33_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_50),
.B(n_48),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_42),
.Y(n_48)
);

OAI32xp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_36),
.A3(n_39),
.B1(n_30),
.B2(n_35),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_50),
.B1(n_45),
.B2(n_43),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_51),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_57),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_54),
.B(n_57),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_56),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_64),
.B1(n_60),
.B2(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_59),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_62),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_66),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_67),
.Y(n_69)
);


endmodule