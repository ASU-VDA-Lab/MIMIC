module fake_jpeg_21330_n_280 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_280);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_32),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_36),
.Y(n_42)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_35),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_16),
.B1(n_29),
.B2(n_35),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_23),
.C(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_30),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_22),
.B(n_26),
.Y(n_87)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_63),
.Y(n_69)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_34),
.B1(n_29),
.B2(n_27),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_59),
.B1(n_64),
.B2(n_36),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_66),
.B1(n_67),
.B2(n_37),
.Y(n_71)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_29),
.B1(n_34),
.B2(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_49),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_23),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_44),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_34),
.B1(n_29),
.B2(n_14),
.Y(n_64)
);

AO22x1_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_36),
.B1(n_35),
.B2(n_32),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_16),
.B1(n_15),
.B2(n_35),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_71),
.A2(n_88),
.B1(n_85),
.B2(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_27),
.C(n_44),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_54),
.C(n_68),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_87),
.B(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_81),
.A2(n_55),
.B1(n_63),
.B2(n_62),
.Y(n_90)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_79),
.B1(n_62),
.B2(n_70),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_100),
.B(n_102),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_103),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_98),
.C(n_28),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_64),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_51),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_57),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_71),
.B1(n_53),
.B2(n_76),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_109),
.A2(n_125),
.B1(n_58),
.B2(n_56),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_66),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_110),
.A2(n_124),
.B(n_122),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_111),
.A2(n_118),
.B1(n_36),
.B2(n_45),
.Y(n_142)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_83),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_113),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_102),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_106),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_79),
.B1(n_62),
.B2(n_53),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_96),
.B(n_67),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_122),
.C(n_45),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_70),
.B(n_22),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_26),
.B(n_18),
.Y(n_141)
);

BUFx4f_ASAP7_75t_SL g123 ( 
.A(n_89),
.Y(n_123)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_36),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_124),
.A2(n_60),
.B(n_94),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_95),
.A2(n_76),
.B1(n_83),
.B2(n_77),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_130),
.A2(n_138),
.B(n_145),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_90),
.B1(n_97),
.B2(n_100),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_132),
.A2(n_140),
.B1(n_141),
.B2(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

OAI22x1_ASAP7_75t_SL g137 ( 
.A1(n_127),
.A2(n_97),
.B1(n_91),
.B2(n_94),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_31),
.B1(n_46),
.B2(n_65),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_60),
.B(n_32),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_28),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_107),
.B1(n_86),
.B2(n_72),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_144),
.B1(n_151),
.B2(n_126),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_110),
.A2(n_107),
.B1(n_72),
.B2(n_61),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_108),
.A2(n_18),
.B(n_13),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_23),
.Y(n_146)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_0),
.B(n_1),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_24),
.B1(n_25),
.B2(n_21),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_150),
.A2(n_153),
.B1(n_38),
.B2(n_40),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_61),
.B1(n_56),
.B2(n_38),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_26),
.B(n_18),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_120),
.C(n_128),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_156),
.C(n_174),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_129),
.C(n_115),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_159),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_148),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_160),
.A2(n_162),
.B1(n_166),
.B2(n_172),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_126),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_146),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_121),
.B1(n_116),
.B2(n_115),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_116),
.C(n_121),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_177),
.C(n_138),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_24),
.C(n_25),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_164),
.A2(n_141),
.B(n_147),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_112),
.B1(n_123),
.B2(n_38),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_167),
.B(n_170),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_123),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_132),
.A2(n_40),
.B1(n_15),
.B2(n_13),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_173),
.B1(n_178),
.B2(n_151),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_40),
.B1(n_15),
.B2(n_43),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_175),
.Y(n_179)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_140),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_182),
.C(n_187),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_184),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_162),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_130),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_188),
.A2(n_190),
.B1(n_194),
.B2(n_197),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_189),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_135),
.B1(n_152),
.B2(n_143),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_131),
.C(n_152),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_199),
.C(n_28),
.Y(n_212)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_174),
.B(n_161),
.CI(n_163),
.CON(n_192),
.SN(n_192)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_153),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_170),
.A2(n_178),
.B1(n_168),
.B2(n_160),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_196),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_149),
.B1(n_136),
.B2(n_134),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_195),
.A2(n_171),
.B1(n_157),
.B2(n_172),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_202),
.A2(n_209),
.B1(n_216),
.B2(n_217),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_205),
.B(n_206),
.Y(n_227)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_181),
.B(n_153),
.CI(n_136),
.CON(n_206),
.SN(n_206)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_210),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_213),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_1),
.B(n_2),
.Y(n_213)
);

O2A1O1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_186),
.A2(n_25),
.B(n_24),
.C(n_31),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_214),
.A2(n_21),
.B1(n_4),
.B2(n_5),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_180),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_190),
.A2(n_31),
.B1(n_19),
.B2(n_43),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_187),
.B1(n_194),
.B2(n_192),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_220),
.A2(n_229),
.B1(n_209),
.B2(n_202),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_182),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_223),
.Y(n_243)
);

NOR2x1_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_188),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_199),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_193),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_226),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_179),
.C(n_43),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_205),
.C(n_206),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_231),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_201),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_3),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_215),
.C(n_204),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_236),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_201),
.C(n_216),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_245),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_206),
.Y(n_238)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_219),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_244),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_228),
.B(n_214),
.Y(n_241)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_21),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_226),
.Y(n_248)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_230),
.C(n_220),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_245),
.C(n_43),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_218),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_250),
.B(n_254),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_238),
.B(n_229),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_17),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_233),
.A2(n_239),
.B(n_222),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_250),
.C(n_247),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_261),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_256),
.B(n_19),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_253),
.A2(n_46),
.B1(n_19),
.B2(n_17),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_263),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_23),
.C(n_17),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_4),
.B(n_5),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_264),
.B(n_265),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_255),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_271),
.B(n_11),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_258),
.C(n_259),
.Y(n_272)
);

NAND2xp33_ASAP7_75t_SL g271 ( 
.A(n_260),
.B(n_247),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_272),
.A2(n_273),
.B(n_274),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_5),
.C(n_6),
.Y(n_274)
);

AOI321xp33_ASAP7_75t_L g276 ( 
.A1(n_273),
.A2(n_267),
.A3(n_269),
.B1(n_266),
.B2(n_9),
.C(n_6),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_6),
.B(n_7),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_275),
.C(n_8),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_279),
.A2(n_7),
.B(n_9),
.Y(n_280)
);


endmodule