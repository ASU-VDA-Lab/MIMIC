module fake_jpeg_20977_n_377 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_377);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_377;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx6p67_ASAP7_75t_R g93 ( 
.A(n_59),
.Y(n_93)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_27),
.B(n_8),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_62),
.B(n_19),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_8),
.C(n_15),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_33),
.C(n_43),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_37),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_75),
.Y(n_106)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_27),
.B(n_8),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_77),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_35),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_80),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_28),
.B(n_16),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_34),
.B1(n_28),
.B2(n_29),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_82),
.A2(n_84),
.B1(n_105),
.B2(n_110),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_64),
.B1(n_34),
.B2(n_55),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_87),
.B(n_35),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_29),
.B(n_40),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_88),
.A2(n_0),
.B(n_2),
.Y(n_153)
);

OR2x4_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_89),
.B(n_102),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_94),
.B(n_114),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_43),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_52),
.A2(n_34),
.B1(n_40),
.B2(n_26),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_24),
.B1(n_30),
.B2(n_40),
.Y(n_107)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_65),
.A3(n_63),
.B1(n_39),
.B2(n_36),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_45),
.A2(n_30),
.B1(n_41),
.B2(n_38),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_48),
.A2(n_35),
.B1(n_19),
.B2(n_33),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_112),
.A2(n_126),
.B1(n_3),
.B2(n_5),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_81),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_115),
.B(n_117),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_31),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_122),
.B(n_123),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_69),
.B(n_31),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_66),
.A2(n_26),
.B1(n_25),
.B2(n_38),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_128),
.B1(n_35),
.B2(n_59),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_56),
.A2(n_25),
.B1(n_41),
.B2(n_38),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_58),
.A2(n_41),
.B1(n_25),
.B2(n_32),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_72),
.B(n_44),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_130),
.Y(n_151)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_50),
.Y(n_131)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_SL g132 ( 
.A(n_61),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_71),
.C(n_77),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_137),
.B(n_133),
.C(n_91),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_138),
.A2(n_161),
.B1(n_168),
.B2(n_172),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_39),
.B(n_2),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_139),
.A2(n_153),
.B(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_142),
.B(n_7),
.Y(n_200)
);

BUFx2_ASAP7_75t_SL g143 ( 
.A(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_143),
.Y(n_207)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_157),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_111),
.A2(n_79),
.B1(n_36),
.B2(n_32),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_147),
.B1(n_150),
.B2(n_152),
.Y(n_178)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_39),
.B1(n_35),
.B2(n_44),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_107),
.B(n_83),
.C(n_124),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_149),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_35),
.B1(n_9),
.B2(n_10),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_107),
.A2(n_0),
.B(n_2),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_154),
.A2(n_155),
.B(n_116),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_100),
.A2(n_0),
.B(n_2),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_86),
.A2(n_9),
.B1(n_14),
.B2(n_12),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_112),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_164),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_97),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_166),
.B(n_169),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_98),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_97),
.Y(n_169)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

O2A1O1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_110),
.A2(n_103),
.B(n_120),
.C(n_98),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_96),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_173),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_99),
.A2(n_16),
.B1(n_6),
.B2(n_7),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_6),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_85),
.B(n_5),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_174),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_176),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_SL g182 ( 
.A1(n_149),
.A2(n_108),
.B(n_103),
.C(n_120),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_182),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_157),
.A2(n_125),
.B1(n_101),
.B2(n_108),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_SL g222 ( 
.A1(n_183),
.A2(n_160),
.B(n_176),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_137),
.B(n_101),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_192),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_116),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_189),
.A2(n_159),
.B1(n_158),
.B2(n_134),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_164),
.B1(n_166),
.B2(n_169),
.Y(n_220)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_145),
.B(n_133),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_195),
.C(n_197),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_154),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_139),
.B(n_138),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_196),
.B(n_201),
.Y(n_246)
);

AND2x2_ASAP7_75t_SL g197 ( 
.A(n_142),
.B(n_92),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_205),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_170),
.B(n_92),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_204),
.B(n_211),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_155),
.B(n_129),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_129),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_213),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_142),
.B(n_104),
.C(n_95),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_151),
.C(n_171),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_170),
.B(n_162),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_212),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_93),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_93),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_148),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_196),
.A2(n_136),
.B1(n_172),
.B2(n_163),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_243),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_214),
.A2(n_136),
.B1(n_135),
.B2(n_141),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_191),
.A2(n_173),
.B1(n_151),
.B2(n_165),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_220),
.B(n_191),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_222),
.A2(n_230),
.B(n_236),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_240),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_229),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_180),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_228),
.B(n_198),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_167),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_144),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_140),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_233),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_140),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_205),
.A2(n_184),
.B(n_192),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_238),
.A2(n_244),
.B(n_188),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_158),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_228),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_187),
.B(n_134),
.C(n_210),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_182),
.A2(n_134),
.B1(n_209),
.B2(n_191),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_189),
.A2(n_182),
.B1(n_212),
.B2(n_195),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_260),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_177),
.B1(n_178),
.B2(n_193),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_253),
.A2(n_267),
.B1(n_217),
.B2(n_230),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_201),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_258),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_234),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_235),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_257),
.A2(n_259),
.B(n_265),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_200),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_226),
.A2(n_184),
.B(n_189),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_197),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_270),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_226),
.A2(n_213),
.B(n_208),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_224),
.A2(n_178),
.B1(n_193),
.B2(n_209),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_236),
.A2(n_197),
.B(n_190),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_269),
.A2(n_225),
.B(n_230),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_197),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_198),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_240),
.Y(n_280)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_272),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_273),
.A2(n_275),
.B1(n_281),
.B2(n_288),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_277),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_268),
.A2(n_246),
.B(n_245),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_SL g299 ( 
.A1(n_278),
.A2(n_264),
.B(n_253),
.C(n_265),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_286),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_247),
.B(n_221),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_282),
.B(n_251),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_239),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_283),
.Y(n_303)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_264),
.A2(n_227),
.B1(n_216),
.B2(n_244),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_267),
.B1(n_248),
.B2(n_263),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_260),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_290),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_252),
.B(n_218),
.C(n_223),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_293),
.C(n_295),
.Y(n_297)
);

AOI221xp5_ASAP7_75t_L g292 ( 
.A1(n_269),
.A2(n_215),
.B1(n_221),
.B2(n_225),
.C(n_230),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_292),
.A2(n_270),
.B1(n_247),
.B2(n_259),
.Y(n_307)
);

OAI322xp33_ASAP7_75t_L g293 ( 
.A1(n_261),
.A2(n_215),
.A3(n_218),
.B1(n_229),
.B2(n_232),
.C1(n_222),
.C2(n_237),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_233),
.Y(n_294)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_252),
.B(n_238),
.C(n_220),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_294),
.Y(n_296)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_296),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_268),
.B(n_257),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_298),
.A2(n_305),
.B1(n_311),
.B2(n_313),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g315 ( 
.A1(n_299),
.A2(n_289),
.B(n_276),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_271),
.C(n_255),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_310),
.C(n_295),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_307),
.B(n_288),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_258),
.C(n_262),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_285),
.A2(n_262),
.B1(n_261),
.B2(n_254),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_287),
.Y(n_312)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_312),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_287),
.A2(n_254),
.B1(n_251),
.B2(n_249),
.Y(n_313)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_314),
.Y(n_327)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_315),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_274),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_318),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_274),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_321),
.C(n_322),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_286),
.C(n_293),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_278),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_278),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_323),
.B(n_326),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_292),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_328),
.C(n_300),
.Y(n_342)
);

OA21x2_ASAP7_75t_SL g326 ( 
.A1(n_298),
.A2(n_282),
.B(n_290),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_305),
.Y(n_328)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_329),
.Y(n_333)
);

NOR3xp33_ASAP7_75t_SL g330 ( 
.A(n_299),
.B(n_277),
.C(n_283),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_330),
.B(n_303),
.Y(n_337)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_320),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_335),
.B(n_338),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_330),
.A2(n_309),
.B(n_299),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_336),
.A2(n_322),
.B1(n_249),
.B2(n_319),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_337),
.B(n_279),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_315),
.A2(n_311),
.B1(n_308),
.B2(n_276),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_327),
.A2(n_300),
.B1(n_308),
.B2(n_284),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_340),
.Y(n_349)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_317),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_341),
.B(n_343),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_342),
.B(n_331),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_324),
.A2(n_299),
.B1(n_306),
.B2(n_279),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_342),
.B(n_329),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_345),
.B(n_353),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_332),
.C(n_316),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_335),
.B(n_328),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_350),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_334),
.B(n_306),
.Y(n_350)
);

NAND4xp25_ASAP7_75t_L g351 ( 
.A(n_343),
.B(n_313),
.C(n_321),
.D(n_325),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_351),
.A2(n_339),
.B(n_331),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_352),
.Y(n_357)
);

NAND4xp25_ASAP7_75t_SL g353 ( 
.A(n_336),
.B(n_203),
.C(n_186),
.D(n_202),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_354),
.B(n_207),
.Y(n_362)
);

OAI221xp5_ASAP7_75t_L g355 ( 
.A1(n_352),
.A2(n_353),
.B1(n_339),
.B2(n_333),
.C(n_349),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_355),
.B(n_346),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_358),
.B(n_360),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_359),
.B(n_347),
.C(n_345),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_344),
.B(n_338),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_350),
.A2(n_318),
.B1(n_332),
.B2(n_186),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_361),
.B(n_362),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_364),
.B(n_367),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_362),
.B(n_349),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_368),
.B(n_369),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_363),
.B(n_199),
.Y(n_369)
);

AOI321xp33_ASAP7_75t_L g370 ( 
.A1(n_365),
.A2(n_357),
.A3(n_356),
.B1(n_360),
.B2(n_199),
.C(n_203),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_370),
.B(n_372),
.Y(n_374)
);

A2O1A1Ixp33_ASAP7_75t_L g372 ( 
.A1(n_366),
.A2(n_206),
.B(n_207),
.C(n_367),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_373),
.A2(n_371),
.B(n_206),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_375),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_376),
.B(n_374),
.Y(n_377)
);


endmodule