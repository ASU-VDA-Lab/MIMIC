module fake_jpeg_13443_n_187 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_187);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_11),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_27),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_23),
.B(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_21),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_40),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_14),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_0),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_1),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_87),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_2),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_60),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_75),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_103),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_56),
.B1(n_64),
.B2(n_73),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_53),
.B1(n_67),
.B2(n_52),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_79),
.B1(n_77),
.B2(n_57),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_73),
.C(n_74),
.Y(n_122)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_100),
.B(n_62),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_110),
.Y(n_128)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_109),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_100),
.B(n_58),
.CI(n_4),
.CON(n_110),
.SN(n_110)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_63),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_121),
.Y(n_139)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_76),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_122),
.A2(n_9),
.B(n_13),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_67),
.B1(n_79),
.B2(n_77),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_89),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_71),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_126),
.C(n_55),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_68),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_72),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_120),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_145),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_131),
.B(n_136),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_118),
.B(n_26),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_17),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_55),
.B1(n_58),
.B2(n_5),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_137),
.A2(n_144),
.B1(n_28),
.B2(n_31),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_146),
.B1(n_48),
.B2(n_30),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_3),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_141),
.B(n_130),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_6),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_146)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_15),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_139),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_152),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_139),
.Y(n_152)
);

A2O1A1O1Ixp25_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_126),
.B(n_125),
.C(n_18),
.D(n_20),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_155),
.A2(n_166),
.B(n_32),
.Y(n_173)
);

AOI21x1_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_141),
.B(n_132),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_164),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_145),
.B1(n_134),
.B2(n_128),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_143),
.B1(n_140),
.B2(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_24),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_165),
.Y(n_168)
);

NOR2xp67_ASAP7_75t_R g175 ( 
.A(n_167),
.B(n_173),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_158),
.A2(n_36),
.B(n_38),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_157),
.Y(n_178)
);

NAND4xp25_ASAP7_75t_SL g177 ( 
.A(n_170),
.B(n_158),
.C(n_161),
.D(n_154),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_178),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_153),
.C(n_168),
.Y(n_179)
);

OA21x2_ASAP7_75t_SL g181 ( 
.A1(n_179),
.A2(n_155),
.B(n_175),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_180),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_182),
.A2(n_168),
.B1(n_176),
.B2(n_172),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_166),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

OAI311xp33_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_171),
.A3(n_156),
.B1(n_43),
.C1(n_44),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_39),
.Y(n_187)
);


endmodule