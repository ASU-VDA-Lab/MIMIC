module fake_jpeg_1349_n_182 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_182);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_36),
.Y(n_48)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_39),
.B(n_43),
.Y(n_71)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_13),
.B(n_11),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_25),
.B1(n_22),
.B2(n_27),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_53),
.B1(n_54),
.B2(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_25),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_54),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_22),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_59),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_13),
.B1(n_16),
.B2(n_14),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_26),
.B1(n_21),
.B2(n_15),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_29),
.A2(n_14),
.B1(n_16),
.B2(n_28),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_35),
.B1(n_38),
.B2(n_30),
.Y(n_73)
);

CKINVDCx12_ASAP7_75t_R g58 ( 
.A(n_30),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_31),
.A2(n_20),
.B1(n_19),
.B2(n_17),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_60),
.A2(n_63),
.B1(n_8),
.B2(n_9),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_29),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_66),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_31),
.A2(n_20),
.B1(n_19),
.B2(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_1),
.Y(n_66)
);

NAND2xp67_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_26),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_44),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_38),
.B1(n_37),
.B2(n_42),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_76),
.B1(n_84),
.B2(n_91),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_99),
.B1(n_68),
.B2(n_52),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_75),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_42),
.B1(n_35),
.B2(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_81),
.Y(n_114)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_85),
.B(n_52),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_61),
.B(n_1),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_88),
.B(n_90),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_2),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_53),
.A2(n_21),
.B1(n_3),
.B2(n_5),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_65),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_70),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_67),
.A2(n_10),
.B1(n_3),
.B2(n_6),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_45),
.B1(n_69),
.B2(n_91),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_2),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_94),
.B(n_95),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_57),
.B(n_7),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_7),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_8),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_47),
.B(n_8),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_89),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_69),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_115),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_108),
.B(n_78),
.Y(n_126)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_82),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_84),
.A2(n_45),
.B1(n_72),
.B2(n_76),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_117),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_73),
.A2(n_97),
.B1(n_79),
.B2(n_86),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_77),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_114),
.C(n_106),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_93),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_96),
.Y(n_125)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_127),
.C(n_120),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_104),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_80),
.B(n_74),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_128),
.A2(n_131),
.B(n_103),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_129),
.B(n_132),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_82),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_130),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_114),
.B(n_110),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_92),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_135),
.C(n_113),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_81),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_111),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_121),
.B(n_128),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_140),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_102),
.B1(n_116),
.B2(n_115),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_145),
.Y(n_149)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_102),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_146),
.B(n_135),
.Y(n_150)
);

XOR2x1_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_151),
.C(n_142),
.Y(n_162)
);

XOR2x2_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_131),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_137),
.Y(n_153)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

OAI22x1_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_121),
.B1(n_122),
.B2(n_127),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_157),
.B1(n_145),
.B2(n_147),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_152),
.Y(n_158)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_158),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_154),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_151),
.C(n_156),
.Y(n_166)
);

XNOR2x1_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_148),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_141),
.B1(n_122),
.B2(n_145),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_164),
.A2(n_149),
.B(n_152),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_139),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_169),
.C(n_158),
.Y(n_173)
);

AOI31xp33_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_162),
.A3(n_159),
.B(n_160),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_171),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_159),
.B(n_139),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_172),
.B(n_155),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_160),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_176),
.Y(n_177)
);

OAI321xp33_ASAP7_75t_L g178 ( 
.A1(n_175),
.A2(n_173),
.A3(n_143),
.B1(n_100),
.B2(n_112),
.C(n_113),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_179),
.Y(n_180)
);

AOI211xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_177),
.B(n_112),
.C(n_101),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_111),
.Y(n_182)
);


endmodule