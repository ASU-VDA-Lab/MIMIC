module fake_ariane_731_n_27 (n_8, n_3, n_2, n_7, n_5, n_1, n_0, n_6, n_9, n_4, n_27);

input n_8;
input n_3;
input n_2;
input n_7;
input n_5;
input n_1;
input n_0;
input n_6;
input n_9;
input n_4;

output n_27;

wire n_24;
wire n_22;
wire n_13;
wire n_20;
wire n_17;
wire n_18;
wire n_11;
wire n_26;
wire n_14;
wire n_19;
wire n_16;
wire n_12;
wire n_15;
wire n_21;
wire n_23;
wire n_10;
wire n_25;

INVx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

OR2x6_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_L g13 ( 
.A1(n_8),
.A2(n_4),
.B1(n_6),
.B2(n_2),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_10),
.A2(n_0),
.B(n_1),
.Y(n_16)
);

AND3x4_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_3),
.C(n_4),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_15),
.B(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_19),
.B(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_18),
.Y(n_22)
);

NOR4xp25_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_17),
.C(n_16),
.D(n_7),
.Y(n_23)
);

AOI32xp33_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_24)
);

NAND4xp75_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_9),
.C(n_22),
.D(n_23),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_25),
.Y(n_26)
);

OR2x6_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_25),
.Y(n_27)
);


endmodule