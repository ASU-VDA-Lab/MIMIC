module fake_jpeg_5344_n_264 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_264);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_SL g14 ( 
.A(n_10),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_6),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_35),
.B(n_37),
.Y(n_64)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_40),
.Y(n_70)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_21),
.B(n_0),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_17),
.B(n_7),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_44),
.B(n_20),
.Y(n_77)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_17),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_49),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_15),
.B1(n_20),
.B2(n_23),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_50),
.A2(n_56),
.B1(n_75),
.B2(n_87),
.Y(n_96)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_62),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_55),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_15),
.B1(n_20),
.B2(n_23),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_68),
.Y(n_107)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_71),
.Y(n_111)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_74),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_41),
.A2(n_15),
.B1(n_21),
.B2(n_26),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_38),
.B(n_14),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_77),
.Y(n_117)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_88),
.Y(n_118)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_36),
.A2(n_16),
.B1(n_22),
.B2(n_28),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_90),
.B1(n_31),
.B2(n_30),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_41),
.B(n_14),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_8),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

BUFx4f_ASAP7_75t_SL g106 ( 
.A(n_85),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_45),
.A2(n_14),
.B(n_28),
.C(n_26),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_8),
.B(n_13),
.C(n_2),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_45),
.A2(n_21),
.B1(n_16),
.B2(n_24),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_38),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_19),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_102),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_19),
.B1(n_18),
.B2(n_31),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_95),
.B(n_119),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_51),
.A2(n_19),
.B1(n_18),
.B2(n_30),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_99),
.A2(n_113),
.B1(n_82),
.B2(n_73),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_87),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_104),
.B(n_109),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_75),
.A2(n_70),
.B1(n_50),
.B2(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_73),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_51),
.A2(n_30),
.B1(n_1),
.B2(n_0),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_111),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_123),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_64),
.B(n_55),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_SL g172 ( 
.A(n_126),
.B(n_148),
.C(n_3),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_128),
.A2(n_138),
.B1(n_118),
.B2(n_120),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_79),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_129),
.B(n_130),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_101),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_135),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_48),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_140),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_134),
.Y(n_175)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_136),
.A2(n_150),
.B1(n_108),
.B2(n_105),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_57),
.Y(n_137)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_96),
.A2(n_82),
.B1(n_52),
.B2(n_74),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_97),
.B(n_47),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_101),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_143),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_97),
.B(n_0),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_66),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_103),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_59),
.Y(n_146)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_57),
.Y(n_147)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_66),
.B(n_59),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_61),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_149),
.Y(n_160)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_112),
.B(n_1),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_123),
.A2(n_113),
.B1(n_119),
.B2(n_100),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_SL g197 ( 
.A(n_154),
.B(n_161),
.C(n_172),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_155),
.B(n_143),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_116),
.C(n_106),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_163),
.C(n_132),
.Y(n_184)
);

AND2x6_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_124),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_58),
.C(n_118),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_166),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_139),
.A2(n_120),
.B1(n_91),
.B2(n_60),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_58),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_144),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_127),
.A2(n_137),
.B(n_129),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_171),
.A2(n_176),
.B(n_142),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_173),
.B(n_136),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_63),
.B1(n_114),
.B2(n_103),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_174),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_127),
.A2(n_3),
.B(n_4),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_144),
.A2(n_114),
.B1(n_103),
.B2(n_121),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_181),
.A2(n_185),
.B(n_195),
.Y(n_201)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_183),
.B(n_186),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_191),
.C(n_196),
.Y(n_208)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_132),
.Y(n_187)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_141),
.Y(n_188)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_151),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_189),
.A2(n_192),
.B(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_193),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_138),
.C(n_140),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_157),
.B(n_125),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_168),
.B(n_147),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_194),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_149),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_131),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_198),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_172),
.C(n_170),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_204),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_163),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_205),
.Y(n_222)
);

AO21x1_ASAP7_75t_L g217 ( 
.A1(n_203),
.A2(n_210),
.B(n_182),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_179),
.A2(n_157),
.B1(n_173),
.B2(n_168),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_179),
.A2(n_162),
.B(n_173),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_165),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_181),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_164),
.B(n_169),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_159),
.C(n_154),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_213),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_193),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_180),
.A2(n_174),
.B1(n_166),
.B2(n_177),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_216),
.A2(n_187),
.B1(n_189),
.B2(n_183),
.Y(n_221)
);

AOI321xp33_ASAP7_75t_L g239 ( 
.A1(n_217),
.A2(n_225),
.A3(n_209),
.B1(n_211),
.B2(n_208),
.C(n_202),
.Y(n_239)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_221),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_214),
.A2(n_186),
.B1(n_197),
.B2(n_195),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_219),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_216),
.A2(n_190),
.B1(n_159),
.B2(n_176),
.Y(n_223)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_169),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_226),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_212),
.B(n_175),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_227),
.B(n_229),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_175),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_228),
.A2(n_205),
.B(n_201),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_232),
.A2(n_236),
.B(n_225),
.Y(n_242)
);

O2A1O1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_204),
.B(n_203),
.C(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_221),
.B(n_215),
.Y(n_235)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_208),
.B(n_207),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_239),
.A2(n_226),
.B(n_153),
.Y(n_247)
);

OAI21x1_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_225),
.B(n_222),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_240),
.A2(n_242),
.B(n_246),
.Y(n_252)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_247),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_223),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_245),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_222),
.C(n_218),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_243),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_145),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_241),
.A2(n_237),
.B1(n_233),
.B2(n_153),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_253),
.B1(n_245),
.B2(n_150),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_246),
.A2(n_230),
.B1(n_232),
.B2(n_239),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_252),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_135),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_255),
.A2(n_257),
.B(n_4),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_4),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_145),
.Y(n_257)
);

AO21x1_ASAP7_75t_L g261 ( 
.A1(n_258),
.A2(n_260),
.B(n_254),
.Y(n_261)
);

NAND4xp25_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_5),
.C(n_9),
.D(n_11),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_261),
.B(n_262),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_9),
.Y(n_264)
);


endmodule