module fake_netlist_1_12024_n_764 (n_117, n_44, n_133, n_149, n_81, n_69, n_185, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_9, n_161, n_10, n_177, n_130, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_184, n_46, n_31, n_58, n_122, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_182, n_166, n_162, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_764);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_185;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_184;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_764;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_227;
wire n_384;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_489;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_602;
wire n_198;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_698;
wire n_555;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g186 ( .A(n_172), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_99), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_159), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_49), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_181), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_17), .Y(n_191) );
INVxp33_ASAP7_75t_SL g192 ( .A(n_109), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_184), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_126), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_81), .Y(n_195) );
BUFx2_ASAP7_75t_L g196 ( .A(n_85), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_149), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_173), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_94), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_111), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_24), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_12), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_32), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_168), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_133), .Y(n_205) );
BUFx5_ASAP7_75t_L g206 ( .A(n_82), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g207 ( .A(n_167), .Y(n_207) );
CKINVDCx14_ASAP7_75t_R g208 ( .A(n_14), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_74), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_83), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_43), .Y(n_211) );
INVx2_ASAP7_75t_SL g212 ( .A(n_3), .Y(n_212) );
OR2x2_ASAP7_75t_L g213 ( .A(n_8), .B(n_169), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_166), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_132), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_112), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_174), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_182), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_158), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_48), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_155), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_171), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_164), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_122), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_177), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_160), .Y(n_226) );
INVxp33_ASAP7_75t_SL g227 ( .A(n_63), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_92), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_80), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_139), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_84), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_170), .Y(n_232) );
INVx1_ASAP7_75t_SL g233 ( .A(n_121), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_30), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_183), .Y(n_235) );
CKINVDCx16_ASAP7_75t_R g236 ( .A(n_47), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_77), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_137), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_178), .Y(n_239) );
BUFx3_ASAP7_75t_L g240 ( .A(n_68), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_145), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_105), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_97), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_141), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_31), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_116), .Y(n_246) );
INVx2_ASAP7_75t_SL g247 ( .A(n_59), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_1), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_118), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_165), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_67), .Y(n_251) );
BUFx2_ASAP7_75t_L g252 ( .A(n_13), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_143), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_86), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_98), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_71), .Y(n_256) );
INVx2_ASAP7_75t_SL g257 ( .A(n_45), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_106), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_12), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_7), .Y(n_260) );
BUFx3_ASAP7_75t_L g261 ( .A(n_138), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_60), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_66), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_123), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_153), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_135), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_154), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_175), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_101), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_117), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_107), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_52), .Y(n_272) );
INVx1_ASAP7_75t_SL g273 ( .A(n_76), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_56), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_113), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_0), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_120), .Y(n_277) );
CKINVDCx14_ASAP7_75t_R g278 ( .A(n_37), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_157), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_40), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_62), .Y(n_281) );
INVxp67_ASAP7_75t_SL g282 ( .A(n_3), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_57), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_44), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_144), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_198), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_198), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_212), .B(n_0), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_190), .B(n_1), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_253), .Y(n_290) );
INVx1_ASAP7_75t_SL g291 ( .A(n_252), .Y(n_291) );
AND2x6_ASAP7_75t_L g292 ( .A(n_190), .B(n_185), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_210), .Y(n_293) );
BUFx6f_ASAP7_75t_L g294 ( .A(n_198), .Y(n_294) );
INVxp67_ASAP7_75t_L g295 ( .A(n_196), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_199), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_202), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_199), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_208), .A2(n_2), .B1(n_4), .B2(n_5), .Y(n_299) );
OA21x2_ASAP7_75t_L g300 ( .A1(n_187), .A2(n_19), .B(n_18), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_199), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_220), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_247), .B(n_2), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_210), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_257), .B(n_4), .Y(n_305) );
INVxp33_ASAP7_75t_SL g306 ( .A(n_248), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_259), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_207), .B(n_5), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_236), .B(n_6), .Y(n_309) );
INVx5_ASAP7_75t_L g310 ( .A(n_220), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_260), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_289), .B(n_206), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_289), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_293), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_288), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_295), .B(n_278), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_286), .Y(n_317) );
INVx1_ASAP7_75t_SL g318 ( .A(n_291), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_286), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_290), .Y(n_320) );
INVx1_ASAP7_75t_SL g321 ( .A(n_291), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_306), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_307), .A2(n_276), .B1(n_227), .B2(n_192), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_299), .A2(n_203), .B1(n_221), .B2(n_193), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_311), .A2(n_282), .B1(n_213), .B2(n_188), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_297), .B(n_233), .Y(n_326) );
BUFx4f_ASAP7_75t_L g327 ( .A(n_292), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_304), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_297), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_287), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_303), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_327), .B(n_308), .Y(n_332) );
INVxp67_ASAP7_75t_L g333 ( .A(n_318), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_327), .Y(n_334) );
OAI22xp33_ASAP7_75t_L g335 ( .A1(n_321), .A2(n_299), .B1(n_309), .B2(n_272), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_331), .B(n_303), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_315), .A2(n_292), .B1(n_305), .B2(n_195), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_327), .A2(n_300), .B(n_305), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_326), .B(n_292), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_320), .B(n_189), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_312), .A2(n_300), .B(n_197), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_320), .B(n_191), .Y(n_342) );
INVxp67_ASAP7_75t_L g343 ( .A(n_316), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_316), .B(n_194), .Y(n_344) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_313), .B(n_233), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_329), .Y(n_346) );
INVxp67_ASAP7_75t_L g347 ( .A(n_322), .Y(n_347) );
INVx2_ASAP7_75t_SL g348 ( .A(n_322), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_328), .Y(n_349) );
NOR2xp67_ASAP7_75t_L g350 ( .A(n_314), .B(n_310), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_312), .B(n_200), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_314), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_323), .B(n_273), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_325), .A2(n_205), .B(n_204), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_336), .B(n_314), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_333), .B(n_201), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_343), .B(n_324), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_333), .A2(n_281), .B1(n_234), .B2(n_214), .Y(n_358) );
O2A1O1Ixp33_ASAP7_75t_L g359 ( .A1(n_343), .A2(n_211), .B(n_218), .C(n_215), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_346), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_339), .A2(n_223), .B(n_222), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_338), .A2(n_341), .B(n_337), .Y(n_362) );
A2O1A1Ixp33_ASAP7_75t_L g363 ( .A1(n_354), .A2(n_225), .B(n_226), .C(n_224), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_334), .Y(n_364) );
INVx2_ASAP7_75t_SL g365 ( .A(n_345), .Y(n_365) );
A2O1A1Ixp33_ASAP7_75t_L g366 ( .A1(n_353), .A2(n_231), .B(n_232), .C(n_228), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_344), .B(n_209), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_332), .A2(n_238), .B(n_237), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_345), .B(n_216), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_349), .B(n_217), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_340), .A2(n_242), .B(n_241), .Y(n_371) );
BUFx8_ASAP7_75t_L g372 ( .A(n_348), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_334), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_342), .A2(n_244), .B(n_243), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_352), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_335), .A2(n_254), .B1(n_263), .B2(n_256), .C(n_267), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_347), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_351), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_360), .Y(n_379) );
BUFx3_ASAP7_75t_L g380 ( .A(n_372), .Y(n_380) );
OAI21x1_ASAP7_75t_L g381 ( .A1(n_362), .A2(n_249), .B(n_246), .Y(n_381) );
AOI221x1_ASAP7_75t_L g382 ( .A1(n_366), .A2(n_283), .B1(n_250), .B2(n_251), .C(n_270), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_357), .B(n_350), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_361), .A2(n_277), .B(n_275), .Y(n_384) );
INVxp67_ASAP7_75t_L g385 ( .A(n_372), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_375), .Y(n_386) );
A2O1A1Ixp33_ASAP7_75t_L g387 ( .A1(n_378), .A2(n_371), .B(n_374), .C(n_359), .Y(n_387) );
NAND3xp33_ASAP7_75t_L g388 ( .A(n_376), .B(n_294), .C(n_287), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_358), .B(n_219), .Y(n_389) );
A2O1A1Ixp33_ASAP7_75t_L g390 ( .A1(n_363), .A2(n_284), .B(n_186), .C(n_258), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_355), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_377), .B(n_229), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_365), .B(n_230), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_367), .B(n_369), .Y(n_394) );
AOI21x1_ASAP7_75t_L g395 ( .A1(n_368), .A2(n_268), .B(n_264), .Y(n_395) );
CKINVDCx6p67_ASAP7_75t_R g396 ( .A(n_356), .Y(n_396) );
AOI221xp5_ASAP7_75t_SL g397 ( .A1(n_370), .A2(n_285), .B1(n_280), .B2(n_279), .C(n_220), .Y(n_397) );
A2O1A1Ixp33_ASAP7_75t_L g398 ( .A1(n_373), .A2(n_261), .B(n_240), .C(n_280), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_364), .A2(n_274), .B1(n_235), .B2(n_239), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_364), .A2(n_280), .B1(n_279), .B2(n_255), .Y(n_400) );
OAI21x1_ASAP7_75t_L g401 ( .A1(n_362), .A2(n_330), .B(n_206), .Y(n_401) );
OAI21xp5_ASAP7_75t_L g402 ( .A1(n_362), .A2(n_262), .B(n_245), .Y(n_402) );
OAI22xp33_ASAP7_75t_L g403 ( .A1(n_358), .A2(n_265), .B1(n_266), .B2(n_269), .Y(n_403) );
AO31x2_ASAP7_75t_L g404 ( .A1(n_362), .A2(n_206), .A3(n_298), .B(n_294), .Y(n_404) );
BUFx8_ASAP7_75t_L g405 ( .A(n_380), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_379), .Y(n_406) );
A2O1A1Ixp33_ASAP7_75t_L g407 ( .A1(n_387), .A2(n_279), .B(n_271), .C(n_310), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_391), .B(n_7), .Y(n_408) );
AO21x2_ASAP7_75t_L g409 ( .A1(n_381), .A2(n_296), .B(n_294), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_386), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_383), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_394), .B(n_9), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_389), .B(n_9), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_404), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_404), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_403), .B(n_10), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_395), .Y(n_417) );
BUFx12f_ASAP7_75t_L g418 ( .A(n_385), .Y(n_418) );
AO21x1_ASAP7_75t_L g419 ( .A1(n_402), .A2(n_10), .B(n_11), .Y(n_419) );
OA21x2_ASAP7_75t_L g420 ( .A1(n_397), .A2(n_302), .B(n_301), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_404), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_388), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_396), .Y(n_423) );
OA21x2_ASAP7_75t_L g424 ( .A1(n_397), .A2(n_302), .B(n_301), .Y(n_424) );
AO31x2_ASAP7_75t_L g425 ( .A1(n_382), .A2(n_301), .A3(n_302), .B(n_310), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_390), .B(n_11), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_393), .Y(n_427) );
AO22x2_ASAP7_75t_L g428 ( .A1(n_388), .A2(n_400), .B1(n_384), .B2(n_398), .Y(n_428) );
OAI21x1_ASAP7_75t_L g429 ( .A1(n_400), .A2(n_104), .B(n_180), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_392), .B(n_15), .Y(n_430) );
OAI21x1_ASAP7_75t_L g431 ( .A1(n_399), .A2(n_103), .B(n_179), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_394), .B(n_15), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_379), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_391), .A2(n_16), .B1(n_319), .B2(n_317), .Y(n_434) );
OAI21x1_ASAP7_75t_L g435 ( .A1(n_401), .A2(n_108), .B(n_20), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_389), .A2(n_319), .B1(n_317), .B2(n_16), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_391), .B(n_21), .Y(n_437) );
OAI21x1_ASAP7_75t_SL g438 ( .A1(n_402), .A2(n_22), .B(n_23), .Y(n_438) );
OAI21x1_ASAP7_75t_L g439 ( .A1(n_401), .A2(n_25), .B(n_26), .Y(n_439) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_380), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_380), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_391), .B(n_27), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_387), .A2(n_319), .B(n_28), .Y(n_443) );
OAI21x1_ASAP7_75t_L g444 ( .A1(n_401), .A2(n_29), .B(n_33), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_379), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_387), .A2(n_34), .B(n_35), .Y(n_446) );
OA21x2_ASAP7_75t_L g447 ( .A1(n_397), .A2(n_36), .B(n_38), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_391), .B(n_39), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_414), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_410), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_433), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_442), .B(n_41), .Y(n_452) );
OR2x6_ASAP7_75t_L g453 ( .A(n_442), .B(n_42), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_415), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_406), .B(n_46), .Y(n_455) );
OA21x2_ASAP7_75t_L g456 ( .A1(n_421), .A2(n_50), .B(n_51), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_411), .A2(n_53), .B1(n_54), .B2(n_55), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_445), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_445), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_421), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_427), .B(n_58), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_432), .B(n_61), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_408), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_412), .A2(n_64), .B(n_65), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_425), .Y(n_465) );
INVx3_ASAP7_75t_L g466 ( .A(n_440), .Y(n_466) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_417), .A2(n_69), .B(n_70), .Y(n_467) );
BUFx2_ASAP7_75t_L g468 ( .A(n_441), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_416), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_419), .B(n_72), .Y(n_470) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_407), .A2(n_73), .B(n_75), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_425), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_426), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_409), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_435), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_430), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_439), .Y(n_477) );
INVx2_ASAP7_75t_SL g478 ( .A(n_405), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_413), .Y(n_479) );
BUFx2_ASAP7_75t_L g480 ( .A(n_440), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_437), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_405), .Y(n_482) );
OR2x6_ASAP7_75t_L g483 ( .A(n_440), .B(n_78), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_444), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_448), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_420), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_420), .Y(n_487) );
AOI21x1_ASAP7_75t_L g488 ( .A1(n_424), .A2(n_447), .B(n_443), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_425), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_423), .B(n_79), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_424), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_436), .B(n_176), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_418), .B(n_87), .Y(n_493) );
INVx3_ASAP7_75t_L g494 ( .A(n_429), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_434), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_438), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_422), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_431), .B(n_88), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_428), .Y(n_499) );
OR2x6_ASAP7_75t_L g500 ( .A(n_446), .B(n_89), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_428), .Y(n_501) );
BUFx3_ASAP7_75t_L g502 ( .A(n_405), .Y(n_502) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_421), .A2(n_90), .B(n_91), .Y(n_503) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_440), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_410), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_410), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_410), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_414), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_410), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_410), .Y(n_510) );
AOI21xp5_ASAP7_75t_SL g511 ( .A1(n_442), .A2(n_93), .B(n_95), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_410), .Y(n_512) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_421), .A2(n_96), .B(n_100), .Y(n_513) );
NAND2x1p5_ASAP7_75t_L g514 ( .A(n_442), .B(n_102), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_414), .Y(n_515) );
BUFx3_ASAP7_75t_L g516 ( .A(n_405), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_406), .B(n_110), .Y(n_517) );
BUFx2_ASAP7_75t_L g518 ( .A(n_504), .Y(n_518) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_449), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_449), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_454), .Y(n_521) );
BUFx2_ASAP7_75t_L g522 ( .A(n_504), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_450), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_451), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_480), .B(n_114), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_505), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_506), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_507), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_454), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_468), .B(n_115), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_509), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_510), .Y(n_532) );
INVxp67_ASAP7_75t_SL g533 ( .A(n_508), .Y(n_533) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_514), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_512), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_508), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_515), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_458), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_466), .B(n_119), .Y(n_539) );
INVx2_ASAP7_75t_SL g540 ( .A(n_482), .Y(n_540) );
INVxp67_ASAP7_75t_SL g541 ( .A(n_515), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_460), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_476), .B(n_124), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_453), .B(n_125), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_460), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_459), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_517), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_517), .Y(n_548) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_514), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_479), .B(n_127), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_499), .B(n_128), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_463), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_486), .Y(n_553) );
BUFx2_ASAP7_75t_L g554 ( .A(n_453), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_493), .B(n_129), .Y(n_555) );
INVx3_ASAP7_75t_L g556 ( .A(n_453), .Y(n_556) );
OR2x6_ASAP7_75t_L g557 ( .A(n_483), .B(n_130), .Y(n_557) );
AO22x1_ASAP7_75t_L g558 ( .A1(n_482), .A2(n_131), .B1(n_134), .B2(n_136), .Y(n_558) );
BUFx2_ASAP7_75t_L g559 ( .A(n_483), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_501), .B(n_140), .Y(n_560) );
INVx4_ASAP7_75t_L g561 ( .A(n_502), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_452), .B(n_142), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_455), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_461), .B(n_146), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_497), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_461), .B(n_147), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_469), .B(n_148), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_486), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_452), .B(n_150), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_483), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_497), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_490), .B(n_151), .Y(n_572) );
INVx5_ASAP7_75t_L g573 ( .A(n_502), .Y(n_573) );
BUFx2_ASAP7_75t_L g574 ( .A(n_516), .Y(n_574) );
NAND2xp33_ASAP7_75t_SL g575 ( .A(n_462), .B(n_152), .Y(n_575) );
INVx4_ASAP7_75t_L g576 ( .A(n_516), .Y(n_576) );
BUFx3_ASAP7_75t_L g577 ( .A(n_478), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_473), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_495), .Y(n_579) );
BUFx2_ASAP7_75t_L g580 ( .A(n_498), .Y(n_580) );
AND2x4_ASAP7_75t_L g581 ( .A(n_496), .B(n_156), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_481), .Y(n_582) );
CKINVDCx8_ASAP7_75t_R g583 ( .A(n_498), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_487), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_487), .Y(n_585) );
BUFx2_ASAP7_75t_L g586 ( .A(n_464), .Y(n_586) );
INVx2_ASAP7_75t_SL g587 ( .A(n_492), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_485), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_491), .Y(n_589) );
BUFx2_ASAP7_75t_L g590 ( .A(n_464), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_465), .Y(n_591) );
AND2x4_ASAP7_75t_SL g592 ( .A(n_561), .B(n_457), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_542), .Y(n_593) );
INVxp67_ASAP7_75t_L g594 ( .A(n_574), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_552), .B(n_465), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_523), .B(n_472), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_542), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_524), .B(n_472), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_582), .B(n_513), .Y(n_599) );
AND2x2_ASAP7_75t_SL g600 ( .A(n_554), .B(n_456), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_526), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_588), .B(n_470), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_527), .B(n_470), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_561), .B(n_511), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_580), .B(n_489), .Y(n_605) );
AND2x4_ASAP7_75t_L g606 ( .A(n_556), .B(n_494), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_528), .B(n_474), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_531), .B(n_503), .Y(n_608) );
AND3x2_ASAP7_75t_L g609 ( .A(n_559), .B(n_491), .C(n_475), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_532), .B(n_513), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_520), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_535), .B(n_474), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_538), .B(n_494), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_546), .Y(n_614) );
BUFx3_ASAP7_75t_L g615 ( .A(n_576), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_578), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_545), .Y(n_617) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_521), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_521), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_583), .B(n_456), .Y(n_620) );
AND2x4_ASAP7_75t_L g621 ( .A(n_556), .B(n_477), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_563), .B(n_484), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_529), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_587), .B(n_484), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_565), .Y(n_625) );
INVx2_ASAP7_75t_SL g626 ( .A(n_576), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_579), .B(n_457), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_536), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_571), .B(n_475), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_537), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_545), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_530), .B(n_467), .Y(n_632) );
INVxp67_ASAP7_75t_L g633 ( .A(n_577), .Y(n_633) );
NOR3xp33_ASAP7_75t_L g634 ( .A(n_540), .B(n_488), .C(n_500), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_547), .B(n_471), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_548), .B(n_471), .Y(n_636) );
AND2x4_ASAP7_75t_L g637 ( .A(n_570), .B(n_500), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_518), .B(n_500), .Y(n_638) );
BUFx2_ASAP7_75t_L g639 ( .A(n_573), .Y(n_639) );
AND2x4_ASAP7_75t_L g640 ( .A(n_570), .B(n_161), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_519), .Y(n_641) );
AND2x4_ASAP7_75t_L g642 ( .A(n_573), .B(n_162), .Y(n_642) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_522), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_551), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_551), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_560), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_519), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_573), .B(n_163), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_577), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_625), .B(n_590), .Y(n_650) );
BUFx2_ASAP7_75t_SL g651 ( .A(n_615), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_643), .B(n_533), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_601), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_594), .B(n_533), .Y(n_654) );
NAND2x1_ASAP7_75t_L g655 ( .A(n_626), .B(n_557), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_613), .B(n_541), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_622), .B(n_541), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_616), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_599), .B(n_591), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_614), .B(n_586), .Y(n_660) );
BUFx2_ASAP7_75t_L g661 ( .A(n_639), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_606), .B(n_591), .Y(n_662) );
OR2x2_ASAP7_75t_L g663 ( .A(n_618), .B(n_568), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_598), .Y(n_664) );
INVx2_ASAP7_75t_SL g665 ( .A(n_611), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_595), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_607), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_644), .B(n_560), .Y(n_668) );
NAND2x1p5_ASAP7_75t_L g669 ( .A(n_642), .B(n_544), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_593), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_612), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_596), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_597), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_608), .B(n_553), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_610), .B(n_553), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_645), .B(n_568), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_624), .B(n_584), .Y(n_677) );
OR2x2_ASAP7_75t_L g678 ( .A(n_619), .B(n_623), .Y(n_678) );
BUFx2_ASAP7_75t_L g679 ( .A(n_633), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_649), .B(n_544), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_597), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_617), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_628), .B(n_589), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_629), .B(n_589), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_646), .B(n_585), .Y(n_685) );
AND2x4_ASAP7_75t_L g686 ( .A(n_606), .B(n_585), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_637), .A2(n_575), .B1(n_562), .B2(n_557), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_638), .B(n_581), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_631), .B(n_584), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_630), .B(n_581), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_653), .Y(n_691) );
OAI22xp33_ASAP7_75t_L g692 ( .A1(n_655), .A2(n_557), .B1(n_534), .B2(n_549), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_658), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_657), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_688), .B(n_637), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_661), .B(n_605), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_657), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_664), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_667), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_671), .Y(n_700) );
OR2x2_ASAP7_75t_L g701 ( .A(n_672), .B(n_641), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_666), .B(n_631), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_679), .B(n_605), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_676), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_652), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_685), .Y(n_706) );
OAI21xp33_ASAP7_75t_L g707 ( .A1(n_687), .A2(n_592), .B(n_620), .Y(n_707) );
NAND2x1p5_ASAP7_75t_L g708 ( .A(n_669), .B(n_642), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_660), .Y(n_709) );
INVxp67_ASAP7_75t_SL g710 ( .A(n_669), .Y(n_710) );
OR2x2_ASAP7_75t_L g711 ( .A(n_678), .B(n_641), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_650), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_681), .Y(n_713) );
INVx1_ASAP7_75t_SL g714 ( .A(n_651), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_665), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_702), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_702), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_691), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_693), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_704), .Y(n_720) );
O2A1O1Ixp33_ASAP7_75t_L g721 ( .A1(n_714), .A2(n_668), .B(n_604), .C(n_634), .Y(n_721) );
NAND3xp33_ASAP7_75t_L g722 ( .A(n_707), .B(n_687), .C(n_654), .Y(n_722) );
INVx2_ASAP7_75t_SL g723 ( .A(n_714), .Y(n_723) );
OAI21xp33_ASAP7_75t_L g724 ( .A1(n_707), .A2(n_665), .B(n_659), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_706), .Y(n_725) );
INVx1_ASAP7_75t_SL g726 ( .A(n_696), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_701), .Y(n_727) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_709), .A2(n_680), .B1(n_659), .B2(n_677), .C(n_656), .Y(n_728) );
OAI22xp33_ASAP7_75t_L g729 ( .A1(n_710), .A2(n_549), .B1(n_534), .B2(n_690), .Y(n_729) );
OAI21xp5_ASAP7_75t_L g730 ( .A1(n_710), .A2(n_562), .B(n_600), .Y(n_730) );
AOI211xp5_ASAP7_75t_L g731 ( .A1(n_724), .A2(n_692), .B(n_712), .C(n_703), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_723), .B(n_698), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_722), .A2(n_699), .B1(n_700), .B2(n_715), .Y(n_733) );
AOI221xp5_ASAP7_75t_L g734 ( .A1(n_728), .A2(n_713), .B1(n_697), .B2(n_694), .C(n_705), .Y(n_734) );
AOI31xp33_ASAP7_75t_L g735 ( .A1(n_730), .A2(n_708), .A3(n_575), .B(n_569), .Y(n_735) );
AOI31xp33_ASAP7_75t_SL g736 ( .A1(n_721), .A2(n_711), .A3(n_708), .B(n_648), .Y(n_736) );
AOI321xp33_ASAP7_75t_L g737 ( .A1(n_720), .A2(n_656), .A3(n_695), .B1(n_662), .B2(n_677), .C(n_686), .Y(n_737) );
AOI221xp5_ASAP7_75t_SL g738 ( .A1(n_726), .A2(n_555), .B1(n_674), .B2(n_675), .C(n_684), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_716), .Y(n_739) );
O2A1O1Ixp33_ASAP7_75t_L g740 ( .A1(n_725), .A2(n_627), .B(n_602), .C(n_603), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g741 ( .A1(n_726), .A2(n_640), .B(n_572), .Y(n_741) );
NOR3xp33_ASAP7_75t_L g742 ( .A(n_729), .B(n_558), .C(n_640), .Y(n_742) );
A2O1A1Ixp33_ASAP7_75t_L g743 ( .A1(n_727), .A2(n_662), .B(n_686), .C(n_684), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g744 ( .A1(n_717), .A2(n_674), .B1(n_675), .B2(n_662), .C(n_686), .Y(n_744) );
NOR3xp33_ASAP7_75t_SL g745 ( .A(n_718), .B(n_636), .C(n_635), .Y(n_745) );
AOI322xp5_ASAP7_75t_L g746 ( .A1(n_719), .A2(n_632), .A3(n_647), .B1(n_689), .B2(n_673), .C1(n_670), .C2(n_682), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g747 ( .A(n_738), .B(n_737), .Y(n_747) );
A2O1A1Ixp33_ASAP7_75t_L g748 ( .A1(n_735), .A2(n_731), .B(n_733), .C(n_734), .Y(n_748) );
AOI211xp5_ASAP7_75t_SL g749 ( .A1(n_742), .A2(n_732), .B(n_743), .C(n_744), .Y(n_749) );
O2A1O1Ixp33_ASAP7_75t_L g750 ( .A1(n_736), .A2(n_740), .B(n_739), .C(n_741), .Y(n_750) );
OR2x2_ASAP7_75t_L g751 ( .A(n_747), .B(n_663), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_749), .B(n_746), .Y(n_752) );
NAND4xp75_ASAP7_75t_L g753 ( .A(n_748), .B(n_745), .C(n_564), .D(n_566), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_751), .B(n_750), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_752), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_753), .B(n_670), .Y(n_756) );
BUFx6f_ASAP7_75t_L g757 ( .A(n_755), .Y(n_757) );
INVx5_ASAP7_75t_L g758 ( .A(n_754), .Y(n_758) );
AO22x2_ASAP7_75t_SL g759 ( .A1(n_758), .A2(n_756), .B1(n_550), .B2(n_543), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_759), .A2(n_758), .B1(n_757), .B2(n_534), .Y(n_760) );
OA22x2_ASAP7_75t_L g761 ( .A1(n_760), .A2(n_609), .B1(n_525), .B2(n_567), .Y(n_761) );
OR2x2_ASAP7_75t_L g762 ( .A(n_761), .B(n_683), .Y(n_762) );
OR2x6_ASAP7_75t_L g763 ( .A(n_762), .B(n_539), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_763), .A2(n_621), .B1(n_549), .B2(n_534), .Y(n_764) );
endmodule