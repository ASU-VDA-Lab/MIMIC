module fake_jpeg_1105_n_204 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_204);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_SL g53 ( 
.A(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_4),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_14),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_31),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_3),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_78),
.B(n_73),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_72),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_47),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_63),
.Y(n_85)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_90),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_70),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_76),
.B1(n_79),
.B2(n_82),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_94),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_53),
.B1(n_50),
.B2(n_56),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_54),
.B1(n_59),
.B2(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_64),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_101),
.Y(n_120)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_99),
.Y(n_133)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_64),
.B(n_68),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_62),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_110),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_69),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_69),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_111),
.B(n_113),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_112),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_49),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_83),
.Y(n_114)
);

OAI32xp33_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_65),
.A3(n_66),
.B1(n_52),
.B2(n_60),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_1),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_52),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_117),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_60),
.Y(n_117)
);

NOR2xp67_ASAP7_75t_SL g118 ( 
.A(n_106),
.B(n_51),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_9),
.B(n_10),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_112),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_129),
.Y(n_143)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_102),
.A2(n_65),
.B1(n_48),
.B2(n_61),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_128),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_108),
.B(n_0),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_107),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_131),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_61),
.B1(n_65),
.B2(n_55),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_134),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_0),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_137),
.Y(n_161)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_145),
.B1(n_154),
.B2(n_155),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_5),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_141),
.Y(n_163)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_25),
.B(n_43),
.Y(n_144)
);

OA21x2_ASAP7_75t_SL g157 ( 
.A1(n_144),
.A2(n_148),
.B(n_149),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_SL g146 ( 
.A1(n_122),
.A2(n_27),
.B(n_42),
.C(n_39),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_146),
.A2(n_147),
.B(n_152),
.Y(n_166)
);

NAND2x1_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_23),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_7),
.B(n_9),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_10),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_35),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_115),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_162),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_133),
.B(n_121),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_160),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_135),
.A2(n_121),
.B(n_18),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_139),
.A2(n_15),
.B1(n_19),
.B2(n_20),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_143),
.A2(n_24),
.B(n_30),
.Y(n_164)
);

NOR2x1_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_166),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_165),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_147),
.A2(n_46),
.B(n_32),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_38),
.Y(n_169)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_153),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_171),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_179),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_183),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_178),
.Y(n_183)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_163),
.C(n_166),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_186),
.C(n_187),
.Y(n_190)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_161),
.C(n_164),
.Y(n_186)
);

BUFx12_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_159),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_182),
.A2(n_172),
.B1(n_170),
.B2(n_167),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_193),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_160),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_157),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_193),
.A2(n_188),
.B1(n_180),
.B2(n_177),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_197),
.Y(n_199)
);

OR2x6_ASAP7_75t_SL g198 ( 
.A(n_195),
.B(n_190),
.Y(n_198)
);

AOI321xp33_ASAP7_75t_SL g200 ( 
.A1(n_198),
.A2(n_196),
.A3(n_188),
.B1(n_189),
.B2(n_177),
.C(n_168),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_199),
.B(n_192),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_203),
.Y(n_204)
);


endmodule