module fake_netlist_6_2187_n_71 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_7, n_2, n_5, n_71);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_7;
input n_2;
input n_5;

output n_71;

wire n_41;
wire n_52;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_70;
wire n_24;
wire n_21;
wire n_37;
wire n_33;
wire n_54;
wire n_67;
wire n_27;
wire n_38;
wire n_61;
wire n_39;
wire n_63;
wire n_60;
wire n_59;
wire n_32;
wire n_66;
wire n_36;
wire n_22;
wire n_26;
wire n_68;
wire n_55;
wire n_35;
wire n_28;
wire n_23;
wire n_58;
wire n_69;
wire n_20;
wire n_50;
wire n_49;
wire n_30;
wire n_64;
wire n_43;
wire n_19;
wire n_47;
wire n_48;
wire n_29;
wire n_62;
wire n_31;
wire n_65;
wire n_25;
wire n_40;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

AND2x6_ASAP7_75t_L g27 ( 
.A(n_2),
.B(n_1),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

OAI21x1_ASAP7_75t_L g29 ( 
.A1(n_12),
.A2(n_11),
.B(n_5),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_7),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

NOR2x2_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_3),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_5),
.Y(n_38)
);

AO31x2_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_28),
.A3(n_30),
.B(n_32),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_29),
.B(n_31),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_25),
.B(n_32),
.C(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_28),
.Y(n_42)
);

AO31x2_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_23),
.A3(n_26),
.B(n_22),
.Y(n_43)
);

AO31x2_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_23),
.A3(n_26),
.B(n_22),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

OR2x6_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_34),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_20),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_39),
.Y(n_53)
);

AND2x4_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_44),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_44),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_49),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_53),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_47),
.B1(n_56),
.B2(n_55),
.Y(n_61)
);

OAI31xp33_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_55),
.A3(n_41),
.B(n_54),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_56),
.B(n_47),
.Y(n_63)
);

AOI221xp5_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_24),
.B1(n_46),
.B2(n_21),
.C(n_45),
.Y(n_64)
);

OAI211xp5_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_24),
.B(n_45),
.C(n_56),
.Y(n_65)
);

NOR2xp67_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_61),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_24),
.B(n_27),
.C(n_10),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

OAI22x1_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_67),
.B1(n_27),
.B2(n_16),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_27),
.Y(n_70)
);

AO21x2_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_40),
.B(n_66),
.Y(n_71)
);


endmodule