module fake_jpeg_13501_n_610 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_610);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_610;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_12),
.B(n_13),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_59),
.B(n_89),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_10),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_63),
.B(n_69),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_65),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_20),
.B(n_10),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_71),
.Y(n_155)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_73),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_74),
.Y(n_194)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_75),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_76),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_77),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_78),
.Y(n_213)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_10),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_80),
.B(n_83),
.Y(n_145)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_81),
.Y(n_176)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_82),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_40),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_84),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_85),
.Y(n_205)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_86),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_88),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_24),
.B(n_18),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_24),
.B(n_10),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_90),
.B(n_92),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_27),
.B(n_11),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

INVx6_ASAP7_75t_SL g94 ( 
.A(n_30),
.Y(n_94)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_94),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_21),
.B(n_8),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_19),
.C(n_48),
.Y(n_136)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

BUFx4f_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_27),
.B(n_12),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_100),
.B(n_101),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_22),
.B(n_7),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_102),
.Y(n_178)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_22),
.Y(n_104)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_105),
.Y(n_217)
);

CKINVDCx9p33_ASAP7_75t_R g106 ( 
.A(n_30),
.Y(n_106)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

INVx6_ASAP7_75t_SL g107 ( 
.A(n_55),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g216 ( 
.A(n_107),
.Y(n_216)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_109),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_18),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_110),
.B(n_17),
.Y(n_160)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_22),
.Y(n_112)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_112),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_113),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_114),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_115),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_116),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_55),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_118),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_119),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_120),
.Y(n_208)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_121),
.Y(n_204)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_122),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_123),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_28),
.Y(n_124)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_124),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_28),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_49),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_41),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_47),
.Y(n_128)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_128),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_63),
.A2(n_42),
.B1(n_52),
.B2(n_25),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_130),
.A2(n_143),
.B1(n_150),
.B2(n_159),
.Y(n_230)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_95),
.B(n_45),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_133),
.B(n_136),
.Y(n_270)
);

AO22x1_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_40),
.B1(n_51),
.B2(n_45),
.Y(n_139)
);

AO22x1_ASAP7_75t_L g260 ( 
.A1(n_139),
.A2(n_142),
.B1(n_151),
.B2(n_181),
.Y(n_260)
);

AO22x1_ASAP7_75t_SL g142 ( 
.A1(n_80),
.A2(n_51),
.B1(n_45),
.B2(n_40),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_69),
.A2(n_42),
.B1(n_25),
.B2(n_40),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_90),
.A2(n_51),
.B1(n_45),
.B2(n_19),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_92),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_157),
.B(n_186),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_100),
.A2(n_51),
.B1(n_58),
.B2(n_56),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_160),
.B(n_193),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_124),
.A2(n_128),
.B1(n_126),
.B2(n_125),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_161),
.A2(n_163),
.B1(n_207),
.B2(n_218),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_64),
.A2(n_67),
.B1(n_119),
.B2(n_117),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_66),
.A2(n_123),
.B1(n_115),
.B2(n_113),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_166),
.A2(n_183),
.B1(n_209),
.B2(n_0),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_82),
.A2(n_57),
.B1(n_49),
.B2(n_56),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_169),
.A2(n_171),
.B(n_175),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_62),
.A2(n_57),
.B1(n_58),
.B2(n_29),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_72),
.A2(n_57),
.B1(n_48),
.B2(n_41),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_177),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_71),
.A2(n_57),
.B1(n_41),
.B2(n_34),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_97),
.Y(n_185)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_85),
.B(n_61),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_76),
.B(n_7),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_73),
.Y(n_196)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_75),
.B(n_7),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_199),
.B(n_203),
.Y(n_257)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_74),
.Y(n_202)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_77),
.B(n_6),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_78),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_84),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_91),
.B(n_6),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_167),
.Y(n_242)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_219),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_133),
.B(n_0),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_220),
.B(n_226),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_129),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_221),
.B(n_228),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_137),
.B(n_105),
.C(n_93),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_223),
.B(n_281),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_224),
.A2(n_239),
.B1(n_241),
.B2(n_272),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_161),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g320 ( 
.A1(n_225),
.A2(n_233),
.B1(n_236),
.B2(n_246),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_153),
.B(n_0),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_129),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_152),
.Y(n_231)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_231),
.Y(n_328)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_146),
.Y(n_232)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_232),
.Y(n_341)
);

OA22x2_ASAP7_75t_L g233 ( 
.A1(n_166),
.A2(n_0),
.B1(n_13),
.B2(n_15),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_149),
.Y(n_234)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_234),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_187),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_235),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_163),
.A2(n_13),
.B1(n_15),
.B2(n_184),
.Y(n_236)
);

BUFx16f_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_237),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_238),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_173),
.A2(n_209),
.B1(n_134),
.B2(n_139),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_180),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_240),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_164),
.A2(n_145),
.B1(n_175),
.B2(n_142),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_242),
.B(n_280),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_135),
.B(n_172),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_243),
.B(n_262),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_162),
.Y(n_244)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_244),
.Y(n_310)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_156),
.Y(n_245)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_245),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_168),
.A2(n_190),
.B1(n_204),
.B2(n_206),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_176),
.Y(n_247)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_247),
.Y(n_316)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_248),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_138),
.A2(n_141),
.B1(n_165),
.B2(n_131),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_249),
.A2(n_278),
.B1(n_289),
.B2(n_191),
.Y(n_297)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_174),
.Y(n_250)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_250),
.Y(n_324)
);

BUFx12_ASAP7_75t_L g251 ( 
.A(n_192),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_251),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_216),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_253),
.B(n_263),
.Y(n_318)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_162),
.Y(n_254)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_254),
.Y(n_300)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_188),
.Y(n_255)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_255),
.Y(n_329)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_197),
.Y(n_258)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_258),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_205),
.Y(n_259)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_259),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_260),
.A2(n_194),
.B(n_198),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_205),
.Y(n_261)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_261),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_147),
.B(n_208),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_216),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_151),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_264),
.Y(n_332)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_178),
.Y(n_265)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_265),
.Y(n_338)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_197),
.Y(n_266)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_266),
.Y(n_322)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_210),
.Y(n_267)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_267),
.Y(n_344)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_154),
.Y(n_268)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_268),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_165),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_271),
.B(n_273),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_171),
.A2(n_195),
.B1(n_169),
.B2(n_189),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_212),
.Y(n_273)
);

INVx3_ASAP7_75t_SL g274 ( 
.A(n_195),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_274),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_189),
.A2(n_132),
.B1(n_213),
.B2(n_140),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_275),
.A2(n_213),
.B1(n_194),
.B2(n_198),
.Y(n_303)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_158),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_281),
.Y(n_302)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_158),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_277),
.B(n_293),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_132),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_179),
.B(n_214),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_279),
.B(n_264),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_148),
.B(n_182),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_148),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_283),
.B(n_284),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_182),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_138),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_285),
.B(n_286),
.Y(n_330)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_170),
.Y(n_286)
);

BUFx2_ASAP7_75t_SL g287 ( 
.A(n_201),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_287),
.B(n_288),
.Y(n_339)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_170),
.Y(n_288)
);

INVx11_ASAP7_75t_L g289 ( 
.A(n_217),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_217),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_290),
.B(n_291),
.Y(n_352)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_218),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_140),
.B(n_144),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_233),
.Y(n_311)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_144),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_155),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_294),
.B(n_278),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_239),
.A2(n_155),
.B(n_191),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_296),
.A2(n_309),
.B(n_350),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_297),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_299),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_303),
.A2(n_294),
.B1(n_258),
.B2(n_266),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_304),
.B(n_311),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_269),
.A2(n_270),
.B(n_280),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_230),
.A2(n_269),
.B1(n_260),
.B2(n_257),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_312),
.A2(n_237),
.B1(n_304),
.B2(n_296),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_251),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_313),
.B(n_317),
.Y(n_366)
);

FAx1_ASAP7_75t_SL g317 ( 
.A(n_220),
.B(n_226),
.CI(n_270),
.CON(n_317),
.SN(n_317)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_252),
.A2(n_244),
.B1(n_274),
.B2(n_219),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_323),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_256),
.B(n_270),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_326),
.B(n_345),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_251),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_331),
.B(n_335),
.Y(n_368)
);

AOI21xp33_ASAP7_75t_L g335 ( 
.A1(n_264),
.A2(n_282),
.B(n_292),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_343),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_223),
.B(n_230),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_346),
.B(n_307),
.Y(n_389)
);

AOI22x1_ASAP7_75t_L g348 ( 
.A1(n_233),
.A2(n_238),
.B1(n_264),
.B2(n_267),
.Y(n_348)
);

AO22x1_ASAP7_75t_SL g367 ( 
.A1(n_348),
.A2(n_283),
.B1(n_284),
.B2(n_289),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_222),
.A2(n_227),
.B(n_229),
.Y(n_350)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_305),
.Y(n_353)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_353),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_318),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_354),
.B(n_363),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_355),
.A2(n_357),
.B1(n_358),
.B2(n_374),
.Y(n_418)
);

OAI21xp33_ASAP7_75t_SL g356 ( 
.A1(n_309),
.A2(n_233),
.B(n_285),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_356),
.A2(n_339),
.B(n_352),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_301),
.A2(n_254),
.B1(n_265),
.B2(n_276),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_301),
.A2(n_234),
.B1(n_245),
.B2(n_247),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_326),
.B(n_232),
.C(n_290),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_359),
.B(n_352),
.C(n_330),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_302),
.A2(n_288),
.B1(n_286),
.B2(n_291),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_361),
.A2(n_383),
.B1(n_386),
.B2(n_393),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_342),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_325),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_364),
.Y(n_414)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_321),
.Y(n_365)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_365),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_367),
.B(n_369),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_306),
.B(n_268),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_321),
.Y(n_370)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_370),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_336),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_371),
.B(n_385),
.Y(n_411)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_338),
.Y(n_373)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_373),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_345),
.A2(n_259),
.B1(n_261),
.B2(n_237),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_322),
.Y(n_375)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_375),
.Y(n_428)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_338),
.Y(n_376)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_376),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_347),
.Y(n_377)
);

INVx5_ASAP7_75t_L g407 ( 
.A(n_377),
.Y(n_407)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_381),
.Y(n_431)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_344),
.Y(n_382)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_382),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_306),
.B(n_312),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_302),
.A2(n_311),
.B1(n_299),
.B2(n_348),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_327),
.B(n_315),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_387),
.B(n_389),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_317),
.B(n_302),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_394),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_348),
.A2(n_320),
.B1(n_303),
.B2(n_319),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g409 ( 
.A1(n_390),
.A2(n_396),
.B1(n_320),
.B2(n_330),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_319),
.A2(n_307),
.B(n_325),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_391),
.A2(n_330),
.B(n_339),
.Y(n_406)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_324),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_392),
.B(n_395),
.Y(n_398)
);

OAI22x1_ASAP7_75t_SL g393 ( 
.A1(n_320),
.A2(n_317),
.B1(n_308),
.B2(n_333),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_350),
.B(n_349),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_324),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_320),
.A2(n_349),
.B1(n_328),
.B2(n_351),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_329),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_397),
.B(n_341),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_399),
.B(n_402),
.C(n_425),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_362),
.B(n_298),
.C(n_329),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_372),
.B(n_325),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_404),
.B(n_367),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_406),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_409),
.A2(n_390),
.B1(n_366),
.B2(n_367),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_386),
.A2(n_332),
.B1(n_337),
.B2(n_322),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_410),
.A2(n_419),
.B1(n_355),
.B2(n_396),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_413),
.B(n_422),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_394),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_415),
.B(n_426),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_379),
.A2(n_339),
.B(n_351),
.Y(n_417)
);

AO21x1_ASAP7_75t_L g458 ( 
.A1(n_417),
.A2(n_420),
.B(n_421),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_383),
.A2(n_333),
.B1(n_300),
.B2(n_310),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_378),
.A2(n_340),
.B(n_334),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_384),
.A2(n_340),
.B(n_334),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_379),
.A2(n_352),
.B(n_310),
.Y(n_422)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_423),
.Y(n_437)
);

INVx8_ASAP7_75t_L g424 ( 
.A(n_380),
.Y(n_424)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_424),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_362),
.B(n_372),
.C(n_385),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_374),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_379),
.B(n_308),
.Y(n_427)
);

AO21x1_ASAP7_75t_L g468 ( 
.A1(n_427),
.A2(n_391),
.B(n_376),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_388),
.B(n_295),
.C(n_314),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_433),
.B(n_359),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_411),
.B(n_369),
.Y(n_435)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_435),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_411),
.B(n_393),
.Y(n_436)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_436),
.Y(n_470)
);

OAI32xp33_ASAP7_75t_L g438 ( 
.A1(n_408),
.A2(n_366),
.A3(n_368),
.B1(n_387),
.B2(n_353),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_438),
.B(n_444),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_398),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_439),
.B(n_455),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_442),
.A2(n_448),
.B1(n_452),
.B2(n_462),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_398),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_398),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_445),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_446),
.A2(n_456),
.B1(n_400),
.B2(n_424),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_408),
.B(n_415),
.Y(n_447)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_447),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_426),
.A2(n_368),
.B1(n_360),
.B2(n_357),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_403),
.B(n_354),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_449),
.B(n_401),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_451),
.B(n_453),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_418),
.A2(n_367),
.B1(n_358),
.B2(n_364),
.Y(n_452)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_405),
.Y(n_454)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_454),
.Y(n_482)
);

INVxp33_ASAP7_75t_L g455 ( 
.A(n_434),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_418),
.A2(n_371),
.B1(n_363),
.B2(n_389),
.Y(n_456)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_405),
.Y(n_459)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_459),
.Y(n_497)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_416),
.Y(n_460)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_460),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_423),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_461),
.Y(n_494)
);

OAI22xp33_ASAP7_75t_SL g462 ( 
.A1(n_400),
.A2(n_414),
.B1(n_403),
.B2(n_413),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_412),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_463),
.Y(n_474)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_412),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_465),
.Y(n_472)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_416),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_423),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_466),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_427),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_467),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_468),
.A2(n_422),
.B(n_406),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_476),
.A2(n_496),
.B1(n_442),
.B2(n_448),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_478),
.B(n_483),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_425),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_479),
.B(n_480),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_450),
.B(n_402),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_441),
.B(n_377),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_446),
.A2(n_421),
.B1(n_420),
.B2(n_417),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_485),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_451),
.B(n_401),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_486),
.B(n_490),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_456),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_491),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_440),
.A2(n_427),
.B(n_443),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_489),
.A2(n_492),
.B(n_458),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_453),
.B(n_404),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_441),
.B(n_407),
.Y(n_491)
);

CKINVDCx14_ASAP7_75t_R g493 ( 
.A(n_457),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_493),
.B(n_445),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_457),
.A2(n_430),
.B1(n_433),
.B2(n_414),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_436),
.A2(n_432),
.B1(n_431),
.B2(n_429),
.Y(n_499)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_499),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_440),
.Y(n_501)
);

MAJx2_ASAP7_75t_L g530 ( 
.A(n_501),
.B(n_515),
.C(n_477),
.Y(n_530)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_504),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_505),
.A2(n_507),
.B1(n_509),
.B2(n_521),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_496),
.A2(n_452),
.B1(n_447),
.B2(n_467),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_472),
.Y(n_508)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_508),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_475),
.A2(n_444),
.B1(n_419),
.B2(n_435),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_475),
.B(n_466),
.Y(n_510)
);

INVxp33_ASAP7_75t_L g539 ( 
.A(n_510),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_471),
.A2(n_458),
.B1(n_468),
.B2(n_439),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_511),
.A2(n_470),
.B1(n_481),
.B2(n_489),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_498),
.B(n_495),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_513),
.B(n_518),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_479),
.B(n_399),
.C(n_468),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_514),
.B(n_512),
.C(n_502),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_486),
.B(n_458),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_472),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_516),
.B(n_523),
.Y(n_526)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_472),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_517),
.A2(n_524),
.B1(n_474),
.B2(n_508),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_498),
.B(n_461),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_519),
.B(n_520),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_477),
.B(n_438),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_494),
.A2(n_410),
.B1(n_437),
.B2(n_463),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_494),
.B(n_437),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_522),
.B(n_459),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_473),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_495),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_527),
.A2(n_429),
.B1(n_407),
.B2(n_428),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_503),
.A2(n_470),
.B1(n_481),
.B2(n_484),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_528),
.A2(n_533),
.B1(n_507),
.B2(n_521),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_530),
.B(n_532),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_524),
.A2(n_484),
.B(n_492),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_531),
.B(n_540),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_506),
.A2(n_469),
.B1(n_471),
.B2(n_478),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_513),
.A2(n_469),
.B(n_474),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_535),
.A2(n_500),
.B(n_454),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_SL g536 ( 
.A(n_515),
.B(n_490),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_536),
.B(n_512),
.Y(n_554)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_537),
.Y(n_550)
);

INVxp33_ASAP7_75t_SL g540 ( 
.A(n_525),
.Y(n_540)
);

FAx1_ASAP7_75t_SL g542 ( 
.A(n_519),
.B(n_497),
.CI(n_482),
.CON(n_542),
.SN(n_542)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_542),
.B(n_504),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_505),
.A2(n_497),
.B1(n_482),
.B2(n_464),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_544),
.A2(n_518),
.B1(n_511),
.B2(n_506),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_502),
.B(n_488),
.C(n_465),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_545),
.B(n_517),
.C(n_522),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_546),
.B(n_510),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_547),
.B(n_552),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_548),
.B(n_556),
.Y(n_567)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_549),
.Y(n_564)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_551),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_541),
.B(n_509),
.Y(n_552)
);

XNOR2x1_ASAP7_75t_L g574 ( 
.A(n_554),
.B(n_557),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_545),
.B(n_514),
.C(n_501),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_558),
.A2(n_559),
.B1(n_561),
.B2(n_527),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_529),
.A2(n_544),
.B1(n_534),
.B2(n_539),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_532),
.B(n_520),
.C(n_488),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_560),
.B(n_538),
.C(n_541),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_529),
.A2(n_460),
.B1(n_432),
.B2(n_431),
.Y(n_561)
);

CKINVDCx14_ASAP7_75t_R g562 ( 
.A(n_526),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_562),
.B(n_533),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_563),
.A2(n_542),
.B1(n_535),
.B2(n_428),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_565),
.B(n_571),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_550),
.A2(n_543),
.B1(n_539),
.B2(n_542),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_568),
.A2(n_558),
.B1(n_551),
.B2(n_547),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_554),
.B(n_560),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_570),
.B(n_577),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_556),
.B(n_538),
.C(n_530),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_572),
.B(n_573),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_548),
.B(n_528),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_575),
.A2(n_569),
.B1(n_555),
.B2(n_563),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_553),
.B(n_536),
.C(n_546),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_576),
.B(n_373),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_578),
.B(n_579),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_567),
.B(n_553),
.C(n_559),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_571),
.B(n_552),
.C(n_561),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_581),
.B(n_584),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_582),
.B(n_587),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_564),
.B(n_375),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_572),
.A2(n_382),
.B(n_381),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_SL g589 ( 
.A1(n_586),
.A2(n_576),
.B(n_566),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_577),
.A2(n_370),
.B1(n_365),
.B2(n_395),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_588),
.B(n_397),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_589),
.B(n_596),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_583),
.B(n_566),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_592),
.A2(n_581),
.B(n_585),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_580),
.B(n_570),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_593),
.B(n_594),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_579),
.B(n_574),
.C(n_575),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_SL g602 ( 
.A(n_598),
.B(n_601),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_591),
.B(n_585),
.C(n_578),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_600),
.B(n_595),
.Y(n_603)
);

MAJx2_ASAP7_75t_L g601 ( 
.A(n_592),
.B(n_574),
.C(n_392),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_603),
.B(n_341),
.C(n_316),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_597),
.B(n_590),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_604),
.A2(n_599),
.B(n_314),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_605),
.B(n_606),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_607),
.A2(n_602),
.B1(n_347),
.B2(n_316),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_608),
.A2(n_300),
.B(n_295),
.Y(n_609)
);

BUFx24_ASAP7_75t_SL g610 ( 
.A(n_609),
.Y(n_610)
);


endmodule