module fake_jpeg_15319_n_8 (n_3, n_2, n_1, n_0, n_4, n_8);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_8;

wire n_6;
wire n_5;
wire n_7;

NAND2xp5_ASAP7_75t_SL g5 ( 
.A(n_1),
.B(n_2),
.Y(n_5)
);

XOR2xp5_ASAP7_75t_L g6 ( 
.A(n_3),
.B(n_1),
.Y(n_6)
);

OAI21xp5_ASAP7_75t_SL g7 ( 
.A1(n_0),
.A2(n_2),
.B(n_4),
.Y(n_7)
);

NAND4xp25_ASAP7_75t_SL g8 ( 
.A(n_7),
.B(n_0),
.C(n_5),
.D(n_6),
.Y(n_8)
);


endmodule