module real_jpeg_26872_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_300;
wire n_292;
wire n_221;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_131;
wire n_47;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_127;
wire n_53;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_0),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_0),
.Y(n_92)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_0),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_1),
.A2(n_77),
.B1(n_78),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_1),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_174),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_174),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_1),
.A2(n_48),
.B1(n_51),
.B2(n_174),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_2),
.A2(n_45),
.B1(n_48),
.B2(n_51),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_2),
.A2(n_45),
.B1(n_77),
.B2(n_78),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_45),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_3),
.A2(n_58),
.B1(n_77),
.B2(n_78),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_3),
.A2(n_48),
.B1(n_51),
.B2(n_58),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_6),
.A2(n_77),
.B1(n_78),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_6),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_153),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_153),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_6),
.A2(n_48),
.B1(n_51),
.B2(n_153),
.Y(n_251)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_8),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_8),
.B(n_73),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_8),
.B(n_29),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g215 ( 
.A1(n_8),
.A2(n_29),
.B(n_211),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_172),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_8),
.A2(n_48),
.B(n_52),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_8),
.B(n_121),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_8),
.A2(n_89),
.B1(n_92),
.B2(n_259),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_9),
.A2(n_39),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_9),
.A2(n_39),
.B1(n_48),
.B2(n_51),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_41),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_10),
.A2(n_41),
.B1(n_48),
.B2(n_51),
.Y(n_143)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_12),
.A2(n_77),
.B1(n_78),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_12),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_127),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_127),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_12),
.A2(n_48),
.B1(n_51),
.B2(n_127),
.Y(n_246)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_14),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_15),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_131),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_102),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_19),
.B(n_102),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_86),
.B2(n_87),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_59),
.B2(n_60),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_23),
.A2(n_24),
.B(n_42),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_42),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_24)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_25),
.B(n_70),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_25),
.A2(n_33),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_25),
.A2(n_33),
.B1(n_168),
.B2(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_25),
.A2(n_33),
.B1(n_197),
.B2(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_33),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_26)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_27),
.Y(n_210)
);

NAND2xp33_ASAP7_75t_SL g212 ( 
.A(n_27),
.B(n_35),
.Y(n_212)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_29),
.A2(n_30),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_29),
.B(n_74),
.Y(n_186)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_30),
.A2(n_81),
.B1(n_171),
.B2(n_186),
.Y(n_185)
);

AOI32xp33_ASAP7_75t_L g209 ( 
.A1(n_30),
.A2(n_34),
.A3(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_209)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_33),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_33),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_33),
.B(n_149),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_35),
.B1(n_50),
.B2(n_52),
.Y(n_56)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_35),
.A2(n_50),
.B(n_172),
.C(n_238),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_38),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_53),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_43),
.A2(n_55),
.B(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_46),
.B(n_57),
.Y(n_98)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_55),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_47),
.A2(n_55),
.B1(n_97),
.B2(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_47),
.A2(n_53),
.B(n_119),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_47),
.A2(n_55),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_47),
.A2(n_55),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_47),
.A2(n_55),
.B1(n_218),
.B2(n_236),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_47),
.B(n_172),
.Y(n_257)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_51),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_55),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_55),
.A2(n_64),
.B(n_98),
.Y(n_165)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_71),
.B1(n_84),
.B2(n_85),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B(n_69),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_67),
.A2(n_69),
.B(n_148),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_67),
.A2(n_182),
.B(n_183),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_71),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_76),
.B(n_79),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_83),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_72),
.A2(n_125),
.B1(n_126),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_72),
.A2(n_125),
.B1(n_152),
.B2(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_74),
.B(n_78),
.C(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_73),
.B(n_100),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_73),
.A2(n_80),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_78),
.Y(n_81)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g171 ( 
.A(n_78),
.B(n_172),
.CON(n_171),
.SN(n_171)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_95),
.B(n_99),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_88),
.A2(n_99),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_88),
.A2(n_96),
.B1(n_106),
.B2(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_92),
.B(n_93),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_89),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_89),
.A2(n_117),
.B1(n_143),
.B2(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_89),
.A2(n_115),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_89),
.A2(n_92),
.B1(n_251),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_90),
.A2(n_94),
.B(n_145),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_90),
.A2(n_116),
.B1(n_250),
.B2(n_252),
.Y(n_249)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_91),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_92),
.B(n_114),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_92),
.A2(n_112),
.B(n_188),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_96),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_99),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.C(n_108),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_103),
.B(n_107),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_108),
.A2(n_109),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_120),
.C(n_123),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_118),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_111),
.B(n_118),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_120),
.A2(n_123),
.B1(n_124),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B(n_128),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_157),
.B(n_303),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_154),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_133),
.B(n_154),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.C(n_140),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_134),
.A2(n_135),
.B1(n_138),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_138),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_140),
.B(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_147),
.C(n_150),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_141),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_146),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_147),
.A2(n_150),
.B1(n_151),
.B2(n_293),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_147),
.Y(n_293)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_297),
.B(n_302),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_201),
.B(n_283),
.C(n_296),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_189),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_160),
.B(n_189),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_175),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_162),
.B(n_163),
.C(n_175),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_170),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_170),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_172),
.B(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_173),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_184),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_177),
.B(n_181),
.C(n_184),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_187),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.C(n_195),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_190),
.A2(n_191),
.B1(n_278),
.B2(n_280),
.Y(n_277)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_195),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.C(n_200),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_200),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_282),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_275),
.B(n_281),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_229),
.B(n_274),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_220),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_205),
.B(n_220),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_213),
.C(n_216),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_206),
.A2(n_207),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_209),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_221),
.B(n_227),
.C(n_228),
.Y(n_276)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_268),
.B(n_273),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_247),
.B(n_267),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_239),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_232),
.B(n_239),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_233),
.A2(n_234),
.B1(n_237),
.B2(n_254),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_245),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_244),
.C(n_245),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_246),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_255),
.B(n_266),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_249),
.B(n_253),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_260),
.B(n_265),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_257),
.B(n_258),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_276),
.B(n_277),
.Y(n_281)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_278),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_285),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_294),
.B2(n_295),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_291),
.C(n_295),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);


endmodule