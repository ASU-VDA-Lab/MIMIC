module fake_jpeg_26887_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_7),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_43),
.B(n_18),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_55),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_18),
.B(n_31),
.C(n_30),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_30),
.B(n_20),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_17),
.C(n_32),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_41),
.C(n_40),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_25),
.B1(n_24),
.B2(n_26),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_41),
.B1(n_37),
.B2(n_25),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_42),
.B(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_33),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_43),
.B(n_20),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_43),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_65),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_66),
.A2(n_74),
.B1(n_87),
.B2(n_61),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_37),
.B1(n_41),
.B2(n_34),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_68),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_76),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_19),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_81),
.C(n_86),
.Y(n_108)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_89),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_37),
.B1(n_41),
.B2(n_34),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_34),
.B1(n_51),
.B2(n_64),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_64),
.A2(n_34),
.B1(n_39),
.B2(n_36),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_86),
.B(n_91),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_63),
.A2(n_25),
.B1(n_23),
.B2(n_33),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_47),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_64),
.A2(n_39),
.B1(n_36),
.B2(n_38),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_83),
.B1(n_84),
.B2(n_46),
.Y(n_98)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_92),
.B(n_22),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_49),
.B1(n_46),
.B2(n_54),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_88),
.B1(n_47),
.B2(n_82),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_63),
.B(n_46),
.C(n_55),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_117),
.B(n_77),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_98),
.A2(n_85),
.B1(n_72),
.B2(n_88),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_76),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_99),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_79),
.A2(n_22),
.B1(n_30),
.B2(n_20),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_101),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_56),
.B(n_50),
.C(n_57),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_91),
.B(n_22),
.Y(n_130)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_106),
.B(n_114),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_43),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_112),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_80),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_110),
.B(n_29),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_70),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_86),
.B(n_43),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_70),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

OAI21x1_ASAP7_75t_SL g117 ( 
.A1(n_75),
.A2(n_38),
.B(n_32),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_38),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_120),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_40),
.Y(n_120)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_130),
.B(n_131),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_81),
.C(n_77),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_122),
.B(n_123),
.C(n_124),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_79),
.C(n_80),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_126),
.B(n_135),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_115),
.A2(n_109),
.B1(n_97),
.B2(n_112),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_97),
.B1(n_98),
.B2(n_96),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_67),
.B(n_27),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_137),
.Y(n_163)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_141),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_67),
.Y(n_139)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_143),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_144),
.B(n_149),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_145),
.A2(n_117),
.B1(n_99),
.B2(n_106),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_94),
.B(n_29),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_104),
.A2(n_27),
.B(n_16),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_150),
.A2(n_96),
.B(n_110),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_SL g198 ( 
.A1(n_151),
.A2(n_175),
.B(n_54),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_119),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_153),
.A2(n_174),
.B(n_177),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_94),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_166),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_156),
.A2(n_158),
.B1(n_143),
.B2(n_140),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g159 ( 
.A(n_132),
.B(n_104),
.CI(n_19),
.CON(n_159),
.SN(n_159)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_164),
.Y(n_199)
);

AOI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_127),
.A2(n_105),
.B(n_102),
.Y(n_162)
);

XNOR2x1_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_180),
.Y(n_194)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_127),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_165),
.Y(n_184)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_167),
.B(n_172),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_116),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_141),
.Y(n_202)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_122),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_123),
.Y(n_187)
);

BUFx12f_ASAP7_75t_SL g174 ( 
.A(n_133),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_114),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_111),
.B1(n_102),
.B2(n_45),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_179),
.A2(n_138),
.B1(n_147),
.B2(n_45),
.Y(n_189)
);

AND2x6_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_14),
.Y(n_180)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_131),
.B(n_40),
.Y(n_182)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_186),
.A2(n_189),
.B1(n_196),
.B2(n_158),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_188),
.C(n_191),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_130),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_176),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_160),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_150),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_156),
.A2(n_149),
.B1(n_135),
.B2(n_45),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_211),
.B1(n_152),
.B2(n_163),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_166),
.A2(n_54),
.B1(n_61),
.B2(n_39),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_201),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_182),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_28),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_207),
.C(n_212),
.Y(n_224)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_205),
.Y(n_223)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_155),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_210),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_154),
.B(n_129),
.C(n_40),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_153),
.B(n_129),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_157),
.A2(n_27),
.B1(n_39),
.B2(n_36),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_153),
.B(n_40),
.C(n_36),
.Y(n_212)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_214),
.B(n_217),
.Y(n_238)
);

AND2x4_ASAP7_75t_SL g215 ( 
.A(n_194),
.B(n_174),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_215),
.A2(n_231),
.B(n_159),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_161),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_235),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_180),
.C(n_178),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_209),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_225),
.A2(n_232),
.B1(n_237),
.B2(n_212),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_184),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_227),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_160),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_230),
.Y(n_255)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_179),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_199),
.B1(n_208),
.B2(n_197),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_185),
.B(n_161),
.Y(n_233)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_185),
.B(n_181),
.Y(n_234)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_193),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_189),
.B1(n_205),
.B2(n_201),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_239),
.A2(n_245),
.B1(n_247),
.B2(n_250),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_191),
.C(n_200),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_251),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_231),
.A2(n_195),
.B1(n_182),
.B2(n_193),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_215),
.A2(n_195),
.B1(n_159),
.B2(n_151),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_248),
.A2(n_254),
.B1(n_226),
.B2(n_237),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_235),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_215),
.A2(n_207),
.B1(n_171),
.B2(n_32),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_224),
.C(n_216),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_225),
.A2(n_171),
.B1(n_16),
.B2(n_11),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_40),
.C(n_28),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_223),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_267),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_257),
.C(n_243),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_233),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_263),
.Y(n_275)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_226),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_268),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_253),
.A2(n_221),
.B1(n_223),
.B2(n_28),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_266),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_244),
.A2(n_221),
.B1(n_10),
.B2(n_11),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_271),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_256),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_8),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_272),
.Y(n_282)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_250),
.Y(n_273)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_238),
.A2(n_9),
.B(n_15),
.Y(n_274)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_274),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_256),
.B1(n_272),
.B2(n_252),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_280),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_246),
.B1(n_241),
.B2(n_263),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_245),
.B1(n_247),
.B2(n_240),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_286),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_4),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_259),
.A2(n_240),
.B1(n_258),
.B2(n_40),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_261),
.B1(n_267),
.B2(n_269),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_296),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_6),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_292),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_284),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_6),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_297),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_277),
.A2(n_5),
.B(n_13),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_294),
.A2(n_12),
.B(n_15),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_279),
.A2(n_5),
.B1(n_12),
.B2(n_10),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_4),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_298),
.B(n_300),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_283),
.C(n_286),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_10),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_0),
.Y(n_316)
);

AOI211xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_281),
.B(n_276),
.C(n_280),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_305),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_295),
.B(n_285),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_3),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_290),
.A2(n_12),
.B(n_2),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_307),
.A2(n_3),
.B(n_0),
.Y(n_314)
);

AOI211x1_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_295),
.B(n_299),
.C(n_3),
.Y(n_311)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_0),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_312),
.B(n_313),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_314),
.A2(n_315),
.B(n_316),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_0),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_318),
.A2(n_310),
.B(n_308),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_321),
.C(n_303),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_312),
.B1(n_319),
.B2(n_302),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_2),
.Y(n_324)
);


endmodule