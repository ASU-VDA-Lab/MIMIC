module fake_netlist_1_9294_n_672 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_672);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_672;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_638;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_33), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_34), .Y(n_78) );
INVx1_ASAP7_75t_SL g79 ( .A(n_6), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_59), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_76), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_23), .Y(n_82) );
INVxp33_ASAP7_75t_L g83 ( .A(n_41), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_42), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_73), .Y(n_85) );
BUFx2_ASAP7_75t_L g86 ( .A(n_25), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_8), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_52), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_35), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_71), .Y(n_90) );
CKINVDCx16_ASAP7_75t_R g91 ( .A(n_68), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_67), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_15), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_2), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_45), .Y(n_95) );
INVxp67_ASAP7_75t_L g96 ( .A(n_65), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_31), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_37), .Y(n_98) );
BUFx3_ASAP7_75t_L g99 ( .A(n_75), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_66), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_16), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_30), .Y(n_102) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_46), .Y(n_103) );
INVxp33_ASAP7_75t_SL g104 ( .A(n_49), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_51), .Y(n_105) );
NOR2xp67_ASAP7_75t_L g106 ( .A(n_9), .B(n_12), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_8), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_63), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_43), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_53), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_20), .Y(n_111) );
INVx1_ASAP7_75t_SL g112 ( .A(n_54), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_12), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_40), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_38), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_5), .Y(n_116) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_69), .Y(n_117) );
INVx4_ASAP7_75t_R g118 ( .A(n_44), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_55), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_36), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_14), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_70), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_86), .B(n_0), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_83), .B(n_0), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_107), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_99), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_99), .Y(n_127) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_81), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_94), .Y(n_129) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_82), .A2(n_26), .B(n_72), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_107), .B(n_1), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_85), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_116), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_116), .B(n_3), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_88), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_89), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_83), .B(n_4), .Y(n_137) );
INVx5_ASAP7_75t_L g138 ( .A(n_103), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_103), .B(n_4), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_103), .B(n_5), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_113), .Y(n_141) );
INVx6_ASAP7_75t_L g142 ( .A(n_103), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_90), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_121), .B(n_6), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_92), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_91), .B(n_7), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_117), .B(n_7), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_93), .Y(n_148) );
AND2x2_ASAP7_75t_SL g149 ( .A(n_95), .B(n_122), .Y(n_149) );
INVxp67_ASAP7_75t_L g150 ( .A(n_94), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_100), .B(n_9), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_102), .Y(n_152) );
AND2x6_ASAP7_75t_L g153 ( .A(n_105), .B(n_32), .Y(n_153) );
INVx6_ASAP7_75t_L g154 ( .A(n_96), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_108), .B(n_10), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_110), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_111), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_77), .B(n_10), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_114), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g160 ( .A1(n_104), .A2(n_11), .B1(n_13), .B2(n_14), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_120), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_119), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_112), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_98), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_164), .B(n_97), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_164), .B(n_97), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_154), .B(n_104), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_131), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_131), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_131), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_154), .B(n_77), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_154), .B(n_84), .Y(n_172) );
OR2x2_ASAP7_75t_L g173 ( .A(n_129), .B(n_79), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_154), .B(n_80), .Y(n_174) );
AO22x2_ASAP7_75t_L g175 ( .A1(n_155), .A2(n_87), .B1(n_78), .B2(n_118), .Y(n_175) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_150), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
INVx4_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_135), .B(n_115), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_149), .B(n_109), .Y(n_180) );
BUFx4f_ASAP7_75t_L g181 ( .A(n_134), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_149), .B(n_115), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_155), .B(n_109), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_134), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_135), .B(n_84), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_144), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_144), .A2(n_143), .B1(n_148), .B2(n_136), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_138), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_136), .B(n_80), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_143), .B(n_101), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_144), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_155), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_138), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_145), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_141), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_148), .B(n_106), .Y(n_196) );
INVx1_ASAP7_75t_SL g197 ( .A(n_147), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_159), .B(n_78), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_138), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_138), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_153), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_141), .Y(n_202) );
INVx4_ASAP7_75t_SL g203 ( .A(n_153), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_138), .Y(n_204) );
AND2x6_ASAP7_75t_L g205 ( .A(n_158), .B(n_47), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_159), .B(n_87), .Y(n_206) );
AOI22xp33_ASAP7_75t_SL g207 ( .A1(n_147), .A2(n_11), .B1(n_13), .B2(n_17), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_141), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_145), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_163), .B(n_18), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_163), .B(n_19), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_132), .B(n_21), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_132), .B(n_162), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_145), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_145), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_145), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_179), .B(n_158), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_194), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_195), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_179), .B(n_124), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_167), .B(n_123), .Y(n_221) );
NOR2xp67_ASAP7_75t_L g222 ( .A(n_176), .B(n_128), .Y(n_222) );
BUFx2_ASAP7_75t_L g223 ( .A(n_197), .Y(n_223) );
INVx5_ASAP7_75t_L g224 ( .A(n_205), .Y(n_224) );
OR2x2_ASAP7_75t_L g225 ( .A(n_173), .B(n_137), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_185), .B(n_162), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_189), .B(n_157), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_169), .A2(n_153), .B1(n_157), .B2(n_156), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_206), .B(n_175), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_202), .Y(n_230) );
NOR2x2_ASAP7_75t_L g231 ( .A(n_175), .B(n_152), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_172), .B(n_152), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_172), .B(n_156), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_178), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_198), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_187), .A2(n_181), .B1(n_192), .B2(n_186), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_178), .B(n_151), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_187), .A2(n_160), .B1(n_146), .B2(n_126), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_190), .B(n_153), .Y(n_239) );
AND2x2_ASAP7_75t_SL g240 ( .A(n_181), .B(n_130), .Y(n_240) );
NOR2xp33_ASAP7_75t_SL g241 ( .A(n_178), .B(n_153), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_205), .Y(n_242) );
INVx1_ASAP7_75t_SL g243 ( .A(n_171), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_201), .B(n_161), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_167), .B(n_126), .Y(n_245) );
INVxp67_ASAP7_75t_L g246 ( .A(n_213), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_208), .Y(n_247) );
OR2x2_ASAP7_75t_L g248 ( .A(n_198), .B(n_133), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_174), .B(n_127), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_169), .A2(n_161), .B1(n_127), .B2(n_133), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_183), .B(n_125), .Y(n_251) );
BUFx3_ASAP7_75t_L g252 ( .A(n_205), .Y(n_252) );
BUFx6f_ASAP7_75t_SL g253 ( .A(n_205), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_175), .B(n_125), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_183), .B(n_161), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_191), .B(n_161), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_177), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g258 ( .A1(n_182), .A2(n_180), .B1(n_168), .B2(n_170), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_165), .B(n_161), .Y(n_259) );
INVxp67_ASAP7_75t_L g260 ( .A(n_166), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_177), .B(n_140), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_182), .A2(n_130), .B(n_139), .Y(n_262) );
AND3x1_ASAP7_75t_L g263 ( .A(n_184), .B(n_169), .C(n_211), .Y(n_263) );
INVx4_ASAP7_75t_L g264 ( .A(n_205), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_184), .A2(n_130), .B1(n_142), .B2(n_27), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_196), .B(n_142), .Y(n_266) );
BUFx2_ASAP7_75t_SL g267 ( .A(n_201), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_201), .A2(n_142), .B1(n_24), .B2(n_28), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_194), .Y(n_269) );
INVx8_ASAP7_75t_L g270 ( .A(n_203), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_196), .B(n_142), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_207), .B(n_22), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_203), .B(n_29), .Y(n_273) );
INVx8_ASAP7_75t_L g274 ( .A(n_203), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_210), .B(n_39), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_212), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_246), .B(n_200), .Y(n_277) );
OAI22x1_ASAP7_75t_L g278 ( .A1(n_223), .A2(n_194), .B1(n_215), .B2(n_209), .Y(n_278) );
BUFx2_ASAP7_75t_L g279 ( .A(n_246), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_234), .B(n_200), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_235), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_257), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_234), .B(n_264), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_241), .A2(n_216), .B(n_214), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_258), .B(n_204), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_239), .A2(n_214), .B(n_204), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_237), .A2(n_199), .B(n_193), .Y(n_287) );
INVx2_ASAP7_75t_SL g288 ( .A(n_225), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_219), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_260), .B(n_199), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_244), .A2(n_193), .B(n_188), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_230), .Y(n_292) );
HAxp5_ASAP7_75t_L g293 ( .A(n_222), .B(n_48), .CON(n_293), .SN(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_247), .Y(n_294) );
BUFx2_ASAP7_75t_L g295 ( .A(n_231), .Y(n_295) );
A2O1A1Ixp33_ASAP7_75t_L g296 ( .A1(n_221), .A2(n_188), .B(n_200), .C(n_57), .Y(n_296) );
INVx4_ASAP7_75t_L g297 ( .A(n_270), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_260), .Y(n_298) );
INVx2_ASAP7_75t_SL g299 ( .A(n_248), .Y(n_299) );
OA22x2_ASAP7_75t_L g300 ( .A1(n_229), .A2(n_50), .B1(n_56), .B2(n_58), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_244), .A2(n_200), .B(n_61), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_262), .A2(n_60), .B(n_62), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_256), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_262), .A2(n_64), .B(n_74), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_251), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_255), .Y(n_306) );
A2O1A1Ixp33_ASAP7_75t_L g307 ( .A1(n_221), .A2(n_220), .B(n_217), .C(n_227), .Y(n_307) );
OAI22x1_ASAP7_75t_L g308 ( .A1(n_254), .A2(n_272), .B1(n_264), .B2(n_224), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_226), .A2(n_249), .B(n_240), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_238), .B(n_243), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_234), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_266), .Y(n_312) );
BUFx2_ASAP7_75t_SL g313 ( .A(n_253), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_234), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_261), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_271), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_236), .A2(n_228), .B1(n_253), .B2(n_242), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_232), .B(n_233), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_270), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_224), .B(n_263), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g321 ( .A1(n_245), .A2(n_259), .B(n_252), .C(n_250), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_228), .A2(n_224), .B1(n_276), .B2(n_250), .Y(n_322) );
O2A1O1Ixp33_ASAP7_75t_L g323 ( .A1(n_273), .A2(n_275), .B(n_268), .C(n_269), .Y(n_323) );
INVxp67_ASAP7_75t_SL g324 ( .A(n_267), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_265), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_224), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_268), .A2(n_240), .B1(n_270), .B2(n_274), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_279), .Y(n_328) );
OAI21xp5_ASAP7_75t_L g329 ( .A1(n_309), .A2(n_218), .B(n_274), .Y(n_329) );
NOR2x1_ASAP7_75t_R g330 ( .A(n_281), .B(n_274), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_288), .A2(n_298), .B1(n_295), .B2(n_310), .Y(n_331) );
BUFx12f_ASAP7_75t_L g332 ( .A(n_297), .Y(n_332) );
A2O1A1Ixp33_ASAP7_75t_L g333 ( .A1(n_307), .A2(n_325), .B(n_318), .C(n_315), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_311), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_319), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_299), .B(n_318), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_323), .A2(n_286), .B(n_285), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_313), .Y(n_338) );
NOR2xp67_ASAP7_75t_SL g339 ( .A(n_297), .B(n_319), .Y(n_339) );
OAI22xp33_ASAP7_75t_L g340 ( .A1(n_290), .A2(n_300), .B1(n_292), .B2(n_294), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_290), .Y(n_341) );
BUFx2_ASAP7_75t_R g342 ( .A(n_320), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_285), .A2(n_287), .B(n_321), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_324), .Y(n_344) );
AOI21x1_ASAP7_75t_L g345 ( .A1(n_302), .A2(n_304), .B(n_327), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_305), .A2(n_322), .B1(n_289), .B2(n_317), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_282), .B(n_322), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_SL g348 ( .A1(n_296), .A2(n_283), .B(n_326), .C(n_327), .Y(n_348) );
AOI221x1_ASAP7_75t_L g349 ( .A1(n_308), .A2(n_317), .B1(n_278), .B2(n_301), .C(n_293), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_316), .Y(n_350) );
INVx2_ASAP7_75t_SL g351 ( .A(n_319), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_311), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_303), .Y(n_353) );
AOI21x1_ASAP7_75t_L g354 ( .A1(n_300), .A2(n_284), .B(n_280), .Y(n_354) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_306), .A2(n_291), .B(n_277), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_311), .Y(n_356) );
BUFx3_ASAP7_75t_L g357 ( .A(n_314), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_312), .Y(n_358) );
AO21x1_ASAP7_75t_L g359 ( .A1(n_314), .A2(n_325), .B(n_327), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_314), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_353), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_333), .B(n_341), .Y(n_362) );
AOI21xp33_ASAP7_75t_L g363 ( .A1(n_340), .A2(n_347), .B(n_346), .Y(n_363) );
OA21x2_ASAP7_75t_L g364 ( .A1(n_337), .A2(n_359), .B(n_343), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_350), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_341), .Y(n_366) );
BUFx12f_ASAP7_75t_L g367 ( .A(n_332), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_336), .B(n_344), .Y(n_368) );
OA21x2_ASAP7_75t_L g369 ( .A1(n_359), .A2(n_349), .B(n_345), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_348), .A2(n_355), .B(n_349), .Y(n_370) );
OR2x6_ASAP7_75t_L g371 ( .A(n_344), .B(n_352), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_334), .Y(n_372) );
OA21x2_ASAP7_75t_L g373 ( .A1(n_345), .A2(n_354), .B(n_329), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_334), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_331), .B(n_328), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g376 ( .A1(n_354), .A2(n_360), .B(n_358), .Y(n_376) );
OAI21xp5_ASAP7_75t_L g377 ( .A1(n_357), .A2(n_351), .B(n_328), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_332), .B(n_330), .Y(n_378) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_352), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_351), .B(n_357), .Y(n_380) );
OAI21x1_ASAP7_75t_L g381 ( .A1(n_352), .A2(n_356), .B(n_342), .Y(n_381) );
OAI21x1_ASAP7_75t_L g382 ( .A1(n_352), .A2(n_356), .B(n_339), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_338), .A2(n_339), .B1(n_335), .B2(n_352), .C(n_356), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_356), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_356), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_335), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_338), .B(n_336), .Y(n_387) );
OA21x2_ASAP7_75t_L g388 ( .A1(n_370), .A2(n_376), .B(n_363), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_362), .B(n_363), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_372), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_385), .B(n_371), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_372), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_374), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_362), .B(n_365), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_366), .B(n_375), .Y(n_395) );
INVxp67_ASAP7_75t_SL g396 ( .A(n_366), .Y(n_396) );
OA21x2_ASAP7_75t_L g397 ( .A1(n_370), .A2(n_376), .B(n_382), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_368), .B(n_374), .Y(n_398) );
BUFx3_ASAP7_75t_L g399 ( .A(n_371), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_384), .Y(n_400) );
OA21x2_ASAP7_75t_L g401 ( .A1(n_382), .A2(n_381), .B(n_384), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_367), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_368), .B(n_361), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_365), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_364), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_361), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_385), .B(n_371), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_384), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_371), .Y(n_409) );
OA21x2_ASAP7_75t_L g410 ( .A1(n_382), .A2(n_381), .B(n_383), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_371), .B(n_369), .Y(n_411) );
BUFx2_ASAP7_75t_L g412 ( .A(n_379), .Y(n_412) );
BUFx3_ASAP7_75t_L g413 ( .A(n_379), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_385), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_375), .A2(n_383), .B1(n_377), .B2(n_387), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_379), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_379), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_379), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_364), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_404), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_400), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_403), .A2(n_387), .B1(n_367), .B2(n_378), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_400), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_404), .Y(n_424) );
INVx1_ASAP7_75t_SL g425 ( .A(n_402), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_403), .B(n_367), .Y(n_426) );
INVx2_ASAP7_75t_SL g427 ( .A(n_399), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_406), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_406), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g430 ( .A1(n_415), .A2(n_377), .B1(n_381), .B2(n_369), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_400), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_403), .B(n_386), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_398), .B(n_369), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_390), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_415), .A2(n_386), .B1(n_380), .B2(n_369), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_408), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_398), .B(n_393), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_408), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_398), .B(n_364), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_408), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_405), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_390), .B(n_386), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_399), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_392), .Y(n_444) );
INVx2_ASAP7_75t_SL g445 ( .A(n_399), .Y(n_445) );
INVxp67_ASAP7_75t_L g446 ( .A(n_396), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_411), .B(n_364), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_405), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_395), .B(n_373), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_392), .Y(n_450) );
NOR2x1_ASAP7_75t_L g451 ( .A(n_399), .B(n_385), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_411), .B(n_373), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_396), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_393), .B(n_380), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_394), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_411), .B(n_373), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_394), .B(n_373), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_405), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_405), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_395), .B(n_379), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_391), .B(n_407), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_419), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_395), .B(n_409), .Y(n_463) );
NOR2x1p5_ASAP7_75t_L g464 ( .A(n_409), .B(n_389), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_419), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_437), .B(n_391), .Y(n_466) );
INVx3_ASAP7_75t_L g467 ( .A(n_465), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_432), .B(n_391), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_433), .B(n_419), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_422), .B(n_389), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_433), .B(n_419), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_453), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_461), .B(n_391), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_422), .B(n_414), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_425), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_451), .A2(n_412), .B(n_410), .Y(n_476) );
AOI22xp33_ASAP7_75t_SL g477 ( .A1(n_426), .A2(n_391), .B1(n_407), .B2(n_410), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_455), .B(n_407), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_439), .B(n_388), .Y(n_479) );
NOR3xp33_ASAP7_75t_SL g480 ( .A(n_454), .B(n_424), .C(n_428), .Y(n_480) );
NAND2x1_ASAP7_75t_L g481 ( .A(n_453), .B(n_410), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_441), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_441), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_448), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_420), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_463), .B(n_407), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_420), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_439), .B(n_388), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_424), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_447), .B(n_388), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_448), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_447), .B(n_388), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_459), .Y(n_493) );
NAND2x1_ASAP7_75t_SL g494 ( .A(n_451), .B(n_410), .Y(n_494) );
INVxp67_ASAP7_75t_L g495 ( .A(n_434), .Y(n_495) );
INVxp67_ASAP7_75t_L g496 ( .A(n_434), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_463), .B(n_407), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_428), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_461), .B(n_412), .Y(n_499) );
BUFx2_ASAP7_75t_SL g500 ( .A(n_427), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_446), .B(n_414), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_459), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_452), .B(n_388), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_452), .B(n_388), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_455), .B(n_412), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_465), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_429), .B(n_410), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_429), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_456), .B(n_413), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_464), .B(n_410), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_456), .B(n_397), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_444), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_444), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_427), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_450), .Y(n_515) );
INVx2_ASAP7_75t_SL g516 ( .A(n_443), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_442), .B(n_416), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_458), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_460), .B(n_416), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_450), .B(n_401), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_457), .B(n_397), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_511), .B(n_457), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_485), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_511), .B(n_449), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_521), .B(n_449), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_521), .B(n_462), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_503), .B(n_462), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_503), .B(n_458), .Y(n_528) );
INVx2_ASAP7_75t_SL g529 ( .A(n_514), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_472), .Y(n_530) );
INVx1_ASAP7_75t_SL g531 ( .A(n_475), .Y(n_531) );
INVx2_ASAP7_75t_SL g532 ( .A(n_514), .Y(n_532) );
INVxp67_ASAP7_75t_L g533 ( .A(n_500), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_469), .B(n_460), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_504), .B(n_464), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_469), .B(n_471), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_473), .B(n_499), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_487), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_471), .B(n_436), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_489), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_504), .B(n_397), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_498), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_490), .B(n_397), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_470), .B(n_435), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_508), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_490), .B(n_397), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_475), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_512), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_513), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_470), .B(n_445), .Y(n_550) );
OAI21xp5_ASAP7_75t_L g551 ( .A1(n_480), .A2(n_430), .B(n_445), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_495), .B(n_443), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_492), .B(n_397), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_492), .B(n_421), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_519), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_518), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_496), .B(n_421), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_479), .B(n_423), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_516), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_515), .B(n_423), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_478), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_501), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_479), .B(n_440), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_505), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_488), .B(n_440), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_466), .B(n_438), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_518), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_520), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_520), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_467), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_473), .B(n_438), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_488), .B(n_509), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_509), .B(n_431), .Y(n_573) );
OAI21xp5_ASAP7_75t_L g574 ( .A1(n_533), .A2(n_477), .B(n_474), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_568), .B(n_510), .Y(n_575) );
INVx2_ASAP7_75t_SL g576 ( .A(n_529), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_568), .B(n_474), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_529), .B(n_516), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_530), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_556), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_536), .B(n_468), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_572), .B(n_473), .Y(n_582) );
INVx2_ASAP7_75t_SL g583 ( .A(n_532), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_536), .B(n_497), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_523), .Y(n_585) );
OAI22xp33_ASAP7_75t_R g586 ( .A1(n_531), .A2(n_486), .B1(n_517), .B2(n_483), .Y(n_586) );
NAND2xp33_ASAP7_75t_SL g587 ( .A(n_532), .B(n_481), .Y(n_587) );
OAI32xp33_ASAP7_75t_L g588 ( .A1(n_547), .A2(n_507), .A3(n_467), .B1(n_502), .B2(n_483), .Y(n_588) );
NAND2xp33_ASAP7_75t_L g589 ( .A(n_551), .B(n_467), .Y(n_589) );
OAI221xp5_ASAP7_75t_L g590 ( .A1(n_544), .A2(n_494), .B1(n_476), .B2(n_502), .C(n_506), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_569), .B(n_499), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_569), .B(n_499), .Y(n_592) );
OAI32xp33_ASAP7_75t_L g593 ( .A1(n_559), .A2(n_493), .A3(n_491), .B1(n_484), .B2(n_482), .Y(n_593) );
NOR2x1p5_ASAP7_75t_L g594 ( .A(n_537), .B(n_509), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_572), .B(n_506), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_523), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_524), .B(n_493), .Y(n_597) );
INVx1_ASAP7_75t_SL g598 ( .A(n_555), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_540), .Y(n_599) );
NAND3xp33_ASAP7_75t_SL g600 ( .A(n_550), .B(n_491), .C(n_484), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_522), .B(n_482), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_522), .B(n_401), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_540), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_571), .B(n_431), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_524), .B(n_436), .Y(n_605) );
INVx2_ASAP7_75t_SL g606 ( .A(n_537), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_539), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_561), .B(n_401), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_535), .B(n_525), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_562), .B(n_401), .Y(n_610) );
OAI21xp33_ASAP7_75t_L g611 ( .A1(n_535), .A2(n_413), .B(n_416), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_610), .B(n_528), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_585), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_596), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_586), .A2(n_553), .B1(n_543), .B2(n_541), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_610), .B(n_553), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_605), .B(n_525), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_599), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_603), .Y(n_619) );
AOI21xp33_ASAP7_75t_L g620 ( .A1(n_589), .A2(n_548), .B(n_538), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_581), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_597), .Y(n_622) );
AOI211x1_ASAP7_75t_SL g623 ( .A1(n_574), .A2(n_552), .B(n_557), .C(n_570), .Y(n_623) );
INVxp67_ASAP7_75t_L g624 ( .A(n_578), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_579), .Y(n_625) );
INVx3_ASAP7_75t_L g626 ( .A(n_606), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_584), .Y(n_627) );
OAI32xp33_ASAP7_75t_L g628 ( .A1(n_587), .A2(n_534), .A3(n_539), .B1(n_526), .B2(n_527), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_598), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_580), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_607), .B(n_526), .Y(n_631) );
OAI211xp5_ASAP7_75t_SL g632 ( .A1(n_589), .A2(n_564), .B(n_549), .C(n_542), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_587), .B(n_578), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_577), .A2(n_527), .B1(n_528), .B2(n_543), .C(n_541), .Y(n_634) );
OAI221xp5_ASAP7_75t_SL g635 ( .A1(n_615), .A2(n_590), .B1(n_576), .B2(n_583), .C(n_611), .Y(n_635) );
OAI21xp33_ASAP7_75t_L g636 ( .A1(n_628), .A2(n_592), .B(n_591), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_613), .Y(n_637) );
OAI211xp5_ASAP7_75t_SL g638 ( .A1(n_623), .A2(n_575), .B(n_606), .C(n_604), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_634), .B(n_602), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_616), .B(n_609), .Y(n_640) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_629), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_614), .Y(n_642) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_629), .A2(n_588), .B1(n_593), .B2(n_537), .Y(n_643) );
OAI322xp33_ASAP7_75t_SL g644 ( .A1(n_612), .A2(n_608), .A3(n_604), .B1(n_549), .B2(n_542), .C1(n_545), .C2(n_580), .Y(n_644) );
AOI222xp33_ASAP7_75t_L g645 ( .A1(n_633), .A2(n_600), .B1(n_546), .B2(n_601), .C1(n_594), .C2(n_595), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_620), .A2(n_600), .B(n_571), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g647 ( .A1(n_624), .A2(n_582), .B(n_546), .Y(n_647) );
OAI21xp5_ASAP7_75t_SL g648 ( .A1(n_620), .A2(n_571), .B(n_573), .Y(n_648) );
OAI211xp5_ASAP7_75t_L g649 ( .A1(n_645), .A2(n_632), .B(n_626), .C(n_625), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_638), .B(n_618), .C(n_619), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_644), .A2(n_612), .B1(n_621), .B2(n_627), .C(n_626), .Y(n_651) );
A2O1A1Ixp33_ASAP7_75t_L g652 ( .A1(n_635), .A2(n_631), .B(n_617), .C(n_622), .Y(n_652) );
NAND2xp33_ASAP7_75t_R g653 ( .A(n_646), .B(n_630), .Y(n_653) );
A2O1A1Ixp33_ASAP7_75t_L g654 ( .A1(n_648), .A2(n_566), .B(n_534), .C(n_565), .Y(n_654) );
NAND3xp33_ASAP7_75t_L g655 ( .A(n_643), .B(n_545), .C(n_567), .Y(n_655) );
OAI211xp5_ASAP7_75t_L g656 ( .A1(n_643), .A2(n_573), .B(n_558), .C(n_554), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_650), .Y(n_657) );
OAI21xp33_ASAP7_75t_SL g658 ( .A1(n_651), .A2(n_639), .B(n_641), .Y(n_658) );
NOR3xp33_ASAP7_75t_L g659 ( .A(n_655), .B(n_636), .C(n_647), .Y(n_659) );
AOI211xp5_ASAP7_75t_SL g660 ( .A1(n_656), .A2(n_642), .B(n_637), .C(n_640), .Y(n_660) );
AOI221xp5_ASAP7_75t_L g661 ( .A1(n_652), .A2(n_565), .B1(n_563), .B2(n_554), .C(n_558), .Y(n_661) );
NOR2x1p5_ASAP7_75t_L g662 ( .A(n_657), .B(n_653), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_660), .B(n_654), .Y(n_663) );
NOR3xp33_ASAP7_75t_L g664 ( .A(n_658), .B(n_649), .C(n_560), .Y(n_664) );
NOR3xp33_ASAP7_75t_SL g665 ( .A(n_662), .B(n_661), .C(n_659), .Y(n_665) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_663), .Y(n_666) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_666), .Y(n_667) );
OAI22xp5_ASAP7_75t_SL g668 ( .A1(n_667), .A2(n_665), .B1(n_664), .B2(n_570), .Y(n_668) );
AOI222xp33_ASAP7_75t_L g669 ( .A1(n_668), .A2(n_556), .B1(n_563), .B2(n_418), .C1(n_417), .C2(n_413), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_669), .B(n_418), .Y(n_670) );
OAI21xp5_ASAP7_75t_L g671 ( .A1(n_670), .A2(n_418), .B(n_417), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_671), .A2(n_401), .B1(n_413), .B2(n_418), .Y(n_672) );
endmodule