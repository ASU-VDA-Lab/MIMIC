module real_jpeg_12471_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx2_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_2),
.A2(n_35),
.B1(n_39),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_2),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_3),
.A2(n_28),
.B1(n_31),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_71),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_3),
.A2(n_35),
.B1(n_39),
.B2(n_71),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_5),
.A2(n_35),
.B1(n_39),
.B2(n_56),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_6),
.A2(n_28),
.B1(n_31),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_64),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_6),
.A2(n_35),
.B1(n_39),
.B2(n_64),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_9),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_10),
.A2(n_35),
.B1(n_39),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_11),
.B(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_11),
.A2(n_43),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_11),
.B(n_88),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_12),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_38),
.Y(n_59)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_92),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_91),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_85),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_18),
.B(n_85),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_60),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_46),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_21),
.B(n_33),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B(n_26),
.C(n_30),
.Y(n_21)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

OA22x2_ASAP7_75t_SL g67 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_32),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_22),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_23),
.A2(n_24),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_23),
.B(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NOR3xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_31),
.C(n_32),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_27),
.A2(n_63),
.B1(n_66),
.B2(n_88),
.Y(n_87)
);

HAxp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_29),
.CON(n_27),
.SN(n_27)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_28),
.A2(n_31),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_29),
.B(n_39),
.C(n_51),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_29),
.B(n_43),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_29),
.B(n_53),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_40),
.B(n_42),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_34),
.B(n_41),
.Y(n_125)
);

CKINVDCx6p67_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_39),
.B1(n_50),
.B2(n_51),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_39),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_40),
.B(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_40),
.A2(n_41),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_40),
.Y(n_115)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_43),
.A2(n_81),
.B(n_83),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_43),
.A2(n_106),
.B1(n_114),
.B2(n_115),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_54),
.B(n_57),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_48),
.A2(n_55),
.B1(n_58),
.B2(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_58),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_48),
.A2(n_58),
.B1(n_90),
.B2(n_101),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_72),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_65),
.B1(n_67),
.B2(n_69),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_79),
.B2(n_80),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.C(n_89),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_86),
.B(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_89),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_132),
.B(n_136),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_121),
.B(n_131),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_109),
.B(n_120),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_104),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_104),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_96)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_102),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_115),
.B(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_116),
.B(n_119),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_118),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_123),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_127),
.C(n_130),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_135),
.Y(n_136)
);


endmodule