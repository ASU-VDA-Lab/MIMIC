module fake_jpeg_5109_n_31 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_31);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_31;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_24;
wire n_28;
wire n_26;
wire n_25;
wire n_17;
wire n_29;

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_12),
.A2(n_0),
.B1(n_5),
.B2(n_15),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_3),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_9),
.B(n_2),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_21),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_24)
);

AOI21x1_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_25),
.B(n_26),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_17),
.A2(n_1),
.B(n_2),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_18),
.A2(n_1),
.B1(n_16),
.B2(n_23),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_28),
.A2(n_24),
.B1(n_27),
.B2(n_20),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_29),
.A2(n_17),
.B(n_22),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_19),
.Y(n_31)
);


endmodule