module fake_ariane_2020_n_774 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_774);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_774;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_116),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_10),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_66),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_21),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

BUFx8_ASAP7_75t_SL g160 ( 
.A(n_43),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_31),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_0),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_4),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_8),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_15),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_11),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_4),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_20),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_107),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_118),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_54),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_37),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_32),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_10),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_152),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_97),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_83),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_44),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_56),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_36),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_17),
.Y(n_185)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_153),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_120),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_29),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_60),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_65),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_52),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_76),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_112),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_69),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_98),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_47),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_90),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_1),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_136),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_18),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_109),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_67),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_102),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_75),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_70),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_127),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_53),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_0),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_166),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_213)
);

AOI22x1_ASAP7_75t_SL g214 ( 
.A1(n_173),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_159),
.B(n_5),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

BUFx8_ASAP7_75t_SL g222 ( 
.A(n_160),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_164),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

XNOR2x2_ASAP7_75t_L g227 ( 
.A(n_155),
.B(n_6),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_168),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_157),
.Y(n_229)
);

OAI21x1_ASAP7_75t_L g230 ( 
.A1(n_157),
.A2(n_82),
.B(n_150),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_165),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_174),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_160),
.Y(n_237)
);

AOI22x1_ASAP7_75t_SL g238 ( 
.A1(n_173),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_196),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_179),
.Y(n_242)
);

OAI21x1_ASAP7_75t_L g243 ( 
.A1(n_205),
.A2(n_84),
.B(n_148),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_176),
.B(n_7),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_184),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_169),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_189),
.Y(n_249)
);

AND3x2_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_158),
.C(n_183),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_210),
.Y(n_251)
);

OR2x6_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_178),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_210),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_235),
.B(n_202),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_210),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_235),
.B(n_203),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_225),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_218),
.B(n_203),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_210),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_221),
.Y(n_271)
);

AO22x2_ASAP7_75t_L g272 ( 
.A1(n_214),
.A2(n_198),
.B1(n_192),
.B2(n_207),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_221),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_234),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_225),
.B(n_190),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_234),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_234),
.Y(n_277)
);

AOI21x1_ASAP7_75t_L g278 ( 
.A1(n_229),
.A2(n_194),
.B(n_186),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_239),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_225),
.B(n_161),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_225),
.B(n_199),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_221),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_208),
.B(n_154),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_208),
.B(n_156),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_239),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_221),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_239),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_221),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_239),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_224),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_224),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_244),
.B(n_167),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_246),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_240),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_240),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_288),
.Y(n_297)
);

NOR2xp67_ASAP7_75t_L g298 ( 
.A(n_261),
.B(n_215),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_240),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_249),
.B(n_240),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_215),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_240),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_283),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_261),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_291),
.Y(n_307)
);

BUFx6f_ASAP7_75t_SL g308 ( 
.A(n_259),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_256),
.B(n_217),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_248),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_256),
.B(n_217),
.Y(n_311)
);

INVx8_ASAP7_75t_L g312 ( 
.A(n_252),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_261),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_262),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_266),
.B(n_219),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_259),
.Y(n_316)
);

OR2x2_ASAP7_75t_SL g317 ( 
.A(n_272),
.B(n_222),
.Y(n_317)
);

NOR3xp33_ASAP7_75t_L g318 ( 
.A(n_269),
.B(n_242),
.C(n_211),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_248),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_252),
.B(n_242),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_266),
.B(n_216),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_262),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_259),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_284),
.B(n_219),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_263),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_293),
.B(n_216),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_269),
.B(n_220),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_262),
.B(n_220),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_291),
.B(n_245),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_253),
.B(n_240),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_253),
.B(n_246),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_278),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_257),
.B(n_258),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_257),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_248),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_245),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_258),
.B(n_246),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_264),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_252),
.A2(n_193),
.B1(n_188),
.B2(n_179),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_263),
.B(n_245),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_264),
.B(n_265),
.Y(n_341)
);

OR2x6_ASAP7_75t_L g342 ( 
.A(n_272),
.B(n_227),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_250),
.B(n_232),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_265),
.B(n_268),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_263),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_268),
.A2(n_236),
.B1(n_241),
.B2(n_232),
.Y(n_346)
);

NOR2xp67_ASAP7_75t_L g347 ( 
.A(n_294),
.B(n_236),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_274),
.B(n_241),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_274),
.B(n_229),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_251),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_294),
.B(n_212),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_254),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_255),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_260),
.Y(n_354)
);

BUFx6f_ASAP7_75t_SL g355 ( 
.A(n_270),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_271),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_276),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_248),
.B(n_188),
.Y(n_358)
);

NAND2x1p5_ASAP7_75t_L g359 ( 
.A(n_340),
.B(n_273),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_351),
.Y(n_360)
);

O2A1O1Ixp33_ASAP7_75t_L g361 ( 
.A1(n_309),
.A2(n_247),
.B(n_228),
.C(n_292),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_334),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_305),
.B(n_282),
.Y(n_364)
);

NAND2x1p5_ASAP7_75t_L g365 ( 
.A(n_323),
.B(n_286),
.Y(n_365)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_325),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_299),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_295),
.A2(n_243),
.B(n_230),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_295),
.A2(n_290),
.B(n_289),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_301),
.A2(n_290),
.B(n_289),
.Y(n_370)
);

NAND3xp33_ASAP7_75t_L g371 ( 
.A(n_303),
.B(n_238),
.C(n_214),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_324),
.B(n_276),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_301),
.A2(n_300),
.B(n_296),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_327),
.B(n_329),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_345),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_332),
.A2(n_230),
.B(n_243),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_336),
.B(n_277),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_326),
.B(n_298),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_296),
.A2(n_287),
.B(n_285),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_316),
.B(n_212),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_311),
.B(n_277),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_300),
.A2(n_287),
.B(n_285),
.Y(n_382)
);

O2A1O1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_315),
.A2(n_228),
.B(n_247),
.C(n_279),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_307),
.B(n_279),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_350),
.A2(n_233),
.B(n_204),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_308),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_339),
.B(n_212),
.Y(n_387)
);

OAI21xp33_ASAP7_75t_L g388 ( 
.A1(n_318),
.A2(n_247),
.B(n_228),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_307),
.B(n_233),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_304),
.B(n_224),
.Y(n_390)
);

O2A1O1Ixp33_ASAP7_75t_L g391 ( 
.A1(n_321),
.A2(n_209),
.B(n_226),
.C(n_223),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_304),
.A2(n_197),
.B(n_171),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_354),
.B(n_193),
.Y(n_393)
);

AOI33xp33_ASAP7_75t_L g394 ( 
.A1(n_313),
.A2(n_209),
.A3(n_226),
.B1(n_227),
.B2(n_346),
.B3(n_238),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_312),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_328),
.B(n_224),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_343),
.Y(n_397)
);

OAI321xp33_ASAP7_75t_L g398 ( 
.A1(n_342),
.A2(n_224),
.A3(n_272),
.B1(n_223),
.B2(n_13),
.C(n_14),
.Y(n_398)
);

A2O1A1Ixp33_ASAP7_75t_L g399 ( 
.A1(n_306),
.A2(n_223),
.B(n_206),
.C(n_200),
.Y(n_399)
);

NOR3xp33_ASAP7_75t_L g400 ( 
.A(n_320),
.B(n_195),
.C(n_187),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_338),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_314),
.B(n_170),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_319),
.A2(n_180),
.B(n_85),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_358),
.B(n_9),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_322),
.A2(n_81),
.B(n_147),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_353),
.B(n_9),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_342),
.A2(n_297),
.B1(n_302),
.B2(n_312),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_333),
.A2(n_80),
.B(n_146),
.Y(n_408)
);

A2O1A1Ixp33_ASAP7_75t_L g409 ( 
.A1(n_352),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_333),
.A2(n_86),
.B(n_145),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_310),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_348),
.B(n_356),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_341),
.A2(n_79),
.B(n_143),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_341),
.A2(n_78),
.B(n_142),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_344),
.B(n_12),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_349),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_344),
.A2(n_87),
.B(n_141),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_L g418 ( 
.A(n_349),
.B(n_19),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_331),
.A2(n_77),
.B(n_140),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_347),
.B(n_14),
.Y(n_420)
);

OAI21xp33_ASAP7_75t_L g421 ( 
.A1(n_342),
.A2(n_15),
.B(n_16),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_357),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_331),
.B(n_16),
.Y(n_423)
);

O2A1O1Ixp5_ASAP7_75t_L g424 ( 
.A1(n_337),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_337),
.A2(n_25),
.B(n_26),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_387),
.B(n_312),
.Y(n_426)
);

AOI21x1_ASAP7_75t_L g427 ( 
.A1(n_373),
.A2(n_330),
.B(n_335),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_363),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_367),
.B(n_308),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_368),
.A2(n_330),
.B(n_335),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_369),
.A2(n_335),
.B(n_310),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_360),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_384),
.A2(n_310),
.B(n_355),
.Y(n_433)
);

OAI21x1_ASAP7_75t_L g434 ( 
.A1(n_376),
.A2(n_355),
.B(n_28),
.Y(n_434)
);

OAI21x1_ASAP7_75t_L g435 ( 
.A1(n_379),
.A2(n_27),
.B(n_30),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_401),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_380),
.Y(n_437)
);

AND2x2_ASAP7_75t_SL g438 ( 
.A(n_394),
.B(n_398),
.Y(n_438)
);

AOI21xp33_ASAP7_75t_L g439 ( 
.A1(n_397),
.A2(n_317),
.B(n_34),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_374),
.A2(n_33),
.B(n_35),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_389),
.A2(n_38),
.B(n_39),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_416),
.B(n_40),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_412),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_422),
.Y(n_444)
);

AO21x1_ASAP7_75t_L g445 ( 
.A1(n_390),
.A2(n_41),
.B(n_42),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_382),
.A2(n_45),
.B(n_46),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_370),
.A2(n_48),
.B(n_49),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_362),
.B(n_50),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_364),
.B(n_51),
.Y(n_449)
);

AOI21x1_ASAP7_75t_L g450 ( 
.A1(n_381),
.A2(n_377),
.B(n_372),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_415),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_375),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_392),
.A2(n_55),
.B(n_57),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_388),
.B(n_58),
.Y(n_454)
);

O2A1O1Ixp5_ASAP7_75t_L g455 ( 
.A1(n_423),
.A2(n_59),
.B(n_61),
.C(n_62),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_378),
.B(n_63),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_383),
.A2(n_64),
.B(n_68),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_361),
.A2(n_385),
.B(n_424),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_396),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_406),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_402),
.A2(n_71),
.B(n_72),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_403),
.A2(n_73),
.B(n_74),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_408),
.A2(n_88),
.B(n_89),
.Y(n_463)
);

OAI21x1_ASAP7_75t_L g464 ( 
.A1(n_410),
.A2(n_91),
.B(n_92),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_375),
.B(n_93),
.Y(n_465)
);

AOI21x1_ASAP7_75t_L g466 ( 
.A1(n_418),
.A2(n_94),
.B(n_95),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_413),
.A2(n_414),
.B(n_417),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_359),
.B(n_96),
.Y(n_468)
);

OAI21x1_ASAP7_75t_SL g469 ( 
.A1(n_366),
.A2(n_151),
.B(n_100),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_399),
.A2(n_99),
.B(n_104),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_419),
.A2(n_105),
.B(n_106),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_425),
.A2(n_108),
.B(n_110),
.Y(n_472)
);

NAND3xp33_ASAP7_75t_L g473 ( 
.A(n_371),
.B(n_421),
.C(n_393),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_359),
.A2(n_111),
.B(n_113),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_420),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_391),
.A2(n_405),
.B(n_404),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_407),
.B(n_114),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_395),
.B(n_115),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_411),
.A2(n_119),
.B(n_122),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_366),
.Y(n_480)
);

OAI21xp33_ASAP7_75t_L g481 ( 
.A1(n_409),
.A2(n_123),
.B(n_124),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_365),
.A2(n_125),
.B(n_126),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_467),
.A2(n_411),
.B(n_365),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_452),
.Y(n_484)
);

NAND3xp33_ASAP7_75t_L g485 ( 
.A(n_481),
.B(n_400),
.C(n_460),
.Y(n_485)
);

OAI21x1_ASAP7_75t_L g486 ( 
.A1(n_434),
.A2(n_411),
.B(n_398),
.Y(n_486)
);

OA21x2_ASAP7_75t_L g487 ( 
.A1(n_430),
.A2(n_386),
.B(n_129),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_434),
.A2(n_128),
.B(n_130),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_482),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_429),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_427),
.A2(n_131),
.B(n_132),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_480),
.Y(n_492)
);

AO21x2_ASAP7_75t_L g493 ( 
.A1(n_458),
.A2(n_133),
.B(n_134),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_426),
.B(n_135),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_428),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_443),
.A2(n_137),
.B(n_138),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_450),
.A2(n_139),
.B(n_431),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_435),
.A2(n_447),
.B(n_464),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_437),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_435),
.A2(n_464),
.B(n_446),
.Y(n_500)
);

OR2x6_ASAP7_75t_L g501 ( 
.A(n_473),
.B(n_437),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_482),
.A2(n_466),
.B(n_457),
.Y(n_502)
);

AOI21x1_ASAP7_75t_L g503 ( 
.A1(n_454),
.A2(n_449),
.B(n_477),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_438),
.B(n_432),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_444),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_451),
.A2(n_442),
.B(n_448),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_428),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_436),
.Y(n_508)
);

CKINVDCx11_ASAP7_75t_R g509 ( 
.A(n_475),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_436),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_459),
.Y(n_511)
);

OA21x2_ASAP7_75t_L g512 ( 
.A1(n_470),
.A2(n_455),
.B(n_459),
.Y(n_512)
);

OAI22x1_ASAP7_75t_L g513 ( 
.A1(n_438),
.A2(n_439),
.B1(n_478),
.B2(n_465),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_456),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_468),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_478),
.Y(n_516)
);

O2A1O1Ixp33_ASAP7_75t_L g517 ( 
.A1(n_476),
.A2(n_455),
.B(n_440),
.C(n_463),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_433),
.Y(n_518)
);

AO21x2_ASAP7_75t_L g519 ( 
.A1(n_445),
.A2(n_469),
.B(n_474),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_462),
.A2(n_453),
.B1(n_471),
.B2(n_472),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_479),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_461),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g523 ( 
.A1(n_441),
.A2(n_434),
.B(n_430),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_426),
.B(n_387),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_443),
.B(n_438),
.Y(n_525)
);

NAND2x1p5_ASAP7_75t_L g526 ( 
.A(n_452),
.B(n_395),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_452),
.Y(n_527)
);

BUFx2_ASAP7_75t_R g528 ( 
.A(n_516),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_509),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_507),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_492),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_494),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_495),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_524),
.A2(n_516),
.B1(n_509),
.B2(n_511),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_499),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_495),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_508),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_501),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_525),
.B(n_494),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_511),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_508),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_492),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_504),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_510),
.Y(n_544)
);

AO21x2_ASAP7_75t_L g545 ( 
.A1(n_500),
.A2(n_503),
.B(n_502),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_510),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_505),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_491),
.Y(n_548)
);

OA21x2_ASAP7_75t_L g549 ( 
.A1(n_500),
.A2(n_523),
.B(n_502),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_501),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_494),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_501),
.Y(n_552)
);

NAND2x1p5_ASAP7_75t_L g553 ( 
.A(n_521),
.B(n_489),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_486),
.B(n_527),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_518),
.B(n_484),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_526),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_526),
.Y(n_557)
);

OAI22xp33_ASAP7_75t_SL g558 ( 
.A1(n_490),
.A2(n_515),
.B1(n_514),
.B2(n_496),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_491),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_486),
.B(n_513),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_497),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_518),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_485),
.Y(n_563)
);

AO21x1_ASAP7_75t_L g564 ( 
.A1(n_517),
.A2(n_520),
.B(n_521),
.Y(n_564)
);

AOI21x1_ASAP7_75t_L g565 ( 
.A1(n_483),
.A2(n_498),
.B(n_522),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_497),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_488),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_535),
.B(n_506),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g569 ( 
.A(n_543),
.B(n_487),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_554),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_554),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_539),
.B(n_487),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_539),
.B(n_487),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_543),
.B(n_493),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_542),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_533),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_562),
.A2(n_493),
.B1(n_512),
.B2(n_519),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_551),
.B(n_512),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_533),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_555),
.B(n_512),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_555),
.B(n_521),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_555),
.B(n_522),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_551),
.B(n_489),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_551),
.B(n_489),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_553),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_542),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_541),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_528),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_553),
.Y(n_589)
);

AO22x1_ASAP7_75t_L g590 ( 
.A1(n_563),
.A2(n_489),
.B1(n_488),
.B2(n_519),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_531),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_529),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_541),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_532),
.B(n_523),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_553),
.Y(n_595)
);

BUFx2_ASAP7_75t_SL g596 ( 
.A(n_532),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_540),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_532),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_540),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_538),
.B(n_498),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_536),
.Y(n_601)
);

INVxp67_ASAP7_75t_SL g602 ( 
.A(n_531),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_536),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_547),
.B(n_530),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_558),
.A2(n_538),
.B1(n_552),
.B2(n_550),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_560),
.B(n_544),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_560),
.B(n_544),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_546),
.B(n_537),
.Y(n_608)
);

AO31x2_ASAP7_75t_L g609 ( 
.A1(n_564),
.A2(n_566),
.A3(n_567),
.B(n_548),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_559),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_565),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_565),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_568),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_570),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_604),
.B(n_556),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_587),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_605),
.A2(n_534),
.B1(n_537),
.B2(n_546),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_587),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_593),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_575),
.B(n_557),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_R g621 ( 
.A(n_592),
.B(n_529),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_593),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_606),
.B(n_567),
.Y(n_623)
);

OAI221xp5_ASAP7_75t_SL g624 ( 
.A1(n_577),
.A2(n_566),
.B1(n_548),
.B2(n_561),
.C(n_559),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_597),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_597),
.Y(n_626)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_580),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_599),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_586),
.B(n_564),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_586),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_586),
.B(n_545),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_599),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_591),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_588),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_602),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_570),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_571),
.B(n_549),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_581),
.A2(n_561),
.B1(n_545),
.B2(n_549),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_585),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_606),
.B(n_549),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_576),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_608),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_576),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_607),
.B(n_549),
.Y(n_644)
);

NOR2xp67_ASAP7_75t_L g645 ( 
.A(n_582),
.B(n_545),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_591),
.B(n_608),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_571),
.B(n_607),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_579),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_579),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_600),
.B(n_572),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_618),
.Y(n_651)
);

INVxp67_ASAP7_75t_SL g652 ( 
.A(n_629),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_613),
.B(n_591),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_616),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_630),
.B(n_600),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_650),
.B(n_594),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_618),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_630),
.B(n_595),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_650),
.B(n_594),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_614),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_623),
.B(n_595),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_627),
.B(n_598),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_647),
.B(n_609),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_635),
.B(n_598),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_640),
.B(n_572),
.Y(n_665)
);

NAND2x1p5_ASAP7_75t_L g666 ( 
.A(n_639),
.B(n_585),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_619),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_623),
.B(n_585),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_623),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_640),
.B(n_573),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_615),
.B(n_642),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_619),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_614),
.B(n_585),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_633),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_644),
.B(n_573),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_622),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_646),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_622),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_654),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_656),
.B(n_644),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_674),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_677),
.B(n_647),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_652),
.A2(n_617),
.B1(n_634),
.B2(n_645),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_651),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_653),
.B(n_660),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_669),
.B(n_636),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_671),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_657),
.Y(n_688)
);

INVxp33_ASAP7_75t_L g689 ( 
.A(n_661),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_664),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_663),
.B(n_636),
.Y(n_691)
);

OAI32xp33_ASAP7_75t_L g692 ( 
.A1(n_663),
.A2(n_620),
.A3(n_631),
.B1(n_632),
.B2(n_625),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_665),
.B(n_637),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_667),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_665),
.B(n_632),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_670),
.B(n_628),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_681),
.B(n_669),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_684),
.Y(n_698)
);

AOI222xp33_ASAP7_75t_L g699 ( 
.A1(n_692),
.A2(n_590),
.B1(n_675),
.B2(n_670),
.C1(n_654),
.C2(n_676),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_688),
.Y(n_700)
);

OAI22xp33_ASAP7_75t_SL g701 ( 
.A1(n_683),
.A2(n_687),
.B1(n_691),
.B2(n_693),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_694),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_691),
.B(n_675),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_696),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_696),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_695),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_695),
.Y(n_707)
);

AOI31xp33_ASAP7_75t_L g708 ( 
.A1(n_699),
.A2(n_690),
.A3(n_697),
.B(n_689),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_703),
.B(n_682),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_703),
.A2(n_669),
.B1(n_685),
.B2(n_661),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_698),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_701),
.A2(n_705),
.B1(n_704),
.B2(n_707),
.Y(n_712)
);

OAI21xp33_ASAP7_75t_L g713 ( 
.A1(n_708),
.A2(n_706),
.B(n_702),
.Y(n_713)
);

AOI221xp5_ASAP7_75t_L g714 ( 
.A1(n_712),
.A2(n_700),
.B1(n_624),
.B2(n_590),
.C(n_678),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_711),
.Y(n_715)
);

AOI21xp33_ASAP7_75t_L g716 ( 
.A1(n_710),
.A2(n_662),
.B(n_672),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_709),
.A2(n_655),
.B1(n_686),
.B2(n_680),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_715),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_714),
.A2(n_668),
.B1(n_661),
.B2(n_655),
.Y(n_719)
);

AOI211xp5_ASAP7_75t_L g720 ( 
.A1(n_713),
.A2(n_621),
.B(n_664),
.C(n_686),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_716),
.B(n_659),
.Y(n_721)
);

NOR2x1_ASAP7_75t_L g722 ( 
.A(n_718),
.B(n_717),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_719),
.A2(n_668),
.B1(n_655),
.B2(n_679),
.Y(n_723)
);

NOR3x1_ASAP7_75t_L g724 ( 
.A(n_720),
.B(n_637),
.C(n_574),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_722),
.B(n_721),
.C(n_638),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_724),
.B(n_723),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_722),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_722),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_727),
.B(n_659),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_728),
.Y(n_730)
);

NOR2x1p5_ASAP7_75t_L g731 ( 
.A(n_725),
.B(n_673),
.Y(n_731)
);

NAND4xp75_ASAP7_75t_L g732 ( 
.A(n_726),
.B(n_656),
.C(n_584),
.D(n_583),
.Y(n_732)
);

NOR2x1_ASAP7_75t_L g733 ( 
.A(n_727),
.B(n_673),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_727),
.B(n_673),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_727),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_730),
.B(n_668),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_735),
.Y(n_737)
);

OAI21xp5_ASAP7_75t_L g738 ( 
.A1(n_733),
.A2(n_666),
.B(n_658),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_732),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_729),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_731),
.Y(n_741)
);

NOR2x1_ASAP7_75t_L g742 ( 
.A(n_734),
.B(n_658),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_730),
.B(n_658),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_740),
.A2(n_666),
.B(n_611),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_739),
.A2(n_574),
.B1(n_583),
.B2(n_584),
.Y(n_745)
);

CKINVDCx20_ASAP7_75t_R g746 ( 
.A(n_740),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_741),
.A2(n_666),
.B1(n_616),
.B2(n_626),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_737),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_736),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_743),
.Y(n_750)
);

NAND3xp33_ASAP7_75t_L g751 ( 
.A(n_742),
.B(n_738),
.C(n_639),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_746),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_751),
.A2(n_626),
.B1(n_628),
.B2(n_639),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_748),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_749),
.A2(n_596),
.B1(n_610),
.B2(n_598),
.Y(n_755)
);

AO22x1_ASAP7_75t_L g756 ( 
.A1(n_750),
.A2(n_598),
.B1(n_578),
.B2(n_610),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_745),
.A2(n_596),
.B1(n_569),
.B2(n_578),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_SL g758 ( 
.A1(n_747),
.A2(n_569),
.B1(n_610),
.B2(n_611),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_744),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_752),
.Y(n_760)
);

NAND4xp75_ASAP7_75t_L g761 ( 
.A(n_754),
.B(n_611),
.C(n_612),
.D(n_649),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_759),
.A2(n_612),
.B(n_610),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_757),
.A2(n_612),
.B1(n_589),
.B2(n_595),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_755),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_758),
.A2(n_589),
.B1(n_595),
.B2(n_610),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_SL g766 ( 
.A1(n_760),
.A2(n_753),
.B1(n_756),
.B2(n_610),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_764),
.A2(n_589),
.B1(n_648),
.B2(n_643),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_762),
.A2(n_589),
.B(n_648),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_761),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_769),
.B(n_763),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_766),
.A2(n_765),
.B(n_643),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_770),
.A2(n_771),
.B(n_767),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_772),
.B(n_768),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_773),
.A2(n_641),
.B1(n_601),
.B2(n_603),
.Y(n_774)
);


endmodule