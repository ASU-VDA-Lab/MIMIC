module fake_jpeg_22791_n_50 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_50);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_50;

wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_40;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_4),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_29),
.B(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_26),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_23),
.B(n_27),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_28),
.B1(n_14),
.B2(n_5),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_1),
.B1(n_2),
.B2(n_26),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_38),
.B1(n_18),
.B2(n_19),
.Y(n_43)
);

NAND3xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.C(n_37),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_10),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_39),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_43),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_48),
.A2(n_36),
.B1(n_44),
.B2(n_21),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_20),
.Y(n_50)
);


endmodule