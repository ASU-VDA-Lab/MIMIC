module fake_jpeg_10715_n_125 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_125);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_7),
.B(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_21),
.A2(n_28),
.B1(n_18),
.B2(n_12),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_39),
.B1(n_43),
.B2(n_30),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_21),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_35),
.A2(n_21),
.B1(n_43),
.B2(n_11),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_36),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_2),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_4),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_48),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_18),
.A2(n_5),
.B1(n_11),
.B2(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_20),
.B(n_5),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_11),
.A2(n_27),
.B1(n_24),
.B2(n_16),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_13),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_29),
.Y(n_54)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_49),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_24),
.A2(n_27),
.B(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_22),
.B(n_14),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_23),
.B(n_11),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_54),
.B(n_60),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_52),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_49),
.B1(n_48),
.B2(n_32),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_33),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_64),
.B(n_65),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_37),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_74),
.C(n_51),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_52),
.B(n_56),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_58),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_29),
.B(n_37),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_55),
.B1(n_53),
.B2(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_80),
.B1(n_81),
.B2(n_87),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_73),
.Y(n_92)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_53),
.A2(n_67),
.B1(n_74),
.B2(n_51),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_69),
.B1(n_75),
.B2(n_68),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_88),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_86),
.B(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_72),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_57),
.C(n_85),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_72),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_93),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_75),
.C(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_97),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_99),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_76),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_78),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_96),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_95),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_86),
.B1(n_91),
.B2(n_81),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_105),
.B1(n_108),
.B2(n_93),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_89),
.B1(n_79),
.B2(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_113),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_110),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_115),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_107),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_104),
.C(n_106),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_122),
.A2(n_111),
.B1(n_117),
.B2(n_120),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_119),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_123),
.Y(n_125)
);


endmodule