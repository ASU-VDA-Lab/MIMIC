module fake_ariane_2142_n_2119 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2119);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2119;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_274;
wire n_1083;
wire n_337;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_2016;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_253;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_363;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_2012;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g215 ( 
.A(n_48),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_68),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_56),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_55),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_126),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_213),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_103),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_150),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_135),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_185),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_51),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_91),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_32),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_74),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_31),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_59),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_99),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_44),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_22),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_58),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_75),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_112),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_64),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_166),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_89),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_37),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_168),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_190),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_8),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_6),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_163),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_134),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_85),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_132),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_88),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_101),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_100),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_64),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_55),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_86),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_113),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_95),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_111),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_106),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_206),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_17),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_82),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_195),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_200),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_70),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_131),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_36),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_115),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_20),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_11),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_60),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_73),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_165),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_143),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_154),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_20),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_188),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_198),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_24),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_110),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_5),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_98),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_40),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_167),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_199),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_66),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_49),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_4),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_42),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_186),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_170),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_121),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_162),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_70),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_61),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_33),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_209),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_81),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_48),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_79),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_182),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_0),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_24),
.Y(n_305)
);

BUFx5_ASAP7_75t_L g306 ( 
.A(n_116),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_30),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_105),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_80),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_10),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_43),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_152),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_147),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_16),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_124),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_180),
.Y(n_316)
);

BUFx10_ASAP7_75t_L g317 ( 
.A(n_203),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_35),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_61),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_83),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_65),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_18),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_16),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_158),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_78),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_26),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_53),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_211),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_117),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_92),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_19),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_33),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_184),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_25),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_84),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_205),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_208),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_193),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_201),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_169),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_119),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_9),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_212),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_175),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_120),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_22),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_196),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_108),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_58),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_176),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_10),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_153),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_74),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_26),
.Y(n_354)
);

BUFx10_ASAP7_75t_L g355 ( 
.A(n_42),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_189),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_77),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_181),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_63),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_93),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_207),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_15),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_122),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_15),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_27),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_5),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_107),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_142),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_109),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_8),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_191),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_21),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_25),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_69),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_73),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_37),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_87),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_2),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_151),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_13),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_36),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_51),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_145),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_141),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_50),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_41),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_140),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_65),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_96),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_63),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_67),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_60),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_19),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_155),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_146),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_183),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_38),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_54),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_43),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_72),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_23),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_104),
.Y(n_402)
);

CKINVDCx14_ASAP7_75t_R g403 ( 
.A(n_128),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_90),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_54),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_149),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_59),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_17),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_50),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_171),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_187),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_97),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_30),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_164),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_179),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_192),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_125),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_44),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_39),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_3),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_18),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_23),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_194),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_133),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_220),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_220),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_242),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_258),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_222),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_222),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_274),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_361),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_402),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_229),
.Y(n_434)
);

INVxp33_ASAP7_75t_SL g435 ( 
.A(n_217),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_215),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_215),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_419),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_310),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_228),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_240),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_419),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_218),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_240),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_229),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_226),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_348),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_302),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_302),
.B(n_0),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_231),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_231),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_296),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_232),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_248),
.Y(n_454)
);

NOR2xp67_ASAP7_75t_L g455 ( 
.A(n_230),
.B(n_1),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_248),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_288),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_254),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_254),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_237),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_259),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_259),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_348),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_334),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_380),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_266),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_238),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_266),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_391),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_403),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_277),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_243),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_317),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_277),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_279),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_279),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_282),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_288),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_282),
.B(n_1),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_247),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_286),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_390),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_286),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_299),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_317),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_317),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_255),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_299),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_317),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_300),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_300),
.B(n_2),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_309),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_256),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_267),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_271),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_309),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_234),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_234),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_273),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_249),
.Y(n_500)
);

INVxp67_ASAP7_75t_SL g501 ( 
.A(n_390),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_316),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_316),
.B(n_3),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_278),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_324),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_249),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_358),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_324),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_281),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_325),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_283),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_325),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_290),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_358),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_297),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_269),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_328),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_269),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_269),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_310),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_244),
.B(n_4),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_304),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_310),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_328),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_305),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_392),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_329),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_310),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_307),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_311),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_R g531 ( 
.A(n_221),
.B(n_223),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_318),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_269),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_329),
.B(n_6),
.Y(n_534)
);

INVxp33_ASAP7_75t_L g535 ( 
.A(n_233),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_425),
.B(n_341),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_523),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_523),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_425),
.B(n_341),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_523),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_439),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_439),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_507),
.B(n_350),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_426),
.B(n_392),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_520),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_520),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_428),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_528),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_426),
.B(n_216),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_528),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_429),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_429),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_430),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_430),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_434),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_434),
.B(n_216),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_521),
.B(n_310),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_SL g558 ( 
.A(n_535),
.B(n_230),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_445),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_438),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_445),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_450),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_450),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_451),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_451),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_442),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_454),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_444),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_454),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_456),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_456),
.B(n_350),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_458),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_458),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_459),
.B(n_235),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_459),
.B(n_356),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_461),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_507),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_461),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_462),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_462),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_466),
.B(n_235),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_466),
.B(n_356),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_468),
.B(n_471),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_457),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_468),
.Y(n_585)
);

AND2x2_ASAP7_75t_SL g586 ( 
.A(n_449),
.B(n_219),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_471),
.B(n_360),
.Y(n_587)
);

AND2x6_ASAP7_75t_L g588 ( 
.A(n_474),
.B(n_219),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_474),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_475),
.B(n_360),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_475),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_476),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_476),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_477),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_477),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_481),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_481),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_483),
.B(n_379),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_432),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_483),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_443),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_484),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_484),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_488),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_488),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_490),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_490),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_492),
.B(n_364),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_492),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_496),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_496),
.B(n_379),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_502),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_531),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_502),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_505),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_505),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_440),
.B(n_319),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_508),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_508),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_441),
.B(n_416),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_510),
.B(n_416),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_448),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_510),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_573),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_537),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_573),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_586),
.A2(n_558),
.B1(n_620),
.B2(n_448),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_537),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_573),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_586),
.B(n_447),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_573),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_537),
.Y(n_632)
);

INVx5_ASAP7_75t_L g633 ( 
.A(n_573),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_613),
.B(n_463),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_573),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_613),
.B(n_435),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_573),
.Y(n_637)
);

AO22x2_ASAP7_75t_L g638 ( 
.A1(n_557),
.A2(n_469),
.B1(n_431),
.B2(n_512),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_586),
.B(n_512),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_622),
.Y(n_640)
);

NAND2xp33_ASAP7_75t_SL g641 ( 
.A(n_601),
.B(n_446),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_577),
.B(n_453),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_573),
.Y(n_643)
);

AOI21x1_ASAP7_75t_L g644 ( 
.A1(n_557),
.A2(n_524),
.B(n_517),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_586),
.B(n_517),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_596),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_583),
.B(n_478),
.Y(n_647)
);

AND2x6_ASAP7_75t_L g648 ( 
.A(n_583),
.B(n_239),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_551),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_537),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_596),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_622),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_547),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_558),
.A2(n_479),
.B1(n_503),
.B2(n_491),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_547),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_577),
.B(n_460),
.Y(n_656)
);

OR2x6_ASAP7_75t_L g657 ( 
.A(n_601),
.B(n_455),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_577),
.B(n_524),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_599),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_537),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_596),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_596),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_596),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_601),
.B(n_467),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_596),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_622),
.B(n_482),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_596),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_577),
.Y(n_668)
);

INVxp33_ASAP7_75t_SL g669 ( 
.A(n_599),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_596),
.Y(n_670)
);

INVx5_ASAP7_75t_L g671 ( 
.A(n_551),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_620),
.A2(n_534),
.B1(n_527),
.B2(n_485),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_548),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_622),
.B(n_472),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_551),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_548),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_551),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_568),
.Y(n_678)
);

INVx4_ASAP7_75t_SL g679 ( 
.A(n_588),
.Y(n_679)
);

AND2x6_ASAP7_75t_L g680 ( 
.A(n_583),
.B(n_239),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_589),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_551),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_622),
.B(n_501),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_551),
.Y(n_684)
);

BUFx4f_ASAP7_75t_L g685 ( 
.A(n_551),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_552),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_622),
.B(n_480),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_552),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_552),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_552),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_608),
.A2(n_527),
.B1(n_486),
.B2(n_489),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_622),
.B(n_487),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_560),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_589),
.B(n_493),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_622),
.B(n_494),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_553),
.B(n_495),
.Y(n_696)
);

AND2x6_ASAP7_75t_L g697 ( 
.A(n_555),
.B(n_340),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_568),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_560),
.B(n_499),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_566),
.B(n_504),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_544),
.B(n_436),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_552),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_552),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_552),
.Y(n_704)
);

INVx5_ASAP7_75t_L g705 ( 
.A(n_565),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_566),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_549),
.B(n_526),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_553),
.B(n_509),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_565),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_589),
.B(n_511),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_565),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_589),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_549),
.B(n_437),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_565),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_565),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_608),
.A2(n_473),
.B1(n_498),
.B2(n_497),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_589),
.B(n_513),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_565),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_544),
.B(n_500),
.Y(n_719)
);

AND3x2_ASAP7_75t_L g720 ( 
.A(n_584),
.B(n_400),
.C(n_298),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_594),
.B(n_515),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_565),
.Y(n_722)
);

AO22x2_ASAP7_75t_L g723 ( 
.A1(n_617),
.A2(n_353),
.B1(n_418),
.B2(n_397),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_594),
.B(n_522),
.Y(n_724)
);

INVx5_ASAP7_75t_L g725 ( 
.A(n_578),
.Y(n_725)
);

OR2x6_ASAP7_75t_L g726 ( 
.A(n_549),
.B(n_364),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_578),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_578),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_578),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_578),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_617),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_578),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_594),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_556),
.B(n_525),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_594),
.B(n_529),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_578),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_604),
.Y(n_737)
);

CKINVDCx6p67_ASAP7_75t_R g738 ( 
.A(n_584),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_604),
.Y(n_739)
);

INVx4_ASAP7_75t_L g740 ( 
.A(n_604),
.Y(n_740)
);

AO22x2_ASAP7_75t_L g741 ( 
.A1(n_617),
.A2(n_377),
.B1(n_315),
.B2(n_236),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_594),
.B(n_530),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_604),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_604),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_554),
.B(n_532),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_604),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_544),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_604),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_554),
.B(n_470),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_606),
.Y(n_750)
);

OAI22xp33_ASAP7_75t_L g751 ( 
.A1(n_536),
.A2(n_571),
.B1(n_575),
.B2(n_539),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_606),
.Y(n_752)
);

INVx4_ASAP7_75t_L g753 ( 
.A(n_606),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_606),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_556),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_543),
.A2(n_322),
.B1(n_327),
.B2(n_321),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_606),
.Y(n_757)
);

OR2x6_ASAP7_75t_L g758 ( 
.A(n_556),
.B(n_378),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_605),
.B(n_506),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_606),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_606),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_614),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_605),
.B(n_514),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_614),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_605),
.B(n_607),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_614),
.Y(n_766)
);

INVx5_ASAP7_75t_L g767 ( 
.A(n_614),
.Y(n_767)
);

OR2x2_ASAP7_75t_L g768 ( 
.A(n_536),
.B(n_233),
.Y(n_768)
);

NAND3xp33_ASAP7_75t_L g769 ( 
.A(n_543),
.B(n_349),
.C(n_331),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_614),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_614),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_605),
.B(n_355),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_614),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_538),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_605),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_608),
.A2(n_373),
.B1(n_351),
.B2(n_354),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_630),
.B(n_607),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_678),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_696),
.B(n_607),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_673),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_678),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_774),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_751),
.B(n_607),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_698),
.B(n_516),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_673),
.Y(n_785)
);

AO221x1_ASAP7_75t_L g786 ( 
.A1(n_741),
.A2(n_399),
.B1(n_291),
.B2(n_285),
.C(n_301),
.Y(n_786)
);

OAI22xp33_ASAP7_75t_SL g787 ( 
.A1(n_657),
.A2(n_571),
.B1(n_575),
.B2(n_539),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_708),
.B(n_607),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_774),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_763),
.B(n_559),
.Y(n_790)
);

INVx8_ASAP7_75t_L g791 ( 
.A(n_648),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_745),
.B(n_642),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_676),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_656),
.B(n_559),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_775),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_648),
.A2(n_608),
.B1(n_561),
.B2(n_562),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_775),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_648),
.A2(n_623),
.B1(n_564),
.B2(n_567),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_694),
.B(n_563),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_676),
.Y(n_800)
);

NAND2xp33_ASAP7_75t_L g801 ( 
.A(n_648),
.B(n_563),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_639),
.B(n_564),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_657),
.B(n_574),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_775),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_625),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_645),
.B(n_627),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_681),
.B(n_567),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_717),
.A2(n_724),
.B(n_721),
.Y(n_808)
);

INVxp67_ASAP7_75t_SL g809 ( 
.A(n_668),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_648),
.A2(n_608),
.B1(n_561),
.B2(n_562),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_742),
.B(n_569),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_625),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_698),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_681),
.B(n_570),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_647),
.B(n_574),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_693),
.B(n_518),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_759),
.B(n_710),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_755),
.B(n_647),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_706),
.B(n_519),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_628),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_SL g821 ( 
.A1(n_731),
.A2(n_464),
.B1(n_465),
.B2(n_452),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_628),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_712),
.B(n_570),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_632),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_768),
.B(n_572),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_768),
.B(n_572),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_632),
.Y(n_827)
);

NOR2x1p5_ASAP7_75t_L g828 ( 
.A(n_655),
.B(n_582),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_712),
.B(n_576),
.Y(n_829)
);

OAI22xp33_ASAP7_75t_L g830 ( 
.A1(n_756),
.A2(n_587),
.B1(n_590),
.B2(n_582),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_650),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_650),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_734),
.B(n_576),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_660),
.Y(n_834)
);

AND2x2_ASAP7_75t_SL g835 ( 
.A(n_654),
.B(n_587),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_668),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_660),
.Y(n_837)
);

INVx4_ASAP7_75t_L g838 ( 
.A(n_648),
.Y(n_838)
);

NAND2xp33_ASAP7_75t_L g839 ( 
.A(n_648),
.B(n_580),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_661),
.Y(n_840)
);

OAI21xp33_ASAP7_75t_L g841 ( 
.A1(n_756),
.A2(n_585),
.B(n_580),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_733),
.Y(n_842)
);

NOR2xp67_ASAP7_75t_L g843 ( 
.A(n_655),
.B(n_659),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_659),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_735),
.B(n_585),
.Y(n_845)
);

INVx8_ASAP7_75t_L g846 ( 
.A(n_680),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_734),
.B(n_636),
.Y(n_847)
);

NAND2xp33_ASAP7_75t_L g848 ( 
.A(n_680),
.B(n_686),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_733),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_726),
.B(n_574),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_661),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_663),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_747),
.A2(n_623),
.B(n_591),
.C(n_597),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_SL g854 ( 
.A(n_653),
.B(n_427),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_701),
.B(n_591),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_SL g856 ( 
.A(n_669),
.B(n_433),
.Y(n_856)
);

BUFx6f_ASAP7_75t_SL g857 ( 
.A(n_719),
.Y(n_857)
);

NAND2x1p5_ASAP7_75t_L g858 ( 
.A(n_666),
.B(n_555),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_701),
.B(n_595),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_701),
.B(n_595),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_663),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_772),
.B(n_597),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_765),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_726),
.B(n_600),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_686),
.B(n_600),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_658),
.Y(n_866)
);

INVxp67_ASAP7_75t_L g867 ( 
.A(n_749),
.Y(n_867)
);

BUFx6f_ASAP7_75t_SL g868 ( 
.A(n_719),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_667),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_680),
.A2(n_615),
.B1(n_618),
.B2(n_612),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_686),
.B(n_612),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_726),
.B(n_581),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_644),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_686),
.B(n_729),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_701),
.B(n_672),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_726),
.B(n_615),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_667),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_758),
.B(n_581),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_713),
.B(n_618),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_686),
.B(n_619),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_713),
.B(n_619),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_666),
.B(n_555),
.Y(n_882)
);

OR2x6_ASAP7_75t_L g883 ( 
.A(n_657),
.B(n_581),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_644),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_680),
.A2(n_562),
.B1(n_579),
.B2(n_561),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_675),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_690),
.Y(n_887)
);

NAND3xp33_ASAP7_75t_L g888 ( 
.A(n_634),
.B(n_598),
.C(n_590),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_675),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_703),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_703),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_666),
.B(n_579),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_677),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_722),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_722),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_719),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_677),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_683),
.B(n_579),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_683),
.B(n_592),
.Y(n_899)
);

OR2x6_ASAP7_75t_L g900 ( 
.A(n_657),
.B(n_598),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_683),
.B(n_592),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_729),
.B(n_592),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_728),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_680),
.B(n_593),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_680),
.B(n_593),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_707),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_728),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_688),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_729),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_664),
.A2(n_621),
.B(n_611),
.C(n_616),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_680),
.B(n_593),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_758),
.B(n_602),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_707),
.B(n_533),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_729),
.B(n_602),
.Y(n_914)
);

INVxp67_ASAP7_75t_L g915 ( 
.A(n_641),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_688),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_638),
.B(n_758),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_729),
.B(n_602),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_699),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_758),
.B(n_769),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_638),
.B(n_603),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_685),
.B(n_649),
.Y(n_922)
);

INVx8_ASAP7_75t_L g923 ( 
.A(n_697),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_638),
.B(n_603),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_674),
.B(n_609),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_689),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_692),
.B(n_609),
.Y(n_927)
);

AO22x2_ASAP7_75t_L g928 ( 
.A1(n_741),
.A2(n_374),
.B1(n_246),
.B2(n_263),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_689),
.Y(n_929)
);

NAND2xp33_ASAP7_75t_L g930 ( 
.A(n_624),
.B(n_609),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_679),
.B(n_610),
.Y(n_931)
);

INVxp67_ASAP7_75t_L g932 ( 
.A(n_700),
.Y(n_932)
);

NAND2xp33_ASAP7_75t_L g933 ( 
.A(n_624),
.B(n_610),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_732),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_685),
.B(n_610),
.Y(n_935)
);

NAND3xp33_ASAP7_75t_L g936 ( 
.A(n_776),
.B(n_621),
.C(n_611),
.Y(n_936)
);

NAND2xp33_ASAP7_75t_L g937 ( 
.A(n_629),
.B(n_616),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_629),
.A2(n_616),
.B(n_540),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_732),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_685),
.B(n_315),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_741),
.A2(n_588),
.B1(n_378),
.B2(n_405),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_739),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_776),
.B(n_359),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_649),
.Y(n_944)
);

NAND2xp33_ASAP7_75t_L g945 ( 
.A(n_792),
.B(n_682),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_943),
.A2(n_684),
.B(n_702),
.C(n_682),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_808),
.A2(n_709),
.B(n_704),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_838),
.B(n_835),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_925),
.A2(n_709),
.B(n_704),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_927),
.A2(n_715),
.B(n_711),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_847),
.B(n_867),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_777),
.A2(n_715),
.B(n_711),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_813),
.B(n_669),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_790),
.B(n_691),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_909),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_922),
.A2(n_730),
.B(n_718),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_844),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_794),
.A2(n_730),
.B(n_718),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_790),
.B(n_738),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_778),
.Y(n_960)
);

CKINVDCx8_ASAP7_75t_R g961 ( 
.A(n_803),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_777),
.A2(n_743),
.B(n_736),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_874),
.A2(n_743),
.B(n_736),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_782),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_830),
.B(n_738),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_830),
.B(n_716),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_835),
.B(n_682),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_815),
.B(n_679),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_874),
.A2(n_762),
.B(n_752),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_779),
.A2(n_762),
.B(n_752),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_789),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_805),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_838),
.B(n_649),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_780),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_788),
.A2(n_766),
.B(n_764),
.Y(n_975)
);

OR2x6_ASAP7_75t_L g976 ( 
.A(n_803),
.B(n_741),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_818),
.B(n_684),
.Y(n_977)
);

NOR3xp33_ASAP7_75t_L g978 ( 
.A(n_943),
.B(n_246),
.C(n_236),
.Y(n_978)
);

AOI21x1_ASAP7_75t_L g979 ( 
.A1(n_922),
.A2(n_766),
.B(n_764),
.Y(n_979)
);

INVx4_ASAP7_75t_L g980 ( 
.A(n_791),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_780),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_781),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_802),
.A2(n_773),
.B(n_770),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_815),
.B(n_679),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_802),
.A2(n_773),
.B(n_770),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_783),
.A2(n_811),
.B(n_799),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_863),
.A2(n_635),
.B(n_631),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_896),
.B(n_740),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_822),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_799),
.A2(n_702),
.B(n_714),
.C(n_684),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_783),
.A2(n_635),
.B(n_631),
.Y(n_991)
);

BUFx4f_ASAP7_75t_L g992 ( 
.A(n_803),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_833),
.B(n_702),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_906),
.B(n_740),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_787),
.B(n_740),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_825),
.B(n_714),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_827),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_785),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_826),
.B(n_714),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_811),
.A2(n_651),
.B(n_637),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_935),
.A2(n_651),
.B(n_637),
.Y(n_1001)
);

OAI21xp33_ASAP7_75t_L g1002 ( 
.A1(n_845),
.A2(n_365),
.B(n_362),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_938),
.A2(n_670),
.B(n_662),
.Y(n_1003)
);

NOR2xp67_ASAP7_75t_L g1004 ( 
.A(n_843),
.B(n_731),
.Y(n_1004)
);

AO21x1_ASAP7_75t_L g1005 ( 
.A1(n_806),
.A2(n_753),
.B(n_670),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_935),
.A2(n_662),
.B(n_687),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_888),
.B(n_753),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_902),
.A2(n_695),
.B(n_739),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_785),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_831),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_821),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_796),
.B(n_753),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_795),
.A2(n_746),
.B(n_744),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_875),
.B(n_727),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_797),
.A2(n_746),
.B(n_744),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_845),
.A2(n_737),
.B(n_727),
.C(n_748),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_879),
.B(n_727),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_902),
.A2(n_750),
.B(n_748),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_837),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_816),
.B(n_723),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_881),
.B(n_737),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_819),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_855),
.B(n_737),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_909),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_909),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_796),
.B(n_671),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_864),
.A2(n_754),
.B(n_757),
.C(n_750),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_914),
.A2(n_757),
.B(n_754),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_859),
.B(n_626),
.Y(n_1029)
);

BUFx12f_ASAP7_75t_L g1030 ( 
.A(n_784),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_914),
.A2(n_761),
.B(n_760),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_918),
.A2(n_820),
.B(n_812),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_918),
.A2(n_824),
.B(n_820),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_824),
.A2(n_761),
.B(n_760),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_930),
.A2(n_771),
.B(n_643),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_860),
.B(n_626),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_909),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_933),
.A2(n_937),
.B(n_871),
.Y(n_1038)
);

CKINVDCx20_ASAP7_75t_R g1039 ( 
.A(n_913),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_850),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_864),
.B(n_626),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_919),
.B(n_643),
.Y(n_1042)
);

OAI21xp33_ASAP7_75t_L g1043 ( 
.A1(n_856),
.A2(n_370),
.B(n_366),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_876),
.B(n_643),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_804),
.A2(n_885),
.B(n_936),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_876),
.B(n_646),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_810),
.B(n_817),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_865),
.A2(n_771),
.B(n_665),
.Y(n_1048)
);

NAND2xp33_ASAP7_75t_L g1049 ( 
.A(n_791),
.B(n_646),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_912),
.B(n_646),
.Y(n_1050)
);

NOR2xp67_ASAP7_75t_L g1051 ( 
.A(n_915),
.B(n_538),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_912),
.B(n_665),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_865),
.A2(n_665),
.B(n_652),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_871),
.A2(n_652),
.B(n_640),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_880),
.A2(n_834),
.B(n_832),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_807),
.A2(n_640),
.B(n_633),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_807),
.A2(n_823),
.B(n_814),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_853),
.A2(n_263),
.B(n_272),
.C(n_285),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_880),
.A2(n_633),
.B(n_671),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_814),
.A2(n_633),
.B(n_671),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_817),
.B(n_540),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_932),
.B(n_720),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_866),
.B(n_671),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_850),
.B(n_671),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_810),
.A2(n_767),
.B1(n_725),
.B2(n_705),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_887),
.Y(n_1066)
);

NAND2x1p5_ASAP7_75t_L g1067 ( 
.A(n_931),
.B(n_872),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_931),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_872),
.B(n_671),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_920),
.B(n_767),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_878),
.B(n_705),
.Y(n_1071)
);

CKINVDCx10_ASAP7_75t_R g1072 ( 
.A(n_857),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_862),
.A2(n_910),
.B(n_841),
.C(n_920),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_798),
.B(n_767),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_823),
.A2(n_272),
.B(n_289),
.C(n_291),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_829),
.A2(n_633),
.B(n_705),
.Y(n_1076)
);

OAI321xp33_ASAP7_75t_L g1077 ( 
.A1(n_941),
.A2(n_342),
.A3(n_289),
.B1(n_301),
.B2(n_314),
.C(n_323),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_887),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_878),
.B(n_705),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_891),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_849),
.B(n_767),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_862),
.B(n_705),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_857),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_870),
.A2(n_314),
.B(n_323),
.C(n_326),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_882),
.B(n_892),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_886),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_889),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_829),
.A2(n_633),
.B(n_705),
.Y(n_1088)
);

AOI21x1_ASAP7_75t_L g1089 ( 
.A1(n_904),
.A2(n_542),
.B(n_541),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_851),
.A2(n_633),
.B(n_725),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_851),
.A2(n_767),
.B(n_725),
.Y(n_1091)
);

OAI21xp33_ASAP7_75t_L g1092 ( 
.A1(n_854),
.A2(n_375),
.B(n_372),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_898),
.B(n_725),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_917),
.B(n_767),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_852),
.A2(n_725),
.B(n_225),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_791),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_944),
.B(n_725),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_852),
.A2(n_227),
.B(n_224),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_899),
.B(n_697),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_883),
.B(n_376),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_842),
.A2(n_409),
.B1(n_388),
.B2(n_386),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_883),
.B(n_382),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_901),
.B(n_697),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_842),
.B(n_697),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_846),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_858),
.B(n_679),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_883),
.B(n_723),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_893),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_891),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_897),
.A2(n_697),
.B(n_588),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_944),
.B(n_377),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_908),
.A2(n_697),
.B(n_588),
.Y(n_1112)
);

AOI21xp33_ASAP7_75t_L g1113 ( 
.A1(n_905),
.A2(n_723),
.B(n_398),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_900),
.B(n_393),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_900),
.B(n_326),
.Y(n_1115)
);

INVx4_ASAP7_75t_L g1116 ( 
.A(n_846),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_861),
.A2(n_245),
.B(n_241),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_916),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_801),
.A2(n_421),
.B(n_385),
.C(n_332),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_858),
.B(n_809),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_926),
.A2(n_346),
.B(n_421),
.C(n_332),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_929),
.A2(n_346),
.B(n_413),
.C(n_374),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_900),
.B(n_697),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_941),
.B(n_342),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_861),
.A2(n_251),
.B(n_250),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_895),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_895),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_903),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_SL g1129 ( 
.A(n_868),
.B(n_355),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_836),
.B(n_381),
.Y(n_1130)
);

NAND2x1p5_ASAP7_75t_L g1131 ( 
.A(n_1068),
.B(n_836),
.Y(n_1131)
);

NAND3xp33_ASAP7_75t_SL g1132 ( 
.A(n_978),
.B(n_959),
.C(n_965),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_951),
.B(n_828),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_986),
.A2(n_848),
.B(n_839),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_953),
.B(n_944),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_945),
.A2(n_846),
.B(n_940),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1086),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_953),
.B(n_944),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1000),
.A2(n_940),
.B(n_911),
.Y(n_1139)
);

NAND2x1p5_ASAP7_75t_L g1140 ( 
.A(n_1068),
.B(n_903),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_978),
.A2(n_928),
.B1(n_786),
.B2(n_723),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_1022),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1049),
.A2(n_877),
.B(n_907),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_951),
.A2(n_877),
.B1(n_928),
.B2(n_939),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_952),
.A2(n_939),
.B(n_907),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_954),
.B(n_928),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1087),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1039),
.A2(n_868),
.B1(n_923),
.B2(n_401),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_974),
.Y(n_1149)
);

BUFx2_ASAP7_75t_L g1150 ( 
.A(n_1030),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_966),
.B(n_921),
.Y(n_1151)
);

O2A1O1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1073),
.A2(n_413),
.B(n_385),
.C(n_381),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1047),
.B(n_924),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1108),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_948),
.A2(n_923),
.B1(n_420),
.B2(n_408),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1007),
.A2(n_923),
.B(n_934),
.C(n_942),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_960),
.Y(n_1157)
);

INVx1_ASAP7_75t_SL g1158 ( 
.A(n_960),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1040),
.B(n_793),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_1043),
.B(n_890),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1118),
.Y(n_1161)
);

NOR2xp67_ASAP7_75t_SL g1162 ( 
.A(n_957),
.B(n_407),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_R g1163 ( 
.A(n_1072),
.B(n_873),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_982),
.B(n_894),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_982),
.B(n_840),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_1096),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_994),
.A2(n_869),
.B1(n_884),
.B2(n_800),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_967),
.A2(n_1052),
.B(n_1050),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_1083),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1040),
.B(n_422),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_962),
.A2(n_340),
.B(n_303),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_994),
.B(n_405),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_1096),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_964),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_948),
.B(n_1067),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1067),
.B(n_355),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_992),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1082),
.A2(n_294),
.B(n_253),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_976),
.A2(n_355),
.B1(n_588),
.B2(n_399),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1041),
.A2(n_399),
.B1(n_352),
.B2(n_347),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1042),
.B(n_588),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_976),
.A2(n_588),
.B1(n_399),
.B2(n_542),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_1011),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_968),
.B(n_541),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_1107),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_976),
.B(n_545),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_971),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1100),
.B(n_252),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_981),
.Y(n_1189)
);

NAND2xp33_ASAP7_75t_SL g1190 ( 
.A(n_980),
.B(n_399),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_972),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_SL g1192 ( 
.A1(n_990),
.A2(n_545),
.B(n_550),
.C(n_11),
.Y(n_1192)
);

NAND3xp33_ASAP7_75t_L g1193 ( 
.A(n_1002),
.B(n_550),
.C(n_546),
.Y(n_1193)
);

O2A1O1Ixp5_ASAP7_75t_L g1194 ( 
.A1(n_1005),
.A2(n_588),
.B(n_546),
.C(n_306),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1044),
.A2(n_406),
.B1(n_337),
.B2(n_336),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1058),
.A2(n_7),
.B(n_9),
.C(n_12),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1046),
.A2(n_410),
.B1(n_333),
.B2(n_330),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_998),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1007),
.A2(n_546),
.B(n_343),
.C(n_424),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1038),
.A2(n_344),
.B(n_260),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1096),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1100),
.B(n_257),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_947),
.A2(n_357),
.B(n_262),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_991),
.A2(n_363),
.B(n_264),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1096),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_989),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_SL g1207 ( 
.A1(n_1045),
.A2(n_588),
.B(n_12),
.C(n_13),
.Y(n_1207)
);

INVx4_ASAP7_75t_L g1208 ( 
.A(n_1105),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1042),
.B(n_588),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1085),
.B(n_7),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_970),
.A2(n_345),
.B(n_423),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1062),
.A2(n_338),
.B1(n_417),
.B2(n_415),
.Y(n_1212)
);

AOI22x1_ASAP7_75t_L g1213 ( 
.A1(n_958),
.A2(n_975),
.B1(n_1053),
.B2(n_950),
.Y(n_1213)
);

CKINVDCx8_ASAP7_75t_R g1214 ( 
.A(n_1115),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1105),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_997),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_968),
.Y(n_1217)
);

OR2x2_ASAP7_75t_L g1218 ( 
.A(n_1020),
.B(n_546),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_949),
.A2(n_339),
.B(n_414),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_996),
.A2(n_335),
.B1(n_412),
.B2(n_411),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_992),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1004),
.B(n_261),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1115),
.B(n_14),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1105),
.Y(n_1224)
);

AOI21x1_ASAP7_75t_L g1225 ( 
.A1(n_995),
.A2(n_546),
.B(n_270),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_SL g1226 ( 
.A1(n_1081),
.A2(n_14),
.B(n_21),
.C(n_27),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1102),
.B(n_265),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1009),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1061),
.B(n_28),
.Y(n_1229)
);

OA22x2_ASAP7_75t_L g1230 ( 
.A1(n_1092),
.A2(n_404),
.B1(n_275),
.B2(n_276),
.Y(n_1230)
);

O2A1O1Ixp5_ASAP7_75t_L g1231 ( 
.A1(n_995),
.A2(n_1111),
.B(n_946),
.C(n_1016),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1121),
.A2(n_1122),
.B(n_1130),
.C(n_1101),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_999),
.A2(n_367),
.B1(n_396),
.B2(n_395),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_987),
.A2(n_313),
.B(n_394),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1006),
.A2(n_1008),
.B(n_1035),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1010),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1014),
.A2(n_546),
.B(n_389),
.C(n_387),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1084),
.A2(n_28),
.B(n_29),
.C(n_31),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1124),
.B(n_29),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_984),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1019),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_984),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1102),
.B(n_32),
.Y(n_1243)
);

NAND3xp33_ASAP7_75t_SL g1244 ( 
.A(n_1114),
.B(n_268),
.C(n_280),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1062),
.Y(n_1245)
);

NAND3xp33_ASAP7_75t_L g1246 ( 
.A(n_988),
.B(n_546),
.C(n_384),
.Y(n_1246)
);

INVxp67_ASAP7_75t_SL g1247 ( 
.A(n_955),
.Y(n_1247)
);

O2A1O1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1119),
.A2(n_34),
.B(n_35),
.C(n_38),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1014),
.B(n_34),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1001),
.A2(n_312),
.B(n_383),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1003),
.A2(n_308),
.B(n_371),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1063),
.A2(n_295),
.B(n_369),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1129),
.B(n_293),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1113),
.A2(n_546),
.B1(n_270),
.B2(n_306),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1114),
.B(n_368),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_963),
.A2(n_969),
.B(n_983),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_961),
.B(n_320),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1064),
.B(n_284),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_988),
.B(n_39),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_985),
.A2(n_287),
.B(n_292),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1017),
.B(n_40),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1077),
.A2(n_306),
.B1(n_270),
.B2(n_46),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1105),
.B(n_306),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1120),
.B(n_306),
.Y(n_1264)
);

AND2x6_ASAP7_75t_L g1265 ( 
.A(n_955),
.B(n_306),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1012),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1069),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_993),
.A2(n_127),
.B(n_214),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1051),
.B(n_41),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1018),
.A2(n_123),
.B(n_204),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1070),
.B(n_306),
.Y(n_1271)
);

NOR2xp67_ASAP7_75t_L g1272 ( 
.A(n_980),
.B(n_1116),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1021),
.B(n_45),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1028),
.A2(n_118),
.B(n_197),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1071),
.B(n_45),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1031),
.A2(n_1090),
.B(n_1048),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1070),
.A2(n_306),
.B(n_270),
.C(n_49),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1023),
.A2(n_46),
.B1(n_47),
.B2(n_52),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_977),
.B(n_47),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1079),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_955),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1116),
.B(n_306),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1024),
.B(n_270),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1024),
.Y(n_1284)
);

A2O1A1Ixp33_ASAP7_75t_SL g1285 ( 
.A1(n_1081),
.A2(n_52),
.B(n_53),
.C(n_56),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1012),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_1123),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1029),
.A2(n_57),
.B1(n_62),
.B2(n_66),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1134),
.A2(n_1074),
.B(n_1097),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1183),
.B(n_1066),
.Y(n_1290)
);

OAI22x1_ASAP7_75t_L g1291 ( 
.A1(n_1188),
.A2(n_1111),
.B1(n_1094),
.B2(n_1026),
.Y(n_1291)
);

AOI211x1_ASAP7_75t_L g1292 ( 
.A1(n_1278),
.A2(n_1057),
.B(n_1036),
.C(n_1110),
.Y(n_1292)
);

OA21x2_ASAP7_75t_L g1293 ( 
.A1(n_1235),
.A2(n_1027),
.B(n_1015),
.Y(n_1293)
);

NAND3x1_ASAP7_75t_L g1294 ( 
.A(n_1243),
.B(n_1094),
.C(n_1112),
.Y(n_1294)
);

INVx4_ASAP7_75t_L g1295 ( 
.A(n_1169),
.Y(n_1295)
);

NAND3xp33_ASAP7_75t_SL g1296 ( 
.A(n_1202),
.B(n_1075),
.C(n_1098),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1157),
.B(n_1128),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1150),
.Y(n_1298)
);

AOI211x1_ASAP7_75t_L g1299 ( 
.A1(n_1288),
.A2(n_1013),
.B(n_1125),
.C(n_1117),
.Y(n_1299)
);

BUFx10_ASAP7_75t_L g1300 ( 
.A(n_1170),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1276),
.A2(n_956),
.B(n_979),
.Y(n_1301)
);

AOI221x1_ASAP7_75t_L g1302 ( 
.A1(n_1277),
.A2(n_1032),
.B1(n_1033),
.B2(n_1055),
.C(n_1034),
.Y(n_1302)
);

BUFx4f_ASAP7_75t_SL g1303 ( 
.A(n_1158),
.Y(n_1303)
);

CKINVDCx11_ASAP7_75t_R g1304 ( 
.A(n_1214),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1256),
.A2(n_1074),
.B(n_1097),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1231),
.A2(n_1099),
.B(n_1103),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1136),
.A2(n_973),
.B(n_1091),
.Y(n_1307)
);

CKINVDCx16_ASAP7_75t_R g1308 ( 
.A(n_1163),
.Y(n_1308)
);

AO32x2_ASAP7_75t_L g1309 ( 
.A1(n_1144),
.A2(n_1065),
.A3(n_1089),
.B1(n_1109),
.B2(n_1127),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1227),
.A2(n_1026),
.B(n_1056),
.Y(n_1310)
);

AO32x2_ASAP7_75t_L g1311 ( 
.A1(n_1167),
.A2(n_1126),
.A3(n_1078),
.B1(n_1080),
.B2(n_1037),
.Y(n_1311)
);

OR2x6_ASAP7_75t_L g1312 ( 
.A(n_1177),
.B(n_1221),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1139),
.A2(n_973),
.B(n_1093),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1245),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1242),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1149),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1217),
.B(n_1024),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1133),
.B(n_1037),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1185),
.B(n_1037),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1190),
.A2(n_1024),
.B(n_1025),
.Y(n_1320)
);

AO31x2_ASAP7_75t_L g1321 ( 
.A1(n_1145),
.A2(n_1104),
.A3(n_1095),
.B(n_1088),
.Y(n_1321)
);

AO31x2_ASAP7_75t_L g1322 ( 
.A1(n_1156),
.A2(n_1076),
.A3(n_1059),
.B(n_1054),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1255),
.B(n_1037),
.Y(n_1323)
);

O2A1O1Ixp33_ASAP7_75t_SL g1324 ( 
.A1(n_1259),
.A2(n_1106),
.B(n_1060),
.C(n_1025),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1147),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1132),
.B(n_1025),
.Y(n_1326)
);

NAND2xp33_ASAP7_75t_L g1327 ( 
.A(n_1249),
.B(n_1025),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1143),
.A2(n_137),
.B(n_178),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1165),
.B(n_1164),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1217),
.B(n_136),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1213),
.A2(n_130),
.B(n_177),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1225),
.A2(n_270),
.B(n_129),
.Y(n_1332)
);

AO31x2_ASAP7_75t_L g1333 ( 
.A1(n_1151),
.A2(n_270),
.A3(n_138),
.B(n_139),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_SL g1334 ( 
.A(n_1132),
.B(n_270),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1240),
.B(n_1146),
.Y(n_1335)
);

NAND3x1_ASAP7_75t_L g1336 ( 
.A(n_1148),
.B(n_57),
.C(n_62),
.Y(n_1336)
);

NAND3xp33_ASAP7_75t_L g1337 ( 
.A(n_1152),
.B(n_67),
.C(n_68),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1154),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1232),
.A2(n_1171),
.B(n_1275),
.C(n_1229),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1161),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1240),
.B(n_69),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1189),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1174),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1168),
.A2(n_148),
.B(n_173),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_SL g1345 ( 
.A1(n_1210),
.A2(n_144),
.B(n_172),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1231),
.A2(n_114),
.B(n_161),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1187),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1184),
.B(n_102),
.Y(n_1348)
);

AOI221x1_ASAP7_75t_L g1349 ( 
.A1(n_1199),
.A2(n_270),
.B1(n_72),
.B2(n_75),
.C(n_76),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1281),
.Y(n_1350)
);

NOR2xp67_ASAP7_75t_SL g1351 ( 
.A(n_1281),
.B(n_71),
.Y(n_1351)
);

O2A1O1Ixp33_ASAP7_75t_SL g1352 ( 
.A1(n_1135),
.A2(n_71),
.B(n_76),
.C(n_94),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1194),
.A2(n_156),
.B(n_157),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1184),
.Y(n_1354)
);

AO31x2_ASAP7_75t_L g1355 ( 
.A1(n_1153),
.A2(n_159),
.A3(n_160),
.B(n_1237),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1281),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1257),
.B(n_1267),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1280),
.B(n_1191),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1194),
.A2(n_1274),
.B(n_1270),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1206),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1281),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1268),
.A2(n_1271),
.B(n_1264),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1283),
.A2(n_1140),
.B(n_1181),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1198),
.Y(n_1364)
);

BUFx10_ASAP7_75t_L g1365 ( 
.A(n_1258),
.Y(n_1365)
);

CKINVDCx11_ASAP7_75t_R g1366 ( 
.A(n_1284),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1216),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1228),
.Y(n_1368)
);

AOI221xp5_ASAP7_75t_SL g1369 ( 
.A1(n_1196),
.A2(n_1238),
.B1(n_1248),
.B2(n_1273),
.C(n_1261),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1166),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1172),
.A2(n_1247),
.B(n_1209),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1239),
.A2(n_1279),
.B(n_1193),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1236),
.B(n_1241),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1140),
.A2(n_1263),
.B(n_1282),
.Y(n_1374)
);

NOR3xp33_ASAP7_75t_SL g1375 ( 
.A(n_1244),
.B(n_1222),
.C(n_1138),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1166),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1247),
.A2(n_1254),
.B(n_1286),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1254),
.A2(n_1266),
.B(n_1286),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1141),
.B(n_1186),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1266),
.A2(n_1160),
.B(n_1131),
.Y(n_1380)
);

NAND3xp33_ASAP7_75t_L g1381 ( 
.A(n_1262),
.B(n_1141),
.C(n_1180),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1223),
.B(n_1212),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1159),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1244),
.B(n_1253),
.Y(n_1384)
);

O2A1O1Ixp5_ASAP7_75t_SL g1385 ( 
.A1(n_1176),
.A2(n_1197),
.B(n_1195),
.C(n_1220),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1218),
.Y(n_1386)
);

O2A1O1Ixp33_ASAP7_75t_SL g1387 ( 
.A1(n_1207),
.A2(n_1285),
.B(n_1226),
.C(n_1252),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1192),
.A2(n_1233),
.B(n_1251),
.C(n_1269),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1179),
.A2(n_1262),
.B1(n_1182),
.B2(n_1155),
.Y(n_1389)
);

NOR2x1_ASAP7_75t_SL g1390 ( 
.A(n_1166),
.B(n_1173),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1230),
.A2(n_1175),
.B1(n_1131),
.B2(n_1287),
.Y(n_1391)
);

AO31x2_ASAP7_75t_L g1392 ( 
.A1(n_1175),
.A2(n_1178),
.A3(n_1234),
.B(n_1203),
.Y(n_1392)
);

AO31x2_ASAP7_75t_L g1393 ( 
.A1(n_1219),
.A2(n_1211),
.A3(n_1204),
.B(n_1200),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_SL g1394 ( 
.A(n_1162),
.B(n_1208),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1246),
.A2(n_1260),
.B(n_1250),
.Y(n_1395)
);

A2O1A1Ixp33_ASAP7_75t_L g1396 ( 
.A1(n_1179),
.A2(n_1182),
.B(n_1272),
.C(n_1215),
.Y(n_1396)
);

BUFx10_ASAP7_75t_L g1397 ( 
.A(n_1284),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1284),
.A2(n_1205),
.B(n_1224),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1230),
.B(n_1284),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1173),
.A2(n_1201),
.B(n_1208),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1265),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1173),
.B(n_1201),
.Y(n_1402)
);

AO31x2_ASAP7_75t_L g1403 ( 
.A1(n_1265),
.A2(n_1005),
.A3(n_1144),
.B(n_1145),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1265),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1265),
.A2(n_986),
.B(n_1073),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1265),
.A2(n_792),
.B(n_951),
.Y(n_1406)
);

NAND2xp33_ASAP7_75t_L g1407 ( 
.A(n_1201),
.B(n_792),
.Y(n_1407)
);

NOR2x1_ASAP7_75t_SL g1408 ( 
.A(n_1201),
.B(n_1132),
.Y(n_1408)
);

CKINVDCx8_ASAP7_75t_R g1409 ( 
.A(n_1169),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1137),
.Y(n_1410)
);

AO21x2_ASAP7_75t_L g1411 ( 
.A1(n_1145),
.A2(n_1005),
.B(n_1168),
.Y(n_1411)
);

OR2x6_ASAP7_75t_L g1412 ( 
.A(n_1177),
.B(n_1221),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1276),
.A2(n_1235),
.B(n_1256),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1134),
.A2(n_986),
.B(n_792),
.Y(n_1414)
);

OAI22x1_ASAP7_75t_L g1415 ( 
.A1(n_1188),
.A2(n_966),
.B1(n_617),
.B2(n_943),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1276),
.A2(n_1235),
.B(n_1256),
.Y(n_1416)
);

NOR2x1_ASAP7_75t_R g1417 ( 
.A(n_1169),
.B(n_844),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_SL g1418 ( 
.A1(n_1243),
.A2(n_792),
.B(n_867),
.Y(n_1418)
);

BUFx12f_ASAP7_75t_L g1419 ( 
.A(n_1169),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1158),
.B(n_959),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1231),
.A2(n_986),
.B(n_1073),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1157),
.B(n_951),
.Y(n_1422)
);

A2O1A1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1152),
.A2(n_792),
.B(n_978),
.C(n_986),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1276),
.A2(n_1235),
.B(n_1256),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1134),
.A2(n_986),
.B(n_792),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1133),
.A2(n_792),
.B1(n_867),
.B2(n_951),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1183),
.B(n_669),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1134),
.A2(n_986),
.B(n_792),
.Y(n_1428)
);

AOI21xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1188),
.A2(n_669),
.B(n_792),
.Y(n_1429)
);

INVx3_ASAP7_75t_SL g1430 ( 
.A(n_1169),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1134),
.A2(n_986),
.B(n_792),
.Y(n_1431)
);

AOI221xp5_ASAP7_75t_L g1432 ( 
.A1(n_1132),
.A2(n_978),
.B1(n_867),
.B2(n_943),
.C(n_966),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1276),
.A2(n_1235),
.B(n_1256),
.Y(n_1433)
);

NAND2x1_ASAP7_75t_L g1434 ( 
.A(n_1281),
.B(n_1284),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1134),
.A2(n_986),
.B(n_792),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1137),
.Y(n_1436)
);

NAND3xp33_ASAP7_75t_SL g1437 ( 
.A(n_1188),
.B(n_659),
.C(n_655),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1276),
.A2(n_1235),
.B(n_1256),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1169),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1134),
.A2(n_986),
.B(n_792),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1208),
.Y(n_1441)
);

AO31x2_ASAP7_75t_L g1442 ( 
.A1(n_1144),
.A2(n_1005),
.A3(n_1145),
.B(n_1276),
.Y(n_1442)
);

NOR2xp67_ASAP7_75t_L g1443 ( 
.A(n_1208),
.B(n_1205),
.Y(n_1443)
);

A2O1A1Ixp33_ASAP7_75t_L g1444 ( 
.A1(n_1152),
.A2(n_792),
.B(n_978),
.C(n_986),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1137),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1141),
.A2(n_978),
.B1(n_723),
.B2(n_741),
.Y(n_1446)
);

AO31x2_ASAP7_75t_L g1447 ( 
.A1(n_1144),
.A2(n_1005),
.A3(n_1145),
.B(n_1276),
.Y(n_1447)
);

O2A1O1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1132),
.A2(n_867),
.B(n_792),
.C(n_847),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1158),
.B(n_959),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_L g1450 ( 
.A(n_1188),
.B(n_792),
.C(n_978),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1137),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1142),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1276),
.A2(n_1235),
.B(n_1256),
.Y(n_1453)
);

AO31x2_ASAP7_75t_L g1454 ( 
.A1(n_1144),
.A2(n_1005),
.A3(n_1145),
.B(n_1276),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1133),
.A2(n_792),
.B1(n_867),
.B2(n_951),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1132),
.A2(n_978),
.B1(n_966),
.B2(n_951),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1397),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1373),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1446),
.A2(n_1415),
.B1(n_1381),
.B2(n_1432),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1381),
.A2(n_1450),
.B1(n_1389),
.B2(n_1456),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1450),
.A2(n_1456),
.B1(n_1379),
.B2(n_1382),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1422),
.B(n_1314),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1337),
.A2(n_1384),
.B1(n_1406),
.B2(n_1334),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1337),
.A2(n_1334),
.B1(n_1329),
.B2(n_1391),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1350),
.Y(n_1465)
);

INVx4_ASAP7_75t_L g1466 ( 
.A(n_1303),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1421),
.A2(n_1455),
.B1(n_1426),
.B2(n_1296),
.Y(n_1467)
);

OAI22xp33_ASAP7_75t_SL g1468 ( 
.A1(n_1420),
.A2(n_1449),
.B1(n_1357),
.B2(n_1323),
.Y(n_1468)
);

AOI22xp5_ASAP7_75t_SL g1469 ( 
.A1(n_1308),
.A2(n_1427),
.B1(n_1330),
.B2(n_1348),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_SL g1470 ( 
.A1(n_1330),
.A2(n_1348),
.B1(n_1354),
.B2(n_1452),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1397),
.Y(n_1471)
);

INVx6_ASAP7_75t_L g1472 ( 
.A(n_1317),
.Y(n_1472)
);

CKINVDCx6p67_ASAP7_75t_R g1473 ( 
.A(n_1430),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1350),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1383),
.B(n_1418),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1325),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1418),
.A2(n_1429),
.B1(n_1444),
.B2(n_1423),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1338),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1340),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_SL g1480 ( 
.A1(n_1405),
.A2(n_1365),
.B1(n_1421),
.B2(n_1300),
.Y(n_1480)
);

OAI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1310),
.A2(n_1349),
.B1(n_1405),
.B2(n_1429),
.Y(n_1481)
);

CKINVDCx11_ASAP7_75t_R g1482 ( 
.A(n_1409),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_SL g1483 ( 
.A1(n_1439),
.A2(n_1315),
.B1(n_1358),
.B2(n_1360),
.Y(n_1483)
);

CKINVDCx6p67_ASAP7_75t_R g1484 ( 
.A(n_1419),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1437),
.A2(n_1290),
.B1(n_1365),
.B2(n_1300),
.Y(n_1485)
);

BUFx12f_ASAP7_75t_L g1486 ( 
.A(n_1304),
.Y(n_1486)
);

INVxp67_ASAP7_75t_SL g1487 ( 
.A(n_1297),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_SL g1488 ( 
.A1(n_1399),
.A2(n_1408),
.B1(n_1353),
.B2(n_1394),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1318),
.Y(n_1489)
);

INVx6_ASAP7_75t_L g1490 ( 
.A(n_1317),
.Y(n_1490)
);

BUFx10_ASAP7_75t_L g1491 ( 
.A(n_1298),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1343),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1347),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1386),
.A2(n_1335),
.B1(n_1451),
.B2(n_1367),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1353),
.A2(n_1394),
.B1(n_1336),
.B2(n_1326),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1410),
.A2(n_1445),
.B1(n_1436),
.B2(n_1291),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_SL g1497 ( 
.A1(n_1372),
.A2(n_1341),
.B1(n_1344),
.B2(n_1346),
.Y(n_1497)
);

INVxp67_ASAP7_75t_SL g1498 ( 
.A(n_1327),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1350),
.Y(n_1499)
);

BUFx12f_ASAP7_75t_L g1500 ( 
.A(n_1295),
.Y(n_1500)
);

INVx6_ASAP7_75t_L g1501 ( 
.A(n_1312),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1311),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1361),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_SL g1504 ( 
.A1(n_1372),
.A2(n_1407),
.B1(n_1310),
.B2(n_1378),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1356),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1316),
.A2(n_1364),
.B1(n_1368),
.B2(n_1342),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1319),
.Y(n_1507)
);

INVx3_ASAP7_75t_SL g1508 ( 
.A(n_1295),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1380),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1312),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1361),
.Y(n_1511)
);

INVx2_ASAP7_75t_SL g1512 ( 
.A(n_1312),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1339),
.A2(n_1448),
.B1(n_1292),
.B2(n_1375),
.Y(n_1513)
);

BUFx12f_ASAP7_75t_L g1514 ( 
.A(n_1412),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1292),
.A2(n_1294),
.B1(n_1388),
.B2(n_1396),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1370),
.Y(n_1516)
);

BUFx10_ASAP7_75t_L g1517 ( 
.A(n_1361),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1376),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1412),
.B(n_1441),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_1402),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1311),
.Y(n_1521)
);

BUFx8_ASAP7_75t_L g1522 ( 
.A(n_1417),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1311),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1414),
.A2(n_1431),
.B1(n_1425),
.B2(n_1428),
.Y(n_1524)
);

CKINVDCx11_ASAP7_75t_R g1525 ( 
.A(n_1417),
.Y(n_1525)
);

CKINVDCx20_ASAP7_75t_R g1526 ( 
.A(n_1400),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1333),
.Y(n_1527)
);

CKINVDCx11_ASAP7_75t_R g1528 ( 
.A(n_1401),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1369),
.B(n_1443),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1369),
.B(n_1443),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1333),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1398),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1333),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1351),
.Y(n_1534)
);

CKINVDCx11_ASAP7_75t_R g1535 ( 
.A(n_1404),
.Y(n_1535)
);

NAND2x1p5_ASAP7_75t_L g1536 ( 
.A(n_1434),
.B(n_1374),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1377),
.Y(n_1537)
);

INVx6_ASAP7_75t_L g1538 ( 
.A(n_1390),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1352),
.Y(n_1539)
);

BUFx12f_ASAP7_75t_L g1540 ( 
.A(n_1345),
.Y(n_1540)
);

BUFx12f_ASAP7_75t_L g1541 ( 
.A(n_1385),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1363),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1306),
.A2(n_1371),
.B1(n_1395),
.B2(n_1411),
.Y(n_1543)
);

BUFx12f_ASAP7_75t_L g1544 ( 
.A(n_1387),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1306),
.A2(n_1395),
.B1(n_1440),
.B2(n_1435),
.Y(n_1545)
);

CKINVDCx6p67_ASAP7_75t_R g1546 ( 
.A(n_1392),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1293),
.A2(n_1331),
.B1(n_1305),
.B2(n_1289),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1309),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1392),
.B(n_1320),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1392),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1293),
.A2(n_1328),
.B1(n_1362),
.B2(n_1313),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1403),
.Y(n_1552)
);

OAI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1302),
.A2(n_1307),
.B1(n_1309),
.B2(n_1355),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1309),
.Y(n_1554)
);

INVx4_ASAP7_75t_L g1555 ( 
.A(n_1324),
.Y(n_1555)
);

BUFx12f_ASAP7_75t_L g1556 ( 
.A(n_1299),
.Y(n_1556)
);

BUFx12f_ASAP7_75t_L g1557 ( 
.A(n_1299),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1332),
.Y(n_1558)
);

INVxp67_ASAP7_75t_L g1559 ( 
.A(n_1301),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_SL g1560 ( 
.A1(n_1355),
.A2(n_1359),
.B1(n_1403),
.B2(n_1393),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1413),
.A2(n_1433),
.B1(n_1453),
.B2(n_1416),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1393),
.Y(n_1562)
);

BUFx4_ASAP7_75t_SL g1563 ( 
.A(n_1393),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1424),
.A2(n_1438),
.B1(n_1442),
.B2(n_1447),
.Y(n_1564)
);

BUFx2_ASAP7_75t_SL g1565 ( 
.A(n_1447),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1447),
.A2(n_1454),
.B1(n_1321),
.B2(n_1322),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1321),
.A2(n_1446),
.B1(n_978),
.B2(n_741),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_SL g1568 ( 
.A1(n_1322),
.A2(n_928),
.B1(n_741),
.B2(n_723),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_SL g1569 ( 
.A1(n_1381),
.A2(n_928),
.B1(n_741),
.B2(n_723),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1373),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1419),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1450),
.A2(n_792),
.B1(n_1456),
.B2(n_1418),
.Y(n_1572)
);

NAND2x1p5_ASAP7_75t_L g1573 ( 
.A(n_1330),
.B(n_992),
.Y(n_1573)
);

INVx6_ASAP7_75t_L g1574 ( 
.A(n_1397),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_SL g1575 ( 
.A1(n_1381),
.A2(n_928),
.B1(n_741),
.B2(n_723),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1366),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1419),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1450),
.A2(n_792),
.B1(n_1456),
.B2(n_1418),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_SL g1579 ( 
.A1(n_1381),
.A2(n_928),
.B1(n_741),
.B2(n_723),
.Y(n_1579)
);

BUFx12f_ASAP7_75t_L g1580 ( 
.A(n_1304),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1450),
.A2(n_792),
.B1(n_1456),
.B2(n_1418),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1450),
.A2(n_792),
.B1(n_1456),
.B2(n_1418),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1366),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_SL g1584 ( 
.A1(n_1381),
.A2(n_928),
.B1(n_741),
.B2(n_723),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1303),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_SL g1586 ( 
.A1(n_1381),
.A2(n_928),
.B1(n_741),
.B2(n_723),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1450),
.A2(n_792),
.B1(n_1456),
.B2(n_1418),
.Y(n_1587)
);

OAI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1456),
.A2(n_966),
.B1(n_965),
.B2(n_1450),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1446),
.A2(n_978),
.B1(n_741),
.B2(n_1415),
.Y(n_1589)
);

INVx4_ASAP7_75t_L g1590 ( 
.A(n_1303),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1366),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_1366),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_SL g1593 ( 
.A1(n_1381),
.A2(n_928),
.B1(n_741),
.B2(n_723),
.Y(n_1593)
);

INVx11_ASAP7_75t_L g1594 ( 
.A(n_1419),
.Y(n_1594)
);

CKINVDCx11_ASAP7_75t_R g1595 ( 
.A(n_1409),
.Y(n_1595)
);

CKINVDCx11_ASAP7_75t_R g1596 ( 
.A(n_1409),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1446),
.A2(n_978),
.B1(n_741),
.B2(n_1415),
.Y(n_1597)
);

CKINVDCx11_ASAP7_75t_R g1598 ( 
.A(n_1409),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1373),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1446),
.A2(n_978),
.B1(n_741),
.B2(n_1415),
.Y(n_1600)
);

CKINVDCx11_ASAP7_75t_R g1601 ( 
.A(n_1409),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1303),
.Y(n_1602)
);

CKINVDCx20_ASAP7_75t_R g1603 ( 
.A(n_1304),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1450),
.A2(n_792),
.B1(n_1456),
.B2(n_1418),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1366),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_SL g1606 ( 
.A1(n_1381),
.A2(n_928),
.B1(n_741),
.B2(n_723),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1373),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_SL g1608 ( 
.A1(n_1381),
.A2(n_928),
.B1(n_741),
.B2(n_723),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1373),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1460),
.A2(n_1459),
.B1(n_1461),
.B2(n_1606),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1505),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1489),
.Y(n_1612)
);

OAI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1572),
.A2(n_1581),
.B(n_1578),
.Y(n_1613)
);

OAI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1524),
.A2(n_1561),
.B(n_1549),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1556),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1509),
.Y(n_1616)
);

AO21x2_ASAP7_75t_L g1617 ( 
.A1(n_1553),
.A2(n_1531),
.B(n_1527),
.Y(n_1617)
);

BUFx2_ASAP7_75t_SL g1618 ( 
.A(n_1498),
.Y(n_1618)
);

BUFx3_ASAP7_75t_L g1619 ( 
.A(n_1501),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1476),
.B(n_1478),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1602),
.B(n_1466),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1502),
.Y(n_1622)
);

OAI22xp33_ASAP7_75t_SL g1623 ( 
.A1(n_1475),
.A2(n_1587),
.B1(n_1582),
.B2(n_1604),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1542),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1482),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1458),
.B(n_1570),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1561),
.A2(n_1550),
.B(n_1547),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1521),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1523),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1523),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_SL g1631 ( 
.A1(n_1573),
.A2(n_1513),
.B(n_1477),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1542),
.Y(n_1632)
);

OA21x2_ASAP7_75t_L g1633 ( 
.A1(n_1533),
.A2(n_1564),
.B(n_1545),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1479),
.B(n_1492),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1501),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1493),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1461),
.B(n_1548),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1547),
.A2(n_1545),
.B(n_1551),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1554),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1507),
.Y(n_1640)
);

AOI21xp33_ASAP7_75t_SL g1641 ( 
.A1(n_1481),
.A2(n_1588),
.B(n_1508),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1562),
.Y(n_1642)
);

OAI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1551),
.A2(n_1564),
.B(n_1543),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1537),
.Y(n_1644)
);

INVx2_ASAP7_75t_SL g1645 ( 
.A(n_1501),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1552),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1563),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1595),
.Y(n_1648)
);

INVx3_ASAP7_75t_L g1649 ( 
.A(n_1557),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1540),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1546),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_L g1652 ( 
.A1(n_1543),
.A2(n_1536),
.B(n_1566),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1555),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1565),
.Y(n_1654)
);

AO31x2_ASAP7_75t_L g1655 ( 
.A1(n_1515),
.A2(n_1555),
.A3(n_1529),
.B(n_1530),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1559),
.Y(n_1656)
);

INVx3_ASAP7_75t_L g1657 ( 
.A(n_1536),
.Y(n_1657)
);

INVx4_ASAP7_75t_L g1658 ( 
.A(n_1573),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1487),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1599),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1607),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1566),
.A2(n_1496),
.B(n_1467),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1460),
.B(n_1609),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1496),
.Y(n_1664)
);

BUFx6f_ASAP7_75t_L g1665 ( 
.A(n_1540),
.Y(n_1665)
);

INVx3_ASAP7_75t_L g1666 ( 
.A(n_1558),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1459),
.A2(n_1608),
.B1(n_1569),
.B2(n_1575),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1553),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1504),
.B(n_1462),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1535),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1494),
.Y(n_1671)
);

INVx2_ASAP7_75t_SL g1672 ( 
.A(n_1576),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1494),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1560),
.Y(n_1674)
);

INVxp33_ASAP7_75t_L g1675 ( 
.A(n_1483),
.Y(n_1675)
);

OA21x2_ASAP7_75t_L g1676 ( 
.A1(n_1467),
.A2(n_1463),
.B(n_1464),
.Y(n_1676)
);

AO21x2_ASAP7_75t_L g1677 ( 
.A1(n_1481),
.A2(n_1588),
.B(n_1539),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1532),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1576),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1472),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1480),
.B(n_1463),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_1465),
.Y(n_1682)
);

AOI21x1_ASAP7_75t_L g1683 ( 
.A1(n_1519),
.A2(n_1534),
.B(n_1516),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1579),
.A2(n_1586),
.B1(n_1584),
.B2(n_1593),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1541),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1576),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1490),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1541),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1520),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1506),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1506),
.Y(n_1691)
);

OAI221xp5_ASAP7_75t_L g1692 ( 
.A1(n_1495),
.A2(n_1597),
.B1(n_1589),
.B2(n_1600),
.C(n_1464),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1465),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1596),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1465),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1512),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1465),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1503),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1468),
.B(n_1470),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1503),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1503),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1469),
.B(n_1568),
.Y(n_1702)
);

OAI21x1_ASAP7_75t_L g1703 ( 
.A1(n_1474),
.A2(n_1499),
.B(n_1457),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1503),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1567),
.B(n_1518),
.Y(n_1705)
);

OAI21x1_ASAP7_75t_L g1706 ( 
.A1(n_1474),
.A2(n_1499),
.B(n_1457),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1526),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1488),
.Y(n_1708)
);

INVx3_ASAP7_75t_L g1709 ( 
.A(n_1544),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1544),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1497),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1538),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1511),
.Y(n_1713)
);

OAI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1485),
.A2(n_1567),
.B(n_1600),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_1528),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1485),
.A2(n_1511),
.B(n_1471),
.Y(n_1716)
);

AO21x2_ASAP7_75t_L g1717 ( 
.A1(n_1589),
.A2(n_1597),
.B(n_1514),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1471),
.Y(n_1718)
);

INVxp67_ASAP7_75t_L g1719 ( 
.A(n_1611),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1612),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1703),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1640),
.B(n_1605),
.Y(n_1722)
);

OAI21x1_ASAP7_75t_L g1723 ( 
.A1(n_1638),
.A2(n_1514),
.B(n_1517),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1647),
.B(n_1592),
.Y(n_1724)
);

AND4x1_ASAP7_75t_L g1725 ( 
.A(n_1613),
.B(n_1522),
.C(n_1525),
.D(n_1576),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1622),
.Y(n_1726)
);

NOR2x1_ASAP7_75t_SL g1727 ( 
.A(n_1618),
.B(n_1592),
.Y(n_1727)
);

A2O1A1Ixp33_ASAP7_75t_L g1728 ( 
.A1(n_1610),
.A2(n_1591),
.B(n_1583),
.C(n_1510),
.Y(n_1728)
);

AOI221xp5_ASAP7_75t_L g1729 ( 
.A1(n_1623),
.A2(n_1585),
.B1(n_1583),
.B2(n_1591),
.C(n_1518),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1610),
.A2(n_1580),
.B1(n_1486),
.B2(n_1603),
.Y(n_1730)
);

AOI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1631),
.A2(n_1517),
.B(n_1590),
.Y(n_1731)
);

A2O1A1Ixp33_ASAP7_75t_L g1732 ( 
.A1(n_1681),
.A2(n_1571),
.B(n_1577),
.C(n_1486),
.Y(n_1732)
);

NOR2x1_ASAP7_75t_SL g1733 ( 
.A(n_1618),
.B(n_1500),
.Y(n_1733)
);

AOI221xp5_ASAP7_75t_L g1734 ( 
.A1(n_1668),
.A2(n_1466),
.B1(n_1590),
.B2(n_1508),
.C(n_1580),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1647),
.B(n_1473),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1676),
.A2(n_1641),
.B1(n_1681),
.B2(n_1631),
.Y(n_1736)
);

O2A1O1Ixp33_ASAP7_75t_L g1737 ( 
.A1(n_1641),
.A2(n_1522),
.B(n_1491),
.C(n_1500),
.Y(n_1737)
);

OAI21xp33_ASAP7_75t_L g1738 ( 
.A1(n_1711),
.A2(n_1484),
.B(n_1574),
.Y(n_1738)
);

INVx8_ASAP7_75t_L g1739 ( 
.A(n_1625),
.Y(n_1739)
);

AO32x2_ASAP7_75t_L g1740 ( 
.A1(n_1635),
.A2(n_1594),
.A3(n_1598),
.B1(n_1601),
.B2(n_1645),
.Y(n_1740)
);

CKINVDCx20_ASAP7_75t_R g1741 ( 
.A(n_1648),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1622),
.Y(n_1742)
);

O2A1O1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1711),
.A2(n_1677),
.B(n_1685),
.C(n_1688),
.Y(n_1743)
);

NAND2xp33_ASAP7_75t_R g1744 ( 
.A(n_1694),
.B(n_1676),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1621),
.B(n_1689),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1707),
.B(n_1669),
.Y(n_1746)
);

AO32x2_ASAP7_75t_L g1747 ( 
.A1(n_1635),
.A2(n_1645),
.A3(n_1672),
.B1(n_1686),
.B2(n_1679),
.Y(n_1747)
);

OA21x2_ASAP7_75t_L g1748 ( 
.A1(n_1614),
.A2(n_1688),
.B(n_1685),
.Y(n_1748)
);

OAI221xp5_ASAP7_75t_L g1749 ( 
.A1(n_1692),
.A2(n_1714),
.B1(n_1668),
.B2(n_1678),
.C(n_1699),
.Y(n_1749)
);

A2O1A1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1667),
.A2(n_1675),
.B(n_1669),
.C(n_1708),
.Y(n_1750)
);

AOI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1702),
.A2(n_1708),
.B(n_1663),
.C(n_1662),
.Y(n_1751)
);

OAI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1676),
.A2(n_1667),
.B1(n_1674),
.B2(n_1664),
.C(n_1684),
.Y(n_1752)
);

OA21x2_ASAP7_75t_L g1753 ( 
.A1(n_1614),
.A2(n_1627),
.B(n_1643),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1636),
.B(n_1659),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1620),
.B(n_1634),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1715),
.B(n_1670),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1659),
.B(n_1660),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1651),
.B(n_1619),
.Y(n_1758)
);

BUFx3_ASAP7_75t_L g1759 ( 
.A(n_1715),
.Y(n_1759)
);

INVx5_ASAP7_75t_SL g1760 ( 
.A(n_1715),
.Y(n_1760)
);

OA21x2_ASAP7_75t_L g1761 ( 
.A1(n_1627),
.A2(n_1643),
.B(n_1652),
.Y(n_1761)
);

AO21x1_ASAP7_75t_L g1762 ( 
.A1(n_1674),
.A2(n_1683),
.B(n_1662),
.Y(n_1762)
);

OA21x2_ASAP7_75t_L g1763 ( 
.A1(n_1652),
.A2(n_1638),
.B(n_1654),
.Y(n_1763)
);

OAI221xp5_ASAP7_75t_L g1764 ( 
.A1(n_1676),
.A2(n_1664),
.B1(n_1671),
.B2(n_1673),
.C(n_1716),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1637),
.B(n_1696),
.Y(n_1765)
);

O2A1O1Ixp33_ASAP7_75t_SL g1766 ( 
.A1(n_1709),
.A2(n_1710),
.B(n_1713),
.C(n_1718),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1660),
.B(n_1661),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1693),
.B(n_1695),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1693),
.B(n_1695),
.Y(n_1769)
);

AO21x1_ASAP7_75t_L g1770 ( 
.A1(n_1683),
.A2(n_1661),
.B(n_1626),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1615),
.B(n_1649),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1697),
.B(n_1698),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1709),
.B(n_1710),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1697),
.B(n_1698),
.Y(n_1774)
);

AOI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1677),
.A2(n_1671),
.B1(n_1673),
.B2(n_1616),
.C(n_1705),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1709),
.B(n_1710),
.Y(n_1776)
);

OAI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1633),
.A2(n_1706),
.B(n_1653),
.Y(n_1777)
);

O2A1O1Ixp33_ASAP7_75t_L g1778 ( 
.A1(n_1709),
.A2(n_1710),
.B(n_1713),
.C(n_1700),
.Y(n_1778)
);

A2O1A1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1615),
.A2(n_1649),
.B(n_1642),
.C(n_1650),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1658),
.B(n_1649),
.Y(n_1780)
);

OAI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1706),
.A2(n_1718),
.B(n_1656),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1701),
.B(n_1704),
.Y(n_1782)
);

A2O1A1Ixp33_ASAP7_75t_L g1783 ( 
.A1(n_1642),
.A2(n_1650),
.B(n_1665),
.C(n_1691),
.Y(n_1783)
);

OAI211xp5_ASAP7_75t_L g1784 ( 
.A1(n_1656),
.A2(n_1704),
.B(n_1701),
.C(n_1616),
.Y(n_1784)
);

A2O1A1Ixp33_ASAP7_75t_L g1785 ( 
.A1(n_1650),
.A2(n_1665),
.B(n_1691),
.C(n_1690),
.Y(n_1785)
);

AO32x2_ASAP7_75t_L g1786 ( 
.A1(n_1658),
.A2(n_1655),
.A3(n_1690),
.B1(n_1639),
.B2(n_1629),
.Y(n_1786)
);

A2O1A1Ixp33_ASAP7_75t_L g1787 ( 
.A1(n_1665),
.A2(n_1632),
.B(n_1624),
.C(n_1657),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1624),
.B(n_1632),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1655),
.B(n_1682),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1789),
.B(n_1777),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1720),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1726),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1726),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1755),
.B(n_1628),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1765),
.B(n_1666),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1742),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1719),
.Y(n_1797)
);

NOR2xp67_ASAP7_75t_L g1798 ( 
.A(n_1721),
.B(n_1653),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1788),
.B(n_1666),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1746),
.B(n_1655),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1754),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1768),
.B(n_1633),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1769),
.B(n_1772),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1757),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1774),
.B(n_1633),
.Y(n_1805)
);

CKINVDCx8_ASAP7_75t_R g1806 ( 
.A(n_1739),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1767),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1770),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1782),
.B(n_1633),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1777),
.B(n_1644),
.Y(n_1810)
);

BUFx2_ASAP7_75t_L g1811 ( 
.A(n_1747),
.Y(n_1811)
);

INVx4_ASAP7_75t_R g1812 ( 
.A(n_1759),
.Y(n_1812)
);

AOI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1736),
.A2(n_1717),
.B1(n_1658),
.B2(n_1712),
.Y(n_1813)
);

INVx2_ASAP7_75t_SL g1814 ( 
.A(n_1722),
.Y(n_1814)
);

NOR2x1_ASAP7_75t_L g1815 ( 
.A(n_1784),
.B(n_1653),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1786),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1747),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1747),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1748),
.B(n_1630),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1786),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1763),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1752),
.A2(n_1717),
.B1(n_1687),
.B2(n_1680),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1721),
.B(n_1646),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1781),
.Y(n_1824)
);

NOR2x1_ASAP7_75t_L g1825 ( 
.A(n_1778),
.B(n_1657),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1762),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1763),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1764),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1811),
.B(n_1753),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1811),
.B(n_1761),
.Y(n_1830)
);

INVxp67_ASAP7_75t_SL g1831 ( 
.A(n_1821),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1815),
.B(n_1787),
.Y(n_1832)
);

BUFx2_ASAP7_75t_L g1833 ( 
.A(n_1815),
.Y(n_1833)
);

AOI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1828),
.A2(n_1749),
.B1(n_1775),
.B2(n_1750),
.C(n_1730),
.Y(n_1834)
);

BUFx2_ASAP7_75t_L g1835 ( 
.A(n_1810),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_SL g1836 ( 
.A1(n_1806),
.A2(n_1730),
.B1(n_1756),
.B2(n_1735),
.Y(n_1836)
);

OAI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1822),
.A2(n_1751),
.B1(n_1728),
.B2(n_1729),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1792),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1800),
.B(n_1761),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1792),
.Y(n_1840)
);

OAI221xp5_ASAP7_75t_L g1841 ( 
.A1(n_1828),
.A2(n_1751),
.B1(n_1744),
.B2(n_1743),
.C(n_1725),
.Y(n_1841)
);

BUFx2_ASAP7_75t_L g1842 ( 
.A(n_1810),
.Y(n_1842)
);

AND2x4_ASAP7_75t_L g1843 ( 
.A(n_1790),
.B(n_1727),
.Y(n_1843)
);

INVx2_ASAP7_75t_SL g1844 ( 
.A(n_1812),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1824),
.B(n_1617),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1793),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1824),
.A2(n_1732),
.B1(n_1738),
.B2(n_1734),
.C(n_1737),
.Y(n_1847)
);

AND2x2_ASAP7_75t_SL g1848 ( 
.A(n_1790),
.B(n_1725),
.Y(n_1848)
);

AND2x4_ASAP7_75t_L g1849 ( 
.A(n_1790),
.B(n_1771),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1806),
.B(n_1739),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1793),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1802),
.B(n_1758),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1803),
.B(n_1724),
.Y(n_1853)
);

BUFx2_ASAP7_75t_L g1854 ( 
.A(n_1817),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1819),
.Y(n_1855)
);

INVxp67_ASAP7_75t_SL g1856 ( 
.A(n_1821),
.Y(n_1856)
);

BUFx2_ASAP7_75t_L g1857 ( 
.A(n_1817),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1819),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1827),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1796),
.Y(n_1860)
);

AOI221xp5_ASAP7_75t_L g1861 ( 
.A1(n_1808),
.A2(n_1738),
.B1(n_1717),
.B2(n_1783),
.C(n_1785),
.Y(n_1861)
);

AOI221xp5_ASAP7_75t_L g1862 ( 
.A1(n_1808),
.A2(n_1779),
.B1(n_1745),
.B2(n_1766),
.C(n_1735),
.Y(n_1862)
);

OAI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1826),
.A2(n_1731),
.B(n_1723),
.Y(n_1863)
);

INVx5_ASAP7_75t_L g1864 ( 
.A(n_1823),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1805),
.B(n_1740),
.Y(n_1865)
);

AND3x1_ASAP7_75t_L g1866 ( 
.A(n_1818),
.B(n_1773),
.C(n_1776),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1865),
.B(n_1791),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1838),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1854),
.B(n_1794),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1864),
.B(n_1825),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1838),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1865),
.B(n_1814),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1840),
.Y(n_1873)
);

INVx4_ASAP7_75t_L g1874 ( 
.A(n_1832),
.Y(n_1874)
);

HB1xp67_ASAP7_75t_L g1875 ( 
.A(n_1854),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1840),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1857),
.B(n_1818),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1865),
.B(n_1814),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1857),
.B(n_1801),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1846),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1864),
.B(n_1825),
.Y(n_1881)
);

INVxp67_ASAP7_75t_L g1882 ( 
.A(n_1833),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1846),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1864),
.B(n_1798),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1835),
.B(n_1799),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1835),
.B(n_1799),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1834),
.A2(n_1826),
.B1(n_1820),
.B2(n_1816),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1842),
.B(n_1805),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1851),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1851),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1833),
.B(n_1807),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1842),
.B(n_1809),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1855),
.B(n_1858),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1829),
.Y(n_1894)
);

AND4x1_ASAP7_75t_L g1895 ( 
.A(n_1862),
.B(n_1740),
.C(n_1813),
.D(n_1780),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1858),
.B(n_1801),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1860),
.B(n_1807),
.Y(n_1897)
);

NOR2xp67_ASAP7_75t_L g1898 ( 
.A(n_1864),
.B(n_1827),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1860),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1859),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1849),
.B(n_1795),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1849),
.B(n_1795),
.Y(n_1902)
);

INVx3_ASAP7_75t_SL g1903 ( 
.A(n_1848),
.Y(n_1903)
);

INVx2_ASAP7_75t_SL g1904 ( 
.A(n_1864),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1829),
.B(n_1804),
.Y(n_1905)
);

NOR2x1_ASAP7_75t_L g1906 ( 
.A(n_1874),
.B(n_1850),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1869),
.B(n_1829),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1875),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1868),
.Y(n_1909)
);

OAI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1903),
.A2(n_1866),
.B1(n_1862),
.B2(n_1841),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1900),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1868),
.Y(n_1912)
);

NOR2xp33_ASAP7_75t_L g1913 ( 
.A(n_1874),
.B(n_1741),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1874),
.B(n_1866),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1900),
.Y(n_1915)
);

INVxp67_ASAP7_75t_SL g1916 ( 
.A(n_1875),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1869),
.B(n_1830),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1871),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1874),
.B(n_1843),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1891),
.B(n_1832),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1900),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1871),
.Y(n_1922)
);

NOR2x1_ASAP7_75t_L g1923 ( 
.A(n_1870),
.B(n_1832),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1873),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1873),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1893),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1879),
.B(n_1830),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1891),
.B(n_1832),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1876),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1876),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1880),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1879),
.B(n_1830),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1880),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1903),
.B(n_1853),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1888),
.B(n_1843),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1903),
.B(n_1853),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1883),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1895),
.B(n_1839),
.Y(n_1938)
);

OR2x2_ASAP7_75t_L g1939 ( 
.A(n_1905),
.B(n_1877),
.Y(n_1939)
);

BUFx3_ASAP7_75t_L g1940 ( 
.A(n_1870),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1883),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1889),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1905),
.B(n_1845),
.Y(n_1943)
);

INVxp67_ASAP7_75t_SL g1944 ( 
.A(n_1895),
.Y(n_1944)
);

INVxp67_ASAP7_75t_L g1945 ( 
.A(n_1867),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1888),
.B(n_1843),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1867),
.B(n_1839),
.Y(n_1947)
);

INVx1_ASAP7_75t_SL g1948 ( 
.A(n_1872),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1888),
.B(n_1892),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1892),
.B(n_1843),
.Y(n_1950)
);

NAND2x1p5_ASAP7_75t_L g1951 ( 
.A(n_1870),
.B(n_1848),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1889),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1892),
.B(n_1852),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1890),
.Y(n_1954)
);

AOI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1887),
.A2(n_1837),
.B1(n_1841),
.B2(n_1834),
.Y(n_1955)
);

AOI21xp33_ASAP7_75t_SL g1956 ( 
.A1(n_1955),
.A2(n_1836),
.B(n_1882),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1918),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1914),
.B(n_1885),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1944),
.B(n_1887),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1918),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1922),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1911),
.Y(n_1962)
);

INVxp67_ASAP7_75t_SL g1963 ( 
.A(n_1910),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1914),
.B(n_1885),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1916),
.B(n_1882),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1953),
.B(n_1886),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1908),
.B(n_1894),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1922),
.Y(n_1968)
);

OR2x2_ASAP7_75t_L g1969 ( 
.A(n_1939),
.B(n_1877),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1909),
.B(n_1894),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1953),
.B(n_1886),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1939),
.B(n_1897),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1911),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1949),
.B(n_1919),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1949),
.B(n_1901),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1913),
.B(n_1836),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1919),
.B(n_1901),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1915),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1945),
.B(n_1897),
.Y(n_1979)
);

AND2x4_ASAP7_75t_L g1980 ( 
.A(n_1923),
.B(n_1870),
.Y(n_1980)
);

OR2x2_ASAP7_75t_L g1981 ( 
.A(n_1907),
.B(n_1896),
.Y(n_1981)
);

OAI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1938),
.A2(n_1848),
.B1(n_1837),
.B2(n_1847),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1948),
.B(n_1935),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1924),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1920),
.B(n_1872),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1924),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1942),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_L g1988 ( 
.A(n_1951),
.B(n_1849),
.Y(n_1988)
);

HB1xp67_ASAP7_75t_L g1989 ( 
.A(n_1912),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1942),
.Y(n_1990)
);

AND2x2_ASAP7_75t_SL g1991 ( 
.A(n_1928),
.B(n_1881),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1925),
.B(n_1890),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1929),
.B(n_1899),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1954),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1930),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1935),
.B(n_1902),
.Y(n_1996)
);

AND2x2_ASAP7_75t_SL g1997 ( 
.A(n_1959),
.B(n_1881),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1963),
.B(n_1926),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1956),
.B(n_1951),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_R g2000 ( 
.A(n_1965),
.B(n_1934),
.Y(n_2000)
);

AOI21xp5_ASAP7_75t_L g2001 ( 
.A1(n_1982),
.A2(n_1951),
.B(n_1906),
.Y(n_2001)
);

AOI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1982),
.A2(n_1861),
.B1(n_1936),
.B2(n_1820),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1975),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_L g2004 ( 
.A(n_1956),
.B(n_1976),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1957),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1957),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1960),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1960),
.Y(n_2008)
);

NAND3xp33_ASAP7_75t_L g2009 ( 
.A(n_1967),
.B(n_1926),
.C(n_1954),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1983),
.B(n_1946),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1983),
.B(n_1946),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_1991),
.B(n_1940),
.Y(n_2012)
);

OAI22xp5_ASAP7_75t_L g2013 ( 
.A1(n_1988),
.A2(n_1881),
.B1(n_1940),
.B2(n_1947),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1966),
.B(n_1878),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1961),
.Y(n_2015)
);

OAI21xp5_ASAP7_75t_L g2016 ( 
.A1(n_1967),
.A2(n_1863),
.B(n_1881),
.Y(n_2016)
);

A2O1A1Ixp33_ASAP7_75t_L g2017 ( 
.A1(n_1991),
.A2(n_1820),
.B(n_1932),
.C(n_1927),
.Y(n_2017)
);

OAI21xp5_ASAP7_75t_L g2018 ( 
.A1(n_1991),
.A2(n_1863),
.B(n_1927),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1961),
.Y(n_2019)
);

INVx1_ASAP7_75t_SL g2020 ( 
.A(n_1958),
.Y(n_2020)
);

INVxp67_ASAP7_75t_L g2021 ( 
.A(n_1989),
.Y(n_2021)
);

OAI21xp33_ASAP7_75t_L g2022 ( 
.A1(n_1958),
.A2(n_1917),
.B(n_1907),
.Y(n_2022)
);

AOI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1970),
.A2(n_1845),
.B(n_1831),
.Y(n_2023)
);

AOI21xp33_ASAP7_75t_L g2024 ( 
.A1(n_1968),
.A2(n_1921),
.B(n_1915),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1968),
.Y(n_2025)
);

NAND4xp25_ASAP7_75t_L g2026 ( 
.A(n_1964),
.B(n_1847),
.C(n_1917),
.D(n_1932),
.Y(n_2026)
);

NAND2x1_ASAP7_75t_L g2027 ( 
.A(n_2001),
.B(n_1980),
.Y(n_2027)
);

INVx1_ASAP7_75t_SL g2028 ( 
.A(n_2020),
.Y(n_2028)
);

AOI22xp33_ASAP7_75t_SL g2029 ( 
.A1(n_1997),
.A2(n_1964),
.B1(n_1980),
.B2(n_1969),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_2004),
.B(n_1966),
.Y(n_2030)
);

INVxp33_ASAP7_75t_L g2031 ( 
.A(n_2004),
.Y(n_2031)
);

AOI22xp33_ASAP7_75t_L g2032 ( 
.A1(n_2002),
.A2(n_1973),
.B1(n_1962),
.B2(n_1978),
.Y(n_2032)
);

OR2x2_ASAP7_75t_L g2033 ( 
.A(n_2026),
.B(n_1969),
.Y(n_2033)
);

NOR2xp33_ASAP7_75t_L g2034 ( 
.A(n_1999),
.B(n_1972),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2003),
.B(n_1971),
.Y(n_2035)
);

AOI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_1999),
.A2(n_1861),
.B1(n_1978),
.B2(n_1962),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_2010),
.B(n_1974),
.Y(n_2037)
);

AOI21xp5_ASAP7_75t_SL g2038 ( 
.A1(n_1998),
.A2(n_2021),
.B(n_2017),
.Y(n_2038)
);

OAI221xp5_ASAP7_75t_SL g2039 ( 
.A1(n_2022),
.A2(n_1981),
.B1(n_1972),
.B2(n_1970),
.C(n_1979),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_2011),
.B(n_1971),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1997),
.B(n_1975),
.Y(n_2041)
);

AOI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_2018),
.A2(n_1973),
.B1(n_1978),
.B2(n_1962),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_2005),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2005),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2014),
.B(n_1995),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_2012),
.B(n_1974),
.Y(n_2046)
);

INVx3_ASAP7_75t_L g2047 ( 
.A(n_2006),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_2012),
.B(n_1979),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2007),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_2016),
.B(n_1996),
.Y(n_2050)
);

BUFx3_ASAP7_75t_L g2051 ( 
.A(n_2008),
.Y(n_2051)
);

INVxp67_ASAP7_75t_L g2052 ( 
.A(n_2043),
.Y(n_2052)
);

OAI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_2038),
.A2(n_1980),
.B1(n_2009),
.B2(n_1985),
.Y(n_2053)
);

AOI21xp33_ASAP7_75t_SL g2054 ( 
.A1(n_2031),
.A2(n_2013),
.B(n_1980),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2043),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_2037),
.Y(n_2056)
);

AOI211xp5_ASAP7_75t_L g2057 ( 
.A1(n_2038),
.A2(n_2024),
.B(n_2000),
.C(n_2019),
.Y(n_2057)
);

INVxp67_ASAP7_75t_L g2058 ( 
.A(n_2044),
.Y(n_2058)
);

NAND2xp33_ASAP7_75t_SL g2059 ( 
.A(n_2027),
.B(n_2000),
.Y(n_2059)
);

AOI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_2036),
.A2(n_2032),
.B1(n_2033),
.B2(n_2042),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2047),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2037),
.B(n_2046),
.Y(n_2062)
);

A2O1A1Ixp33_ASAP7_75t_L g2063 ( 
.A1(n_2034),
.A2(n_2023),
.B(n_2025),
.C(n_2015),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2046),
.B(n_1996),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_L g2065 ( 
.A(n_2031),
.B(n_2030),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2028),
.B(n_1981),
.Y(n_2066)
);

O2A1O1Ixp33_ASAP7_75t_SL g2067 ( 
.A1(n_2041),
.A2(n_1994),
.B(n_1984),
.C(n_1986),
.Y(n_2067)
);

AOI21xp33_ASAP7_75t_SL g2068 ( 
.A1(n_2029),
.A2(n_1904),
.B(n_1984),
.Y(n_2068)
);

OR2x2_ASAP7_75t_L g2069 ( 
.A(n_2056),
.B(n_2040),
.Y(n_2069)
);

NAND3xp33_ASAP7_75t_L g2070 ( 
.A(n_2057),
.B(n_2051),
.C(n_2048),
.Y(n_2070)
);

AOI221xp5_ASAP7_75t_L g2071 ( 
.A1(n_2060),
.A2(n_2039),
.B1(n_2051),
.B2(n_2050),
.C(n_2047),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2062),
.Y(n_2072)
);

AOI222xp33_ASAP7_75t_L g2073 ( 
.A1(n_2052),
.A2(n_2050),
.B1(n_2049),
.B2(n_2047),
.C1(n_1973),
.C2(n_2045),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2064),
.B(n_2035),
.Y(n_2074)
);

OAI21xp33_ASAP7_75t_SL g2075 ( 
.A1(n_2065),
.A2(n_1977),
.B(n_1994),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2066),
.B(n_1977),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2063),
.B(n_1986),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_2052),
.B(n_1987),
.Y(n_2078)
);

NOR2xp33_ASAP7_75t_SL g2079 ( 
.A(n_2058),
.B(n_1904),
.Y(n_2079)
);

INVxp67_ASAP7_75t_L g2080 ( 
.A(n_2059),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2061),
.B(n_2054),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2072),
.Y(n_2082)
);

OAI221xp5_ASAP7_75t_L g2083 ( 
.A1(n_2071),
.A2(n_2053),
.B1(n_2068),
.B2(n_2055),
.C(n_2058),
.Y(n_2083)
);

AOI21xp33_ASAP7_75t_SL g2084 ( 
.A1(n_2070),
.A2(n_1990),
.B(n_1987),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_R g2085 ( 
.A(n_2080),
.B(n_2067),
.Y(n_2085)
);

XNOR2xp5_ASAP7_75t_L g2086 ( 
.A(n_2074),
.B(n_1990),
.Y(n_2086)
);

O2A1O1Ixp5_ASAP7_75t_SL g2087 ( 
.A1(n_2081),
.A2(n_1993),
.B(n_1992),
.C(n_1952),
.Y(n_2087)
);

AOI211xp5_ASAP7_75t_L g2088 ( 
.A1(n_2077),
.A2(n_1898),
.B(n_1993),
.C(n_1992),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2086),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2082),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2084),
.B(n_2076),
.Y(n_2091)
);

A2O1A1Ixp33_ASAP7_75t_L g2092 ( 
.A1(n_2083),
.A2(n_2075),
.B(n_2078),
.C(n_2079),
.Y(n_2092)
);

BUFx2_ASAP7_75t_L g2093 ( 
.A(n_2085),
.Y(n_2093)
);

BUFx2_ASAP7_75t_L g2094 ( 
.A(n_2088),
.Y(n_2094)
);

AOI21xp33_ASAP7_75t_L g2095 ( 
.A1(n_2087),
.A2(n_2073),
.B(n_2079),
.Y(n_2095)
);

INVx2_ASAP7_75t_SL g2096 ( 
.A(n_2082),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_2093),
.B(n_2096),
.Y(n_2097)
);

XNOR2x1_ASAP7_75t_L g2098 ( 
.A(n_2089),
.B(n_2069),
.Y(n_2098)
);

AND2x4_ASAP7_75t_L g2099 ( 
.A(n_2090),
.B(n_1950),
.Y(n_2099)
);

NAND4xp75_ASAP7_75t_L g2100 ( 
.A(n_2095),
.B(n_1898),
.C(n_1904),
.D(n_1950),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2091),
.B(n_1878),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_2094),
.Y(n_2102)
);

OAI22xp5_ASAP7_75t_L g2103 ( 
.A1(n_2098),
.A2(n_2092),
.B1(n_2095),
.B2(n_1937),
.Y(n_2103)
);

HB1xp67_ASAP7_75t_L g2104 ( 
.A(n_2097),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2101),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2099),
.B(n_1902),
.Y(n_2106)
);

NAND3x1_ASAP7_75t_L g2107 ( 
.A(n_2105),
.B(n_2102),
.C(n_2100),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2104),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2108),
.Y(n_2109)
);

OAI22xp5_ASAP7_75t_L g2110 ( 
.A1(n_2109),
.A2(n_2100),
.B1(n_2103),
.B2(n_2107),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2109),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2111),
.B(n_2106),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_2110),
.Y(n_2113)
);

AOI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_2112),
.A2(n_1921),
.B(n_1943),
.Y(n_2114)
);

AOI22xp33_ASAP7_75t_L g2115 ( 
.A1(n_2114),
.A2(n_2113),
.B1(n_1943),
.B2(n_1831),
.Y(n_2115)
);

AOI22x1_ASAP7_75t_L g2116 ( 
.A1(n_2115),
.A2(n_1941),
.B1(n_1933),
.B2(n_1931),
.Y(n_2116)
);

XOR2xp5_ASAP7_75t_L g2117 ( 
.A(n_2116),
.B(n_1733),
.Y(n_2117)
);

OAI221xp5_ASAP7_75t_R g2118 ( 
.A1(n_2117),
.A2(n_1797),
.B1(n_1760),
.B2(n_1844),
.C(n_1884),
.Y(n_2118)
);

AOI211xp5_ASAP7_75t_L g2119 ( 
.A1(n_2118),
.A2(n_1856),
.B(n_1844),
.C(n_1884),
.Y(n_2119)
);


endmodule