module fake_aes_11572_n_599 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_599);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_599;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g73 ( .A(n_9), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_20), .Y(n_74) );
INVx2_ASAP7_75t_L g75 ( .A(n_13), .Y(n_75) );
INVxp67_ASAP7_75t_SL g76 ( .A(n_25), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_37), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_56), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_57), .Y(n_79) );
INVxp33_ASAP7_75t_L g80 ( .A(n_17), .Y(n_80) );
BUFx3_ASAP7_75t_L g81 ( .A(n_27), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_2), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_33), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_9), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_64), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_32), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_41), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_47), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_52), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_4), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_7), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_34), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_60), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_4), .Y(n_94) );
INVxp67_ASAP7_75t_L g95 ( .A(n_28), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_62), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_18), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_22), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_6), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_49), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_46), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_3), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_30), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_23), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_10), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_69), .Y(n_106) );
AND2x2_ASAP7_75t_L g107 ( .A(n_21), .B(n_15), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_55), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_59), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_54), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_11), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_36), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_68), .Y(n_113) );
CKINVDCx14_ASAP7_75t_R g114 ( .A(n_61), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_11), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_38), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_50), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_73), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_74), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_74), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_77), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_97), .Y(n_122) );
INVxp33_ASAP7_75t_L g123 ( .A(n_82), .Y(n_123) );
BUFx2_ASAP7_75t_L g124 ( .A(n_73), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_97), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_91), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_109), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_77), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_109), .B(n_0), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_78), .B(n_0), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_99), .Y(n_131) );
INVx2_ASAP7_75t_SL g132 ( .A(n_81), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_75), .B(n_84), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_111), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_75), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_78), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_114), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_81), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_98), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_80), .B(n_1), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_81), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_79), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g143 ( .A(n_82), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_79), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_100), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_83), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_90), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_83), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_90), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_85), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_113), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_102), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_85), .Y(n_153) );
NOR2xp33_ASAP7_75t_R g154 ( .A(n_107), .B(n_35), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_87), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_87), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_153), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_153), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_123), .A2(n_102), .B1(n_115), .B2(n_84), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_133), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g161 ( .A1(n_119), .A2(n_117), .B(n_116), .C(n_88), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_137), .B(n_95), .Y(n_162) );
NAND2x1p5_ASAP7_75t_L g163 ( .A(n_119), .B(n_107), .Y(n_163) );
INVxp67_ASAP7_75t_SL g164 ( .A(n_124), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_124), .B(n_117), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_153), .Y(n_166) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_120), .A2(n_115), .B1(n_94), .B2(n_105), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_120), .B(n_116), .Y(n_169) );
INVx4_ASAP7_75t_L g170 ( .A(n_133), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_122), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_121), .B(n_112), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_122), .Y(n_174) );
BUFx4f_ASAP7_75t_L g175 ( .A(n_121), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_125), .Y(n_176) );
INVx4_ASAP7_75t_L g177 ( .A(n_133), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_125), .Y(n_178) );
BUFx2_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_140), .B(n_94), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
BUFx2_ASAP7_75t_L g182 ( .A(n_134), .Y(n_182) );
INVx1_ASAP7_75t_SL g183 ( .A(n_126), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_141), .Y(n_184) );
INVx1_ASAP7_75t_SL g185 ( .A(n_118), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_138), .Y(n_186) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_139), .B(n_112), .Y(n_188) );
INVxp67_ASAP7_75t_L g189 ( .A(n_140), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_127), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_138), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_127), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_146), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_151), .B(n_110), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_128), .B(n_136), .Y(n_195) );
INVxp33_ASAP7_75t_L g196 ( .A(n_133), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_146), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_128), .B(n_110), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_136), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_142), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_142), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_144), .B(n_105), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_144), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_148), .B(n_108), .Y(n_204) );
OR2x2_ASAP7_75t_SL g205 ( .A(n_143), .B(n_108), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_148), .B(n_106), .Y(n_206) );
BUFx2_ASAP7_75t_L g207 ( .A(n_147), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_150), .B(n_106), .Y(n_208) );
AO22x2_ASAP7_75t_L g209 ( .A1(n_150), .A2(n_104), .B1(n_103), .B2(n_101), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_155), .B(n_104), .Y(n_210) );
INVx4_ASAP7_75t_SL g211 ( .A(n_132), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_157), .Y(n_212) );
NOR3xp33_ASAP7_75t_SL g213 ( .A(n_162), .B(n_130), .C(n_129), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_163), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_164), .B(n_152), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_207), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_170), .B(n_156), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_170), .B(n_156), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_170), .B(n_155), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_209), .A2(n_135), .B1(n_88), .B2(n_93), .Y(n_220) );
BUFx10_ASAP7_75t_L g221 ( .A(n_194), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_168), .Y(n_222) );
INVxp67_ASAP7_75t_SL g223 ( .A(n_163), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_163), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_193), .Y(n_225) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_179), .Y(n_226) );
BUFx8_ASAP7_75t_L g227 ( .A(n_179), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_177), .B(n_180), .Y(n_228) );
NAND3xp33_ASAP7_75t_SL g229 ( .A(n_185), .B(n_149), .C(n_154), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_177), .B(n_135), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_193), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_177), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_180), .B(n_135), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_206), .B(n_135), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_168), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_160), .B(n_103), .Y(n_236) );
NAND2x1p5_ASAP7_75t_L g237 ( .A(n_182), .B(n_101), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_189), .B(n_210), .Y(n_238) );
OR2x2_ASAP7_75t_L g239 ( .A(n_183), .B(n_1), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_197), .Y(n_240) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_182), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_206), .B(n_89), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_207), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_197), .Y(n_244) );
INVx3_ASAP7_75t_SL g245 ( .A(n_205), .Y(n_245) );
BUFx2_ASAP7_75t_L g246 ( .A(n_187), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_157), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_158), .Y(n_248) );
BUFx4f_ASAP7_75t_L g249 ( .A(n_206), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_158), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_209), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_166), .Y(n_252) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_166), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_202), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_210), .B(n_96), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_202), .Y(n_256) );
INVx3_ASAP7_75t_L g257 ( .A(n_171), .Y(n_257) );
NAND2xp33_ASAP7_75t_SL g258 ( .A(n_199), .B(n_96), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_208), .B(n_93), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_174), .Y(n_260) );
INVx3_ASAP7_75t_L g261 ( .A(n_171), .Y(n_261) );
BUFx12f_ASAP7_75t_L g262 ( .A(n_205), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_174), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_208), .B(n_86), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_173), .Y(n_265) );
NOR2xp33_ASAP7_75t_R g266 ( .A(n_188), .B(n_2), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_171), .Y(n_267) );
AND2x4_ASAP7_75t_SL g268 ( .A(n_208), .B(n_92), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_227), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_220), .A2(n_209), .B1(n_175), .B2(n_200), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_250), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_252), .Y(n_272) );
HAxp5_ASAP7_75t_L g273 ( .A(n_216), .B(n_196), .CON(n_273), .SN(n_273) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_251), .A2(n_209), .B1(n_175), .B2(n_165), .Y(n_274) );
INVx4_ASAP7_75t_L g275 ( .A(n_249), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_212), .Y(n_276) );
BUFx2_ASAP7_75t_L g277 ( .A(n_249), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_212), .Y(n_278) );
INVx3_ASAP7_75t_SL g279 ( .A(n_216), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_212), .Y(n_280) );
INVx1_ASAP7_75t_SL g281 ( .A(n_268), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_226), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_268), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_249), .Y(n_284) );
NAND2x1p5_ASAP7_75t_L g285 ( .A(n_214), .B(n_175), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_212), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_238), .B(n_159), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_238), .B(n_195), .Y(n_288) );
INVx4_ASAP7_75t_SL g289 ( .A(n_247), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_238), .B(n_199), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_224), .B(n_203), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_247), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_247), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_220), .A2(n_203), .B1(n_201), .B2(n_200), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_247), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_237), .B(n_241), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_248), .Y(n_297) );
AOI22xp33_ASAP7_75t_SL g298 ( .A1(n_227), .A2(n_169), .B1(n_172), .B2(n_198), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_255), .B(n_201), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_248), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_223), .B(n_192), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_248), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_260), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_255), .B(n_167), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_263), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_246), .Y(n_306) );
BUFx12f_ASAP7_75t_L g307 ( .A(n_227), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_225), .Y(n_308) );
INVx2_ASAP7_75t_SL g309 ( .A(n_237), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_243), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_248), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_217), .A2(n_204), .B(n_181), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_271), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_309), .B(n_254), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_271), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_301), .B(n_255), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_287), .A2(n_262), .B1(n_215), .B2(n_245), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_292), .Y(n_318) );
INVx4_ASAP7_75t_L g319 ( .A(n_289), .Y(n_319) );
OAI21x1_ASAP7_75t_L g320 ( .A1(n_270), .A2(n_173), .B(n_184), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_282), .A2(n_262), .B1(n_245), .B2(n_229), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_288), .A2(n_256), .B1(n_233), .B2(n_228), .C(n_161), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_272), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_301), .B(n_259), .Y(n_324) );
NAND3xp33_ASAP7_75t_SL g325 ( .A(n_298), .B(n_266), .C(n_239), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_292), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_304), .A2(n_259), .B1(n_236), .B2(n_258), .Y(n_327) );
NOR2xp33_ASAP7_75t_R g328 ( .A(n_269), .B(n_258), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_306), .B(n_242), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_281), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_281), .Y(n_331) );
AOI21x1_ASAP7_75t_L g332 ( .A1(n_270), .A2(n_184), .B(n_186), .Y(n_332) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_307), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_309), .B(n_232), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_292), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_310), .A2(n_259), .B1(n_232), .B2(n_236), .Y(n_336) );
BUFx3_ASAP7_75t_L g337 ( .A(n_285), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_275), .Y(n_338) );
CKINVDCx8_ASAP7_75t_R g339 ( .A(n_289), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_294), .A2(n_236), .B1(n_231), .B2(n_240), .Y(n_340) );
AND2x4_ASAP7_75t_SL g341 ( .A(n_333), .B(n_275), .Y(n_341) );
OAI22xp33_ASAP7_75t_L g342 ( .A1(n_340), .A2(n_279), .B1(n_283), .B2(n_307), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_325), .A2(n_279), .B1(n_340), .B2(n_316), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_325), .A2(n_279), .B1(n_296), .B2(n_274), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_316), .B(n_291), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_313), .Y(n_346) );
AOI222xp33_ASAP7_75t_L g347 ( .A1(n_316), .A2(n_317), .B1(n_322), .B2(n_324), .C1(n_321), .C2(n_315), .Y(n_347) );
INVx1_ASAP7_75t_SL g348 ( .A(n_331), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_337), .B(n_275), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_324), .B(n_283), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_324), .A2(n_266), .B1(n_221), .B2(n_291), .Y(n_351) );
AOI322xp5_ASAP7_75t_L g352 ( .A1(n_313), .A2(n_273), .A3(n_213), .B1(n_290), .B2(n_192), .C1(n_190), .C2(n_178), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_320), .A2(n_299), .B(n_303), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_315), .B(n_291), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_327), .A2(n_294), .B1(n_291), .B2(n_272), .Y(n_355) );
A2O1A1Ixp33_ASAP7_75t_SL g356 ( .A1(n_338), .A2(n_267), .B(n_261), .C(n_257), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_323), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_327), .A2(n_221), .B1(n_303), .B2(n_308), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_336), .A2(n_308), .B1(n_305), .B2(n_285), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_323), .B(n_305), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_314), .A2(n_285), .B1(n_264), .B2(n_284), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_339), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_322), .A2(n_244), .B1(n_234), .B2(n_277), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_332), .A2(n_276), .B(n_311), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_329), .B(n_277), .Y(n_365) );
AND2x4_ASAP7_75t_SL g366 ( .A(n_349), .B(n_319), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_342), .A2(n_329), .B1(n_314), .B2(n_328), .C(n_330), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_349), .Y(n_368) );
AOI21x1_ASAP7_75t_L g369 ( .A1(n_364), .A2(n_332), .B(n_320), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_354), .B(n_273), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_343), .A2(n_314), .B1(n_331), .B2(n_330), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_347), .A2(n_314), .B1(n_338), .B2(n_337), .Y(n_372) );
INVx2_ASAP7_75t_SL g373 ( .A(n_341), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_348), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_357), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_355), .A2(n_337), .B1(n_338), .B2(n_334), .Y(n_376) );
OAI33xp33_ASAP7_75t_L g377 ( .A1(n_359), .A2(n_92), .A3(n_178), .B1(n_176), .B2(n_190), .B3(n_273), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_348), .Y(n_378) );
AOI21x1_ASAP7_75t_L g379 ( .A1(n_364), .A2(n_320), .B(n_335), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_346), .Y(n_380) );
OAI22xp33_ASAP7_75t_L g381 ( .A1(n_363), .A2(n_339), .B1(n_338), .B2(n_275), .Y(n_381) );
AO21x2_ASAP7_75t_L g382 ( .A1(n_353), .A2(n_335), .B(n_326), .Y(n_382) );
INVxp67_ASAP7_75t_L g383 ( .A(n_365), .Y(n_383) );
BUFx10_ASAP7_75t_L g384 ( .A(n_341), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_354), .B(n_326), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_346), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_345), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_362), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_357), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_360), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_344), .A2(n_230), .B1(n_218), .B2(n_219), .C(n_176), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_360), .B(n_326), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_363), .Y(n_393) );
AOI33xp33_ASAP7_75t_L g394 ( .A1(n_358), .A2(n_334), .A3(n_191), .B1(n_186), .B2(n_7), .B3(n_8), .Y(n_394) );
NAND3xp33_ASAP7_75t_L g395 ( .A(n_352), .B(n_335), .C(n_318), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_345), .A2(n_334), .B1(n_221), .B2(n_284), .Y(n_396) );
NOR2xp33_ASAP7_75t_R g397 ( .A(n_362), .B(n_339), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_362), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_383), .B(n_352), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_370), .B(n_350), .Y(n_400) );
INVx2_ASAP7_75t_SL g401 ( .A(n_384), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_370), .A2(n_351), .B1(n_361), .B2(n_349), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_374), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_375), .Y(n_404) );
OAI33xp33_ASAP7_75t_L g405 ( .A1(n_375), .A2(n_3), .A3(n_5), .B1(n_6), .B2(n_8), .B3(n_10), .Y(n_405) );
NAND3xp33_ASAP7_75t_L g406 ( .A(n_367), .B(n_76), .C(n_356), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_390), .B(n_334), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_377), .A2(n_267), .B1(n_261), .B2(n_257), .C(n_312), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_393), .A2(n_372), .B1(n_381), .B2(n_371), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_380), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_389), .Y(n_411) );
INVx3_ASAP7_75t_L g412 ( .A(n_398), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_376), .A2(n_319), .B1(n_318), .B2(n_311), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_376), .A2(n_319), .B1(n_318), .B2(n_302), .Y(n_414) );
NAND2xp33_ASAP7_75t_R g415 ( .A(n_397), .B(n_5), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_380), .Y(n_416) );
OAI21xp5_ASAP7_75t_L g417 ( .A1(n_394), .A2(n_181), .B(n_191), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_380), .B(n_318), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_390), .B(n_319), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_393), .A2(n_257), .B1(n_261), .B2(n_267), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_386), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_389), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_386), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_386), .B(n_318), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_382), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_390), .Y(n_426) );
INVx6_ASAP7_75t_L g427 ( .A(n_384), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_385), .B(n_318), .Y(n_428) );
INVx5_ASAP7_75t_L g429 ( .A(n_384), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_384), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_382), .Y(n_431) );
INVxp67_ASAP7_75t_L g432 ( .A(n_378), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_387), .B(n_318), .Y(n_433) );
INVx5_ASAP7_75t_L g434 ( .A(n_373), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_385), .B(n_12), .Y(n_435) );
AOI211xp5_ASAP7_75t_SL g436 ( .A1(n_392), .A2(n_302), .B(n_300), .C(n_297), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_382), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_379), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_368), .B(n_12), .Y(n_439) );
OAI21xp5_ASAP7_75t_SL g440 ( .A1(n_373), .A2(n_253), .B(n_14), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_379), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_368), .B(n_13), .Y(n_442) );
INVx4_ASAP7_75t_L g443 ( .A(n_366), .Y(n_443) );
OAI31xp33_ASAP7_75t_L g444 ( .A1(n_395), .A2(n_232), .A3(n_222), .B(n_235), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_369), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_411), .B(n_369), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_410), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_403), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_432), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_411), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_422), .B(n_398), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_422), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_404), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_428), .B(n_398), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_428), .B(n_398), .Y(n_455) );
NAND2x1p5_ASAP7_75t_L g456 ( .A(n_443), .B(n_398), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_426), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_441), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_410), .B(n_395), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_416), .B(n_398), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_416), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_441), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_399), .B(n_388), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_421), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_421), .B(n_366), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_423), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_438), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_423), .B(n_366), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_438), .Y(n_469) );
BUFx2_ASAP7_75t_L g470 ( .A(n_443), .Y(n_470) );
AOI211x1_ASAP7_75t_L g471 ( .A1(n_439), .A2(n_14), .B(n_15), .C(n_16), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_400), .B(n_16), .Y(n_472) );
INVxp67_ASAP7_75t_SL g473 ( .A(n_433), .Y(n_473) );
NAND2xp33_ASAP7_75t_SL g474 ( .A(n_443), .B(n_396), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_429), .B(n_434), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_407), .B(n_431), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_431), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_435), .B(n_391), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_435), .B(n_19), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_418), .B(n_24), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_418), .B(n_26), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_424), .B(n_29), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_424), .B(n_31), .Y(n_483) );
INVx3_ASAP7_75t_L g484 ( .A(n_425), .Y(n_484) );
NAND2xp33_ASAP7_75t_SL g485 ( .A(n_415), .B(n_253), .Y(n_485) );
NOR3xp33_ASAP7_75t_L g486 ( .A(n_440), .B(n_222), .C(n_235), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_437), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_437), .B(n_39), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_425), .B(n_40), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_412), .B(n_42), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_430), .B(n_43), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_445), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_412), .B(n_44), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_409), .B(n_442), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_419), .B(n_253), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_445), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_412), .B(n_45), .Y(n_497) );
OAI33xp33_ASAP7_75t_L g498 ( .A1(n_406), .A2(n_419), .A3(n_413), .B1(n_414), .B2(n_405), .B3(n_402), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_463), .B(n_427), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_448), .B(n_442), .Y(n_500) );
NOR2xp33_ASAP7_75t_SL g501 ( .A(n_470), .B(n_429), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_450), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_449), .B(n_439), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_473), .B(n_401), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_450), .Y(n_505) );
AOI21xp33_ASAP7_75t_L g506 ( .A1(n_472), .A2(n_434), .B(n_444), .Y(n_506) );
OAI22xp33_ASAP7_75t_L g507 ( .A1(n_470), .A2(n_429), .B1(n_427), .B2(n_434), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_453), .B(n_434), .Y(n_508) );
NOR2x1_ASAP7_75t_L g509 ( .A(n_475), .B(n_429), .Y(n_509) );
CKINVDCx16_ASAP7_75t_R g510 ( .A(n_485), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_452), .Y(n_511) );
OAI221xp5_ASAP7_75t_L g512 ( .A1(n_486), .A2(n_427), .B1(n_420), .B2(n_417), .C(n_434), .Y(n_512) );
OAI211xp5_ASAP7_75t_L g513 ( .A1(n_471), .A2(n_429), .B(n_436), .C(n_408), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_471), .A2(n_427), .B1(n_300), .B2(n_297), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_457), .Y(n_515) );
NAND3x1_ASAP7_75t_L g516 ( .A(n_494), .B(n_48), .C(n_51), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_454), .B(n_53), .Y(n_517) );
OAI321xp33_ASAP7_75t_L g518 ( .A1(n_456), .A2(n_295), .A3(n_293), .B1(n_286), .B2(n_280), .C(n_278), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_476), .B(n_58), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_465), .B(n_289), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_SL g521 ( .A1(n_472), .A2(n_63), .B(n_65), .C(n_66), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_474), .A2(n_289), .B1(n_295), .B2(n_278), .Y(n_522) );
O2A1O1Ixp5_ASAP7_75t_L g523 ( .A1(n_498), .A2(n_293), .B(n_286), .C(n_280), .Y(n_523) );
OAI221xp5_ASAP7_75t_L g524 ( .A1(n_478), .A2(n_265), .B1(n_276), .B2(n_71), .C(n_72), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_457), .B(n_265), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_479), .A2(n_67), .B(n_70), .C(n_211), .Y(n_526) );
INVxp67_ASAP7_75t_SL g527 ( .A(n_484), .Y(n_527) );
NAND4xp25_ASAP7_75t_L g528 ( .A(n_477), .B(n_211), .C(n_487), .D(n_446), .Y(n_528) );
INVxp67_ASAP7_75t_L g529 ( .A(n_468), .Y(n_529) );
NOR3xp33_ASAP7_75t_SL g530 ( .A(n_491), .B(n_211), .C(n_477), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_495), .A2(n_211), .B(n_488), .C(n_481), .Y(n_531) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_446), .A2(n_451), .B1(n_484), .B2(n_469), .C(n_467), .Y(n_532) );
OAI221xp5_ASAP7_75t_L g533 ( .A1(n_456), .A2(n_469), .B1(n_467), .B2(n_484), .C(n_459), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_465), .B(n_468), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_467), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_495), .A2(n_488), .B(n_481), .C(n_482), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_502), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_505), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_529), .B(n_454), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_511), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_515), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_535), .Y(n_542) );
OAI22xp33_ASAP7_75t_L g543 ( .A1(n_501), .A2(n_456), .B1(n_459), .B2(n_465), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_500), .B(n_464), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_503), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_504), .B(n_455), .Y(n_546) );
NOR4xp25_ASAP7_75t_SL g547 ( .A(n_512), .B(n_496), .C(n_492), .D(n_461), .Y(n_547) );
INVxp67_ASAP7_75t_L g548 ( .A(n_533), .Y(n_548) );
XOR2xp5_ASAP7_75t_L g549 ( .A(n_510), .B(n_455), .Y(n_549) );
NOR2xp33_ASAP7_75t_R g550 ( .A(n_499), .B(n_483), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_534), .B(n_483), .Y(n_551) );
NOR2xp33_ASAP7_75t_R g552 ( .A(n_508), .B(n_482), .Y(n_552) );
AOI221xp5_ASAP7_75t_SL g553 ( .A1(n_536), .A2(n_480), .B1(n_496), .B2(n_492), .C(n_493), .Y(n_553) );
XNOR2xp5_ASAP7_75t_L g554 ( .A(n_516), .B(n_480), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_532), .B(n_458), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_507), .A2(n_497), .B(n_493), .Y(n_556) );
NOR2xp67_ASAP7_75t_L g557 ( .A(n_528), .B(n_484), .Y(n_557) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_522), .A2(n_447), .B1(n_466), .B2(n_462), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_536), .B(n_458), .Y(n_559) );
OAI21xp33_ASAP7_75t_L g560 ( .A1(n_548), .A2(n_513), .B(n_506), .Y(n_560) );
XNOR2xp5_ASAP7_75t_L g561 ( .A(n_549), .B(n_509), .Y(n_561) );
NOR2x1_ASAP7_75t_L g562 ( .A(n_554), .B(n_513), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_548), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_553), .B(n_523), .C(n_514), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_547), .A2(n_520), .B(n_531), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_545), .B(n_519), .Y(n_566) );
OAI21xp33_ASAP7_75t_L g567 ( .A1(n_559), .A2(n_527), .B(n_517), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_555), .B(n_462), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_543), .B(n_530), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_542), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_557), .B(n_460), .Y(n_571) );
XNOR2x1_ASAP7_75t_L g572 ( .A(n_546), .B(n_525), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_551), .A2(n_531), .B1(n_524), .B2(n_526), .Y(n_573) );
OAI22xp33_ASAP7_75t_L g574 ( .A1(n_556), .A2(n_518), .B1(n_490), .B2(n_497), .Y(n_574) );
XNOR2xp5_ASAP7_75t_L g575 ( .A(n_539), .B(n_523), .Y(n_575) );
AOI221xp5_ASAP7_75t_L g576 ( .A1(n_544), .A2(n_489), .B1(n_490), .B2(n_521), .C(n_543), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_562), .A2(n_542), .B1(n_537), .B2(n_538), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_570), .Y(n_578) );
OAI22xp33_ASAP7_75t_L g579 ( .A1(n_564), .A2(n_550), .B1(n_552), .B2(n_558), .Y(n_579) );
CKINVDCx16_ASAP7_75t_R g580 ( .A(n_561), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_572), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_563), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_575), .B(n_540), .Y(n_583) );
NAND2xp33_ASAP7_75t_SL g584 ( .A(n_569), .B(n_541), .Y(n_584) );
A2O1A1Ixp33_ASAP7_75t_L g585 ( .A1(n_565), .A2(n_489), .B(n_567), .C(n_576), .Y(n_585) );
AOI32xp33_ASAP7_75t_L g586 ( .A1(n_573), .A2(n_562), .A3(n_560), .B1(n_574), .B2(n_576), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_571), .A2(n_562), .B1(n_560), .B2(n_563), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_566), .B(n_568), .Y(n_588) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_582), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_578), .Y(n_590) );
NAND2x1_ASAP7_75t_L g591 ( .A(n_577), .B(n_587), .Y(n_591) );
NOR3xp33_ASAP7_75t_L g592 ( .A(n_584), .B(n_579), .C(n_580), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_590), .Y(n_593) );
AOI22xp33_ASAP7_75t_SL g594 ( .A1(n_592), .A2(n_581), .B1(n_583), .B2(n_586), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_593), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_594), .Y(n_596) );
INVxp67_ASAP7_75t_SL g597 ( .A(n_596), .Y(n_597) );
AOI222xp33_ASAP7_75t_L g598 ( .A1(n_597), .A2(n_595), .B1(n_584), .B2(n_579), .C1(n_589), .C2(n_585), .Y(n_598) );
AOI21xp33_ASAP7_75t_L g599 ( .A1(n_598), .A2(n_591), .B(n_588), .Y(n_599) );
endmodule