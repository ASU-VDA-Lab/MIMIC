module fake_ariane_712_n_1956 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1956);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1956;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_194;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_38),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_8),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_174),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_142),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_80),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_114),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_0),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_88),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_103),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_52),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_189),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_66),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_95),
.Y(n_208)
);

BUFx8_ASAP7_75t_SL g209 ( 
.A(n_73),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_68),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_34),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_102),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_106),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_45),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_162),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_29),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_183),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_168),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_188),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_15),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_147),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_78),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_65),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_37),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_166),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_156),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_65),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_54),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_179),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_75),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_139),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_90),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_4),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_144),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_184),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_25),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_70),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_171),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_89),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_175),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_35),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_2),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_69),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_51),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_173),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_59),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_5),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_119),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_33),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_8),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_172),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_24),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_128),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_68),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_53),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_131),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_86),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_149),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_104),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_50),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_100),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_72),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_62),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_1),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_34),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_93),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_73),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_146),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_124),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_115),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_27),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_22),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_9),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_32),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_31),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_122),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_170),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_111),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_192),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_62),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_81),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_83),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_41),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_17),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_7),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_43),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_181),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_59),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_44),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_126),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_98),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_132),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_3),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_9),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_87),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_31),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_150),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_71),
.Y(n_299)
);

BUFx10_ASAP7_75t_L g300 ( 
.A(n_135),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_72),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_56),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_43),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_158),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_52),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_11),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_76),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_108),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_66),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_29),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_159),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_30),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_143),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_85),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_97),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_38),
.Y(n_316)
);

BUFx10_ASAP7_75t_L g317 ( 
.A(n_141),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_16),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_64),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_48),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_69),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_26),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_32),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_13),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_113),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_0),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_48),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_37),
.Y(n_328)
);

BUFx10_ASAP7_75t_L g329 ( 
.A(n_79),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_190),
.Y(n_330)
);

BUFx10_ASAP7_75t_L g331 ( 
.A(n_44),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_26),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_94),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_110),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_20),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_50),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_19),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_129),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_157),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_39),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_165),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_82),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_63),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_187),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_28),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_191),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_109),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_137),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_57),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_36),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_77),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_121),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_23),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_1),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_10),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_77),
.Y(n_356)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_101),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_84),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_46),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_10),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_41),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_67),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_51),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_92),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_45),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_21),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_22),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_57),
.Y(n_368)
);

INVx4_ASAP7_75t_R g369 ( 
.A(n_178),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_6),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_61),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_140),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_33),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_74),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_64),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_46),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_3),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_76),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_16),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_138),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_35),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_4),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_96),
.Y(n_383)
);

BUFx2_ASAP7_75t_SL g384 ( 
.A(n_169),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_161),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_186),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_209),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_249),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_249),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_204),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_249),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_297),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_249),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_201),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_297),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_300),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_220),
.B(n_2),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_321),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_218),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_300),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_194),
.B(n_5),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_321),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_194),
.B(n_6),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_204),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_227),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_196),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_L g407 ( 
.A(n_261),
.B(n_7),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_196),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_242),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_247),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_300),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_228),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_287),
.Y(n_413)
);

NOR2xp67_ASAP7_75t_L g414 ( 
.A(n_286),
.B(n_327),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_220),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_220),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_220),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_368),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_228),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_300),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_317),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_234),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_374),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_317),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_234),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_357),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_317),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_348),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_317),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_329),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_329),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_245),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_216),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_202),
.B(n_11),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_329),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_201),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_329),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_202),
.B(n_12),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_195),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_206),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_245),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_264),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_232),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_201),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_264),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_274),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_340),
.B(n_12),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_274),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_210),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_211),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_223),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_276),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_276),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_348),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_224),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_281),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_281),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_230),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_203),
.B(n_13),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_237),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_201),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_299),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_238),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_216),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_232),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_299),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_243),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_220),
.B(n_14),
.Y(n_468)
);

INVxp33_ASAP7_75t_SL g469 ( 
.A(n_244),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_203),
.B(n_212),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_302),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_250),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_251),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_302),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_303),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_253),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_303),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_255),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_256),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_306),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_263),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_364),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_306),
.Y(n_483)
);

NOR2xp67_ASAP7_75t_L g484 ( 
.A(n_343),
.B(n_14),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_220),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_L g486 ( 
.A(n_248),
.B(n_15),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_212),
.B(n_17),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_415),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_415),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_416),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_433),
.B(n_220),
.Y(n_491)
);

NAND2x1_ASAP7_75t_L g492 ( 
.A(n_470),
.B(n_369),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_428),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_428),
.Y(n_494)
);

BUFx8_ASAP7_75t_L g495 ( 
.A(n_404),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_428),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_428),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_416),
.Y(n_498)
);

AND2x6_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_358),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_464),
.B(n_220),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_428),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_417),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_485),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_469),
.B(n_221),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_454),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_406),
.B(n_248),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_417),
.B(n_220),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_454),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_399),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_397),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_408),
.B(n_284),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_412),
.B(n_284),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_390),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_468),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_454),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_454),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_394),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_454),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_388),
.B(n_216),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_392),
.B(n_221),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_419),
.Y(n_521)
);

AND3x2_ASAP7_75t_L g522 ( 
.A(n_467),
.B(n_403),
.C(n_401),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_422),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_425),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_432),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_441),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_395),
.B(n_231),
.Y(n_527)
);

AND3x2_ASAP7_75t_L g528 ( 
.A(n_434),
.B(n_381),
.C(n_266),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_442),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_388),
.B(n_389),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_445),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_448),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_452),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_453),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_426),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g536 ( 
.A1(n_456),
.A2(n_358),
.B(n_233),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_439),
.Y(n_537)
);

AND2x6_ASAP7_75t_L g538 ( 
.A(n_438),
.B(n_358),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_405),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_457),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_466),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_471),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_474),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_475),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_477),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_480),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_398),
.B(n_402),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_389),
.B(n_216),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_391),
.B(n_216),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_483),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_459),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_436),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_487),
.Y(n_553)
);

AND3x2_ASAP7_75t_L g554 ( 
.A(n_446),
.B(n_207),
.C(n_324),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_462),
.B(n_231),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_391),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_443),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_486),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_447),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_393),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_393),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_465),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_439),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_484),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_440),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_407),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_440),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_561),
.B(n_396),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_509),
.Y(n_569)
);

INVxp33_ASAP7_75t_L g570 ( 
.A(n_513),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_503),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_503),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_503),
.Y(n_573)
);

OR2x6_ASAP7_75t_L g574 ( 
.A(n_492),
.B(n_324),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_556),
.B(n_396),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_552),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_507),
.Y(n_577)
);

NAND3xp33_ASAP7_75t_L g578 ( 
.A(n_510),
.B(n_514),
.C(n_553),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_561),
.B(n_400),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_503),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_503),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_524),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_488),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_524),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_553),
.B(n_444),
.Y(n_585)
);

CKINVDCx16_ASAP7_75t_R g586 ( 
.A(n_517),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_510),
.B(n_411),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_556),
.B(n_411),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_524),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_507),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_538),
.A2(n_427),
.B1(n_437),
.B2(n_430),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_561),
.B(n_420),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_552),
.B(n_420),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_552),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_L g595 ( 
.A1(n_555),
.A2(n_424),
.B1(n_429),
.B2(n_421),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_556),
.B(n_421),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_491),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_538),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_514),
.B(n_553),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_556),
.B(n_424),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_491),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_SL g602 ( 
.A(n_495),
.B(n_429),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_500),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_488),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_489),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_489),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_504),
.A2(n_435),
.B1(n_431),
.B2(n_449),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_560),
.B(n_431),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_552),
.B(n_435),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_538),
.A2(n_551),
.B1(n_504),
.B2(n_555),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_490),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_552),
.B(n_449),
.Y(n_612)
);

AND2x2_ASAP7_75t_SL g613 ( 
.A(n_538),
.B(n_226),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_490),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_524),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_500),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_538),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_551),
.A2(n_451),
.B1(n_455),
.B2(n_450),
.Y(n_618)
);

BUFx4f_ASAP7_75t_L g619 ( 
.A(n_538),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_498),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_498),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_560),
.B(n_530),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_502),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_539),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_560),
.B(n_461),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_502),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_524),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_538),
.A2(n_379),
.B1(n_289),
.B2(n_265),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_552),
.B(n_450),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_560),
.B(n_451),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_538),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_524),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_524),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_534),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g635 ( 
.A1(n_536),
.A2(n_240),
.B(n_233),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_493),
.Y(n_636)
);

OAI21xp33_ASAP7_75t_SL g637 ( 
.A1(n_519),
.A2(n_320),
.B(n_310),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_519),
.B(n_458),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_534),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_534),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_534),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_548),
.B(n_458),
.Y(n_642)
);

OR2x6_ASAP7_75t_L g643 ( 
.A(n_492),
.B(n_520),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_548),
.B(n_460),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_549),
.B(n_460),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_493),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_493),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_496),
.Y(n_648)
);

INVx5_ASAP7_75t_L g649 ( 
.A(n_499),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_534),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_496),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_530),
.B(n_463),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_534),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_534),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_496),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_529),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_549),
.B(n_463),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_523),
.B(n_472),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_520),
.B(n_384),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_543),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_499),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_552),
.B(n_472),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_SL g663 ( 
.A1(n_495),
.A2(n_482),
.B1(n_409),
.B2(n_413),
.Y(n_663)
);

INVxp67_ASAP7_75t_SL g664 ( 
.A(n_547),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_543),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_543),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_543),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_501),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_529),
.B(n_473),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_543),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_537),
.B(n_473),
.Y(n_671)
);

BUFx6f_ASAP7_75t_SL g672 ( 
.A(n_566),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_537),
.B(n_476),
.Y(n_673)
);

NAND3xp33_ASAP7_75t_L g674 ( 
.A(n_543),
.B(n_252),
.C(n_240),
.Y(n_674)
);

BUFx4f_ASAP7_75t_L g675 ( 
.A(n_543),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_528),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_499),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_499),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_532),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_501),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_523),
.B(n_476),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_532),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_499),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_522),
.A2(n_414),
.B1(n_310),
.B2(n_322),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_563),
.B(n_478),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_499),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_529),
.B(n_478),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_501),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_563),
.B(n_479),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_494),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_532),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_565),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_565),
.B(n_481),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_532),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_567),
.B(n_214),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_567),
.B(n_214),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_540),
.B(n_222),
.Y(n_697)
);

AND3x1_ASAP7_75t_L g698 ( 
.A(n_513),
.B(n_564),
.C(n_559),
.Y(n_698)
);

INVx5_ASAP7_75t_L g699 ( 
.A(n_499),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_517),
.B(n_387),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_558),
.B(n_320),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_559),
.B(n_269),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_528),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_564),
.B(n_270),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_505),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_540),
.B(n_338),
.Y(n_706)
);

AND2x2_ASAP7_75t_SL g707 ( 
.A(n_506),
.B(n_226),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_532),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_499),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_505),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_540),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_541),
.B(n_252),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_525),
.B(n_214),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_541),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_SL g715 ( 
.A(n_566),
.B(n_268),
.Y(n_715)
);

NOR2x1p5_ASAP7_75t_L g716 ( 
.A(n_700),
.B(n_535),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_664),
.B(n_541),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_585),
.B(n_525),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_692),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_583),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_656),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_610),
.B(n_522),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_575),
.B(n_526),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_628),
.A2(n_613),
.B1(n_707),
.B2(n_642),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_630),
.B(n_495),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_588),
.B(n_526),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_596),
.B(n_531),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_625),
.B(n_495),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_600),
.B(n_495),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_605),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_605),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_608),
.B(n_531),
.Y(n_732)
);

NOR3xp33_ASAP7_75t_L g733 ( 
.A(n_692),
.B(n_545),
.C(n_544),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_620),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_622),
.B(n_707),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_604),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_569),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_685),
.B(n_545),
.C(n_544),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_606),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_689),
.B(n_550),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_620),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_638),
.B(n_550),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_676),
.B(n_506),
.Y(n_743)
);

O2A1O1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_599),
.A2(n_533),
.B(n_542),
.C(n_521),
.Y(n_744)
);

OAI22xp33_ASAP7_75t_L g745 ( 
.A1(n_628),
.A2(n_533),
.B1(n_542),
.B2(n_521),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_606),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_644),
.B(n_645),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_676),
.B(n_506),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_585),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_707),
.A2(n_558),
.B1(n_533),
.B2(n_542),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_621),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_597),
.B(n_601),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_621),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_597),
.B(n_521),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_611),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_586),
.B(n_557),
.Y(n_756)
);

AOI221xp5_ASAP7_75t_L g757 ( 
.A1(n_607),
.A2(n_322),
.B1(n_326),
.B2(n_349),
.C(n_350),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_611),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_613),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_587),
.B(n_546),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_619),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_656),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_586),
.B(n_557),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_626),
.Y(n_764)
);

NOR2xp67_ASAP7_75t_L g765 ( 
.A(n_700),
.B(n_557),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_619),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_614),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_L g768 ( 
.A(n_618),
.B(n_554),
.C(n_527),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_614),
.Y(n_769)
);

NOR3xp33_ASAP7_75t_L g770 ( 
.A(n_595),
.B(n_349),
.C(n_326),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_626),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_652),
.B(n_562),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_601),
.B(n_546),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_603),
.B(n_546),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_657),
.B(n_562),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_570),
.B(n_562),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_572),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_L g778 ( 
.A(n_577),
.B(n_499),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_613),
.B(n_506),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_603),
.B(n_527),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_572),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_659),
.A2(n_512),
.B1(n_511),
.B2(n_506),
.Y(n_782)
);

NAND3xp33_ASAP7_75t_L g783 ( 
.A(n_578),
.B(n_554),
.C(n_273),
.Y(n_783)
);

OR2x6_ASAP7_75t_L g784 ( 
.A(n_703),
.B(n_511),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_711),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_711),
.Y(n_786)
);

NAND3xp33_ASAP7_75t_L g787 ( 
.A(n_578),
.B(n_687),
.C(n_669),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_573),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_568),
.B(n_410),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_659),
.A2(n_279),
.B1(n_347),
.B2(n_342),
.Y(n_790)
);

AND2x6_ASAP7_75t_L g791 ( 
.A(n_619),
.B(n_709),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_616),
.B(n_511),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_714),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_713),
.B(n_511),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_658),
.B(n_511),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_573),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_713),
.B(n_512),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_579),
.B(n_418),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_616),
.B(n_512),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_659),
.A2(n_512),
.B1(n_214),
.B2(n_331),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_581),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_577),
.B(n_512),
.Y(n_802)
);

NOR2xp67_ASAP7_75t_L g803 ( 
.A(n_569),
.B(n_217),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_590),
.B(n_536),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_581),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_679),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_658),
.B(n_331),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_624),
.B(n_591),
.Y(n_808)
);

INVx5_ASAP7_75t_L g809 ( 
.A(n_598),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_714),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_590),
.B(n_536),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_702),
.B(n_704),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_592),
.B(n_423),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_681),
.B(n_254),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_681),
.B(n_254),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_679),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_694),
.A2(n_315),
.B(n_271),
.C(n_314),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_694),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_598),
.B(n_617),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_604),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_598),
.B(n_331),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_617),
.Y(n_822)
);

INVxp67_ASAP7_75t_SL g823 ( 
.A(n_617),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_703),
.B(n_350),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_697),
.B(n_271),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_SL g826 ( 
.A(n_602),
.B(n_624),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_708),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_SL g828 ( 
.A(n_602),
.B(n_672),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_708),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_682),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_682),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_659),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_631),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_671),
.B(n_272),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_631),
.B(n_331),
.Y(n_835)
);

NOR3xp33_ASAP7_75t_L g836 ( 
.A(n_693),
.B(n_360),
.C(n_356),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_659),
.A2(n_217),
.B1(n_384),
.B2(n_364),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_698),
.B(n_684),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_631),
.B(n_275),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_SL g840 ( 
.A(n_672),
.B(n_285),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_706),
.B(n_277),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_673),
.B(n_290),
.Y(n_842)
);

NAND2xp33_ASAP7_75t_L g843 ( 
.A(n_635),
.B(n_584),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_584),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_574),
.B(n_356),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_682),
.B(n_277),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_698),
.B(n_294),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_695),
.B(n_295),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_623),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_691),
.B(n_279),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_662),
.B(n_301),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_715),
.Y(n_852)
);

NOR2xp67_ASAP7_75t_L g853 ( 
.A(n_674),
.B(n_701),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_691),
.B(n_280),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_571),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_691),
.B(n_360),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_623),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_571),
.B(n_280),
.Y(n_858)
);

NAND2xp33_ASAP7_75t_L g859 ( 
.A(n_584),
.B(n_305),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_580),
.B(n_282),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_580),
.B(n_282),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_580),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_636),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_637),
.B(n_283),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_637),
.B(n_283),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_701),
.B(n_361),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_636),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_646),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_643),
.B(n_314),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_646),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_677),
.B(n_307),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_709),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_696),
.B(n_309),
.Y(n_873)
);

OAI22xp33_ASAP7_75t_L g874 ( 
.A1(n_643),
.A2(n_366),
.B1(n_361),
.B2(n_362),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_643),
.B(n_315),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_627),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_643),
.B(n_325),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_677),
.B(n_312),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_672),
.B(n_316),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_643),
.B(n_325),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_712),
.B(n_342),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_574),
.A2(n_347),
.B1(n_383),
.B2(n_330),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_574),
.B(n_383),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_752),
.A2(n_629),
.B(n_612),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_719),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_784),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_721),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_804),
.A2(n_632),
.B(n_627),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_844),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_811),
.A2(n_787),
.B(n_780),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_843),
.A2(n_594),
.B(n_576),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_724),
.A2(n_709),
.B(n_653),
.C(n_650),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_771),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_809),
.B(n_677),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_812),
.A2(n_574),
.B1(n_593),
.B2(n_609),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_809),
.B(n_678),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_735),
.A2(n_370),
.B(n_371),
.C(n_377),
.Y(n_897)
);

INVxp67_ASAP7_75t_L g898 ( 
.A(n_776),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_749),
.B(n_663),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_734),
.A2(n_574),
.B1(n_576),
.B2(n_589),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_771),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_772),
.B(n_582),
.Y(n_902)
);

O2A1O1Ixp5_ASAP7_75t_L g903 ( 
.A1(n_723),
.A2(n_675),
.B(n_654),
.C(n_641),
.Y(n_903)
);

NAND3xp33_ASAP7_75t_L g904 ( 
.A(n_757),
.B(n_633),
.C(n_632),
.Y(n_904)
);

AOI21xp33_ASAP7_75t_L g905 ( 
.A1(n_834),
.A2(n_842),
.B(n_808),
.Y(n_905)
);

AND2x6_ASAP7_75t_L g906 ( 
.A(n_822),
.B(n_584),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_718),
.B(n_582),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_718),
.B(n_582),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_747),
.A2(n_653),
.B(n_654),
.C(n_650),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_794),
.B(n_362),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_784),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_722),
.B(n_589),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_806),
.Y(n_913)
);

BUFx8_ASAP7_75t_L g914 ( 
.A(n_756),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_743),
.B(n_678),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_721),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_823),
.A2(n_639),
.B(n_633),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_809),
.B(n_678),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_838),
.A2(n_674),
.B1(n_686),
.B2(n_683),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_809),
.A2(n_773),
.B(n_754),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_775),
.B(n_589),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_794),
.B(n_615),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_797),
.B(n_615),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_809),
.B(n_822),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_737),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_797),
.B(n_615),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_802),
.A2(n_665),
.B(n_641),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_806),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_774),
.A2(n_666),
.B(n_665),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_734),
.Y(n_930)
);

OAI321xp33_ASAP7_75t_L g931 ( 
.A1(n_790),
.A2(n_382),
.A3(n_377),
.B1(n_366),
.B2(n_367),
.C(n_370),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_765),
.B(n_367),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_824),
.B(n_634),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_763),
.B(n_808),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_741),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_763),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_824),
.B(n_634),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_741),
.A2(n_666),
.B(n_670),
.C(n_634),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_726),
.A2(n_670),
.B(n_667),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_751),
.Y(n_940)
);

AND2x4_ASAP7_75t_SL g941 ( 
.A(n_784),
.B(n_683),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_743),
.B(n_683),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_824),
.B(n_640),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_727),
.B(n_640),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_822),
.B(n_833),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_770),
.A2(n_371),
.B(n_382),
.C(n_640),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_866),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_751),
.Y(n_948)
);

AOI21x1_ASAP7_75t_L g949 ( 
.A1(n_839),
.A2(n_648),
.B(n_647),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_732),
.B(n_667),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_816),
.A2(n_667),
.B(n_686),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_743),
.B(n_686),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_818),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_748),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_795),
.A2(n_710),
.B(n_705),
.C(n_688),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_748),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_753),
.A2(n_584),
.B1(n_660),
.B2(n_319),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_844),
.Y(n_958)
);

OAI21xp33_ASAP7_75t_L g959 ( 
.A1(n_814),
.A2(n_323),
.B(n_318),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_818),
.Y(n_960)
);

OR2x6_ASAP7_75t_L g961 ( 
.A(n_784),
.B(n_660),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_748),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_716),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_759),
.A2(n_660),
.B1(n_332),
.B2(n_335),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_826),
.B(n_660),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_717),
.A2(n_690),
.B(n_651),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_760),
.A2(n_819),
.B(n_822),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_822),
.A2(n_690),
.B(n_651),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_764),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_815),
.B(n_647),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_833),
.B(n_690),
.Y(n_971)
);

BUFx12f_ASAP7_75t_L g972 ( 
.A(n_716),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_829),
.Y(n_973)
);

BUFx4f_ASAP7_75t_L g974 ( 
.A(n_845),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_764),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_785),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_853),
.B(n_655),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_SL g978 ( 
.A(n_828),
.B(n_649),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_789),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_838),
.B(n_328),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_833),
.A2(n_690),
.B(n_668),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_740),
.B(n_680),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_833),
.B(n_759),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_792),
.B(n_680),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_799),
.B(n_688),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_856),
.B(n_705),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_827),
.A2(n_661),
.B(n_649),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_857),
.A2(n_260),
.B(n_308),
.C(n_363),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_785),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_762),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_829),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_866),
.B(n_798),
.Y(n_992)
);

AO22x1_ASAP7_75t_L g993 ( 
.A1(n_813),
.A2(n_355),
.B1(n_336),
.B2(n_337),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_827),
.A2(n_793),
.B(n_786),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_845),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_856),
.B(n_345),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_820),
.B(n_351),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_786),
.A2(n_661),
.B(n_649),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_793),
.A2(n_661),
.B(n_649),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_820),
.B(n_353),
.Y(n_1000)
);

AO21x1_ASAP7_75t_L g1001 ( 
.A1(n_729),
.A2(n_308),
.B(n_260),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_733),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_742),
.B(n_354),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_845),
.Y(n_1004)
);

NAND2x1p5_ASAP7_75t_L g1005 ( 
.A(n_736),
.B(n_649),
.Y(n_1005)
);

O2A1O1Ixp5_ASAP7_75t_L g1006 ( 
.A1(n_851),
.A2(n_505),
.B(n_508),
.C(n_515),
.Y(n_1006)
);

OAI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_882),
.A2(n_376),
.B1(n_365),
.B2(n_373),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_810),
.A2(n_699),
.B(n_661),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_750),
.B(n_359),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_810),
.A2(n_699),
.B(n_661),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_817),
.A2(n_508),
.B(n_515),
.C(n_375),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_840),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_768),
.B(n_378),
.Y(n_1013)
);

INVx5_ASAP7_75t_L g1014 ( 
.A(n_791),
.Y(n_1014)
);

AOI21x1_ASAP7_75t_L g1015 ( 
.A1(n_871),
.A2(n_515),
.B(n_508),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_878),
.A2(n_699),
.B(n_661),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_736),
.B(n_649),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_736),
.B(n_849),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_864),
.A2(n_699),
.B(n_348),
.C(n_291),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_849),
.B(n_699),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_846),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_779),
.A2(n_292),
.B1(n_198),
.B2(n_199),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_807),
.B(n_699),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_883),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_782),
.B(n_197),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_874),
.B(n_738),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_832),
.A2(n_296),
.B1(n_205),
.B2(n_208),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_852),
.B(n_18),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_825),
.B(n_200),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_841),
.B(n_213),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_876),
.A2(n_304),
.B(n_219),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_830),
.B(n_21),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_876),
.A2(n_311),
.B(n_225),
.Y(n_1033)
);

O2A1O1Ixp5_ASAP7_75t_L g1034 ( 
.A1(n_881),
.A2(n_518),
.B(n_516),
.C(n_497),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_855),
.A2(n_313),
.B(n_229),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_720),
.B(n_215),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_762),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_879),
.B(n_23),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_831),
.B(n_24),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_730),
.B(n_235),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_872),
.Y(n_1041)
);

AND2x4_ASAP7_75t_SL g1042 ( 
.A(n_836),
.B(n_348),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_855),
.A2(n_334),
.B1(n_239),
.B2(n_241),
.Y(n_1043)
);

INVx11_ASAP7_75t_L g1044 ( 
.A(n_791),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_862),
.A2(n_341),
.B(n_246),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_847),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_832),
.A2(n_344),
.B1(n_257),
.B2(n_258),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_730),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_731),
.B(n_236),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_848),
.B(n_25),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_850),
.A2(n_854),
.B(n_860),
.C(n_861),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_869),
.A2(n_259),
.B(n_262),
.C(n_267),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_739),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_844),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_778),
.A2(n_352),
.B(n_288),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_873),
.B(n_27),
.Y(n_1056)
);

OAI21xp33_ASAP7_75t_L g1057 ( 
.A1(n_837),
.A2(n_278),
.B(n_293),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_858),
.A2(n_28),
.B(n_30),
.C(n_36),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_761),
.B(n_766),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_744),
.A2(n_372),
.B(n_333),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_898),
.B(n_783),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_898),
.B(n_803),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_992),
.B(n_800),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_930),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_935),
.B(n_746),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_979),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_974),
.B(n_761),
.Y(n_1067)
);

AOI221xp5_ASAP7_75t_L g1068 ( 
.A1(n_905),
.A2(n_865),
.B1(n_745),
.B2(n_875),
.C(n_880),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_913),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_914),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_885),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_920),
.A2(n_778),
.B(n_766),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_889),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_940),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_948),
.B(n_755),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_925),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1056),
.A2(n_728),
.B1(n_725),
.B2(n_791),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_1002),
.B(n_877),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_914),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_928),
.Y(n_1080)
);

BUFx12f_ASAP7_75t_L g1081 ( 
.A(n_972),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_1056),
.A2(n_755),
.B1(n_758),
.B2(n_767),
.Y(n_1082)
);

BUFx8_ASAP7_75t_L g1083 ( 
.A(n_963),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_936),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_947),
.B(n_758),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_974),
.B(n_761),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_980),
.B(n_767),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_890),
.A2(n_950),
.B(n_944),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_953),
.Y(n_1089)
);

AO31x2_ASAP7_75t_L g1090 ( 
.A1(n_1001),
.A2(n_769),
.A3(n_870),
.B(n_868),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_1002),
.B(n_769),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1026),
.A2(n_844),
.B1(n_761),
.B2(n_766),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_889),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_1050),
.A2(n_859),
.B(n_835),
.C(n_821),
.Y(n_1094)
);

INVx3_ASAP7_75t_SL g1095 ( 
.A(n_1046),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_902),
.A2(n_761),
.B(n_766),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_1007),
.A2(n_1028),
.B(n_1038),
.C(n_1003),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_969),
.A2(n_844),
.B1(n_766),
.B2(n_777),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_899),
.B(n_777),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_1013),
.A2(n_1028),
.B(n_912),
.C(n_946),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_1004),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_960),
.Y(n_1102)
);

OR2x6_ASAP7_75t_SL g1103 ( 
.A(n_934),
.B(n_298),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_1013),
.A2(n_872),
.B(n_859),
.C(n_781),
.Y(n_1104)
);

INVx2_ASAP7_75t_SL g1105 ( 
.A(n_1012),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_1007),
.A2(n_805),
.B(n_788),
.C(n_796),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_902),
.A2(n_888),
.B(n_1051),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_975),
.A2(n_989),
.B1(n_976),
.B2(n_907),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_915),
.B(n_781),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_915),
.B(n_942),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_908),
.A2(n_796),
.B1(n_788),
.B2(n_801),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1003),
.A2(n_805),
.B(n_801),
.C(n_870),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_897),
.A2(n_868),
.B1(n_867),
.B2(n_863),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_889),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_995),
.B(n_867),
.Y(n_1115)
);

NOR3xp33_ASAP7_75t_L g1116 ( 
.A(n_993),
.B(n_863),
.C(n_386),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_893),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_973),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_942),
.B(n_791),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_901),
.B(n_791),
.Y(n_1120)
);

NAND2xp33_ASAP7_75t_SL g1121 ( 
.A(n_889),
.B(n_339),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_887),
.B(n_385),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_912),
.A2(n_380),
.B(n_346),
.C(n_348),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1024),
.B(n_39),
.Y(n_1124)
);

AOI33xp33_ASAP7_75t_L g1125 ( 
.A1(n_910),
.A2(n_40),
.A3(n_42),
.B1(n_47),
.B2(n_49),
.B3(n_53),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_991),
.B(n_40),
.Y(n_1126)
);

O2A1O1Ixp5_ASAP7_75t_L g1127 ( 
.A1(n_1060),
.A2(n_42),
.B(n_47),
.C(n_49),
.Y(n_1127)
);

AO32x1_ASAP7_75t_L g1128 ( 
.A1(n_957),
.A2(n_54),
.A3(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_958),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_994),
.B(n_55),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_997),
.B(n_58),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_951),
.A2(n_518),
.B(n_516),
.Y(n_1132)
);

AOI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1015),
.A2(n_518),
.B(n_516),
.Y(n_1133)
);

NOR3xp33_ASAP7_75t_SL g1134 ( 
.A(n_959),
.B(n_60),
.C(n_61),
.Y(n_1134)
);

AOI21xp33_ASAP7_75t_L g1135 ( 
.A1(n_931),
.A2(n_60),
.B(n_63),
.Y(n_1135)
);

BUFx2_ASAP7_75t_SL g1136 ( 
.A(n_1014),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1048),
.Y(n_1137)
);

O2A1O1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_996),
.A2(n_67),
.B(n_70),
.C(n_71),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_1000),
.B(n_74),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_954),
.B(n_75),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_887),
.B(n_916),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_921),
.A2(n_518),
.B(n_516),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_956),
.B(n_91),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_962),
.B(n_518),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1053),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_916),
.B(n_518),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_990),
.B(n_516),
.Y(n_1147)
);

BUFx4f_ASAP7_75t_L g1148 ( 
.A(n_961),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_903),
.A2(n_369),
.B(n_516),
.Y(n_1149)
);

BUFx12f_ASAP7_75t_L g1150 ( 
.A(n_961),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_932),
.B(n_494),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_886),
.B(n_497),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_886),
.B(n_497),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1032),
.A2(n_497),
.B(n_494),
.C(n_112),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_990),
.Y(n_1155)
);

INVxp67_ASAP7_75t_L g1156 ( 
.A(n_1032),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_897),
.A2(n_497),
.B(n_494),
.C(n_116),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_911),
.B(n_933),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_961),
.B(n_99),
.Y(n_1159)
);

AOI21x1_ASAP7_75t_L g1160 ( 
.A1(n_949),
.A2(n_494),
.B(n_117),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1039),
.A2(n_494),
.B(n_118),
.C(n_120),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_952),
.B(n_105),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_884),
.A2(n_123),
.B(n_125),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_911),
.B(n_127),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1021),
.A2(n_130),
.B(n_133),
.C(n_134),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_958),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_937),
.B(n_136),
.Y(n_1167)
);

OAI21xp33_ASAP7_75t_L g1168 ( 
.A1(n_1031),
.A2(n_145),
.B(n_148),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1039),
.A2(n_151),
.B(n_152),
.C(n_153),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1037),
.B(n_154),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_943),
.B(n_155),
.Y(n_1171)
);

OAI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1009),
.A2(n_1025),
.B1(n_1047),
.B2(n_1027),
.Y(n_1172)
);

AOI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1059),
.A2(n_891),
.B(n_971),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1037),
.B(n_1029),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_895),
.A2(n_163),
.B(n_164),
.C(n_167),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_958),
.Y(n_1176)
);

CKINVDCx6p67_ASAP7_75t_R g1177 ( 
.A(n_1014),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1058),
.A2(n_177),
.B(n_180),
.C(n_182),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1041),
.B(n_185),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1054),
.Y(n_1180)
);

BUFx12f_ASAP7_75t_L g1181 ( 
.A(n_1054),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1033),
.A2(n_193),
.B(n_1030),
.C(n_1052),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_965),
.B(n_1054),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1044),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_982),
.A2(n_927),
.B(n_965),
.C(n_929),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1041),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_L g1187 ( 
.A(n_988),
.B(n_964),
.C(n_982),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1054),
.B(n_1014),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_900),
.A2(n_941),
.B1(n_919),
.B2(n_1057),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_945),
.A2(n_971),
.B(n_939),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_919),
.B(n_984),
.Y(n_1191)
);

O2A1O1Ixp5_ASAP7_75t_L g1192 ( 
.A1(n_903),
.A2(n_1006),
.B(n_909),
.C(n_1034),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_945),
.A2(n_924),
.B(n_967),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_977),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_922),
.A2(n_926),
.B(n_923),
.C(n_938),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_R g1196 ( 
.A(n_978),
.B(n_1014),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_985),
.B(n_970),
.Y(n_1197)
);

BUFx12f_ASAP7_75t_L g1198 ( 
.A(n_906),
.Y(n_1198)
);

INVx4_ASAP7_75t_L g1199 ( 
.A(n_906),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_986),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1042),
.B(n_1018),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_924),
.A2(n_917),
.B(n_966),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_983),
.B(n_906),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_906),
.Y(n_1204)
);

OAI21xp33_ASAP7_75t_L g1205 ( 
.A1(n_1022),
.A2(n_1043),
.B(n_1040),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_983),
.B(n_906),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_1036),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_892),
.B(n_1017),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_1049),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_968),
.A2(n_981),
.B(n_1020),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1023),
.B(n_904),
.Y(n_1211)
);

NAND2xp33_ASAP7_75t_L g1212 ( 
.A(n_1005),
.B(n_894),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1083),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1078),
.B(n_1023),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1069),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1160),
.A2(n_1034),
.B(n_1006),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1080),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1156),
.A2(n_1055),
.B1(n_1017),
.B2(n_1019),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1066),
.B(n_1035),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1097),
.A2(n_1019),
.B(n_1011),
.C(n_1045),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1064),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1107),
.A2(n_1059),
.B(n_896),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1088),
.A2(n_894),
.B(n_896),
.Y(n_1223)
);

AOI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1207),
.A2(n_918),
.B1(n_1005),
.B2(n_987),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1092),
.A2(n_1016),
.A3(n_998),
.B(n_999),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1099),
.B(n_955),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1074),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1133),
.A2(n_1008),
.B(n_1010),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1065),
.Y(n_1229)
);

NOR2xp67_ASAP7_75t_L g1230 ( 
.A(n_1071),
.B(n_918),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1076),
.Y(n_1231)
);

O2A1O1Ixp5_ASAP7_75t_SL g1232 ( 
.A1(n_1211),
.A2(n_1082),
.B(n_1183),
.C(n_1092),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1208),
.A2(n_1096),
.B(n_1072),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1089),
.Y(n_1234)
);

BUFx5_ASAP7_75t_L g1235 ( 
.A(n_1198),
.Y(n_1235)
);

O2A1O1Ixp5_ASAP7_75t_SL g1236 ( 
.A1(n_1082),
.A2(n_1108),
.B(n_1149),
.C(n_1209),
.Y(n_1236)
);

OAI22x1_ASAP7_75t_L g1237 ( 
.A1(n_1061),
.A2(n_1143),
.B1(n_1095),
.B2(n_1131),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_1084),
.B(n_1105),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1111),
.A2(n_1210),
.A3(n_1104),
.B(n_1113),
.Y(n_1239)
);

OAI22x1_ASAP7_75t_L g1240 ( 
.A1(n_1143),
.A2(n_1139),
.B1(n_1062),
.B2(n_1189),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1102),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1208),
.A2(n_1108),
.B(n_1185),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1065),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1091),
.B(n_1200),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1085),
.B(n_1087),
.Y(n_1245)
);

OA21x2_ASAP7_75t_L g1246 ( 
.A1(n_1192),
.A2(n_1142),
.B(n_1190),
.Y(n_1246)
);

AO32x2_ASAP7_75t_L g1247 ( 
.A1(n_1098),
.A2(n_1111),
.A3(n_1113),
.B1(n_1155),
.B2(n_1128),
.Y(n_1247)
);

NAND2xp33_ASAP7_75t_SL g1248 ( 
.A(n_1196),
.B(n_1199),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1063),
.B(n_1115),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1103),
.B(n_1110),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1075),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1205),
.A2(n_1187),
.B(n_1168),
.C(n_1182),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1202),
.A2(n_1173),
.B(n_1193),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1194),
.B(n_1101),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1077),
.A2(n_1068),
.B(n_1094),
.C(n_1134),
.Y(n_1255)
);

AO21x1_ASAP7_75t_L g1256 ( 
.A1(n_1130),
.A2(n_1172),
.B(n_1191),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1081),
.Y(n_1257)
);

OA21x2_ASAP7_75t_L g1258 ( 
.A1(n_1132),
.A2(n_1191),
.B(n_1154),
.Y(n_1258)
);

INVx5_ASAP7_75t_L g1259 ( 
.A(n_1204),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1098),
.A2(n_1197),
.A3(n_1120),
.B(n_1175),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1116),
.A2(n_1070),
.B1(n_1159),
.B2(n_1079),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1075),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1181),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1138),
.A2(n_1130),
.B(n_1161),
.C(n_1169),
.Y(n_1264)
);

OAI21xp33_ASAP7_75t_L g1265 ( 
.A1(n_1125),
.A2(n_1135),
.B(n_1123),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_SL g1266 ( 
.A1(n_1124),
.A2(n_1140),
.B1(n_1159),
.B2(n_1150),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1127),
.A2(n_1135),
.B(n_1165),
.C(n_1178),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1174),
.A2(n_1140),
.B(n_1157),
.C(n_1195),
.Y(n_1268)
);

BUFx10_ASAP7_75t_L g1269 ( 
.A(n_1170),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1186),
.B(n_1141),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_SL g1271 ( 
.A1(n_1199),
.A2(n_1204),
.B(n_1112),
.Y(n_1271)
);

AO31x2_ASAP7_75t_L g1272 ( 
.A1(n_1162),
.A2(n_1203),
.A3(n_1206),
.B(n_1117),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1137),
.Y(n_1273)
);

INVxp67_ASAP7_75t_SL g1274 ( 
.A(n_1204),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1212),
.A2(n_1162),
.B(n_1163),
.Y(n_1275)
);

BUFx8_ASAP7_75t_SL g1276 ( 
.A(n_1176),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1179),
.A2(n_1188),
.B(n_1106),
.Y(n_1277)
);

BUFx12f_ASAP7_75t_L g1278 ( 
.A(n_1073),
.Y(n_1278)
);

AOI31xp67_ASAP7_75t_L g1279 ( 
.A1(n_1179),
.A2(n_1146),
.A3(n_1147),
.B(n_1126),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1145),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1151),
.A2(n_1171),
.B(n_1167),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1118),
.Y(n_1282)
);

AOI221x1_ASAP7_75t_L g1283 ( 
.A1(n_1126),
.A2(n_1201),
.B1(n_1158),
.B2(n_1121),
.C(n_1164),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1119),
.A2(n_1067),
.B(n_1086),
.Y(n_1284)
);

AO21x2_ASAP7_75t_L g1285 ( 
.A1(n_1109),
.A2(n_1122),
.B(n_1119),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1148),
.A2(n_1109),
.B(n_1180),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1144),
.A2(n_1153),
.B(n_1152),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1090),
.A2(n_1128),
.A3(n_1136),
.B(n_1177),
.Y(n_1288)
);

AOI21x1_ASAP7_75t_SL g1289 ( 
.A1(n_1128),
.A2(n_1073),
.B(n_1180),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_SL g1290 ( 
.A1(n_1184),
.A2(n_1093),
.B(n_1114),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1093),
.A2(n_1114),
.B(n_1129),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1090),
.A2(n_1114),
.A3(n_1129),
.B(n_1166),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1090),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1160),
.A2(n_1133),
.B(n_1210),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1160),
.A2(n_1133),
.B(n_1210),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1107),
.A2(n_619),
.B(n_752),
.Y(n_1296)
);

O2A1O1Ixp5_ASAP7_75t_L g1297 ( 
.A1(n_1107),
.A2(n_1056),
.B(n_1100),
.C(n_905),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1160),
.A2(n_1133),
.B(n_1210),
.Y(n_1298)
);

AO22x2_ASAP7_75t_L g1299 ( 
.A1(n_1082),
.A2(n_808),
.B1(n_980),
.B2(n_1108),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1076),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1065),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1078),
.B(n_992),
.Y(n_1302)
);

INVxp67_ASAP7_75t_SL g1303 ( 
.A(n_1115),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1107),
.A2(n_619),
.B(n_752),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1084),
.B(n_936),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1084),
.B(n_934),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1149),
.A2(n_1107),
.B(n_1160),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1160),
.A2(n_1133),
.B(n_1210),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1156),
.A2(n_724),
.B1(n_1056),
.B2(n_1100),
.Y(n_1309)
);

O2A1O1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1097),
.A2(n_1056),
.B(n_1100),
.C(n_905),
.Y(n_1310)
);

AO21x2_ASAP7_75t_L g1311 ( 
.A1(n_1149),
.A2(n_1107),
.B(n_1160),
.Y(n_1311)
);

OAI22x1_ASAP7_75t_L g1312 ( 
.A1(n_1207),
.A2(n_979),
.B1(n_1056),
.B2(n_808),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1097),
.A2(n_1056),
.B(n_1100),
.C(n_905),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1066),
.Y(n_1314)
);

NAND2xp33_ASAP7_75t_SL g1315 ( 
.A(n_1196),
.B(n_1066),
.Y(n_1315)
);

AO31x2_ASAP7_75t_L g1316 ( 
.A1(n_1092),
.A2(n_1001),
.A3(n_1107),
.B(n_1082),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1065),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1092),
.A2(n_1001),
.A3(n_1107),
.B(n_1082),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1065),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1107),
.A2(n_619),
.B(n_752),
.Y(n_1320)
);

AOI221xp5_ASAP7_75t_L g1321 ( 
.A1(n_1097),
.A2(n_905),
.B1(n_504),
.B2(n_992),
.C(n_757),
.Y(n_1321)
);

AO31x2_ASAP7_75t_L g1322 ( 
.A1(n_1092),
.A2(n_1001),
.A3(n_1107),
.B(n_1082),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1110),
.B(n_1004),
.Y(n_1323)
);

INVxp67_ASAP7_75t_SL g1324 ( 
.A(n_1115),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1100),
.A2(n_1056),
.B(n_812),
.Y(n_1325)
);

BUFx8_ASAP7_75t_L g1326 ( 
.A(n_1079),
.Y(n_1326)
);

INVxp67_ASAP7_75t_SL g1327 ( 
.A(n_1115),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1084),
.B(n_934),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1084),
.B(n_936),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1084),
.B(n_936),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1110),
.B(n_1004),
.Y(n_1331)
);

O2A1O1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1097),
.A2(n_1056),
.B(n_1100),
.C(n_905),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1097),
.A2(n_1056),
.B(n_905),
.C(n_1100),
.Y(n_1333)
);

OR2x6_ASAP7_75t_L g1334 ( 
.A(n_1070),
.B(n_1081),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1107),
.A2(n_619),
.B(n_752),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1107),
.A2(n_619),
.B(n_752),
.Y(n_1336)
);

A2O1A1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1097),
.A2(n_1056),
.B(n_905),
.C(n_1100),
.Y(n_1337)
);

AO32x2_ASAP7_75t_L g1338 ( 
.A1(n_1108),
.A2(n_1092),
.A3(n_1082),
.B1(n_1098),
.B2(n_1111),
.Y(n_1338)
);

OAI22x1_ASAP7_75t_L g1339 ( 
.A1(n_1207),
.A2(n_979),
.B1(n_1056),
.B2(n_808),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1160),
.A2(n_1133),
.B(n_1210),
.Y(n_1340)
);

OR2x6_ASAP7_75t_L g1341 ( 
.A(n_1070),
.B(n_1081),
.Y(n_1341)
);

AO31x2_ASAP7_75t_L g1342 ( 
.A1(n_1092),
.A2(n_1001),
.A3(n_1107),
.B(n_1082),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1100),
.A2(n_1056),
.B(n_812),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1084),
.B(n_934),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1069),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1100),
.A2(n_1056),
.B(n_812),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1078),
.B(n_992),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1107),
.A2(n_619),
.B(n_752),
.Y(n_1348)
);

NOR2x1_ASAP7_75t_SL g1349 ( 
.A(n_1199),
.B(n_1204),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_SL g1350 ( 
.A(n_1066),
.B(n_569),
.Y(n_1350)
);

INVx4_ASAP7_75t_L g1351 ( 
.A(n_1198),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_SL g1352 ( 
.A(n_1066),
.B(n_569),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1107),
.A2(n_619),
.B(n_752),
.Y(n_1353)
);

INVx4_ASAP7_75t_SL g1354 ( 
.A(n_1095),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1100),
.A2(n_1056),
.B(n_812),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1069),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1107),
.A2(n_619),
.B(n_752),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1107),
.A2(n_619),
.B(n_752),
.Y(n_1358)
);

AO32x2_ASAP7_75t_L g1359 ( 
.A1(n_1108),
.A2(n_1092),
.A3(n_1082),
.B1(n_1098),
.B2(n_1111),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1078),
.A2(n_1056),
.B1(n_692),
.B2(n_979),
.Y(n_1360)
);

AO31x2_ASAP7_75t_L g1361 ( 
.A1(n_1092),
.A2(n_1001),
.A3(n_1107),
.B(n_1082),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1156),
.A2(n_724),
.B1(n_1056),
.B2(n_1100),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1066),
.B(n_692),
.Y(n_1363)
);

AOI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1078),
.A2(n_1056),
.B1(n_692),
.B2(n_979),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1160),
.A2(n_1133),
.B(n_1210),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_1066),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1100),
.A2(n_1056),
.B(n_812),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1107),
.A2(n_619),
.B(n_752),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1084),
.B(n_934),
.Y(n_1369)
);

AO31x2_ASAP7_75t_L g1370 ( 
.A1(n_1092),
.A2(n_1001),
.A3(n_1107),
.B(n_1082),
.Y(n_1370)
);

AOI221xp5_ASAP7_75t_SL g1371 ( 
.A1(n_1097),
.A2(n_1056),
.B1(n_1156),
.B2(n_1007),
.C(n_757),
.Y(n_1371)
);

BUFx4f_ASAP7_75t_L g1372 ( 
.A(n_1081),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1198),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_SL g1374 ( 
.A1(n_1299),
.A2(n_1309),
.B1(n_1362),
.B2(n_1266),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1221),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1302),
.B(n_1347),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1321),
.A2(n_1299),
.B1(n_1355),
.B2(n_1367),
.Y(n_1377)
);

INVx6_ASAP7_75t_L g1378 ( 
.A(n_1259),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1276),
.Y(n_1379)
);

BUFx10_ASAP7_75t_L g1380 ( 
.A(n_1363),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1227),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1278),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_SL g1383 ( 
.A1(n_1325),
.A2(n_1343),
.B1(n_1346),
.B2(n_1250),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1303),
.A2(n_1327),
.B1(n_1324),
.B2(n_1214),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1360),
.A2(n_1364),
.B(n_1313),
.Y(n_1385)
);

AOI21xp33_ASAP7_75t_L g1386 ( 
.A1(n_1310),
.A2(n_1332),
.B(n_1264),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1315),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1333),
.A2(n_1337),
.B1(n_1242),
.B2(n_1255),
.Y(n_1388)
);

CKINVDCx11_ASAP7_75t_R g1389 ( 
.A(n_1366),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_SL g1390 ( 
.A1(n_1249),
.A2(n_1244),
.B1(n_1312),
.B2(n_1339),
.Y(n_1390)
);

BUFx12f_ASAP7_75t_L g1391 ( 
.A(n_1314),
.Y(n_1391)
);

BUFx8_ASAP7_75t_L g1392 ( 
.A(n_1213),
.Y(n_1392)
);

CKINVDCx11_ASAP7_75t_R g1393 ( 
.A(n_1354),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1263),
.Y(n_1394)
);

BUFx12f_ASAP7_75t_L g1395 ( 
.A(n_1326),
.Y(n_1395)
);

CKINVDCx11_ASAP7_75t_R g1396 ( 
.A(n_1354),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1273),
.Y(n_1397)
);

INVx6_ASAP7_75t_L g1398 ( 
.A(n_1263),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1240),
.A2(n_1256),
.B1(n_1237),
.B2(n_1265),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1245),
.A2(n_1226),
.B1(n_1328),
.B2(n_1344),
.Y(n_1400)
);

INVx6_ASAP7_75t_L g1401 ( 
.A(n_1351),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1269),
.A2(n_1371),
.B1(n_1219),
.B2(n_1254),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_SL g1403 ( 
.A1(n_1269),
.A2(n_1218),
.B1(n_1331),
.B2(n_1323),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1280),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1306),
.A2(n_1369),
.B1(n_1262),
.B2(n_1251),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1305),
.Y(n_1406)
);

CKINVDCx14_ASAP7_75t_R g1407 ( 
.A(n_1372),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1229),
.A2(n_1262),
.B1(n_1251),
.B2(n_1243),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1351),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1350),
.A2(n_1352),
.B1(n_1261),
.B2(n_1323),
.Y(n_1410)
);

INVx4_ASAP7_75t_L g1411 ( 
.A(n_1372),
.Y(n_1411)
);

INVx3_ASAP7_75t_SL g1412 ( 
.A(n_1334),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1329),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1272),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1331),
.Y(n_1415)
);

INVx8_ASAP7_75t_L g1416 ( 
.A(n_1334),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1229),
.A2(n_1243),
.B1(n_1301),
.B2(n_1317),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1330),
.Y(n_1418)
);

AND2x4_ASAP7_75t_SL g1419 ( 
.A(n_1341),
.B(n_1373),
.Y(n_1419)
);

INVx3_ASAP7_75t_SL g1420 ( 
.A(n_1341),
.Y(n_1420)
);

INVx6_ASAP7_75t_L g1421 ( 
.A(n_1326),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_SL g1422 ( 
.A1(n_1349),
.A2(n_1235),
.B1(n_1373),
.B2(n_1317),
.Y(n_1422)
);

OAI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1238),
.A2(n_1300),
.B1(n_1231),
.B2(n_1319),
.Y(n_1423)
);

INVx6_ASAP7_75t_L g1424 ( 
.A(n_1235),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1235),
.Y(n_1425)
);

CKINVDCx11_ASAP7_75t_R g1426 ( 
.A(n_1235),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1252),
.A2(n_1267),
.B1(n_1268),
.B2(n_1224),
.Y(n_1427)
);

OAI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1301),
.A2(n_1319),
.B1(n_1283),
.B2(n_1230),
.Y(n_1428)
);

CKINVDCx11_ASAP7_75t_R g1429 ( 
.A(n_1257),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1270),
.B(n_1217),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1234),
.A2(n_1345),
.B1(n_1356),
.B2(n_1241),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1282),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1286),
.B(n_1290),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1285),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1248),
.A2(n_1258),
.B1(n_1293),
.B2(n_1304),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1297),
.A2(n_1348),
.B1(n_1368),
.B2(n_1336),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_SL g1437 ( 
.A1(n_1349),
.A2(n_1274),
.B1(n_1258),
.B2(n_1311),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1296),
.A2(n_1357),
.B1(n_1320),
.B2(n_1353),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_1291),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1272),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1335),
.A2(n_1358),
.B1(n_1307),
.B2(n_1275),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1284),
.A2(n_1222),
.B1(n_1277),
.B2(n_1287),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1236),
.A2(n_1220),
.B(n_1232),
.Y(n_1443)
);

NAND2x1p5_ASAP7_75t_L g1444 ( 
.A(n_1228),
.B(n_1233),
.Y(n_1444)
);

BUFx8_ASAP7_75t_L g1445 ( 
.A(n_1338),
.Y(n_1445)
);

BUFx8_ASAP7_75t_L g1446 ( 
.A(n_1338),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1338),
.A2(n_1359),
.B1(n_1281),
.B2(n_1223),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1292),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1271),
.A2(n_1359),
.B1(n_1246),
.B2(n_1289),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1359),
.A2(n_1247),
.B1(n_1246),
.B2(n_1260),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1279),
.A2(n_1247),
.B1(n_1316),
.B2(n_1361),
.Y(n_1451)
);

CKINVDCx11_ASAP7_75t_R g1452 ( 
.A(n_1292),
.Y(n_1452)
);

CKINVDCx11_ASAP7_75t_R g1453 ( 
.A(n_1288),
.Y(n_1453)
);

INVx3_ASAP7_75t_SL g1454 ( 
.A(n_1288),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1260),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1260),
.Y(n_1456)
);

BUFx12f_ASAP7_75t_L g1457 ( 
.A(n_1288),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1316),
.B(n_1370),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1239),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1239),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1247),
.Y(n_1461)
);

CKINVDCx6p67_ASAP7_75t_R g1462 ( 
.A(n_1316),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1318),
.A2(n_1370),
.B1(n_1361),
.B2(n_1342),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1318),
.B(n_1370),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1318),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1253),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1322),
.A2(n_1361),
.B1(n_1342),
.B2(n_1239),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1322),
.A2(n_1216),
.B1(n_1298),
.B2(n_1294),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1295),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1308),
.A2(n_1340),
.B1(n_1365),
.B2(n_1225),
.Y(n_1470)
);

BUFx4f_ASAP7_75t_SL g1471 ( 
.A(n_1225),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1321),
.A2(n_905),
.B1(n_1299),
.B2(n_1325),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1259),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1360),
.A2(n_1364),
.B1(n_979),
.B2(n_1056),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1372),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1272),
.Y(n_1476)
);

BUFx2_ASAP7_75t_SL g1477 ( 
.A(n_1366),
.Y(n_1477)
);

OAI22xp33_ASAP7_75t_R g1478 ( 
.A1(n_1363),
.A2(n_504),
.B1(n_381),
.B2(n_266),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1302),
.B(n_1347),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1276),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1259),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1321),
.A2(n_905),
.B1(n_1299),
.B2(n_1325),
.Y(n_1482)
);

BUFx12f_ASAP7_75t_L g1483 ( 
.A(n_1314),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1215),
.Y(n_1484)
);

CKINVDCx11_ASAP7_75t_R g1485 ( 
.A(n_1366),
.Y(n_1485)
);

BUFx10_ASAP7_75t_L g1486 ( 
.A(n_1363),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1360),
.A2(n_1364),
.B1(n_1056),
.B2(n_1343),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1302),
.B(n_1347),
.Y(n_1488)
);

CKINVDCx11_ASAP7_75t_R g1489 ( 
.A(n_1366),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_SL g1490 ( 
.A1(n_1299),
.A2(n_495),
.B1(n_399),
.B2(n_409),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1321),
.A2(n_905),
.B1(n_1299),
.B2(n_1325),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1321),
.A2(n_905),
.B1(n_1299),
.B2(n_1325),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1276),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1305),
.B(n_1329),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1302),
.B(n_1347),
.Y(n_1495)
);

BUFx10_ASAP7_75t_L g1496 ( 
.A(n_1363),
.Y(n_1496)
);

OAI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1360),
.A2(n_1364),
.B1(n_724),
.B2(n_1343),
.Y(n_1497)
);

BUFx3_ASAP7_75t_L g1498 ( 
.A(n_1276),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1221),
.Y(n_1499)
);

INVx6_ASAP7_75t_L g1500 ( 
.A(n_1259),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1305),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1305),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1276),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1321),
.A2(n_905),
.B1(n_1299),
.B2(n_1325),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1221),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1221),
.Y(n_1506)
);

CKINVDCx11_ASAP7_75t_R g1507 ( 
.A(n_1366),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_SL g1508 ( 
.A1(n_1299),
.A2(n_495),
.B1(n_399),
.B2(n_409),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1360),
.A2(n_1364),
.B1(n_1056),
.B2(n_1343),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1215),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1221),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1221),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1448),
.B(n_1425),
.Y(n_1513)
);

INVx4_ASAP7_75t_SL g1514 ( 
.A(n_1471),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1375),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1381),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1416),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1400),
.B(n_1384),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1440),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1426),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1487),
.A2(n_1509),
.B(n_1474),
.Y(n_1521)
);

INVxp67_ASAP7_75t_L g1522 ( 
.A(n_1418),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1499),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1424),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1424),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1505),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1424),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1506),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1457),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1461),
.B(n_1458),
.Y(n_1530)
);

AOI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1478),
.A2(n_1374),
.B1(n_1385),
.B2(n_1497),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1443),
.A2(n_1441),
.B(n_1464),
.Y(n_1532)
);

AO21x2_ASAP7_75t_L g1533 ( 
.A1(n_1451),
.A2(n_1434),
.B(n_1428),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1414),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1459),
.B(n_1465),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1414),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1476),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1466),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1450),
.B(n_1511),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1476),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1406),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1466),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1380),
.B(n_1486),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1416),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1400),
.B(n_1376),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1512),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1397),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1404),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1388),
.A2(n_1497),
.B(n_1427),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1416),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1444),
.A2(n_1441),
.B(n_1438),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1389),
.Y(n_1552)
);

AO21x2_ASAP7_75t_L g1553 ( 
.A1(n_1428),
.A2(n_1436),
.B(n_1467),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1432),
.Y(n_1554)
);

INVxp33_ASAP7_75t_L g1555 ( 
.A(n_1494),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1430),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1484),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1510),
.Y(n_1558)
);

INVxp67_ASAP7_75t_L g1559 ( 
.A(n_1501),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1423),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1479),
.B(n_1488),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1423),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1405),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1405),
.Y(n_1564)
);

NAND3xp33_ASAP7_75t_L g1565 ( 
.A(n_1383),
.B(n_1504),
.C(n_1472),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1456),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1502),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1408),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1408),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1417),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1417),
.Y(n_1571)
);

INVx4_ASAP7_75t_L g1572 ( 
.A(n_1412),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1445),
.Y(n_1573)
);

OA21x2_ASAP7_75t_L g1574 ( 
.A1(n_1463),
.A2(n_1438),
.B(n_1468),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1445),
.Y(n_1575)
);

AO21x2_ASAP7_75t_L g1576 ( 
.A1(n_1436),
.A2(n_1449),
.B(n_1460),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1455),
.B(n_1463),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1446),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_1485),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1413),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1446),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1433),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1462),
.B(n_1454),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1431),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1387),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1431),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1490),
.A2(n_1508),
.B1(n_1504),
.B2(n_1492),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1454),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1386),
.A2(n_1377),
.B(n_1492),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1472),
.A2(n_1482),
.B1(n_1491),
.B2(n_1377),
.Y(n_1590)
);

AOI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1482),
.A2(n_1491),
.B1(n_1390),
.B2(n_1402),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1495),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1415),
.Y(n_1593)
);

INVx4_ASAP7_75t_L g1594 ( 
.A(n_1412),
.Y(n_1594)
);

AOI21xp33_ASAP7_75t_L g1595 ( 
.A1(n_1399),
.A2(n_1439),
.B(n_1403),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1447),
.B(n_1420),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1415),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1447),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1410),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1419),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1419),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1453),
.A2(n_1452),
.B1(n_1496),
.B2(n_1380),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1442),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1469),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1444),
.A2(n_1468),
.B(n_1442),
.Y(n_1605)
);

INVx4_ASAP7_75t_L g1606 ( 
.A(n_1420),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1469),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1409),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1435),
.B(n_1470),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1437),
.Y(n_1610)
);

BUFx8_ASAP7_75t_L g1611 ( 
.A(n_1395),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1378),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1435),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1409),
.Y(n_1614)
);

OAI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1549),
.A2(n_1422),
.B(n_1407),
.Y(n_1615)
);

AOI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1531),
.A2(n_1486),
.B1(n_1407),
.B2(n_1396),
.Y(n_1616)
);

OA21x2_ASAP7_75t_L g1617 ( 
.A1(n_1551),
.A2(n_1382),
.B(n_1475),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1589),
.A2(n_1473),
.B(n_1411),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1582),
.B(n_1394),
.Y(n_1619)
);

INVxp67_ASAP7_75t_L g1620 ( 
.A(n_1585),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1539),
.B(n_1394),
.Y(n_1621)
);

NAND4xp25_ASAP7_75t_L g1622 ( 
.A(n_1521),
.B(n_1498),
.C(n_1379),
.D(n_1480),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1592),
.B(n_1398),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1580),
.B(n_1477),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1530),
.B(n_1503),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1565),
.A2(n_1473),
.B(n_1493),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1515),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1543),
.B(n_1507),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1604),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1516),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1587),
.A2(n_1393),
.B1(n_1421),
.B2(n_1429),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1539),
.B(n_1421),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1574),
.B(n_1379),
.Y(n_1633)
);

A2O1A1Ixp33_ASAP7_75t_L g1634 ( 
.A1(n_1591),
.A2(n_1590),
.B(n_1518),
.C(n_1595),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1577),
.A2(n_1401),
.B1(n_1392),
.B2(n_1500),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1574),
.B(n_1609),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1574),
.B(n_1498),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1609),
.B(n_1480),
.Y(n_1638)
);

O2A1O1Ixp33_ASAP7_75t_SL g1639 ( 
.A1(n_1552),
.A2(n_1489),
.B(n_1392),
.C(n_1391),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1552),
.B(n_1483),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1530),
.B(n_1481),
.Y(n_1641)
);

AOI221xp5_ASAP7_75t_L g1642 ( 
.A1(n_1560),
.A2(n_1562),
.B1(n_1598),
.B2(n_1545),
.C(n_1570),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1532),
.B(n_1603),
.Y(n_1643)
);

AO32x2_ASAP7_75t_L g1644 ( 
.A1(n_1524),
.A2(n_1527),
.A3(n_1525),
.B1(n_1572),
.B2(n_1606),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1532),
.B(n_1577),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1556),
.B(n_1522),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1576),
.B(n_1598),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1563),
.A2(n_1564),
.B1(n_1584),
.B2(n_1586),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1541),
.B(n_1567),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1534),
.B(n_1536),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1561),
.B(n_1555),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1579),
.B(n_1572),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1576),
.B(n_1553),
.Y(n_1653)
);

A2O1A1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1610),
.A2(n_1599),
.B(n_1613),
.C(n_1596),
.Y(n_1654)
);

CKINVDCx6p67_ASAP7_75t_R g1655 ( 
.A(n_1579),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1553),
.A2(n_1551),
.B(n_1576),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1613),
.A2(n_1533),
.B(n_1605),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1535),
.B(n_1523),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1568),
.A2(n_1569),
.B1(n_1571),
.B2(n_1575),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1526),
.B(n_1528),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1514),
.B(n_1513),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1546),
.B(n_1547),
.Y(n_1662)
);

AO21x1_ASAP7_75t_L g1663 ( 
.A1(n_1596),
.A2(n_1548),
.B(n_1540),
.Y(n_1663)
);

OR2x6_ASAP7_75t_L g1664 ( 
.A(n_1588),
.B(n_1583),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1611),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1633),
.B(n_1637),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1650),
.Y(n_1667)
);

INVx3_ASAP7_75t_SL g1668 ( 
.A(n_1655),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1650),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1645),
.B(n_1537),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1645),
.B(n_1607),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1643),
.B(n_1533),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1658),
.B(n_1607),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1658),
.B(n_1559),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1644),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1622),
.B(n_1594),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1636),
.B(n_1519),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1661),
.B(n_1513),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1627),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1642),
.A2(n_1653),
.B1(n_1647),
.B2(n_1648),
.Y(n_1680)
);

NAND2x1p5_ASAP7_75t_SL g1681 ( 
.A(n_1653),
.B(n_1638),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1660),
.B(n_1566),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_SL g1683 ( 
.A1(n_1647),
.A2(n_1638),
.B1(n_1615),
.B2(n_1581),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1630),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1664),
.B(n_1542),
.Y(n_1685)
);

AND2x2_ASAP7_75t_SL g1686 ( 
.A(n_1661),
.B(n_1513),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1634),
.A2(n_1578),
.B1(n_1573),
.B2(n_1606),
.Y(n_1687)
);

NAND2xp33_ASAP7_75t_SL g1688 ( 
.A(n_1665),
.B(n_1520),
.Y(n_1688)
);

INVxp67_ASAP7_75t_L g1689 ( 
.A(n_1629),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1659),
.A2(n_1529),
.B1(n_1602),
.B2(n_1558),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1662),
.B(n_1651),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1631),
.A2(n_1529),
.B1(n_1632),
.B2(n_1663),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1620),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1663),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1656),
.A2(n_1614),
.B(n_1608),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1649),
.B(n_1538),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1625),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1695),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1675),
.B(n_1644),
.Y(n_1699)
);

INVx3_ASAP7_75t_SL g1700 ( 
.A(n_1668),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1670),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1668),
.B(n_1625),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1668),
.B(n_1655),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1675),
.B(n_1666),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1694),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1667),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1666),
.B(n_1644),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1681),
.B(n_1646),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1667),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1695),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1671),
.B(n_1644),
.Y(n_1711)
);

OAI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1680),
.A2(n_1654),
.B1(n_1616),
.B2(n_1635),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1669),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1686),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1694),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1669),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1681),
.B(n_1657),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1671),
.B(n_1644),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1670),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1689),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1681),
.A2(n_1626),
.B1(n_1619),
.B2(n_1618),
.C(n_1632),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1677),
.B(n_1641),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1673),
.B(n_1617),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1686),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1683),
.A2(n_1692),
.B1(n_1687),
.B2(n_1674),
.Y(n_1725)
);

OAI33xp33_ASAP7_75t_L g1726 ( 
.A1(n_1687),
.A2(n_1623),
.A3(n_1624),
.B1(n_1665),
.B2(n_1554),
.B3(n_1601),
.Y(n_1726)
);

OAI33xp33_ASAP7_75t_L g1727 ( 
.A1(n_1672),
.A2(n_1600),
.A3(n_1597),
.B1(n_1593),
.B2(n_1557),
.B3(n_1612),
.Y(n_1727)
);

INVx4_ASAP7_75t_L g1728 ( 
.A(n_1678),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1707),
.B(n_1689),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1719),
.B(n_1682),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1705),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1706),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1698),
.B(n_1679),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1724),
.B(n_1678),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1707),
.B(n_1697),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1706),
.Y(n_1736)
);

NOR2x1_ASAP7_75t_L g1737 ( 
.A(n_1714),
.B(n_1652),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1699),
.B(n_1693),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1699),
.B(n_1696),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_SL g1740 ( 
.A(n_1726),
.B(n_1594),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1706),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1709),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1720),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1698),
.B(n_1679),
.Y(n_1744)
);

INVx2_ASAP7_75t_SL g1745 ( 
.A(n_1724),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1720),
.Y(n_1746)
);

NAND2xp33_ASAP7_75t_R g1747 ( 
.A(n_1714),
.B(n_1676),
.Y(n_1747)
);

BUFx3_ASAP7_75t_L g1748 ( 
.A(n_1700),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1709),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1699),
.B(n_1696),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1705),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1709),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1710),
.B(n_1684),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1724),
.B(n_1678),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_R g1755 ( 
.A(n_1700),
.B(n_1611),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1711),
.B(n_1718),
.Y(n_1756)
);

NOR2xp67_ASAP7_75t_L g1757 ( 
.A(n_1724),
.B(n_1678),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1712),
.A2(n_1683),
.B1(n_1690),
.B2(n_1621),
.Y(n_1758)
);

OR2x6_ASAP7_75t_SL g1759 ( 
.A(n_1725),
.B(n_1717),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1724),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1710),
.B(n_1674),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1705),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1704),
.B(n_1685),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1705),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1701),
.B(n_1691),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1733),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1733),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1744),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1732),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1732),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1761),
.B(n_1708),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1761),
.B(n_1708),
.Y(n_1772)
);

NAND2x1p5_ASAP7_75t_L g1773 ( 
.A(n_1748),
.B(n_1714),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1737),
.B(n_1728),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1765),
.B(n_1708),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1765),
.B(n_1717),
.Y(n_1776)
);

NAND4xp75_ASAP7_75t_L g1777 ( 
.A(n_1759),
.B(n_1721),
.C(n_1640),
.D(n_1703),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1755),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1737),
.B(n_1728),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_1744),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1731),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1755),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1736),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1756),
.B(n_1728),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1753),
.B(n_1701),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1736),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1756),
.B(n_1763),
.Y(n_1787)
);

AND2x4_ASAP7_75t_SL g1788 ( 
.A(n_1734),
.B(n_1724),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1756),
.B(n_1728),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1753),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1765),
.B(n_1717),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1759),
.B(n_1713),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1743),
.Y(n_1793)
);

INVxp67_ASAP7_75t_L g1794 ( 
.A(n_1740),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1759),
.B(n_1713),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1741),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1743),
.Y(n_1797)
);

AND2x4_ASAP7_75t_SL g1798 ( 
.A(n_1734),
.B(n_1703),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1746),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1746),
.Y(n_1800)
);

INVx2_ASAP7_75t_SL g1801 ( 
.A(n_1748),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1731),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1763),
.B(n_1728),
.Y(n_1803)
);

NOR2x1_ASAP7_75t_L g1804 ( 
.A(n_1748),
.B(n_1628),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1741),
.Y(n_1805)
);

NAND2xp67_ASAP7_75t_L g1806 ( 
.A(n_1731),
.B(n_1715),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1742),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1742),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1738),
.B(n_1716),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1730),
.B(n_1722),
.Y(n_1810)
);

NOR2xp67_ASAP7_75t_SL g1811 ( 
.A(n_1760),
.B(n_1606),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1806),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1787),
.B(n_1734),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1787),
.B(n_1734),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1773),
.B(n_1734),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1769),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1773),
.B(n_1754),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1773),
.B(n_1754),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1766),
.B(n_1738),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1780),
.B(n_1767),
.Y(n_1820)
);

AOI211xp5_ASAP7_75t_L g1821 ( 
.A1(n_1792),
.A2(n_1725),
.B(n_1740),
.C(n_1712),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1768),
.B(n_1738),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1785),
.B(n_1730),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1769),
.Y(n_1824)
);

NOR3x1_ASAP7_75t_L g1825 ( 
.A(n_1777),
.B(n_1745),
.C(n_1700),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1788),
.B(n_1754),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1788),
.B(n_1754),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1784),
.B(n_1754),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1775),
.B(n_1749),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1784),
.B(n_1760),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1789),
.B(n_1760),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1775),
.B(n_1749),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1806),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_SL g1834 ( 
.A(n_1777),
.B(n_1700),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1790),
.B(n_1735),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1794),
.B(n_1700),
.Y(n_1836)
);

INVx3_ASAP7_75t_L g1837 ( 
.A(n_1798),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1797),
.B(n_1793),
.Y(n_1838)
);

NAND2x1_ASAP7_75t_L g1839 ( 
.A(n_1774),
.B(n_1760),
.Y(n_1839)
);

AND2x4_ASAP7_75t_L g1840 ( 
.A(n_1789),
.B(n_1757),
.Y(n_1840)
);

INVxp67_ASAP7_75t_L g1841 ( 
.A(n_1801),
.Y(n_1841)
);

INVx2_ASAP7_75t_SL g1842 ( 
.A(n_1798),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1770),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1781),
.Y(n_1844)
);

OAI221xp5_ASAP7_75t_L g1845 ( 
.A1(n_1795),
.A2(n_1758),
.B1(n_1747),
.B2(n_1721),
.C(n_1715),
.Y(n_1845)
);

INVx3_ASAP7_75t_L g1846 ( 
.A(n_1803),
.Y(n_1846)
);

AOI21x1_ASAP7_75t_L g1847 ( 
.A1(n_1804),
.A2(n_1762),
.B(n_1751),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1774),
.B(n_1760),
.Y(n_1848)
);

AOI222xp33_ASAP7_75t_L g1849 ( 
.A1(n_1845),
.A2(n_1758),
.B1(n_1772),
.B2(n_1771),
.C1(n_1726),
.C2(n_1727),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1834),
.A2(n_1782),
.B(n_1778),
.Y(n_1850)
);

OAI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1845),
.A2(n_1747),
.B1(n_1776),
.B2(n_1791),
.Y(n_1851)
);

INVx2_ASAP7_75t_SL g1852 ( 
.A(n_1837),
.Y(n_1852)
);

AOI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1821),
.A2(n_1727),
.B1(n_1715),
.B2(n_1723),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1816),
.Y(n_1854)
);

AOI211xp5_ASAP7_75t_SL g1855 ( 
.A1(n_1834),
.A2(n_1639),
.B(n_1800),
.C(n_1799),
.Y(n_1855)
);

OAI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1821),
.A2(n_1801),
.B(n_1779),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1816),
.Y(n_1857)
);

INVx2_ASAP7_75t_SL g1858 ( 
.A(n_1837),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1837),
.B(n_1763),
.Y(n_1859)
);

OAI22xp33_ASAP7_75t_SL g1860 ( 
.A1(n_1847),
.A2(n_1812),
.B1(n_1833),
.B2(n_1776),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1824),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1837),
.A2(n_1757),
.B1(n_1728),
.B2(n_1810),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1824),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1819),
.B(n_1810),
.Y(n_1864)
);

OAI32xp33_ASAP7_75t_L g1865 ( 
.A1(n_1819),
.A2(n_1791),
.A3(n_1779),
.B1(n_1809),
.B2(n_1745),
.Y(n_1865)
);

OAI221xp5_ASAP7_75t_L g1866 ( 
.A1(n_1847),
.A2(n_1812),
.B1(n_1833),
.B2(n_1820),
.C(n_1825),
.Y(n_1866)
);

AOI221xp5_ASAP7_75t_L g1867 ( 
.A1(n_1820),
.A2(n_1786),
.B1(n_1770),
.B2(n_1807),
.C(n_1805),
.Y(n_1867)
);

AOI211xp5_ASAP7_75t_L g1868 ( 
.A1(n_1825),
.A2(n_1811),
.B(n_1745),
.C(n_1807),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1841),
.B(n_1739),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1842),
.B(n_1803),
.Y(n_1870)
);

INVxp67_ASAP7_75t_L g1871 ( 
.A(n_1842),
.Y(n_1871)
);

AOI221xp5_ASAP7_75t_L g1872 ( 
.A1(n_1838),
.A2(n_1783),
.B1(n_1805),
.B2(n_1796),
.C(n_1786),
.Y(n_1872)
);

OAI21xp33_ASAP7_75t_SL g1873 ( 
.A1(n_1815),
.A2(n_1729),
.B(n_1735),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1843),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1841),
.B(n_1739),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1854),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1871),
.B(n_1838),
.Y(n_1877)
);

INVx3_ASAP7_75t_L g1878 ( 
.A(n_1859),
.Y(n_1878)
);

AOI221xp5_ASAP7_75t_L g1879 ( 
.A1(n_1851),
.A2(n_1812),
.B1(n_1833),
.B2(n_1822),
.C(n_1843),
.Y(n_1879)
);

AOI21xp33_ASAP7_75t_SL g1880 ( 
.A1(n_1866),
.A2(n_1842),
.B(n_1836),
.Y(n_1880)
);

AOI21xp33_ASAP7_75t_L g1881 ( 
.A1(n_1860),
.A2(n_1844),
.B(n_1832),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1849),
.B(n_1823),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1852),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1866),
.A2(n_1814),
.B1(n_1813),
.B2(n_1822),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1858),
.B(n_1813),
.Y(n_1885)
);

INVxp67_ASAP7_75t_SL g1886 ( 
.A(n_1850),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1857),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1853),
.A2(n_1844),
.B1(n_1818),
.B2(n_1815),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1861),
.Y(n_1889)
);

AOI332xp33_ASAP7_75t_L g1890 ( 
.A1(n_1863),
.A2(n_1846),
.A3(n_1835),
.B1(n_1815),
.B2(n_1817),
.B3(n_1818),
.C1(n_1848),
.C2(n_1840),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1855),
.B(n_1813),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1864),
.B(n_1823),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1874),
.Y(n_1893)
);

OAI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1856),
.A2(n_1873),
.B(n_1868),
.Y(n_1894)
);

OAI21xp5_ASAP7_75t_SL g1895 ( 
.A1(n_1867),
.A2(n_1818),
.B(n_1817),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1869),
.B(n_1829),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1878),
.B(n_1867),
.Y(n_1897)
);

AOI21xp33_ASAP7_75t_L g1898 ( 
.A1(n_1886),
.A2(n_1844),
.B(n_1872),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1880),
.B(n_1872),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1876),
.Y(n_1900)
);

NAND2x1_ASAP7_75t_L g1901 ( 
.A(n_1878),
.B(n_1817),
.Y(n_1901)
);

AOI31xp33_ASAP7_75t_SL g1902 ( 
.A1(n_1882),
.A2(n_1875),
.A3(n_1835),
.B(n_1832),
.Y(n_1902)
);

OAI221xp5_ASAP7_75t_L g1903 ( 
.A1(n_1888),
.A2(n_1862),
.B1(n_1870),
.B2(n_1829),
.C(n_1832),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1876),
.Y(n_1904)
);

AOI222xp33_ASAP7_75t_L g1905 ( 
.A1(n_1879),
.A2(n_1865),
.B1(n_1715),
.B2(n_1802),
.C1(n_1781),
.C2(n_1751),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1887),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1878),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1887),
.Y(n_1908)
);

NAND4xp75_ASAP7_75t_L g1909 ( 
.A(n_1894),
.B(n_1848),
.C(n_1826),
.D(n_1827),
.Y(n_1909)
);

NAND2x1p5_ASAP7_75t_L g1910 ( 
.A(n_1883),
.B(n_1611),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1907),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1907),
.Y(n_1912)
);

NOR3xp33_ASAP7_75t_L g1913 ( 
.A(n_1899),
.B(n_1881),
.C(n_1895),
.Y(n_1913)
);

OAI21xp5_ASAP7_75t_SL g1914 ( 
.A1(n_1899),
.A2(n_1891),
.B(n_1910),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1900),
.Y(n_1915)
);

OAI21xp33_ASAP7_75t_SL g1916 ( 
.A1(n_1905),
.A2(n_1891),
.B(n_1885),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1898),
.A2(n_1884),
.B1(n_1892),
.B2(n_1885),
.Y(n_1917)
);

NAND3xp33_ASAP7_75t_L g1918 ( 
.A(n_1897),
.B(n_1883),
.C(n_1877),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1910),
.B(n_1896),
.Y(n_1919)
);

AO22x1_ASAP7_75t_L g1920 ( 
.A1(n_1904),
.A2(n_1889),
.B1(n_1893),
.B2(n_1890),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1901),
.B(n_1896),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_SL g1922 ( 
.A(n_1913),
.B(n_1906),
.Y(n_1922)
);

OAI21xp33_ASAP7_75t_L g1923 ( 
.A1(n_1913),
.A2(n_1903),
.B(n_1908),
.Y(n_1923)
);

AOI221xp5_ASAP7_75t_L g1924 ( 
.A1(n_1916),
.A2(n_1889),
.B1(n_1902),
.B2(n_1909),
.C(n_1802),
.Y(n_1924)
);

OAI211xp5_ASAP7_75t_L g1925 ( 
.A1(n_1914),
.A2(n_1839),
.B(n_1846),
.C(n_1848),
.Y(n_1925)
);

AOI211xp5_ASAP7_75t_L g1926 ( 
.A1(n_1920),
.A2(n_1829),
.B(n_1826),
.C(n_1827),
.Y(n_1926)
);

AOI221xp5_ASAP7_75t_L g1927 ( 
.A1(n_1918),
.A2(n_1846),
.B1(n_1783),
.B2(n_1796),
.C(n_1751),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1922),
.Y(n_1928)
);

AOI221xp5_ASAP7_75t_L g1929 ( 
.A1(n_1924),
.A2(n_1917),
.B1(n_1921),
.B2(n_1912),
.C(n_1911),
.Y(n_1929)
);

OAI211xp5_ASAP7_75t_L g1930 ( 
.A1(n_1923),
.A2(n_1919),
.B(n_1915),
.C(n_1839),
.Y(n_1930)
);

AOI222xp33_ASAP7_75t_L g1931 ( 
.A1(n_1927),
.A2(n_1762),
.B1(n_1764),
.B2(n_1846),
.C1(n_1808),
.C2(n_1814),
.Y(n_1931)
);

AOI211xp5_ASAP7_75t_L g1932 ( 
.A1(n_1926),
.A2(n_1827),
.B(n_1826),
.C(n_1840),
.Y(n_1932)
);

NAND4xp25_ASAP7_75t_L g1933 ( 
.A(n_1925),
.B(n_1814),
.C(n_1840),
.D(n_1828),
.Y(n_1933)
);

AOI221x1_ASAP7_75t_L g1934 ( 
.A1(n_1923),
.A2(n_1840),
.B1(n_1831),
.B2(n_1830),
.C(n_1828),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1928),
.B(n_1828),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1930),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1929),
.B(n_1830),
.Y(n_1937)
);

NOR2x1_ASAP7_75t_L g1938 ( 
.A(n_1933),
.B(n_1934),
.Y(n_1938)
);

INVxp67_ASAP7_75t_L g1939 ( 
.A(n_1931),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1932),
.Y(n_1940)
);

AND2x4_ASAP7_75t_L g1941 ( 
.A(n_1935),
.B(n_1840),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1938),
.Y(n_1942)
);

INVxp67_ASAP7_75t_L g1943 ( 
.A(n_1937),
.Y(n_1943)
);

INVx3_ASAP7_75t_L g1944 ( 
.A(n_1941),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1944),
.Y(n_1945)
);

OAI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1945),
.A2(n_1942),
.B1(n_1943),
.B2(n_1939),
.Y(n_1946)
);

OR2x2_ASAP7_75t_L g1947 ( 
.A(n_1945),
.B(n_1944),
.Y(n_1947)
);

OAI22xp5_ASAP7_75t_SL g1948 ( 
.A1(n_1947),
.A2(n_1936),
.B1(n_1940),
.B2(n_1702),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1946),
.Y(n_1949)
);

HB1xp67_ASAP7_75t_L g1950 ( 
.A(n_1949),
.Y(n_1950)
);

AO21x1_ASAP7_75t_L g1951 ( 
.A1(n_1948),
.A2(n_1831),
.B(n_1830),
.Y(n_1951)
);

AOI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1950),
.A2(n_1831),
.B(n_1750),
.Y(n_1952)
);

O2A1O1Ixp33_ASAP7_75t_SL g1953 ( 
.A1(n_1952),
.A2(n_1951),
.B(n_1702),
.C(n_1752),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1953),
.A2(n_1739),
.B1(n_1750),
.B2(n_1729),
.Y(n_1954)
);

OAI221xp5_ASAP7_75t_R g1955 ( 
.A1(n_1954),
.A2(n_1811),
.B1(n_1729),
.B2(n_1735),
.C(n_1688),
.Y(n_1955)
);

AOI211xp5_ASAP7_75t_L g1956 ( 
.A1(n_1955),
.A2(n_1517),
.B(n_1544),
.C(n_1550),
.Y(n_1956)
);


endmodule