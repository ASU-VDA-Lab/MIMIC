module fake_jpeg_1319_n_296 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_227;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_270;
wire n_199;
wire n_112;
wire n_260;
wire n_176;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVxp67_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVxp33_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_3),
.B(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_44),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_48),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g130 ( 
.A(n_49),
.Y(n_130)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx4f_ASAP7_75t_SL g51 ( 
.A(n_25),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_51),
.Y(n_104)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_62),
.Y(n_100)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

NAND2x1_ASAP7_75t_SL g64 ( 
.A(n_16),
.B(n_0),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_64),
.B(n_11),
.C(n_12),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_21),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_70),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx2_ASAP7_75t_R g70 ( 
.A(n_22),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_26),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_74),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_19),
.B(n_1),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_79),
.Y(n_118)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_27),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_81),
.Y(n_117)
);

INVx2_ASAP7_75t_R g81 ( 
.A(n_19),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_23),
.B(n_2),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_87),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_41),
.B(n_14),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_41),
.B1(n_28),
.B2(n_29),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_89),
.A2(n_94),
.B1(n_96),
.B2(n_102),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_55),
.A2(n_23),
.B1(n_37),
.B2(n_36),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_28),
.B1(n_37),
.B2(n_36),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_29),
.B1(n_33),
.B2(n_32),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_99),
.A2(n_63),
.B1(n_60),
.B2(n_47),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_50),
.A2(n_33),
.B1(n_32),
.B2(n_30),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_74),
.A2(n_40),
.B1(n_5),
.B2(n_7),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_111),
.A2(n_114),
.B1(n_95),
.B2(n_113),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_52),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_73),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_132),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_81),
.A2(n_13),
.B1(n_15),
.B2(n_75),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_130),
.B(n_97),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_51),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_133),
.B(n_139),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_61),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_150),
.Y(n_167)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_46),
.B1(n_66),
.B2(n_64),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_137),
.B(n_140),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g138 ( 
.A(n_131),
.B(n_70),
.CI(n_53),
.CON(n_138),
.SN(n_138)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_119),
.C(n_110),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_51),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_160),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_147),
.B1(n_151),
.B2(n_127),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_132),
.A2(n_72),
.B1(n_65),
.B2(n_58),
.Y(n_147)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_118),
.B(n_86),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_149),
.B(n_156),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_83),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_99),
.A2(n_76),
.B1(n_49),
.B2(n_53),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_83),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_152),
.B(n_155),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_49),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_157),
.Y(n_169)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_107),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_96),
.B(n_98),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_158),
.B(n_163),
.Y(n_191)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_88),
.B(n_125),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_94),
.B(n_128),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_102),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_105),
.Y(n_162)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_106),
.B(n_129),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_164),
.Y(n_190)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_165),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_173),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_119),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_89),
.B(n_105),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_145),
.B(n_157),
.Y(n_193)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_178),
.B(n_135),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_121),
.C(n_123),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_192),
.C(n_144),
.Y(n_212)
);

AND2x6_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_116),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_186),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_147),
.A2(n_115),
.B1(n_123),
.B2(n_120),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_143),
.B1(n_144),
.B2(n_165),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_150),
.B(n_115),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_193),
.A2(n_175),
.B(n_186),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_191),
.A2(n_158),
.B1(n_142),
.B2(n_137),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_195),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_142),
.B1(n_141),
.B2(n_138),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_192),
.B(n_169),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_196),
.B(n_199),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_167),
.B(n_149),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_156),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_163),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_204),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_159),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_180),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_205),
.B(n_211),
.Y(n_227)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_162),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_209),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_177),
.B1(n_190),
.B2(n_168),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_172),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_212),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_170),
.A2(n_164),
.B1(n_146),
.B2(n_136),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_213),
.A2(n_182),
.B1(n_190),
.B2(n_183),
.Y(n_226)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_215),
.A2(n_218),
.B(n_229),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_193),
.A2(n_186),
.B(n_188),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_209),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_214),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_231),
.B1(n_203),
.B2(n_202),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_200),
.A2(n_187),
.B(n_178),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_200),
.A2(n_202),
.B1(n_205),
.B2(n_199),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_233),
.A2(n_236),
.B1(n_217),
.B2(n_224),
.Y(n_254)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_217),
.A2(n_229),
.B1(n_219),
.B2(n_223),
.Y(n_236)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_228),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_239),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_232),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_211),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_244),
.C(n_245),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_204),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_242),
.Y(n_255)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_212),
.C(n_196),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_195),
.C(n_194),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_247),
.Y(n_260)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

AOI321xp33_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_221),
.A3(n_215),
.B1(n_218),
.B2(n_222),
.C(n_219),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_251),
.B(n_238),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_240),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_257),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_239),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_234),
.A2(n_222),
.B1(n_221),
.B2(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_256),
.B(n_249),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_198),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_233),
.A2(n_208),
.B1(n_213),
.B2(n_210),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_258),
.B(n_246),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_206),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_237),
.Y(n_264)
);

XOR2x2_ASAP7_75t_L g261 ( 
.A(n_259),
.B(n_245),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_268),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_262),
.A2(n_265),
.B1(n_269),
.B2(n_270),
.Y(n_273)
);

XOR2x1_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_234),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_266),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_253),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_255),
.B(n_247),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_176),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_261),
.A2(n_250),
.B(n_251),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_242),
.B(n_226),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_252),
.C(n_253),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_258),
.C(n_172),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_235),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_263),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_189),
.B1(n_176),
.B2(n_181),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_248),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_242),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_279),
.B(n_280),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_271),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_283),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_273),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_286),
.A2(n_272),
.B(n_279),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_289),
.B(n_290),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_278),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_288),
.A2(n_276),
.A3(n_275),
.B1(n_154),
.B2(n_148),
.C1(n_177),
.C2(n_181),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_184),
.C(n_177),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_293),
.B(n_292),
.Y(n_294)
);

AOI221xp5_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_184),
.B1(n_168),
.B2(n_93),
.C(n_126),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_120),
.Y(n_296)
);


endmodule