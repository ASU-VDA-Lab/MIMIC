module fake_jpeg_29756_n_441 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_441);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_441;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_49),
.Y(n_91)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_21),
.B(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_15),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_51),
.B(n_59),
.Y(n_125)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_54),
.Y(n_138)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx2_ASAP7_75t_SL g96 ( 
.A(n_55),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_0),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_61),
.B(n_63),
.Y(n_126)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_17),
.B(n_1),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_64),
.B(n_65),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_69),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_16),
.B(n_1),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_83),
.C(n_25),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_19),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_75),
.B(n_78),
.Y(n_120)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_43),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_43),
.Y(n_82)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_16),
.B(n_1),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_27),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_19),
.B(n_2),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_88),
.B(n_38),
.Y(n_136)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_89),
.A2(n_31),
.B1(n_24),
.B2(n_39),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_47),
.A2(n_22),
.B1(n_41),
.B2(n_45),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_93),
.A2(n_97),
.B1(n_98),
.B2(n_116),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_49),
.A2(n_22),
.B1(n_41),
.B2(n_45),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_41),
.B1(n_45),
.B2(n_40),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_136),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_103),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_83),
.B1(n_87),
.B2(n_86),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_106),
.A2(n_117),
.B1(n_82),
.B2(n_69),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_73),
.A2(n_29),
.B1(n_30),
.B2(n_24),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_66),
.A2(n_29),
.B1(n_30),
.B2(n_24),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_67),
.A2(n_29),
.B1(n_30),
.B2(n_16),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_27),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_122),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_115),
.B(n_10),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_51),
.A2(n_25),
.B1(n_35),
.B2(n_40),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_39),
.B1(n_37),
.B2(n_31),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_50),
.B(n_35),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_55),
.A2(n_39),
.B1(n_37),
.B2(n_31),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_130),
.A2(n_54),
.B1(n_57),
.B2(n_52),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_56),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_133),
.A2(n_70),
.B1(n_62),
.B2(n_7),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_55),
.B(n_36),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_65),
.Y(n_154)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

INVx13_ASAP7_75t_L g201 ( 
.A(n_141),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_91),
.B(n_58),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_142),
.B(n_155),
.Y(n_197)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_143),
.Y(n_202)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_152),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_91),
.A2(n_84),
.B1(n_72),
.B2(n_89),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_148),
.A2(n_157),
.B1(n_172),
.B2(n_173),
.Y(n_209)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_151),
.Y(n_226)
);

OR2x4_ASAP7_75t_L g152 ( 
.A(n_106),
.B(n_80),
.Y(n_152)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_153),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_154),
.B(n_159),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_111),
.B(n_74),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_120),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_156),
.B(n_160),
.Y(n_211)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_102),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_43),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_43),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_161),
.B(n_175),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_126),
.B(n_64),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_162),
.B(n_163),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_60),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_99),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_165),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_112),
.B(n_65),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_64),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_181),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_167),
.A2(n_128),
.B1(n_100),
.B2(n_121),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_117),
.B(n_2),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_168),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_118),
.A2(n_77),
.B1(n_85),
.B2(n_43),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_169),
.A2(n_180),
.B1(n_138),
.B2(n_113),
.Y(n_222)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_107),
.A2(n_85),
.B1(n_77),
.B2(n_44),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_114),
.A2(n_44),
.B1(n_4),
.B2(n_7),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_97),
.B(n_44),
.C(n_4),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_127),
.C(n_100),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_96),
.A2(n_2),
.B(n_4),
.C(n_7),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

INVx3_ASAP7_75t_SL g177 ( 
.A(n_123),
.Y(n_177)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

OR2x2_ASAP7_75t_SL g178 ( 
.A(n_114),
.B(n_44),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_184),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_104),
.A2(n_44),
.B(n_8),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_179),
.A2(n_98),
.B(n_134),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_139),
.A2(n_2),
.B1(n_9),
.B2(n_10),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_10),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_133),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_128),
.Y(n_206)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_104),
.Y(n_183)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_132),
.Y(n_185)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_185),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_105),
.B1(n_121),
.B2(n_139),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_189),
.A2(n_178),
.B1(n_150),
.B2(n_183),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_199),
.A2(n_209),
.B(n_175),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_159),
.B(n_105),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_214),
.Y(n_227)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_203),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_206),
.Y(n_239)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_144),
.Y(n_207)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_207),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_208),
.A2(n_222),
.B1(n_177),
.B2(n_151),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_119),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_220),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_161),
.B(n_92),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_160),
.Y(n_231)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_156),
.B(n_119),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_162),
.B(n_92),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_224),
.Y(n_232)
);

AO22x2_ASAP7_75t_L g223 ( 
.A1(n_147),
.A2(n_123),
.B1(n_127),
.B2(n_113),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_223),
.B(n_167),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_149),
.B(n_95),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_228),
.B(n_235),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_230),
.A2(n_255),
.B(n_262),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_248),
.C(n_253),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_199),
.A2(n_150),
.B1(n_152),
.B2(n_142),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_233),
.A2(n_247),
.B1(n_212),
.B2(n_223),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_140),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_238),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_200),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_149),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_236),
.Y(n_264)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_181),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_168),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_245),
.Y(n_273)
);

INVxp33_ASAP7_75t_L g241 ( 
.A(n_193),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_241),
.B(n_243),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g243 ( 
.A(n_211),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_244),
.A2(n_261),
.B1(n_209),
.B2(n_208),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_190),
.B(n_163),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_186),
.A2(n_174),
.B1(n_140),
.B2(n_148),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_184),
.C(n_155),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_196),
.B(n_154),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_252),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_226),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_251),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_197),
.B(n_146),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_184),
.C(n_179),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_143),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_258),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_226),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_256),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_186),
.B(n_171),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_226),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_259),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_191),
.B(n_212),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_260),
.B(n_223),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_191),
.A2(n_138),
.B(n_185),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_263),
.A2(n_291),
.B1(n_268),
.B2(n_275),
.Y(n_309)
);

FAx1_ASAP7_75t_SL g265 ( 
.A(n_260),
.B(n_212),
.CI(n_191),
.CON(n_265),
.SN(n_265)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_265),
.B(n_234),
.Y(n_302)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_267),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_268),
.B(n_253),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_223),
.B(n_188),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_271),
.A2(n_288),
.B(n_259),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_230),
.A2(n_252),
.B1(n_235),
.B2(n_258),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_272),
.A2(n_294),
.B1(n_244),
.B2(n_254),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_236),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_229),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_281),
.Y(n_300)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_246),
.Y(n_279)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_246),
.Y(n_280)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_280),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_229),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_257),
.Y(n_282)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_231),
.B(n_223),
.C(n_203),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_283),
.B(n_296),
.C(n_250),
.Y(n_314)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_287),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_262),
.A2(n_188),
.B(n_198),
.Y(n_288)
);

OR2x6_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_198),
.Y(n_289)
);

INVx13_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_233),
.A2(n_153),
.B1(n_151),
.B2(n_225),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_227),
.A2(n_153),
.B1(n_210),
.B2(n_219),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_232),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_239),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_248),
.B(n_218),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_278),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_299),
.B(n_307),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_271),
.A2(n_261),
.B1(n_239),
.B2(n_227),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_301),
.A2(n_309),
.B1(n_312),
.B2(n_324),
.Y(n_351)
);

OAI21x1_ASAP7_75t_L g346 ( 
.A1(n_302),
.A2(n_290),
.B(n_289),
.Y(n_346)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_305),
.B(n_314),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_285),
.A2(n_232),
.B(n_247),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_308),
.A2(n_315),
.B1(n_325),
.B2(n_288),
.Y(n_339)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_310),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_264),
.B(n_238),
.Y(n_311)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_311),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_289),
.A2(n_283),
.B1(n_295),
.B2(n_278),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_273),
.B(n_240),
.Y(n_313)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_313),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_289),
.A2(n_270),
.B1(n_293),
.B2(n_292),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_245),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_274),
.C(n_276),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_317),
.B(n_319),
.Y(n_336)
);

FAx1_ASAP7_75t_SL g319 ( 
.A(n_272),
.B(n_207),
.CI(n_256),
.CON(n_319),
.SN(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_269),
.B(n_251),
.Y(n_320)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_320),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_269),
.B(n_237),
.Y(n_322)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_322),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_289),
.A2(n_237),
.B1(n_210),
.B2(n_187),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_289),
.A2(n_225),
.B1(n_195),
.B2(n_204),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_299),
.B(n_273),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_326),
.B(n_267),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_327),
.B(n_330),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_281),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_329),
.B(n_319),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_305),
.B(n_274),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_314),
.B(n_286),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_333),
.Y(n_353)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_300),
.Y(n_332)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_332),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_286),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_265),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_335),
.B(n_340),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_265),
.C(n_285),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_337),
.B(n_348),
.C(n_330),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_339),
.A2(n_270),
.B1(n_303),
.B2(n_298),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_320),
.B(n_290),
.Y(n_340)
);

A2O1A1O1Ixp25_ASAP7_75t_L g355 ( 
.A1(n_346),
.A2(n_311),
.B(n_304),
.C(n_319),
.D(n_306),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_313),
.A2(n_291),
.B1(n_293),
.B2(n_292),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_347),
.A2(n_309),
.B1(n_321),
.B2(n_297),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_322),
.B(n_294),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_301),
.B(n_284),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_308),
.Y(n_359)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_300),
.Y(n_350)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_350),
.Y(n_356)
);

FAx1_ASAP7_75t_SL g352 ( 
.A(n_335),
.B(n_302),
.CI(n_317),
.CON(n_352),
.SN(n_352)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_363),
.Y(n_379)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_355),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_336),
.A2(n_325),
.B(n_306),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_357),
.A2(n_351),
.B(n_338),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_359),
.B(n_371),
.Y(n_386)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_360),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_344),
.A2(n_324),
.B(n_323),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_361),
.B(n_364),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_362),
.A2(n_366),
.B1(n_367),
.B2(n_345),
.Y(n_376)
);

FAx1_ASAP7_75t_SL g363 ( 
.A(n_337),
.B(n_306),
.CI(n_319),
.CON(n_363),
.SN(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_332),
.B(n_321),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_334),
.A2(n_323),
.B(n_318),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_368),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_341),
.A2(n_318),
.B1(n_303),
.B2(n_298),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_343),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_297),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_333),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_336),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_280),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_373),
.A2(n_342),
.B1(n_351),
.B2(n_277),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_372),
.B(n_327),
.C(n_328),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_374),
.B(n_380),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_376),
.B(n_381),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_378),
.A2(n_369),
.B(n_358),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_359),
.A2(n_348),
.B1(n_349),
.B2(n_340),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_385),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_353),
.B(n_328),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_287),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_387),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_356),
.B(n_282),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_388),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_370),
.A2(n_354),
.B1(n_363),
.B2(n_366),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_389),
.A2(n_363),
.B1(n_355),
.B2(n_352),
.Y(n_391)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_390),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_391),
.B(n_385),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_383),
.B(n_352),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_392),
.B(n_395),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_379),
.A2(n_371),
.B(n_367),
.Y(n_394)
);

AO21x1_ASAP7_75t_L g411 ( 
.A1(n_394),
.A2(n_400),
.B(n_187),
.Y(n_411)
);

NOR3xp33_ASAP7_75t_L g395 ( 
.A(n_377),
.B(n_357),
.C(n_279),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_396),
.B(n_249),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_379),
.A2(n_378),
.B(n_389),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_398),
.B(n_402),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_375),
.A2(n_266),
.B(n_353),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_376),
.A2(n_384),
.B(n_381),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_403),
.B(n_386),
.C(n_374),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_406),
.B(n_407),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_393),
.B(n_386),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_399),
.A2(n_358),
.B1(n_266),
.B2(n_387),
.Y(n_408)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_408),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_409),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_402),
.B(n_382),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_410),
.B(n_411),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_398),
.B(n_192),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_414),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_413),
.B(n_396),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_SL g414 ( 
.A1(n_401),
.A2(n_249),
.B1(n_145),
.B2(n_195),
.Y(n_414)
);

BUFx24_ASAP7_75t_SL g416 ( 
.A(n_391),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_416),
.B(n_170),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_415),
.C(n_409),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_419),
.B(n_421),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_414),
.B(n_393),
.C(n_404),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_423),
.A2(n_192),
.B1(n_194),
.B2(n_216),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_407),
.B(n_397),
.C(n_204),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_424),
.A2(n_426),
.B(n_425),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_427),
.B(n_428),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_417),
.A2(n_216),
.B1(n_194),
.B2(n_141),
.Y(n_428)
);

AOI21x1_ASAP7_75t_SL g429 ( 
.A1(n_420),
.A2(n_201),
.B(n_202),
.Y(n_429)
);

MAJx2_ASAP7_75t_L g435 ( 
.A(n_429),
.B(n_430),
.C(n_13),
.Y(n_435)
);

AOI322xp5_ASAP7_75t_L g430 ( 
.A1(n_420),
.A2(n_201),
.A3(n_202),
.B1(n_94),
.B2(n_14),
.C1(n_11),
.C2(n_13),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_432),
.Y(n_436)
);

AO221x1_ASAP7_75t_L g433 ( 
.A1(n_422),
.A2(n_418),
.B1(n_424),
.B2(n_201),
.C(n_202),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_433),
.A2(n_11),
.B(n_13),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_434),
.Y(n_438)
);

O2A1O1Ixp33_ASAP7_75t_SL g439 ( 
.A1(n_435),
.A2(n_430),
.B(n_431),
.C(n_13),
.Y(n_439)
);

NOR4xp25_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_437),
.C(n_14),
.D(n_436),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_438),
.Y(n_441)
);


endmodule