module fake_jpeg_12561_n_271 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_271);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_11),
.B(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_55),
.Y(n_86)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_53),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_52),
.Y(n_71)
);

BUFx4f_ASAP7_75t_SL g53 ( 
.A(n_24),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_0),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_1),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_3),
.B(n_5),
.Y(n_99)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_23),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_62),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_40),
.B(n_2),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_65),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_28),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_24),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_38),
.B1(n_30),
.B2(n_37),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_68),
.A2(n_77),
.B1(n_88),
.B2(n_92),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_29),
.B1(n_37),
.B2(n_31),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_69),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_38),
.C(n_35),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_79),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_37),
.B1(n_31),
.B2(n_26),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_73),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_65),
.B1(n_51),
.B2(n_61),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_18),
.C(n_27),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_27),
.C(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_97),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_87),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_25),
.B1(n_31),
.B2(n_26),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_46),
.A2(n_63),
.B1(n_43),
.B2(n_26),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_25),
.B1(n_39),
.B2(n_32),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_93),
.A2(n_94),
.B1(n_98),
.B2(n_101),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_44),
.A2(n_25),
.B1(n_32),
.B2(n_23),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_95),
.B(n_102),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_39),
.C(n_4),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_62),
.A2(n_39),
.B1(n_4),
.B2(n_5),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_87),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_53),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_56),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_59),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_60),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_14),
.B1(n_16),
.B2(n_89),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_104),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g153 ( 
.A(n_108),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_53),
.B(n_12),
.C(n_13),
.Y(n_109)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_109),
.A2(n_82),
.A3(n_119),
.B1(n_110),
.B2(n_107),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_10),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_117),
.Y(n_139)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_12),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_72),
.B(n_13),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_85),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_116),
.A2(n_83),
.B1(n_90),
.B2(n_67),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_16),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_81),
.B1(n_83),
.B2(n_90),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_126),
.A2(n_131),
.B1(n_128),
.B2(n_125),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_92),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_132),
.Y(n_152)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_134),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_81),
.A2(n_83),
.B1(n_90),
.B2(n_67),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_80),
.B(n_76),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_75),
.B(n_78),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_96),
.Y(n_146)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_132),
.B(n_97),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_158),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_127),
.A2(n_102),
.B(n_67),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_158),
.B(n_113),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_141),
.B(n_146),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_91),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_151),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_111),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_150),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_96),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_155),
.B1(n_104),
.B2(n_150),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_67),
.B1(n_82),
.B2(n_121),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_160),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_106),
.A2(n_82),
.B(n_115),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_105),
.B(n_123),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_159),
.B(n_139),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_109),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_157),
.B1(n_161),
.B2(n_138),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_166),
.C(n_169),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_104),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_114),
.C(n_121),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_182),
.Y(n_208)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_152),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_140),
.A2(n_120),
.B(n_129),
.C(n_133),
.Y(n_170)
);

OA21x2_ASAP7_75t_L g194 ( 
.A1(n_170),
.A2(n_162),
.B(n_145),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_177),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_120),
.B1(n_129),
.B2(n_118),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_129),
.B1(n_130),
.B2(n_134),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_147),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_137),
.A2(n_129),
.B1(n_122),
.B2(n_104),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_163),
.B1(n_155),
.B2(n_149),
.Y(n_189)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_184),
.Y(n_197)
);

OAI221xp5_ASAP7_75t_L g184 ( 
.A1(n_160),
.A2(n_139),
.B1(n_159),
.B2(n_156),
.C(n_151),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_188),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_141),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_186),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_143),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_187),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_147),
.B(n_142),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_189),
.A2(n_194),
.B(n_183),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_164),
.A2(n_154),
.B1(n_142),
.B2(n_144),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_191),
.A2(n_203),
.B1(n_204),
.B2(n_170),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_149),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_176),
.C(n_172),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_145),
.Y(n_200)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_180),
.A2(n_145),
.B1(n_162),
.B2(n_165),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_201),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_173),
.A2(n_178),
.B1(n_174),
.B2(n_177),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_178),
.A2(n_184),
.B1(n_170),
.B2(n_167),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_179),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_206),
.B(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_182),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_210),
.B(n_218),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_170),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_213),
.C(n_219),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_206),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_215),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_170),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_168),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_220),
.B(n_221),
.Y(n_235)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

BUFx12_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_222),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_205),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_223),
.A2(n_224),
.B1(n_199),
.B2(n_192),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_192),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_216),
.A2(n_197),
.B1(n_224),
.B2(n_214),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_212),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_193),
.C(n_204),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_234),
.C(n_236),
.Y(n_240)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_231),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_197),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_215),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_203),
.C(n_190),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_190),
.C(n_198),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_238),
.A2(n_244),
.B(n_235),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_226),
.B(n_198),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_241),
.Y(n_250)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_243),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_229),
.A2(n_214),
.B(n_194),
.Y(n_243)
);

AO21x1_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_202),
.B(n_217),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_200),
.C(n_217),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_232),
.C(n_236),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_220),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_194),
.C(n_191),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_249),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_230),
.C(n_234),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_225),
.C(n_233),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_253),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_248),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_258),
.Y(n_261)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

AOI21x1_ASAP7_75t_SL g259 ( 
.A1(n_257),
.A2(n_243),
.B(n_237),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_260),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_254),
.A2(n_256),
.B(n_245),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_194),
.B1(n_241),
.B2(n_209),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_262),
.A2(n_244),
.B(n_246),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_263),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_250),
.B(n_222),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_264),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_265),
.C(n_259),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_268),
.B(n_267),
.Y(n_269)
);

AOI321xp33_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_189),
.A3(n_207),
.B1(n_221),
.B2(n_222),
.C(n_254),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_207),
.Y(n_271)
);


endmodule