module fake_jpeg_18840_n_30 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_30);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_30;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_29;
wire n_15;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_5),
.A2(n_8),
.B1(n_0),
.B2(n_12),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_6),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_17),
.A2(n_18),
.B1(n_13),
.B2(n_5),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_20),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_2),
.B(n_3),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_4),
.C(n_7),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_4),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_23),
.A2(n_13),
.B(n_6),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_25),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_22),
.B(n_19),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_21),
.C(n_8),
.Y(n_28)
);

AOI21xp33_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_7),
.B(n_9),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_29),
.A2(n_27),
.B(n_9),
.Y(n_30)
);


endmodule