module real_aes_16925_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1034;
wire n_549;
wire n_1328;
wire n_571;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_1301;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_580;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_550;
wire n_966;
wire n_333;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_769;
wire n_434;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_1343;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_340;
wire n_483;
wire n_394;
wire n_1280;
wire n_729;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_SL g1261 ( .A1(n_0), .A2(n_79), .B1(n_734), .B2(n_822), .Y(n_1261) );
AOI22xp33_ASAP7_75t_L g1284 ( .A1(n_0), .A2(n_232), .B1(n_501), .B2(n_933), .Y(n_1284) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_1), .A2(n_6), .B1(n_1058), .B2(n_1061), .Y(n_1100) );
OAI22xp33_ASAP7_75t_SL g878 ( .A1(n_2), .A2(n_113), .B1(n_394), .B2(n_397), .Y(n_878) );
OAI22xp33_ASAP7_75t_L g888 ( .A1(n_2), .A2(n_27), .B1(n_407), .B2(n_408), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_3), .A2(n_28), .B1(n_388), .B2(n_758), .Y(n_1023) );
OAI22xp5_ASAP7_75t_SL g1031 ( .A1(n_3), .A2(n_116), .B1(n_407), .B2(n_429), .Y(n_1031) );
INVx1_ASAP7_75t_L g1270 ( .A(n_4), .Y(n_1270) );
INVx1_ASAP7_75t_L g1347 ( .A(n_5), .Y(n_1347) );
OAI22xp33_ASAP7_75t_L g575 ( .A1(n_7), .A2(n_157), .B1(n_388), .B2(n_397), .Y(n_575) );
OAI22xp33_ASAP7_75t_SL g591 ( .A1(n_7), .A2(n_157), .B1(n_407), .B2(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g692 ( .A(n_8), .Y(n_692) );
OAI211xp5_ASAP7_75t_L g696 ( .A1(n_8), .A2(n_577), .B(n_697), .C(n_698), .Y(n_696) );
CKINVDCx5p33_ASAP7_75t_R g1026 ( .A(n_9), .Y(n_1026) );
INVx1_ASAP7_75t_L g785 ( .A(n_10), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g1004 ( .A(n_11), .Y(n_1004) );
INVx1_ASAP7_75t_L g262 ( .A(n_12), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_12), .B(n_272), .Y(n_341) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_12), .B(n_205), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_12), .B(n_396), .Y(n_1273) );
CKINVDCx5p33_ASAP7_75t_R g864 ( .A(n_13), .Y(n_864) );
OAI22xp33_ASAP7_75t_L g977 ( .A1(n_14), .A2(n_187), .B1(n_264), .B2(n_760), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_14), .A2(n_187), .B1(n_987), .B2(n_989), .Y(n_986) );
CKINVDCx5p33_ASAP7_75t_R g854 ( .A(n_15), .Y(n_854) );
INVx1_ASAP7_75t_L g633 ( .A(n_16), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g858 ( .A(n_17), .Y(n_858) );
AOI221xp5_ASAP7_75t_L g1260 ( .A1(n_18), .A2(n_128), .B1(n_470), .B2(n_894), .C(n_897), .Y(n_1260) );
AOI22xp33_ASAP7_75t_L g1289 ( .A1(n_18), .A2(n_67), .B1(n_501), .B2(n_1290), .Y(n_1289) );
INVx1_ASAP7_75t_L g911 ( .A(n_19), .Y(n_911) );
INVx2_ASAP7_75t_L g1046 ( .A(n_20), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_20), .B(n_101), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_20), .B(n_1060), .Y(n_1062) );
CKINVDCx5p33_ASAP7_75t_R g1252 ( .A(n_21), .Y(n_1252) );
AOI22xp33_ASAP7_75t_SL g810 ( .A1(n_22), .A2(n_239), .B1(n_584), .B2(n_800), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_22), .A2(n_26), .B1(n_816), .B2(n_819), .Y(n_825) );
OAI22xp5_ASAP7_75t_SL g657 ( .A1(n_23), .A2(n_130), .B1(n_658), .B2(n_659), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_23), .A2(n_130), .B1(n_664), .B2(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g835 ( .A(n_24), .Y(n_835) );
AO22x2_ASAP7_75t_L g534 ( .A1(n_25), .A2(n_535), .B1(n_600), .B2(n_601), .Y(n_534) );
INVx1_ASAP7_75t_L g600 ( .A(n_25), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_26), .A2(n_161), .B1(n_501), .B2(n_804), .Y(n_803) );
OAI22xp33_ASAP7_75t_SL g877 ( .A1(n_27), .A2(n_223), .B1(n_388), .B2(n_523), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g1030 ( .A(n_28), .B(n_428), .Y(n_1030) );
AOI22xp5_ASAP7_75t_L g1064 ( .A1(n_29), .A2(n_211), .B1(n_1058), .B2(n_1061), .Y(n_1064) );
INVx1_ASAP7_75t_L g782 ( .A(n_30), .Y(n_782) );
INVx1_ASAP7_75t_L g613 ( .A(n_31), .Y(n_613) );
XOR2xp5_ASAP7_75t_L g849 ( .A(n_32), .B(n_850), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_33), .A2(n_150), .B1(n_264), .B2(n_397), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_33), .A2(n_150), .B1(n_408), .B2(n_839), .Y(n_838) );
OAI22xp33_ASAP7_75t_L g759 ( .A1(n_34), .A2(n_127), .B1(n_388), .B2(n_760), .Y(n_759) );
OAI22xp33_ASAP7_75t_SL g762 ( .A1(n_34), .A2(n_127), .B1(n_407), .B2(n_592), .Y(n_762) );
CKINVDCx5p33_ASAP7_75t_R g1014 ( .A(n_35), .Y(n_1014) );
INVx1_ASAP7_75t_L g542 ( .A(n_36), .Y(n_542) );
OAI22xp33_ASAP7_75t_L g387 ( .A1(n_37), .A2(n_180), .B1(n_388), .B2(n_390), .Y(n_387) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_37), .A2(n_98), .B1(n_407), .B2(n_408), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g1010 ( .A(n_38), .Y(n_1010) );
CKINVDCx5p33_ASAP7_75t_R g862 ( .A(n_39), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g1070 ( .A1(n_40), .A2(n_236), .B1(n_1043), .B2(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g1338 ( .A(n_41), .Y(n_1338) );
OAI22xp33_ASAP7_75t_L g660 ( .A1(n_42), .A2(n_149), .B1(n_264), .B2(n_397), .Y(n_660) );
OAI22xp33_ASAP7_75t_L g674 ( .A1(n_42), .A2(n_149), .B1(n_675), .B2(n_677), .Y(n_674) );
INVx1_ASAP7_75t_L g718 ( .A(n_43), .Y(n_718) );
XOR2x2_ASAP7_75t_L g795 ( .A(n_44), .B(n_796), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g1074 ( .A1(n_44), .A2(n_228), .B1(n_1058), .B2(n_1061), .Y(n_1074) );
XNOR2xp5_ASAP7_75t_L g606 ( .A(n_45), .B(n_607), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_46), .A2(n_160), .B1(n_408), .B2(n_429), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_46), .A2(n_48), .B1(n_587), .B2(n_758), .Y(n_919) );
INVx1_ASAP7_75t_L g831 ( .A(n_47), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_48), .A2(n_245), .B1(n_407), .B2(n_428), .Y(n_905) );
CKINVDCx5p33_ASAP7_75t_R g1011 ( .A(n_49), .Y(n_1011) );
AO22x1_ASAP7_75t_L g1054 ( .A1(n_50), .A2(n_66), .B1(n_1043), .B2(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g756 ( .A(n_51), .Y(n_756) );
INVx1_ASAP7_75t_L g296 ( .A(n_52), .Y(n_296) );
INVx1_ASAP7_75t_L g303 ( .A(n_52), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g1317 ( .A1(n_53), .A2(n_124), .B1(n_677), .B2(n_987), .Y(n_1317) );
OAI22xp33_ASAP7_75t_L g1333 ( .A1(n_53), .A2(n_124), .B1(n_264), .B2(n_397), .Y(n_1333) );
INVx1_ASAP7_75t_L g962 ( .A(n_54), .Y(n_962) );
CKINVDCx5p33_ASAP7_75t_R g1005 ( .A(n_55), .Y(n_1005) );
OAI22xp33_ASAP7_75t_L g586 ( .A1(n_56), .A2(n_102), .B1(n_587), .B2(n_588), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g598 ( .A1(n_56), .A2(n_102), .B1(n_428), .B2(n_429), .Y(n_598) );
INVx1_ASAP7_75t_L g956 ( .A(n_57), .Y(n_956) );
OAI211xp5_ASAP7_75t_L g369 ( .A1(n_58), .A2(n_370), .B(n_371), .C(n_377), .Y(n_369) );
INVx1_ASAP7_75t_L g426 ( .A(n_58), .Y(n_426) );
INVx1_ASAP7_75t_L g255 ( .A(n_59), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_60), .A2(n_178), .B1(n_464), .B2(n_480), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_60), .A2(n_185), .B1(n_504), .B2(n_508), .Y(n_510) );
INVx2_ASAP7_75t_L g289 ( .A(n_61), .Y(n_289) );
INVx1_ASAP7_75t_L g621 ( .A(n_62), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g893 ( .A1(n_63), .A2(n_226), .B1(n_842), .B2(n_894), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_63), .A2(n_164), .B1(n_935), .B2(n_937), .Y(n_938) );
XNOR2x2_ASAP7_75t_L g947 ( .A(n_64), .B(n_948), .Y(n_947) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_65), .A2(n_204), .B1(n_522), .B2(n_659), .Y(n_984) );
OAI22xp33_ASAP7_75t_L g994 ( .A1(n_65), .A2(n_204), .B1(n_685), .B2(n_995), .Y(n_994) );
AOI221xp5_ASAP7_75t_L g1257 ( .A1(n_67), .A2(n_77), .B1(n_332), .B2(n_894), .C(n_1258), .Y(n_1257) );
INVx1_ASAP7_75t_L g910 ( .A(n_68), .Y(n_910) );
INVx1_ASAP7_75t_L g908 ( .A(n_69), .Y(n_908) );
AOI22xp5_ASAP7_75t_L g1075 ( .A1(n_70), .A2(n_162), .B1(n_1043), .B2(n_1055), .Y(n_1075) );
INVx1_ASAP7_75t_L g1246 ( .A(n_71), .Y(n_1246) );
INVx1_ASAP7_75t_L g1236 ( .A(n_72), .Y(n_1236) );
OAI222xp33_ASAP7_75t_L g450 ( .A1(n_73), .A2(n_103), .B1(n_218), .B2(n_451), .C1(n_453), .C2(n_455), .Y(n_450) );
OAI222xp33_ASAP7_75t_L g525 ( .A1(n_73), .A2(n_103), .B1(n_218), .B2(n_526), .C1(n_528), .C2(n_530), .Y(n_525) );
INVx1_ASAP7_75t_L g957 ( .A(n_74), .Y(n_957) );
INVx1_ASAP7_75t_L g725 ( .A(n_75), .Y(n_725) );
AO221x2_ASAP7_75t_L g1101 ( .A1(n_76), .A2(n_195), .B1(n_1058), .B2(n_1061), .C(n_1102), .Y(n_1101) );
AOI221xp5_ASAP7_75t_L g1279 ( .A1(n_77), .A2(n_128), .B1(n_1280), .B2(n_1281), .C(n_1283), .Y(n_1279) );
OAI22xp33_ASAP7_75t_L g393 ( .A1(n_78), .A2(n_98), .B1(n_394), .B2(n_397), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g427 ( .A1(n_78), .A2(n_180), .B1(n_428), .B2(n_429), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g1291 ( .A1(n_79), .A2(n_86), .B1(n_937), .B2(n_1281), .C(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g776 ( .A(n_80), .Y(n_776) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_81), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_82), .A2(n_246), .B1(n_473), .B2(n_475), .Y(n_472) );
AOI22xp33_ASAP7_75t_SL g514 ( .A1(n_82), .A2(n_122), .B1(n_515), .B2(n_516), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_83), .A2(n_122), .B1(n_483), .B2(n_484), .Y(n_482) );
AOI22xp33_ASAP7_75t_SL g503 ( .A1(n_83), .A2(n_246), .B1(n_504), .B2(n_508), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g896 ( .A1(n_84), .A2(n_244), .B1(n_484), .B2(n_640), .C(n_897), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_84), .A2(n_121), .B1(n_516), .B2(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g755 ( .A(n_85), .Y(n_755) );
AOI22xp33_ASAP7_75t_SL g1259 ( .A1(n_86), .A2(n_232), .B1(n_734), .B2(n_822), .Y(n_1259) );
AOI22xp33_ASAP7_75t_SL g808 ( .A1(n_87), .A2(n_193), .B1(n_501), .B2(n_809), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_87), .A2(n_89), .B1(n_565), .B2(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g875 ( .A(n_88), .Y(n_875) );
OAI211xp5_ASAP7_75t_SL g881 ( .A1(n_88), .A2(n_451), .B(n_594), .C(n_882), .Y(n_881) );
AOI22xp33_ASAP7_75t_SL g799 ( .A1(n_89), .A2(n_147), .B1(n_584), .B2(n_800), .Y(n_799) );
XOR2x2_ASAP7_75t_L g749 ( .A(n_90), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g952 ( .A(n_91), .Y(n_952) );
OAI211xp5_ASAP7_75t_L g978 ( .A1(n_92), .A2(n_649), .B(n_979), .C(n_983), .Y(n_978) );
INVx1_ASAP7_75t_L g993 ( .A(n_92), .Y(n_993) );
INVx1_ASAP7_75t_L g626 ( .A(n_93), .Y(n_626) );
INVx1_ASAP7_75t_L g278 ( .A(n_94), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_95), .A2(n_148), .B1(n_587), .B2(n_758), .Y(n_757) );
OAI22xp33_ASAP7_75t_L g769 ( .A1(n_95), .A2(n_148), .B1(n_428), .B2(n_429), .Y(n_769) );
INVx1_ASAP7_75t_L g1343 ( .A(n_96), .Y(n_1343) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_97), .Y(n_257) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_97), .B(n_255), .Y(n_1044) );
CKINVDCx5p33_ASAP7_75t_R g1249 ( .A(n_99), .Y(n_1249) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_100), .A2(n_153), .B1(n_665), .B2(n_685), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_100), .A2(n_153), .B1(n_522), .B2(n_659), .Y(n_701) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_101), .B(n_1046), .Y(n_1045) );
INVx1_ASAP7_75t_L g1060 ( .A(n_101), .Y(n_1060) );
INVx1_ASAP7_75t_L g559 ( .A(n_104), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_105), .A2(n_208), .B1(n_447), .B2(n_448), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_105), .A2(n_208), .B1(n_522), .B2(n_523), .Y(n_521) );
INVx2_ASAP7_75t_L g288 ( .A(n_106), .Y(n_288) );
INVx1_ASAP7_75t_L g336 ( .A(n_106), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_106), .B(n_289), .Y(n_1241) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_107), .Y(n_297) );
INVx1_ASAP7_75t_L g691 ( .A(n_108), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_109), .A2(n_189), .B1(n_1043), .B2(n_1055), .Y(n_1099) );
INVx1_ASAP7_75t_L g774 ( .A(n_110), .Y(n_774) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_111), .Y(n_312) );
INVx1_ASAP7_75t_L g654 ( .A(n_112), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_113), .A2(n_223), .B1(n_428), .B2(n_429), .Y(n_880) );
OAI22xp33_ASAP7_75t_SL g1028 ( .A1(n_114), .A2(n_116), .B1(n_587), .B2(n_760), .Y(n_1028) );
OAI22xp5_ASAP7_75t_L g1035 ( .A1(n_114), .A2(n_120), .B1(n_885), .B2(n_886), .Y(n_1035) );
INVx1_ASAP7_75t_L g441 ( .A(n_115), .Y(n_441) );
INVx1_ASAP7_75t_L g1351 ( .A(n_117), .Y(n_1351) );
INVx1_ASAP7_75t_L g580 ( .A(n_118), .Y(n_580) );
INVx1_ASAP7_75t_L g784 ( .A(n_119), .Y(n_784) );
INVx1_ASAP7_75t_L g1027 ( .A(n_120), .Y(n_1027) );
AOI221xp5_ASAP7_75t_L g898 ( .A1(n_121), .A2(n_197), .B1(n_484), .B2(n_640), .C(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g710 ( .A(n_123), .Y(n_710) );
XOR2xp5_ASAP7_75t_L g437 ( .A(n_125), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g716 ( .A(n_126), .Y(n_716) );
INVx1_ASAP7_75t_L g557 ( .A(n_129), .Y(n_557) );
AOI31xp33_ASAP7_75t_L g891 ( .A1(n_131), .A2(n_892), .A3(n_904), .B(n_913), .Y(n_891) );
NAND2xp33_ASAP7_75t_SL g929 ( .A(n_131), .B(n_930), .Y(n_929) );
INVxp67_ASAP7_75t_SL g942 ( .A(n_131), .Y(n_942) );
AO22x1_ASAP7_75t_L g1057 ( .A1(n_131), .A2(n_209), .B1(n_1058), .B2(n_1061), .Y(n_1057) );
BUFx3_ASAP7_75t_L g294 ( .A(n_132), .Y(n_294) );
OAI211xp5_ASAP7_75t_SL g1024 ( .A1(n_133), .A2(n_371), .B(n_873), .C(n_1025), .Y(n_1024) );
OAI211xp5_ASAP7_75t_SL g1032 ( .A1(n_133), .A2(n_594), .B(n_1033), .C(n_1034), .Y(n_1032) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_134), .Y(n_329) );
INVx1_ASAP7_75t_L g1337 ( .A(n_135), .Y(n_1337) );
INVx1_ASAP7_75t_L g954 ( .A(n_136), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_137), .A2(n_158), .B1(n_1058), .B2(n_1061), .Y(n_1080) );
INVx1_ASAP7_75t_L g656 ( .A(n_138), .Y(n_656) );
OAI211xp5_ASAP7_75t_SL g666 ( .A1(n_138), .A2(n_594), .B(n_667), .C(n_669), .Y(n_666) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_139), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_140), .A2(n_185), .B1(n_464), .B2(n_470), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_140), .A2(n_178), .B1(n_496), .B2(n_500), .Y(n_495) );
OAI22xp33_ASAP7_75t_L g693 ( .A1(n_141), .A2(n_184), .B1(n_675), .B2(n_694), .Y(n_693) );
OAI22xp33_ASAP7_75t_L g702 ( .A1(n_141), .A2(n_184), .B1(n_388), .B2(n_397), .Y(n_702) );
CKINVDCx5p33_ASAP7_75t_R g1008 ( .A(n_142), .Y(n_1008) );
INVx1_ASAP7_75t_L g1274 ( .A(n_143), .Y(n_1274) );
INVx1_ASAP7_75t_L g554 ( .A(n_144), .Y(n_554) );
INVx1_ASAP7_75t_L g1341 ( .A(n_145), .Y(n_1341) );
INVx1_ASAP7_75t_L g545 ( .A(n_146), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_147), .A2(n_193), .B1(n_813), .B2(n_814), .Y(n_812) );
INVx1_ASAP7_75t_L g902 ( .A(n_151), .Y(n_902) );
AOI22xp33_ASAP7_75t_SL g932 ( .A1(n_151), .A2(n_226), .B1(n_501), .B2(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g960 ( .A(n_152), .Y(n_960) );
OAI21xp5_ASAP7_75t_SL g1296 ( .A1(n_154), .A2(n_1297), .B(n_1301), .Y(n_1296) );
INVx1_ASAP7_75t_L g1320 ( .A(n_155), .Y(n_1320) );
OA22x2_ASAP7_75t_L g681 ( .A1(n_156), .A2(n_682), .B1(n_740), .B2(n_741), .Y(n_681) );
INVxp67_ASAP7_75t_L g741 ( .A(n_156), .Y(n_741) );
CKINVDCx5p33_ASAP7_75t_R g857 ( .A(n_159), .Y(n_857) );
INVxp67_ASAP7_75t_SL g917 ( .A(n_160), .Y(n_917) );
AOI22xp33_ASAP7_75t_SL g815 ( .A1(n_161), .A2(n_239), .B1(n_816), .B2(n_819), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g1065 ( .A1(n_163), .A2(n_227), .B1(n_1043), .B2(n_1055), .Y(n_1065) );
INVx1_ASAP7_75t_L g901 ( .A(n_164), .Y(n_901) );
INVx1_ASAP7_75t_L g833 ( .A(n_165), .Y(n_833) );
INVx1_ASAP7_75t_L g631 ( .A(n_166), .Y(n_631) );
INVx1_ASAP7_75t_L g707 ( .A(n_167), .Y(n_707) );
OAI211xp5_ASAP7_75t_SL g1318 ( .A1(n_168), .A2(n_594), .B(n_991), .C(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1329 ( .A(n_168), .Y(n_1329) );
INVx1_ASAP7_75t_L g582 ( .A(n_169), .Y(n_582) );
OAI211xp5_ASAP7_75t_L g686 ( .A1(n_170), .A2(n_415), .B(n_687), .C(n_690), .Y(n_686) );
INVx1_ASAP7_75t_L g699 ( .A(n_170), .Y(n_699) );
CKINVDCx5p33_ASAP7_75t_R g865 ( .A(n_171), .Y(n_865) );
OAI211xp5_ASAP7_75t_L g872 ( .A1(n_172), .A2(n_371), .B(n_873), .C(n_874), .Y(n_872) );
INVx1_ASAP7_75t_L g887 ( .A(n_172), .Y(n_887) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_173), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_174), .A2(n_222), .B1(n_1043), .B2(n_1055), .Y(n_1079) );
OAI22xp33_ASAP7_75t_L g1322 ( .A1(n_175), .A2(n_237), .B1(n_685), .B2(n_995), .Y(n_1322) );
OAI22xp5_ASAP7_75t_L g1330 ( .A1(n_175), .A2(n_237), .B1(n_658), .B2(n_1331), .Y(n_1330) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_176), .Y(n_268) );
INVx1_ASAP7_75t_L g834 ( .A(n_177), .Y(n_834) );
INVx1_ASAP7_75t_L g628 ( .A(n_179), .Y(n_628) );
INVx1_ASAP7_75t_L g546 ( .A(n_181), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g855 ( .A(n_182), .Y(n_855) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_183), .Y(n_291) );
AO22x1_ASAP7_75t_L g1095 ( .A1(n_186), .A2(n_210), .B1(n_1043), .B2(n_1096), .Y(n_1095) );
CKINVDCx16_ASAP7_75t_R g1103 ( .A(n_188), .Y(n_1103) );
OAI211xp5_ASAP7_75t_SL g648 ( .A1(n_190), .A2(n_649), .B(n_652), .C(n_653), .Y(n_648) );
INVx1_ASAP7_75t_L g672 ( .A(n_190), .Y(n_672) );
INVx1_ASAP7_75t_L g780 ( .A(n_191), .Y(n_780) );
INVx1_ASAP7_75t_L g539 ( .A(n_192), .Y(n_539) );
INVx1_ASAP7_75t_L g982 ( .A(n_194), .Y(n_982) );
OAI211xp5_ASAP7_75t_L g990 ( .A1(n_194), .A2(n_594), .B(n_991), .C(n_992), .Y(n_990) );
INVx1_ASAP7_75t_L g552 ( .A(n_196), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_197), .A2(n_244), .B1(n_935), .B2(n_937), .Y(n_934) );
INVx1_ASAP7_75t_L g829 ( .A(n_198), .Y(n_829) );
INVx1_ASAP7_75t_L g724 ( .A(n_199), .Y(n_724) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_200), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g1015 ( .A(n_201), .Y(n_1015) );
INVx1_ASAP7_75t_L g777 ( .A(n_202), .Y(n_777) );
XOR2xp5_ASAP7_75t_L g999 ( .A(n_203), .B(n_1000), .Y(n_999) );
AOI22xp5_ASAP7_75t_L g1069 ( .A1(n_203), .A2(n_230), .B1(n_1058), .B2(n_1061), .Y(n_1069) );
BUFx3_ASAP7_75t_L g272 ( .A(n_205), .Y(n_272) );
INVx1_ASAP7_75t_L g396 ( .A(n_205), .Y(n_396) );
INVx1_ASAP7_75t_L g980 ( .A(n_206), .Y(n_980) );
CKINVDCx20_ASAP7_75t_R g1104 ( .A(n_207), .Y(n_1104) );
CKINVDCx5p33_ASAP7_75t_R g876 ( .A(n_212), .Y(n_876) );
INVx1_ASAP7_75t_L g1348 ( .A(n_213), .Y(n_1348) );
CKINVDCx5p33_ASAP7_75t_R g1007 ( .A(n_214), .Y(n_1007) );
AOI22xp5_ASAP7_75t_L g1311 ( .A1(n_215), .A2(n_1312), .B1(n_1313), .B2(n_1314), .Y(n_1311) );
CKINVDCx5p33_ASAP7_75t_R g1312 ( .A(n_215), .Y(n_1312) );
INVx1_ASAP7_75t_L g719 ( .A(n_216), .Y(n_719) );
INVx1_ASAP7_75t_L g714 ( .A(n_217), .Y(n_714) );
INVx1_ASAP7_75t_L g773 ( .A(n_219), .Y(n_773) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_220), .Y(n_322) );
INVx1_ASAP7_75t_L g585 ( .A(n_221), .Y(n_585) );
OAI211xp5_ASAP7_75t_L g752 ( .A1(n_224), .A2(n_371), .B(n_753), .C(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g765 ( .A(n_224), .Y(n_765) );
INVx1_ASAP7_75t_L g286 ( .A(n_225), .Y(n_286) );
INVx2_ASAP7_75t_L g334 ( .A(n_225), .Y(n_334) );
INVx1_ASAP7_75t_L g490 ( .A(n_225), .Y(n_490) );
AOI222xp33_ASAP7_75t_L g1225 ( .A1(n_227), .A2(n_1226), .B1(n_1307), .B2(n_1310), .C1(n_1362), .C2(n_1364), .Y(n_1225) );
XNOR2x1_ASAP7_75t_L g1227 ( .A(n_227), .B(n_1228), .Y(n_1227) );
AO22x1_ASAP7_75t_L g1097 ( .A1(n_229), .A2(n_240), .B1(n_1058), .B2(n_1061), .Y(n_1097) );
CKINVDCx5p33_ASAP7_75t_R g861 ( .A(n_231), .Y(n_861) );
INVx1_ASAP7_75t_L g611 ( .A(n_233), .Y(n_611) );
INVx1_ASAP7_75t_L g963 ( .A(n_234), .Y(n_963) );
INVx1_ASAP7_75t_L g617 ( .A(n_235), .Y(n_617) );
INVx1_ASAP7_75t_L g1350 ( .A(n_238), .Y(n_1350) );
INVx1_ASAP7_75t_L g1321 ( .A(n_241), .Y(n_1321) );
OAI211xp5_ASAP7_75t_L g1324 ( .A1(n_241), .A2(n_652), .B(n_1325), .C(n_1328), .Y(n_1324) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_242), .Y(n_331) );
INVx1_ASAP7_75t_L g443 ( .A(n_243), .Y(n_443) );
INVx1_ASAP7_75t_L g915 ( .A(n_245), .Y(n_915) );
INVx1_ASAP7_75t_L g959 ( .A(n_247), .Y(n_959) );
INVx1_ASAP7_75t_L g386 ( .A(n_248), .Y(n_386) );
OAI211xp5_ASAP7_75t_L g411 ( .A1(n_248), .A2(n_412), .B(n_415), .C(n_419), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_273), .B(n_1039), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_258), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g1309 ( .A(n_252), .B(n_261), .Y(n_1309) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g1363 ( .A(n_254), .B(n_257), .Y(n_1363) );
INVx1_ASAP7_75t_L g1365 ( .A(n_254), .Y(n_1365) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g1367 ( .A(n_257), .B(n_1365), .Y(n_1367) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g402 ( .A(n_261), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g367 ( .A(n_262), .B(n_272), .Y(n_367) );
AND2x4_ASAP7_75t_L g1293 ( .A(n_262), .B(n_271), .Y(n_1293) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_263), .A2(n_398), .B1(n_441), .B2(n_443), .Y(n_519) );
AND2x4_ASAP7_75t_SL g1308 ( .A(n_263), .B(n_1309), .Y(n_1308) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x6_ASAP7_75t_L g264 ( .A(n_265), .B(n_270), .Y(n_264) );
OR2x6_ASAP7_75t_L g394 ( .A(n_265), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g587 ( .A(n_265), .B(n_395), .Y(n_587) );
INVx1_ASAP7_75t_L g794 ( .A(n_265), .Y(n_794) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
BUFx4f_ASAP7_75t_L g344 ( .A(n_266), .Y(n_344) );
INVx3_ASAP7_75t_L g389 ( .A(n_266), .Y(n_389) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx2_ASAP7_75t_L g350 ( .A(n_268), .Y(n_350) );
INVx2_ASAP7_75t_L g355 ( .A(n_268), .Y(n_355) );
NAND2x1_ASAP7_75t_L g359 ( .A(n_268), .B(n_269), .Y(n_359) );
AND2x2_ASAP7_75t_L g376 ( .A(n_268), .B(n_269), .Y(n_376) );
INVx1_ASAP7_75t_L g385 ( .A(n_268), .Y(n_385) );
AND2x2_ASAP7_75t_L g399 ( .A(n_268), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_269), .B(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g354 ( .A(n_269), .B(n_355), .Y(n_354) );
BUFx2_ASAP7_75t_L g379 ( .A(n_269), .Y(n_379) );
INVx2_ASAP7_75t_L g400 ( .A(n_269), .Y(n_400) );
INVx1_ASAP7_75t_L g499 ( .A(n_269), .Y(n_499) );
AND2x2_ASAP7_75t_L g502 ( .A(n_269), .B(n_350), .Y(n_502) );
OR2x6_ASAP7_75t_L g388 ( .A(n_270), .B(n_389), .Y(n_388) );
INVxp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g373 ( .A(n_271), .Y(n_373) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x4_ASAP7_75t_L g383 ( .A(n_272), .B(n_384), .Y(n_383) );
BUFx2_ASAP7_75t_L g392 ( .A(n_272), .Y(n_392) );
OAI22xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_743), .B1(n_744), .B2(n_1038), .Y(n_273) );
INVx1_ASAP7_75t_L g1038 ( .A(n_274), .Y(n_1038) );
AO22x1_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_276), .B1(n_435), .B2(n_742), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
XNOR2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND3x1_ASAP7_75t_L g279 ( .A(n_280), .B(n_368), .C(n_405), .Y(n_279) );
NOR2xp33_ASAP7_75t_SL g280 ( .A(n_281), .B(n_338), .Y(n_280) );
OAI33xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_290), .A3(n_305), .B1(n_317), .B2(n_326), .B3(n_332), .Y(n_281) );
OAI33xp33_ASAP7_75t_L g771 ( .A1(n_282), .A2(n_332), .A3(n_772), .B1(n_775), .B2(n_778), .B3(n_783), .Y(n_771) );
OAI33xp33_ASAP7_75t_L g852 ( .A1(n_282), .A2(n_332), .A3(n_853), .B1(n_856), .B2(n_859), .B3(n_863), .Y(n_852) );
OAI33xp33_ASAP7_75t_L g1002 ( .A1(n_282), .A2(n_332), .A3(n_1003), .B1(n_1006), .B2(n_1009), .B3(n_1013), .Y(n_1002) );
BUFx4f_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx2_ASAP7_75t_L g561 ( .A(n_283), .Y(n_561) );
BUFx4f_ASAP7_75t_L g965 ( .A(n_283), .Y(n_965) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_287), .Y(n_283) );
AND2x2_ASAP7_75t_SL g366 ( .A(n_284), .B(n_367), .Y(n_366) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_284), .Y(n_434) );
INVx1_ASAP7_75t_L g513 ( .A(n_284), .Y(n_513) );
OR2x2_ASAP7_75t_L g1240 ( .A(n_284), .B(n_1241), .Y(n_1240) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g404 ( .A(n_285), .Y(n_404) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp33_ASAP7_75t_SL g287 ( .A(n_288), .B(n_289), .Y(n_287) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_288), .Y(n_432) );
AND3x4_ASAP7_75t_L g461 ( .A(n_288), .B(n_422), .C(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g1234 ( .A(n_288), .Y(n_1234) );
INVx3_ASAP7_75t_L g337 ( .A(n_289), .Y(n_337) );
BUFx3_ASAP7_75t_L g422 ( .A(n_289), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_292), .B1(n_297), .B2(n_298), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_291), .A2(n_329), .B1(n_343), .B2(n_345), .Y(n_342) );
OAI22xp33_ASAP7_75t_L g562 ( .A1(n_292), .A2(n_298), .B1(n_545), .B2(n_557), .Y(n_562) );
OAI22xp33_ASAP7_75t_L g573 ( .A1(n_292), .A2(n_330), .B1(n_546), .B2(n_559), .Y(n_573) );
OAI22xp33_ASAP7_75t_L g772 ( .A1(n_292), .A2(n_689), .B1(n_773), .B2(n_774), .Y(n_772) );
OAI22xp33_ASAP7_75t_L g783 ( .A1(n_292), .A2(n_330), .B1(n_784), .B2(n_785), .Y(n_783) );
OAI22xp33_ASAP7_75t_L g853 ( .A1(n_292), .A2(n_689), .B1(n_854), .B2(n_855), .Y(n_853) );
OAI22xp33_ASAP7_75t_L g863 ( .A1(n_292), .A2(n_330), .B1(n_864), .B2(n_865), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_292), .A2(n_298), .B1(n_1004), .B2(n_1005), .Y(n_1003) );
OAI22xp5_ASAP7_75t_L g1013 ( .A1(n_292), .A2(n_330), .B1(n_1014), .B2(n_1015), .Y(n_1013) );
BUFx4f_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g328 ( .A(n_293), .Y(n_328) );
OR2x4_ASAP7_75t_L g407 ( .A(n_293), .B(n_337), .Y(n_407) );
OR2x4_ASAP7_75t_L g428 ( .A(n_293), .B(n_410), .Y(n_428) );
BUFx3_ASAP7_75t_L g636 ( .A(n_293), .Y(n_636) );
BUFx3_ASAP7_75t_L g730 ( .A(n_293), .Y(n_730) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_294), .Y(n_304) );
INVx2_ASAP7_75t_L g311 ( .A(n_294), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_294), .B(n_303), .Y(n_316) );
AND2x4_ASAP7_75t_L g417 ( .A(n_294), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g469 ( .A(n_295), .Y(n_469) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVxp67_ASAP7_75t_L g310 ( .A(n_296), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_297), .A2(n_331), .B1(n_361), .B2(n_362), .Y(n_360) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g1339 ( .A(n_299), .Y(n_1339) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx4_ASAP7_75t_L g454 ( .A(n_300), .Y(n_454) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_300), .Y(n_637) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_300), .Y(n_689) );
OR2x2_ASAP7_75t_L g1298 ( .A(n_300), .B(n_1240), .Y(n_1298) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx3_ASAP7_75t_L g330 ( .A(n_301), .Y(n_330) );
BUFx2_ASAP7_75t_L g414 ( .A(n_301), .Y(n_414) );
NAND2x1p5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
BUFx2_ASAP7_75t_L g425 ( .A(n_302), .Y(n_425) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g418 ( .A(n_303), .Y(n_418) );
BUFx2_ASAP7_75t_L g423 ( .A(n_304), .Y(n_423) );
AND2x4_ASAP7_75t_L g477 ( .A(n_304), .B(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g886 ( .A(n_304), .Y(n_886) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B1(n_312), .B2(n_313), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_306), .A2(n_318), .B1(n_352), .B2(n_356), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g1006 ( .A1(n_307), .A2(n_313), .B1(n_1007), .B2(n_1008), .Y(n_1006) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g409 ( .A(n_308), .B(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g444 ( .A(n_308), .B(n_410), .Y(n_444) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_308), .Y(n_640) );
INVx2_ASAP7_75t_L g643 ( .A(n_308), .Y(n_643) );
BUFx6f_ASAP7_75t_L g734 ( .A(n_308), .Y(n_734) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g321 ( .A(n_309), .Y(n_321) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_309), .Y(n_565) );
BUFx8_ASAP7_75t_L g568 ( .A(n_309), .Y(n_568) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
AND2x4_ASAP7_75t_L g468 ( .A(n_311), .B(n_469), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_312), .A2(n_322), .B1(n_343), .B2(n_364), .Y(n_363) );
INVx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
CKINVDCx8_ASAP7_75t_R g735 ( .A(n_314), .Y(n_735) );
INVx3_ASAP7_75t_L g1012 ( .A(n_314), .Y(n_1012) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g571 ( .A(n_315), .Y(n_571) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_L g325 ( .A(n_316), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B1(n_322), .B2(n_323), .Y(n_317) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g737 ( .A(n_320), .Y(n_737) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_320), .B(n_1306), .Y(n_1305) );
INVx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g474 ( .A(n_321), .Y(n_474) );
INVx1_ASAP7_75t_L g483 ( .A(n_321), .Y(n_483) );
OAI22xp33_ASAP7_75t_SL g563 ( .A1(n_323), .A2(n_539), .B1(n_552), .B2(n_564), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_323), .A2(n_567), .B1(n_776), .B2(n_777), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_323), .A2(n_779), .B1(n_857), .B2(n_858), .Y(n_856) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x6_ASAP7_75t_L g429 ( .A(n_325), .B(n_337), .Y(n_429) );
BUFx3_ASAP7_75t_L g641 ( .A(n_325), .Y(n_641) );
OAI22xp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_329), .B1(n_330), .B2(n_331), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g970 ( .A(n_330), .Y(n_970) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
AND2x4_ASAP7_75t_L g340 ( .A(n_333), .B(n_341), .Y(n_340) );
OR2x6_ASAP7_75t_L g572 ( .A(n_333), .B(n_335), .Y(n_572) );
INVx1_ASAP7_75t_L g1267 ( .A(n_333), .Y(n_1267) );
BUFx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g462 ( .A(n_334), .Y(n_462) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
NAND3x1_ASAP7_75t_L g488 ( .A(n_336), .B(n_337), .C(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g410 ( .A(n_337), .Y(n_410) );
AND2x4_ASAP7_75t_L g416 ( .A(n_337), .B(n_417), .Y(n_416) );
AND2x4_ASAP7_75t_L g1233 ( .A(n_337), .B(n_1234), .Y(n_1233) );
OAI33xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_342), .A3(n_351), .B1(n_360), .B2(n_363), .B3(n_365), .Y(n_338) );
OAI33xp33_ASAP7_75t_L g786 ( .A1(n_339), .A2(n_787), .A3(n_789), .B1(n_790), .B2(n_791), .B3(n_792), .Y(n_786) );
OAI33xp33_ASAP7_75t_L g866 ( .A1(n_339), .A2(n_791), .A3(n_867), .B1(n_868), .B2(n_869), .B3(n_870), .Y(n_866) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g494 ( .A(n_340), .Y(n_494) );
INVx4_ASAP7_75t_L g550 ( .A(n_340), .Y(n_550) );
INVx2_ASAP7_75t_L g712 ( .A(n_340), .Y(n_712) );
OAI22xp33_ASAP7_75t_L g544 ( .A1(n_343), .A2(n_545), .B1(n_546), .B2(n_547), .Y(n_544) );
OAI22xp33_ASAP7_75t_L g787 ( .A1(n_343), .A2(n_773), .B1(n_784), .B2(n_788), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_343), .A2(n_364), .B1(n_854), .B2(n_864), .Y(n_867) );
INVx4_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_344), .Y(n_709) );
INVx3_ASAP7_75t_L g953 ( .A(n_344), .Y(n_953) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_345), .A2(n_552), .B1(n_553), .B2(n_554), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_345), .A2(n_553), .B1(n_1004), .B2(n_1014), .Y(n_1017) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx4_ASAP7_75t_L g364 ( .A(n_347), .Y(n_364) );
INVx1_ASAP7_75t_L g547 ( .A(n_347), .Y(n_547) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_347), .Y(n_615) );
INVx1_ASAP7_75t_L g788 ( .A(n_347), .Y(n_788) );
INVx8_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g391 ( .A(n_348), .B(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g758 ( .A(n_348), .B(n_373), .Y(n_758) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g625 ( .A(n_353), .Y(n_625) );
BUFx2_ASAP7_75t_L g1358 ( .A(n_353), .Y(n_1358) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g361 ( .A(n_354), .Y(n_361) );
INVx1_ASAP7_75t_L g541 ( .A(n_354), .Y(n_541) );
BUFx3_ASAP7_75t_L g556 ( .A(n_354), .Y(n_556) );
BUFx2_ASAP7_75t_L g620 ( .A(n_354), .Y(n_620) );
AND2x2_ASAP7_75t_L g498 ( .A(n_355), .B(n_499), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_356), .A2(n_540), .B1(n_776), .B2(n_780), .Y(n_789) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_356), .A2(n_540), .B1(n_857), .B2(n_861), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_356), .A2(n_540), .B1(n_855), .B2(n_865), .Y(n_869) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g370 ( .A(n_357), .Y(n_370) );
INVx1_ASAP7_75t_L g697 ( .A(n_357), .Y(n_697) );
INVx2_ASAP7_75t_L g1020 ( .A(n_357), .Y(n_1020) );
INVx2_ASAP7_75t_L g1359 ( .A(n_357), .Y(n_1359) );
INVx4_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_358), .Y(n_543) );
BUFx4f_ASAP7_75t_L g558 ( .A(n_358), .Y(n_558) );
BUFx4f_ASAP7_75t_L g651 ( .A(n_358), .Y(n_651) );
BUFx4f_ASAP7_75t_L g873 ( .A(n_358), .Y(n_873) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx3_ASAP7_75t_L g362 ( .A(n_359), .Y(n_362) );
INVx2_ASAP7_75t_SL g529 ( .A(n_362), .Y(n_529) );
BUFx2_ASAP7_75t_SL g627 ( .A(n_362), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_362), .A2(n_540), .B1(n_774), .B2(n_785), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_362), .A2(n_625), .B1(n_956), .B2(n_957), .Y(n_955) );
BUFx3_ASAP7_75t_L g1327 ( .A(n_362), .Y(n_1327) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_364), .A2(n_777), .B1(n_782), .B2(n_793), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_364), .A2(n_793), .B1(n_858), .B2(n_862), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g1021 ( .A1(n_364), .A2(n_553), .B1(n_1008), .B2(n_1011), .Y(n_1021) );
OAI33xp33_ASAP7_75t_L g537 ( .A1(n_365), .A2(n_538), .A3(n_544), .B1(n_548), .B2(n_551), .B3(n_555), .Y(n_537) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g791 ( .A(n_366), .Y(n_791) );
NAND3xp33_ASAP7_75t_L g807 ( .A(n_366), .B(n_808), .C(n_810), .Y(n_807) );
AOI33xp33_ASAP7_75t_L g930 ( .A1(n_366), .A2(n_931), .A3(n_932), .B1(n_934), .B2(n_938), .B3(n_939), .Y(n_930) );
AND2x4_ASAP7_75t_L g511 ( .A(n_367), .B(n_512), .Y(n_511) );
INVx4_ASAP7_75t_L g1283 ( .A(n_367), .Y(n_1283) );
OAI31xp33_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_387), .A3(n_393), .B(n_401), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g1360 ( .A1(n_370), .A2(n_1338), .B1(n_1351), .B2(n_1357), .Y(n_1360) );
NAND3xp33_ASAP7_75t_L g827 ( .A(n_371), .B(n_828), .C(n_832), .Y(n_827) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g925 ( .A(n_372), .Y(n_925) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
AND2x2_ASAP7_75t_L g378 ( .A(n_373), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g531 ( .A(n_373), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g924 ( .A(n_374), .Y(n_924) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g509 ( .A(n_375), .Y(n_509) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_376), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_380), .B1(n_381), .B2(n_386), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_378), .A2(n_383), .B1(n_908), .B2(n_910), .Y(n_921) );
AND2x4_ASAP7_75t_L g527 ( .A(n_379), .B(n_392), .Y(n_527) );
AND2x2_ASAP7_75t_L g579 ( .A(n_379), .B(n_392), .Y(n_579) );
BUFx2_ASAP7_75t_L g1295 ( .A(n_379), .Y(n_1295) );
AOI22xp33_ASAP7_75t_SL g419 ( .A1(n_380), .A2(n_420), .B1(n_424), .B2(n_426), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g874 ( .A1(n_381), .A2(n_579), .B1(n_875), .B2(n_876), .Y(n_874) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g530 ( .A(n_383), .Y(n_530) );
BUFx3_ASAP7_75t_L g581 ( .A(n_383), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_384), .B(n_1245), .Y(n_1300) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g916 ( .A(n_388), .Y(n_916) );
BUFx3_ASAP7_75t_L g553 ( .A(n_389), .Y(n_553) );
BUFx3_ASAP7_75t_L g612 ( .A(n_389), .Y(n_612) );
INVx2_ASAP7_75t_SL g723 ( .A(n_389), .Y(n_723) );
INVx2_ASAP7_75t_SL g1332 ( .A(n_390), .Y(n_1332) );
BUFx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g524 ( .A(n_391), .Y(n_524) );
INVx2_ASAP7_75t_L g589 ( .A(n_391), .Y(n_589) );
AND2x2_ASAP7_75t_L g830 ( .A(n_392), .B(n_806), .Y(n_830) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_394), .Y(n_522) );
BUFx2_ASAP7_75t_L g658 ( .A(n_394), .Y(n_658) );
AND2x4_ASAP7_75t_L g398 ( .A(n_395), .B(n_399), .Y(n_398) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
CKINVDCx16_ASAP7_75t_R g397 ( .A(n_398), .Y(n_397) );
INVx4_ASAP7_75t_L g760 ( .A(n_398), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g914 ( .A1(n_398), .A2(n_915), .B1(n_916), .B2(n_917), .Y(n_914) );
INVx2_ASAP7_75t_L g507 ( .A(n_399), .Y(n_507) );
BUFx3_ASAP7_75t_L g802 ( .A(n_399), .Y(n_802) );
BUFx6f_ASAP7_75t_L g936 ( .A(n_399), .Y(n_936) );
OAI31xp33_ASAP7_75t_L g574 ( .A1(n_401), .A2(n_575), .A3(n_576), .B(n_586), .Y(n_574) );
OAI31xp33_ASAP7_75t_L g871 ( .A1(n_401), .A2(n_872), .A3(n_877), .B(n_878), .Y(n_871) );
BUFx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g533 ( .A(n_402), .Y(n_533) );
BUFx3_ASAP7_75t_L g661 ( .A(n_402), .Y(n_661) );
BUFx2_ASAP7_75t_SL g703 ( .A(n_402), .Y(n_703) );
OAI31xp33_ASAP7_75t_L g1022 ( .A1(n_402), .A2(n_1023), .A3(n_1024), .B(n_1028), .Y(n_1022) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g1235 ( .A(n_404), .Y(n_1235) );
OR2x2_ASAP7_75t_L g1299 ( .A(n_404), .B(n_1300), .Y(n_1299) );
OAI31xp33_ASAP7_75t_SL g405 ( .A1(n_406), .A2(n_411), .A3(n_427), .B(n_430), .Y(n_405) );
INVx2_ASAP7_75t_SL g442 ( .A(n_407), .Y(n_442) );
INVx1_ASAP7_75t_L g676 ( .A(n_407), .Y(n_676) );
INVx2_ASAP7_75t_SL g988 ( .A(n_407), .Y(n_988) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI22xp33_ASAP7_75t_L g975 ( .A1(n_412), .A2(n_954), .B1(n_960), .B2(n_967), .Y(n_975) );
OAI22xp33_ASAP7_75t_L g1349 ( .A1(n_412), .A2(n_636), .B1(n_1350), .B2(n_1351), .Y(n_1349) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g646 ( .A(n_414), .Y(n_646) );
INVx1_ASAP7_75t_L g668 ( .A(n_414), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g763 ( .A(n_415), .B(n_764), .C(n_766), .Y(n_763) );
NAND3xp33_ASAP7_75t_SL g906 ( .A(n_415), .B(n_907), .C(n_909), .Y(n_906) );
CKINVDCx8_ASAP7_75t_R g415 ( .A(n_416), .Y(n_415) );
NOR3xp33_ASAP7_75t_L g445 ( .A(n_416), .B(n_446), .C(n_450), .Y(n_445) );
CKINVDCx8_ASAP7_75t_R g594 ( .A(n_416), .Y(n_594) );
INVx2_ASAP7_75t_L g471 ( .A(n_417), .Y(n_471) );
BUFx2_ASAP7_75t_L g481 ( .A(n_417), .Y(n_481) );
BUFx2_ASAP7_75t_L g597 ( .A(n_417), .Y(n_597) );
BUFx3_ASAP7_75t_L g768 ( .A(n_417), .Y(n_768) );
BUFx2_ASAP7_75t_L g842 ( .A(n_417), .Y(n_842) );
BUFx2_ASAP7_75t_L g1258 ( .A(n_417), .Y(n_1258) );
INVx1_ASAP7_75t_L g478 ( .A(n_418), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_420), .A2(n_424), .B1(n_910), .B2(n_911), .Y(n_909) );
AOI22xp5_ASAP7_75t_L g1034 ( .A1(n_420), .A2(n_883), .B1(n_1026), .B2(n_1035), .Y(n_1034) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_423), .Y(n_420) );
AND2x2_ASAP7_75t_L g424 ( .A(n_421), .B(n_425), .Y(n_424) );
AND2x4_ASAP7_75t_L g452 ( .A(n_421), .B(n_423), .Y(n_452) );
AND2x4_ASAP7_75t_L g456 ( .A(n_421), .B(n_425), .Y(n_456) );
AND2x2_ASAP7_75t_L g671 ( .A(n_421), .B(n_423), .Y(n_671) );
INVx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g883 ( .A(n_422), .B(n_884), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_424), .A2(n_452), .B1(n_755), .B2(n_765), .Y(n_764) );
AOI32xp33_ASAP7_75t_L g882 ( .A1(n_424), .A2(n_876), .A3(n_883), .B1(n_885), .B2(n_887), .Y(n_882) );
INVxp67_ASAP7_75t_L g1033 ( .A(n_424), .Y(n_1033) );
BUFx2_ASAP7_75t_L g447 ( .A(n_428), .Y(n_447) );
BUFx2_ASAP7_75t_L g664 ( .A(n_428), .Y(n_664) );
BUFx3_ASAP7_75t_L g685 ( .A(n_428), .Y(n_685) );
INVx2_ASAP7_75t_SL g845 ( .A(n_428), .Y(n_845) );
INVx2_ASAP7_75t_L g449 ( .A(n_429), .Y(n_449) );
BUFx3_ASAP7_75t_L g665 ( .A(n_429), .Y(n_665) );
INVx1_ASAP7_75t_L g996 ( .A(n_429), .Y(n_996) );
OAI31xp33_ASAP7_75t_L g761 ( .A1(n_430), .A2(n_762), .A3(n_763), .B(n_769), .Y(n_761) );
OAI21xp5_ASAP7_75t_L g837 ( .A1(n_430), .A2(n_838), .B(n_840), .Y(n_837) );
OAI31xp33_ASAP7_75t_SL g879 ( .A1(n_430), .A2(n_880), .A3(n_881), .B(n_888), .Y(n_879) );
OAI31xp33_ASAP7_75t_SL g1029 ( .A1(n_430), .A2(n_1030), .A3(n_1031), .B(n_1032), .Y(n_1029) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_433), .Y(n_430) );
AND2x4_ASAP7_75t_L g458 ( .A(n_431), .B(n_433), .Y(n_458) );
AND2x2_ASAP7_75t_L g599 ( .A(n_431), .B(n_433), .Y(n_599) );
AND2x2_ASAP7_75t_SL g679 ( .A(n_431), .B(n_433), .Y(n_679) );
INVx1_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g742 ( .A(n_435), .Y(n_742) );
XNOR2x1_ASAP7_75t_L g435 ( .A(n_436), .B(n_604), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_534), .B1(n_602), .B2(n_603), .Y(n_436) );
INVx1_ASAP7_75t_L g603 ( .A(n_437), .Y(n_603) );
NAND4xp25_ASAP7_75t_SL g438 ( .A(n_439), .B(n_459), .C(n_491), .D(n_518), .Y(n_438) );
AO21x1_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_445), .B(n_457), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .B1(n_443), .B2(n_444), .Y(n_440) );
INVx2_ASAP7_75t_SL g839 ( .A(n_442), .Y(n_839) );
INVx1_ASAP7_75t_L g592 ( .A(n_444), .Y(n_592) );
INVx2_ASAP7_75t_L g677 ( .A(n_444), .Y(n_677) );
INVx1_ASAP7_75t_L g694 ( .A(n_444), .Y(n_694) );
INVx1_ASAP7_75t_L g989 ( .A(n_444), .Y(n_989) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_449), .A2(n_829), .B1(n_831), .B2(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_452), .A2(n_456), .B1(n_580), .B2(n_585), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_452), .A2(n_456), .B1(n_691), .B2(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g991 ( .A(n_454), .Y(n_991) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_456), .Y(n_673) );
AOI222xp33_ASAP7_75t_L g841 ( .A1(n_456), .A2(n_833), .B1(n_834), .B2(n_835), .C1(n_842), .C2(n_843), .Y(n_841) );
CKINVDCx14_ASAP7_75t_R g457 ( .A(n_458), .Y(n_457) );
OAI31xp33_ASAP7_75t_L g683 ( .A1(n_458), .A2(n_684), .A3(n_686), .B(n_693), .Y(n_683) );
AOI33xp33_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_463), .A3(n_472), .B1(n_479), .B2(n_482), .B3(n_485), .Y(n_459) );
BUFx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g811 ( .A(n_461), .B(n_812), .C(n_815), .Y(n_811) );
INVx1_ASAP7_75t_L g897 ( .A(n_461), .Y(n_897) );
BUFx2_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI221xp5_ASAP7_75t_L g899 ( .A1(n_466), .A2(n_900), .B1(n_901), .B2(n_902), .C(n_903), .Y(n_899) );
INVx2_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
BUFx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx3_ASAP7_75t_L g818 ( .A(n_468), .Y(n_818) );
INVx8_ASAP7_75t_L g895 ( .A(n_468), .Y(n_895) );
NAND2x1p5_ASAP7_75t_L g1232 ( .A(n_468), .B(n_1233), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_470), .B(n_908), .Y(n_907) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g819 ( .A(n_471), .Y(n_819) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g484 ( .A(n_476), .Y(n_484) );
INVx5_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx3_ASAP7_75t_L g814 ( .A(n_477), .Y(n_814) );
BUFx12f_ASAP7_75t_L g822 ( .A(n_477), .Y(n_822) );
INVx1_ASAP7_75t_L g884 ( .A(n_478), .Y(n_884) );
BUFx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x4_ASAP7_75t_L g1263 ( .A(n_481), .B(n_1251), .Y(n_1263) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI33xp33_ASAP7_75t_L g634 ( .A1(n_486), .A2(n_561), .A3(n_635), .B1(n_638), .B2(n_642), .B3(n_644), .Y(n_634) );
OAI33xp33_ASAP7_75t_L g1335 ( .A1(n_486), .A2(n_561), .A3(n_1336), .B1(n_1340), .B2(n_1344), .B3(n_1349), .Y(n_1335) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g738 ( .A(n_487), .Y(n_738) );
INVx2_ASAP7_75t_L g974 ( .A(n_487), .Y(n_974) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g824 ( .A(n_488), .Y(n_824) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g1243 ( .A(n_490), .Y(n_1243) );
AOI33xp33_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_495), .A3(n_503), .B1(n_510), .B2(n_511), .B3(n_514), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OAI33xp33_ASAP7_75t_L g609 ( .A1(n_493), .A2(n_610), .A3(n_616), .B1(n_622), .B2(n_629), .B3(n_630), .Y(n_609) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
OAI33xp33_ASAP7_75t_L g1016 ( .A1(n_494), .A2(n_791), .A3(n_1017), .B1(n_1018), .B2(n_1019), .B3(n_1021), .Y(n_1016) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_SL g515 ( .A(n_497), .Y(n_515) );
INVx2_ASAP7_75t_L g933 ( .A(n_497), .Y(n_933) );
INVx1_ASAP7_75t_L g1290 ( .A(n_497), .Y(n_1290) );
INVx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx6f_ASAP7_75t_L g806 ( .A(n_498), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_498), .B(n_1245), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_498), .B(n_1273), .Y(n_1272) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g517 ( .A(n_502), .Y(n_517) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g629 ( .A(n_511), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g720 ( .A(n_511), .Y(n_720) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx3_ASAP7_75t_L g1278 ( .A(n_517), .Y(n_1278) );
AO21x1_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_533), .Y(n_518) );
NOR3xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .C(n_531), .Y(n_520) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g655 ( .A(n_527), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_527), .A2(n_581), .B1(n_755), .B2(n_756), .Y(n_754) );
AOI222xp33_ASAP7_75t_L g832 ( .A1(n_527), .A2(n_581), .B1(n_584), .B2(n_833), .C1(n_834), .C2(n_835), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g1025 ( .A1(n_527), .A2(n_581), .B1(n_1026), .B2(n_1027), .Y(n_1025) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_528), .A2(n_617), .B1(n_618), .B2(n_621), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_528), .A2(n_714), .B1(n_715), .B2(n_716), .Y(n_713) );
INVx5_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g700 ( .A(n_530), .Y(n_700) );
INVx2_ASAP7_75t_L g981 ( .A(n_530), .Y(n_981) );
INVx3_ASAP7_75t_L g577 ( .A(n_531), .Y(n_577) );
INVx1_ASAP7_75t_L g652 ( .A(n_531), .Y(n_652) );
INVx1_ASAP7_75t_L g983 ( .A(n_531), .Y(n_983) );
BUFx3_ASAP7_75t_L g584 ( .A(n_532), .Y(n_584) );
BUFx3_ASAP7_75t_L g937 ( .A(n_532), .Y(n_937) );
BUFx6f_ASAP7_75t_L g1280 ( .A(n_532), .Y(n_1280) );
AND2x6_ASAP7_75t_L g1285 ( .A(n_532), .B(n_1245), .Y(n_1285) );
AND2x4_ASAP7_75t_SL g1288 ( .A(n_532), .B(n_1273), .Y(n_1288) );
AO21x1_ASAP7_75t_L g913 ( .A1(n_533), .A2(n_914), .B(n_918), .Y(n_913) );
INVx3_ASAP7_75t_SL g602 ( .A(n_534), .Y(n_602) );
INVx1_ASAP7_75t_L g601 ( .A(n_535), .Y(n_601) );
NAND3xp33_ASAP7_75t_L g535 ( .A(n_536), .B(n_574), .C(n_590), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_560), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B1(n_542), .B2(n_543), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_540), .A2(n_558), .B1(n_1007), .B2(n_1010), .Y(n_1018) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g715 ( .A(n_541), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_542), .A2(n_554), .B1(n_567), .B2(n_569), .Y(n_566) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_543), .Y(n_753) );
BUFx3_ASAP7_75t_L g632 ( .A(n_547), .Y(n_632) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND3xp33_ASAP7_75t_L g798 ( .A(n_549), .B(n_799), .C(n_803), .Y(n_798) );
INVx2_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_SL g931 ( .A(n_550), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_558), .B2(n_559), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_556), .A2(n_1005), .B1(n_1015), .B2(n_1020), .Y(n_1019) );
OAI33xp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_562), .A3(n_563), .B1(n_566), .B2(n_572), .B3(n_573), .Y(n_560) );
OAI33xp33_ASAP7_75t_L g726 ( .A1(n_561), .A2(n_727), .A3(n_732), .B1(n_736), .B2(n_738), .B3(n_739), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_564), .A2(n_735), .B1(n_956), .B2(n_962), .Y(n_971) );
BUFx3_ASAP7_75t_L g1342 ( .A(n_564), .Y(n_1342) );
INVx5_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_565), .Y(n_813) );
INVx3_ASAP7_75t_L g860 ( .A(n_565), .Y(n_860) );
INVx2_ASAP7_75t_SL g973 ( .A(n_565), .Y(n_973) );
INVx3_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_SL g779 ( .A(n_568), .Y(n_779) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
BUFx3_ASAP7_75t_L g781 ( .A(n_571), .Y(n_781) );
OR2x2_ASAP7_75t_L g1239 ( .A(n_571), .B(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g903 ( .A(n_572), .Y(n_903) );
NAND3xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .C(n_583), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_580), .B1(n_581), .B2(n_582), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_579), .A2(n_691), .B1(n_699), .B2(n_700), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g1328 ( .A1(n_579), .A2(n_981), .B1(n_1320), .B2(n_1329), .Y(n_1328) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_581), .A2(n_654), .B1(n_655), .B2(n_656), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_582), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g659 ( .A(n_589), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_589), .A2(n_829), .B1(n_830), .B2(n_831), .Y(n_828) );
OAI31xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_593), .A3(n_598), .B(n_599), .Y(n_590) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .C(n_596), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g840 ( .A(n_594), .B(n_841), .C(n_844), .Y(n_840) );
OAI31xp33_ASAP7_75t_SL g904 ( .A1(n_599), .A2(n_905), .A3(n_906), .B(n_912), .Y(n_904) );
OA22x2_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B1(n_680), .B2(n_681), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_647), .C(n_662), .Y(n_607) );
NOR2xp33_ASAP7_75t_SL g608 ( .A(n_609), .B(n_634), .Y(n_608) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B1(n_613), .B2(n_614), .Y(n_610) );
OAI22xp33_ASAP7_75t_L g635 ( .A1(n_611), .A2(n_626), .B1(n_636), .B2(n_637), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_612), .A2(n_631), .B1(n_632), .B2(n_633), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_612), .A2(n_614), .B1(n_962), .B2(n_963), .Y(n_961) );
OAI22xp33_ASAP7_75t_L g644 ( .A1(n_613), .A2(n_628), .B1(n_636), .B2(n_645), .Y(n_644) );
OAI22xp5_ASAP7_75t_SL g951 ( .A1(n_614), .A2(n_952), .B1(n_953), .B2(n_954), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g1353 ( .A1(n_614), .A2(n_1337), .B1(n_1350), .B2(n_1354), .Y(n_1353) );
OAI22xp5_ASAP7_75t_L g1361 ( .A1(n_614), .A2(n_1343), .B1(n_1348), .B2(n_1354), .Y(n_1361) );
INVx6_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx5_ASAP7_75t_L g711 ( .A(n_615), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_617), .A2(n_631), .B1(n_639), .B2(n_641), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g958 ( .A1(n_618), .A2(n_627), .B1(n_959), .B2(n_960), .Y(n_958) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx4_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_621), .A2(n_633), .B1(n_641), .B2(n_643), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_626), .B1(n_627), .B2(n_628), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI33xp33_ASAP7_75t_L g950 ( .A1(n_629), .A2(n_712), .A3(n_951), .B1(n_955), .B2(n_958), .B3(n_961), .Y(n_950) );
OAI22xp33_ASAP7_75t_L g1336 ( .A1(n_636), .A2(n_1337), .B1(n_1338), .B2(n_1339), .Y(n_1336) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_641), .A2(n_716), .B1(n_725), .B2(n_737), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g972 ( .A1(n_641), .A2(n_957), .B1(n_963), .B2(n_973), .Y(n_972) );
OAI22xp5_ASAP7_75t_L g1344 ( .A1(n_641), .A2(n_1345), .B1(n_1347), .B2(n_1348), .Y(n_1344) );
INVxp67_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
OAI31xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_657), .A3(n_660), .B(n_661), .Y(n_647) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_651), .A2(n_715), .B1(n_718), .B2(n_719), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_654), .A2(n_670), .B1(n_672), .B2(n_673), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_655), .A2(n_980), .B1(n_981), .B2(n_982), .Y(n_979) );
OAI31xp33_ASAP7_75t_L g976 ( .A1(n_661), .A2(n_977), .A3(n_978), .B(n_984), .Y(n_976) );
OAI31xp33_ASAP7_75t_L g1323 ( .A1(n_661), .A2(n_1324), .A3(n_1330), .B(n_1333), .Y(n_1323) );
OAI31xp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_666), .A3(n_674), .B(n_678), .Y(n_662) );
INVxp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g731 ( .A(n_668), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_670), .A2(n_673), .B1(n_980), .B2(n_993), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1319 ( .A1(n_670), .A2(n_673), .B1(n_1320), .B2(n_1321), .Y(n_1319) );
BUFx3_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
BUFx3_ASAP7_75t_L g843 ( .A(n_671), .Y(n_843) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI31xp33_ASAP7_75t_L g985 ( .A1(n_678), .A2(n_986), .A3(n_990), .B(n_994), .Y(n_985) );
OAI31xp33_ASAP7_75t_L g1316 ( .A1(n_678), .A2(n_1317), .A3(n_1318), .B(n_1322), .Y(n_1316) );
BUFx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g740 ( .A(n_682), .Y(n_740) );
NAND3xp33_ASAP7_75t_L g682 ( .A(n_683), .B(n_695), .C(n_704), .Y(n_682) );
INVx2_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI22xp33_ASAP7_75t_L g739 ( .A1(n_689), .A2(n_710), .B1(n_719), .B2(n_728), .Y(n_739) );
OAI31xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_701), .A3(n_702), .B(n_703), .Y(n_695) );
OAI31xp33_ASAP7_75t_SL g751 ( .A1(n_703), .A2(n_752), .A3(n_757), .B(n_759), .Y(n_751) );
OAI21xp5_ASAP7_75t_L g826 ( .A1(n_703), .A2(n_827), .B(n_836), .Y(n_826) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_726), .Y(n_704) );
OAI33xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_712), .A3(n_713), .B1(n_717), .B2(n_720), .B3(n_721), .Y(n_705) );
OAI22xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B1(n_710), .B2(n_711), .Y(n_706) );
OAI22xp33_ASAP7_75t_L g727 ( .A1(n_707), .A2(n_718), .B1(n_728), .B2(n_731), .Y(n_727) );
INVx3_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_711), .A2(n_722), .B1(n_724), .B2(n_725), .Y(n_721) );
OAI33xp33_ASAP7_75t_L g1352 ( .A1(n_712), .A2(n_720), .A3(n_1353), .B1(n_1356), .B2(n_1360), .B3(n_1361), .Y(n_1352) );
OAI22xp33_ASAP7_75t_L g732 ( .A1(n_714), .A2(n_724), .B1(n_733), .B2(n_735), .Y(n_732) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVxp67_ASAP7_75t_SL g968 ( .A(n_730), .Y(n_968) );
INVx2_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g1340 ( .A1(n_735), .A2(n_1341), .B1(n_1342), .B2(n_1343), .Y(n_1340) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B1(n_946), .B2(n_1037), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AO22x1_ASAP7_75t_SL g746 ( .A1(n_747), .A2(n_748), .B1(n_846), .B2(n_945), .Y(n_746) );
INVx2_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
XNOR2x1_ASAP7_75t_L g748 ( .A(n_749), .B(n_795), .Y(n_748) );
NAND3xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_761), .C(n_770), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_756), .B(n_767), .Y(n_766) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g900 ( .A(n_768), .Y(n_900) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_771), .B(n_786), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_780), .B1(n_781), .B2(n_782), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_781), .A2(n_860), .B1(n_861), .B2(n_862), .Y(n_859) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NAND3xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_826), .C(n_837), .Y(n_796) );
AND4x1_ASAP7_75t_L g797 ( .A(n_798), .B(n_807), .C(n_811), .D(n_820), .Y(n_797) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g940 ( .A(n_805), .Y(n_940) );
INVx3_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
BUFx6f_ASAP7_75t_L g809 ( .A(n_806), .Y(n_809) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
NAND3xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_823), .C(n_825), .Y(n_820) );
BUFx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g945 ( .A(n_846), .Y(n_945) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_848), .B1(n_889), .B2(n_944), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
NAND3xp33_ASAP7_75t_L g850 ( .A(n_851), .B(n_871), .C(n_879), .Y(n_850) );
NOR2xp33_ASAP7_75t_SL g851 ( .A(n_852), .B(n_866), .Y(n_851) );
INVx2_ASAP7_75t_L g1346 ( .A(n_860), .Y(n_1346) );
INVx1_ASAP7_75t_L g1255 ( .A(n_884), .Y(n_1255) );
AND2x4_ASAP7_75t_SL g1250 ( .A(n_885), .B(n_1251), .Y(n_1250) );
INVx3_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVxp67_ASAP7_75t_SL g944 ( .A(n_889), .Y(n_944) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
OR2x2_ASAP7_75t_L g890 ( .A(n_891), .B(n_926), .Y(n_890) );
INVx1_ASAP7_75t_L g928 ( .A(n_892), .Y(n_928) );
AOI21xp5_ASAP7_75t_L g892 ( .A1(n_893), .A2(n_896), .B(n_898), .Y(n_892) );
INVx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx2_ASAP7_75t_L g1303 ( .A(n_895), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_904), .B(n_913), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_911), .B(n_923), .Y(n_922) );
NOR2xp33_ASAP7_75t_L g918 ( .A(n_919), .B(n_920), .Y(n_918) );
NAND3xp33_ASAP7_75t_L g920 ( .A(n_921), .B(n_922), .C(n_925), .Y(n_920) );
INVx2_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
OAI31xp33_ASAP7_75t_L g926 ( .A1(n_927), .A2(n_928), .A3(n_929), .B(n_941), .Y(n_926) );
INVx1_ASAP7_75t_L g943 ( .A(n_930), .Y(n_943) );
BUFx6f_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
AND2x4_ASAP7_75t_L g1275 ( .A(n_936), .B(n_1273), .Y(n_1275) );
INVx2_ASAP7_75t_L g1282 ( .A(n_936), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_942), .B(n_943), .Y(n_941) );
INVx1_ASAP7_75t_L g1037 ( .A(n_946), .Y(n_1037) );
OAI22xp33_ASAP7_75t_L g946 ( .A1(n_947), .A2(n_997), .B1(n_998), .B2(n_1036), .Y(n_946) );
INVx2_ASAP7_75t_SL g1036 ( .A(n_947), .Y(n_1036) );
NAND3xp33_ASAP7_75t_L g948 ( .A(n_949), .B(n_976), .C(n_985), .Y(n_948) );
NOR2xp33_ASAP7_75t_L g949 ( .A(n_950), .B(n_964), .Y(n_949) );
OAI22xp33_ASAP7_75t_L g966 ( .A1(n_952), .A2(n_959), .B1(n_967), .B2(n_969), .Y(n_966) );
INVx2_ASAP7_75t_SL g1355 ( .A(n_953), .Y(n_1355) );
OAI33xp33_ASAP7_75t_L g964 ( .A1(n_965), .A2(n_966), .A3(n_971), .B1(n_972), .B2(n_974), .B3(n_975), .Y(n_964) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx2_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g1009 ( .A1(n_973), .A2(n_1010), .B1(n_1011), .B2(n_1012), .Y(n_1009) );
INVx2_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
NAND3xp33_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1022), .C(n_1029), .Y(n_1000) );
NOR2xp33_ASAP7_75t_SL g1001 ( .A(n_1002), .B(n_1016), .Y(n_1001) );
OAI21xp5_ASAP7_75t_L g1039 ( .A1(n_1040), .A2(n_1047), .B(n_1225), .Y(n_1039) );
CKINVDCx20_ASAP7_75t_R g1040 ( .A(n_1041), .Y(n_1040) );
CKINVDCx20_ASAP7_75t_R g1041 ( .A(n_1042), .Y(n_1041) );
OAI22xp5_ASAP7_75t_SL g1102 ( .A1(n_1042), .A2(n_1103), .B1(n_1104), .B2(n_1105), .Y(n_1102) );
INVx2_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
AND2x6_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1045), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_1044), .B(n_1056), .Y(n_1055) );
AND2x4_ASAP7_75t_L g1058 ( .A(n_1044), .B(n_1059), .Y(n_1058) );
AND2x6_ASAP7_75t_L g1061 ( .A(n_1044), .B(n_1062), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_1044), .B(n_1056), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_1044), .B(n_1056), .Y(n_1096) );
OAI21xp5_ASAP7_75t_L g1364 ( .A1(n_1045), .A2(n_1365), .B(n_1366), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_1046), .B(n_1060), .Y(n_1059) );
AOI221xp5_ASAP7_75t_SL g1047 ( .A1(n_1048), .A2(n_1106), .B1(n_1163), .B2(n_1165), .C(n_1192), .Y(n_1047) );
A2O1A1Ixp33_ASAP7_75t_L g1048 ( .A1(n_1049), .A2(n_1081), .B(n_1092), .C(n_1101), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1076), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1066), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1052), .B(n_1073), .Y(n_1117) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1052), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1052), .B(n_1187), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1063), .Y(n_1052) );
INVx2_ASAP7_75t_L g1088 ( .A(n_1053), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_1053), .B(n_1091), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1053), .B(n_1086), .Y(n_1114) );
OR2x2_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1057), .Y(n_1053) );
INVxp67_ASAP7_75t_L g1105 ( .A(n_1055), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_1063), .B(n_1088), .Y(n_1087) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1063), .Y(n_1091) );
AND3x1_ASAP7_75t_L g1135 ( .A(n_1063), .B(n_1067), .C(n_1088), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1063), .B(n_1086), .Y(n_1137) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1063), .B(n_1067), .Y(n_1144) );
OAI32xp33_ASAP7_75t_L g1221 ( .A1(n_1063), .A2(n_1136), .A3(n_1146), .B1(n_1222), .B2(n_1224), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1065), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1066), .B(n_1151), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1066), .B(n_1087), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1072), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1067), .B(n_1090), .Y(n_1110) );
OR2x2_ASAP7_75t_L g1204 ( .A(n_1067), .B(n_1158), .Y(n_1204) );
INVx2_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
BUFx2_ASAP7_75t_L g1086 ( .A(n_1068), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_1068), .B(n_1090), .Y(n_1089) );
OR2x2_ASAP7_75t_L g1116 ( .A(n_1068), .B(n_1117), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1155 ( .A(n_1068), .B(n_1156), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1068), .B(n_1151), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1070), .Y(n_1068) );
NOR2xp33_ASAP7_75t_L g1113 ( .A(n_1072), .B(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1072), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_1072), .B(n_1137), .Y(n_1136) );
NOR2xp33_ASAP7_75t_L g1139 ( .A(n_1072), .B(n_1140), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1072), .B(n_1132), .Y(n_1191) );
INVx2_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1073), .Y(n_1084) );
OR2x2_ASAP7_75t_L g1142 ( .A(n_1073), .B(n_1078), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1073), .B(n_1151), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1073), .B(n_1098), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1073), .B(n_1078), .Y(n_1172) );
OR2x2_ASAP7_75t_L g1178 ( .A(n_1073), .B(n_1114), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1073), .B(n_1086), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1073), .B(n_1143), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1073), .B(n_1094), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1075), .Y(n_1073) );
INVx2_ASAP7_75t_L g1108 ( .A(n_1076), .Y(n_1108) );
A2O1A1Ixp33_ASAP7_75t_L g1111 ( .A1(n_1076), .A2(n_1112), .B(n_1113), .C(n_1115), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1076), .B(n_1126), .Y(n_1159) );
OR2x2_ASAP7_75t_L g1208 ( .A(n_1076), .B(n_1209), .Y(n_1208) );
INVx2_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1077), .B(n_1098), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1077), .B(n_1126), .Y(n_1199) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
OR2x2_ASAP7_75t_L g1127 ( .A(n_1078), .B(n_1098), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1078), .B(n_1133), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1078), .B(n_1098), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1080), .Y(n_1078) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_1082), .A2(n_1083), .B1(n_1085), .B2(n_1089), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1083), .B(n_1110), .Y(n_1109) );
INVx2_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
NAND2xp5_ASAP7_75t_L g1158 ( .A(n_1084), .B(n_1151), .Y(n_1158) );
O2A1O1Ixp33_ASAP7_75t_SL g1160 ( .A1(n_1084), .A2(n_1088), .B(n_1161), .C(n_1162), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1084), .B(n_1085), .Y(n_1194) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1085), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1087), .Y(n_1085) );
AOI221xp5_ASAP7_75t_L g1118 ( .A1(n_1086), .A2(n_1119), .B1(n_1123), .B2(n_1125), .C(n_1128), .Y(n_1118) );
OR2x2_ASAP7_75t_L g1124 ( .A(n_1086), .B(n_1088), .Y(n_1124) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1087), .Y(n_1140) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1087), .B(n_1090), .Y(n_1168) );
OAI332xp33_ASAP7_75t_L g1128 ( .A1(n_1088), .A2(n_1094), .A3(n_1098), .B1(n_1129), .B2(n_1131), .B3(n_1132), .C1(n_1134), .C2(n_1136), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1088), .B(n_1091), .Y(n_1151) );
O2A1O1Ixp33_ASAP7_75t_L g1173 ( .A1(n_1089), .A2(n_1174), .B(n_1176), .C(n_1177), .Y(n_1173) );
AOI22xp5_ASAP7_75t_L g1166 ( .A1(n_1091), .A2(n_1167), .B1(n_1169), .B2(n_1171), .Y(n_1166) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1098), .Y(n_1093) );
OR2x2_ASAP7_75t_L g1120 ( .A(n_1094), .B(n_1121), .Y(n_1120) );
CKINVDCx6p67_ASAP7_75t_R g1126 ( .A(n_1094), .Y(n_1126) );
CKINVDCx5p33_ASAP7_75t_R g1131 ( .A(n_1094), .Y(n_1131) );
OR2x2_ASAP7_75t_L g1179 ( .A(n_1094), .B(n_1098), .Y(n_1179) );
OR2x6_ASAP7_75t_L g1094 ( .A(n_1095), .B(n_1097), .Y(n_1094) );
OR2x2_ASAP7_75t_L g1112 ( .A(n_1095), .B(n_1097), .Y(n_1112) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1098), .Y(n_1133) );
OR2x2_ASAP7_75t_L g1146 ( .A(n_1098), .B(n_1126), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1098), .B(n_1172), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1098), .B(n_1126), .Y(n_1205) );
AND2x4_ASAP7_75t_L g1098 ( .A(n_1099), .B(n_1100), .Y(n_1098) );
INVx2_ASAP7_75t_SL g1152 ( .A(n_1101), .Y(n_1152) );
INVx2_ASAP7_75t_SL g1164 ( .A(n_1101), .Y(n_1164) );
NAND5xp2_ASAP7_75t_SL g1106 ( .A(n_1107), .B(n_1111), .C(n_1118), .D(n_1138), .E(n_1153), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1109), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_1108), .B(n_1181), .Y(n_1180) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1110), .Y(n_1161) );
OAI211xp5_ASAP7_75t_SL g1165 ( .A1(n_1112), .A2(n_1166), .B(n_1173), .C(n_1182), .Y(n_1165) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1114), .Y(n_1224) );
OAI21xp5_ASAP7_75t_L g1206 ( .A1(n_1115), .A2(n_1131), .B(n_1207), .Y(n_1206) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
NOR2xp33_ASAP7_75t_L g1218 ( .A(n_1120), .B(n_1155), .Y(n_1218) );
CKINVDCx6p67_ASAP7_75t_R g1121 ( .A(n_1122), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1122), .B(n_1130), .Y(n_1129) );
AOI221xp5_ASAP7_75t_L g1138 ( .A1(n_1122), .A2(n_1139), .B1(n_1141), .B2(n_1143), .C(n_1145), .Y(n_1138) );
OAI22xp5_ASAP7_75t_L g1182 ( .A1(n_1122), .A2(n_1183), .B1(n_1188), .B2(n_1191), .Y(n_1182) );
O2A1O1Ixp33_ASAP7_75t_L g1219 ( .A1(n_1122), .A2(n_1181), .B(n_1220), .C(n_1221), .Y(n_1219) );
A2O1A1Ixp33_ASAP7_75t_L g1202 ( .A1(n_1123), .A2(n_1130), .B(n_1203), .C(n_1205), .Y(n_1202) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
AOI221xp5_ASAP7_75t_L g1193 ( .A1(n_1125), .A2(n_1137), .B1(n_1194), .B2(n_1195), .C(n_1200), .Y(n_1193) );
NOR2xp33_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1127), .Y(n_1125) );
NOR2xp33_ASAP7_75t_L g1141 ( .A(n_1126), .B(n_1142), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1175 ( .A(n_1126), .B(n_1149), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1126), .B(n_1132), .Y(n_1217) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1127), .Y(n_1149) );
AOI21xp33_ASAP7_75t_L g1200 ( .A1(n_1127), .A2(n_1178), .B(n_1201), .Y(n_1200) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1132), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1132), .B(n_1223), .Y(n_1222) );
A2O1A1Ixp33_ASAP7_75t_L g1177 ( .A1(n_1134), .A2(n_1178), .B(n_1179), .C(n_1180), .Y(n_1177) );
INVx2_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1137), .Y(n_1147) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1142), .Y(n_1176) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
OAI211xp5_ASAP7_75t_SL g1145 ( .A1(n_1146), .A2(n_1147), .B(n_1148), .C(n_1152), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1149), .B(n_1150), .Y(n_1148) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1151), .Y(n_1211) );
O2A1O1Ixp33_ASAP7_75t_L g1153 ( .A1(n_1154), .A2(n_1157), .B(n_1159), .C(n_1160), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
NAND3xp33_ASAP7_75t_SL g1213 ( .A(n_1158), .B(n_1214), .C(n_1215), .Y(n_1213) );
NOR2xp33_ASAP7_75t_L g1188 ( .A(n_1162), .B(n_1189), .Y(n_1188) );
INVx3_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
AOI21xp33_ASAP7_75t_L g1195 ( .A1(n_1164), .A2(n_1196), .B(n_1198), .Y(n_1195) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
INVxp67_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVxp67_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
NOR2xp33_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1186), .Y(n_1184) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1187), .Y(n_1210) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
NAND5xp2_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1202), .C(n_1206), .D(n_1212), .E(n_1219), .Y(n_1192) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1205), .Y(n_1214) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1209), .Y(n_1220) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_1210), .B(n_1211), .Y(n_1209) );
AOI21xp5_ASAP7_75t_L g1212 ( .A1(n_1213), .A2(n_1217), .B(n_1218), .Y(n_1212) );
INVxp67_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1229), .B(n_1264), .Y(n_1228) );
AOI221xp5_ASAP7_75t_L g1229 ( .A1(n_1230), .A2(n_1236), .B1(n_1237), .B2(n_1246), .C(n_1247), .Y(n_1229) );
INVx3_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
OR2x6_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1235), .Y(n_1231) );
AND2x4_ASAP7_75t_L g1251 ( .A(n_1233), .B(n_1243), .Y(n_1251) );
AOI221xp5_ASAP7_75t_L g1276 ( .A1(n_1236), .A2(n_1277), .B1(n_1279), .B2(n_1284), .C(n_1285), .Y(n_1276) );
INVx8_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
AND2x4_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1242), .Y(n_1238) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1240), .Y(n_1304) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1240), .Y(n_1306) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1244), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1245), .B(n_1295), .Y(n_1294) );
NAND3xp33_ASAP7_75t_SL g1247 ( .A(n_1248), .B(n_1256), .C(n_1262), .Y(n_1247) );
AOI22xp5_ASAP7_75t_L g1248 ( .A1(n_1249), .A2(n_1250), .B1(n_1252), .B2(n_1253), .Y(n_1248) );
AOI222xp33_ASAP7_75t_L g1286 ( .A1(n_1249), .A2(n_1252), .B1(n_1287), .B2(n_1289), .C1(n_1291), .C2(n_1294), .Y(n_1286) );
AND2x4_ASAP7_75t_SL g1253 ( .A(n_1251), .B(n_1254), .Y(n_1253) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
AOI22xp5_ASAP7_75t_L g1256 ( .A1(n_1257), .A2(n_1259), .B1(n_1260), .B2(n_1261), .Y(n_1256) );
INVx3_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
AOI21xp5_ASAP7_75t_L g1264 ( .A1(n_1265), .A2(n_1268), .B(n_1296), .Y(n_1264) );
INVx2_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
BUFx2_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
NAND3xp33_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1276), .C(n_1286), .Y(n_1268) );
AOI22xp5_ASAP7_75t_L g1269 ( .A1(n_1270), .A2(n_1271), .B1(n_1274), .B2(n_1275), .Y(n_1269) );
AOI22xp33_ASAP7_75t_L g1301 ( .A1(n_1270), .A2(n_1274), .B1(n_1302), .B2(n_1305), .Y(n_1301) );
BUFx6f_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1273), .B(n_1278), .Y(n_1277) );
INVx2_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
BUFx3_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
INVx2_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
AND2x4_ASAP7_75t_L g1297 ( .A(n_1298), .B(n_1299), .Y(n_1297) );
AND2x4_ASAP7_75t_L g1302 ( .A(n_1303), .B(n_1304), .Y(n_1302) );
BUFx4f_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
INVxp67_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
HB1xp67_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
NAND3xp33_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1323), .C(n_1334), .Y(n_1315) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
NOR2xp33_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1352), .Y(n_1334) );
OAI22xp5_ASAP7_75t_L g1356 ( .A1(n_1341), .A2(n_1347), .B1(n_1357), .B2(n_1359), .Y(n_1356) );
INVx2_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
INVx2_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
INVx4_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
HB1xp67_ASAP7_75t_SL g1362 ( .A(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
endmodule