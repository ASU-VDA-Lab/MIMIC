module fake_jpeg_2965_n_111 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_22),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_34),
.B1(n_36),
.B2(n_29),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_0),
.B(n_1),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_37),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_12),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_38),
.B1(n_39),
.B2(n_35),
.Y(n_56)
);

AO22x2_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_46),
.B1(n_49),
.B2(n_2),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_38),
.B1(n_33),
.B2(n_40),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_46),
.B1(n_47),
.B2(n_54),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

OR2x4_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_43),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_3),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_63),
.Y(n_73)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_68),
.B1(n_63),
.B2(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_72),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_49),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_71),
.C(n_18),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_13),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_75),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_73),
.B(n_4),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_82),
.Y(n_92)
);

OR2x2_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_6),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_7),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_20),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_86),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_90),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_96),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_15),
.Y(n_96)
);

AOI221xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_82),
.B1(n_77),
.B2(n_7),
.C(n_8),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_99),
.A2(n_101),
.B(n_92),
.Y(n_102)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_103),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_93),
.C(n_87),
.Y(n_103)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_98),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_100),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_87),
.Y(n_108)
);

OAI221xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_99),
.B1(n_93),
.B2(n_14),
.C(n_23),
.Y(n_109)
);

OAI221xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_10),
.B1(n_11),
.B2(n_25),
.C(n_26),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_27),
.Y(n_111)
);


endmodule