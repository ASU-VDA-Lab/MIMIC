module fake_jpeg_20754_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx6_ASAP7_75t_SL g8 ( 
.A(n_7),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_19),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_12),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_7),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_9),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_15),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_22),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_28),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_20),
.B(n_10),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_32),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_21),
.B(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_17),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_14),
.B(n_13),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_8),
.C(n_11),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_13),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_40),
.B(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_30),
.B(n_27),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_34),
.B1(n_40),
.B2(n_39),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_11),
.C(n_8),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_45),
.B(n_6),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_49),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_1),
.C(n_2),
.Y(n_51)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_51),
.B(n_2),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_50),
.B(n_48),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_2),
.B(n_3),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_47),
.B1(n_49),
.B2(n_46),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B(n_3),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_4),
.C(n_5),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_4),
.Y(n_58)
);


endmodule