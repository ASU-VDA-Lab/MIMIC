module fake_netlist_1_9482_n_507 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_507);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_507;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_486;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g65 ( .A(n_35), .Y(n_65) );
INVx1_ASAP7_75t_L g66 ( .A(n_41), .Y(n_66) );
INVx1_ASAP7_75t_L g67 ( .A(n_53), .Y(n_67) );
NOR2xp33_ASAP7_75t_L g68 ( .A(n_56), .B(n_15), .Y(n_68) );
INVx1_ASAP7_75t_L g69 ( .A(n_28), .Y(n_69) );
INVxp67_ASAP7_75t_SL g70 ( .A(n_47), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_37), .Y(n_71) );
INVxp33_ASAP7_75t_SL g72 ( .A(n_4), .Y(n_72) );
CKINVDCx5p33_ASAP7_75t_R g73 ( .A(n_8), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_63), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_5), .Y(n_75) );
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_39), .Y(n_76) );
BUFx6f_ASAP7_75t_L g77 ( .A(n_3), .Y(n_77) );
NOR2xp33_ASAP7_75t_L g78 ( .A(n_49), .B(n_23), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_45), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_10), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_1), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_30), .Y(n_82) );
BUFx5_ASAP7_75t_L g83 ( .A(n_42), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_10), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_32), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_12), .Y(n_86) );
INVx2_ASAP7_75t_SL g87 ( .A(n_11), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_12), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_54), .Y(n_89) );
NOR2xp67_ASAP7_75t_L g90 ( .A(n_5), .B(n_58), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_57), .Y(n_91) );
CKINVDCx16_ASAP7_75t_R g92 ( .A(n_44), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_11), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_25), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_29), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_27), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_52), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_0), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_3), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_31), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_26), .Y(n_101) );
INVx3_ASAP7_75t_L g102 ( .A(n_51), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_48), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_55), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_65), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_93), .Y(n_106) );
AND2x4_ASAP7_75t_L g107 ( .A(n_102), .B(n_0), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_82), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_92), .Y(n_109) );
AND2x4_ASAP7_75t_L g110 ( .A(n_102), .B(n_1), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_87), .B(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_66), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_67), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_73), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_84), .Y(n_115) );
AND2x4_ASAP7_75t_L g116 ( .A(n_75), .B(n_6), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_72), .Y(n_117) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_69), .A2(n_33), .B(n_62), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_76), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_83), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_71), .Y(n_121) );
AND2x4_ASAP7_75t_L g122 ( .A(n_80), .B(n_7), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_70), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_77), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_81), .B(n_9), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_74), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_70), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_79), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_83), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_77), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_86), .B(n_9), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_85), .Y(n_132) );
CKINVDCx8_ASAP7_75t_R g133 ( .A(n_77), .Y(n_133) );
INVxp33_ASAP7_75t_SL g134 ( .A(n_90), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_88), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_77), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_105), .B(n_95), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_107), .B(n_98), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_108), .Y(n_139) );
INVx2_ASAP7_75t_SL g140 ( .A(n_107), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_120), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_107), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_110), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_110), .Y(n_144) );
INVx2_ASAP7_75t_SL g145 ( .A(n_110), .Y(n_145) );
INVx4_ASAP7_75t_L g146 ( .A(n_110), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_134), .B(n_96), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_116), .B(n_99), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_116), .B(n_104), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_116), .Y(n_150) );
OAI22xp5_ASAP7_75t_L g151 ( .A1(n_106), .A2(n_104), .B1(n_103), .B2(n_101), .Y(n_151) );
OR2x6_ASAP7_75t_SL g152 ( .A(n_109), .B(n_97), .Y(n_152) );
OAI22xp5_ASAP7_75t_L g153 ( .A1(n_117), .A2(n_100), .B1(n_94), .B2(n_91), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_116), .B(n_89), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_135), .B(n_83), .Y(n_155) );
BUFx2_ASAP7_75t_L g156 ( .A(n_114), .Y(n_156) );
OR2x6_ASAP7_75t_L g157 ( .A(n_122), .B(n_78), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_120), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_122), .B(n_78), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_120), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_105), .B(n_83), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_122), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_122), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_111), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_129), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_112), .B(n_83), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_112), .B(n_68), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_125), .Y(n_168) );
AND2x6_ASAP7_75t_L g169 ( .A(n_125), .B(n_68), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_119), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_118), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_113), .B(n_13), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_113), .B(n_14), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_131), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_123), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_129), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_121), .B(n_19), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_129), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_118), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_121), .B(n_20), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_127), .B(n_21), .Y(n_181) );
NAND2x1p5_ASAP7_75t_L g182 ( .A(n_131), .B(n_22), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_124), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_126), .B(n_24), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_126), .B(n_34), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_138), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_164), .B(n_128), .Y(n_187) );
CKINVDCx14_ASAP7_75t_R g188 ( .A(n_156), .Y(n_188) );
INVx4_ASAP7_75t_L g189 ( .A(n_146), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_146), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_141), .Y(n_191) );
BUFx4_ASAP7_75t_SL g192 ( .A(n_139), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_149), .B(n_132), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_141), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_182), .Y(n_195) );
BUFx8_ASAP7_75t_L g196 ( .A(n_170), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_138), .Y(n_197) );
INVx4_ASAP7_75t_L g198 ( .A(n_146), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_168), .B(n_115), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_158), .Y(n_200) );
BUFx2_ASAP7_75t_L g201 ( .A(n_170), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_174), .B(n_115), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_151), .A2(n_118), .B1(n_130), .B2(n_124), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_177), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_147), .B(n_133), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_155), .B(n_118), .Y(n_206) );
NOR2xp33_ASAP7_75t_R g207 ( .A(n_142), .B(n_36), .Y(n_207) );
BUFx3_ASAP7_75t_L g208 ( .A(n_182), .Y(n_208) );
NAND2xp33_ASAP7_75t_R g209 ( .A(n_159), .B(n_38), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_158), .Y(n_210) );
OR2x2_ASAP7_75t_L g211 ( .A(n_153), .B(n_136), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_160), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_152), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_160), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_171), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_143), .Y(n_216) );
AOI211xp5_ASAP7_75t_L g217 ( .A1(n_167), .A2(n_130), .B(n_124), .C(n_43), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_165), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_142), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_142), .Y(n_220) );
INVx8_ASAP7_75t_L g221 ( .A(n_157), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_148), .B(n_130), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_165), .Y(n_223) );
BUFx4f_ASAP7_75t_L g224 ( .A(n_177), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_177), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_144), .Y(n_226) );
BUFx2_ASAP7_75t_L g227 ( .A(n_169), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_150), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_162), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_148), .B(n_40), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_224), .A2(n_145), .B(n_140), .Y(n_231) );
BUFx2_ASAP7_75t_L g232 ( .A(n_188), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_191), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_189), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_193), .A2(n_221), .B1(n_227), .B2(n_197), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_204), .A2(n_154), .B1(n_163), .B2(n_148), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_191), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_187), .B(n_137), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_194), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_224), .A2(n_140), .B(n_145), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_186), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_192), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_199), .B(n_201), .Y(n_243) );
NAND2xp33_ASAP7_75t_L g244 ( .A(n_221), .B(n_179), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_194), .Y(n_245) );
BUFx6f_ASAP7_75t_SL g246 ( .A(n_230), .Y(n_246) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_206), .A2(n_184), .B(n_185), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_193), .B(n_154), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_196), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_204), .A2(n_157), .B1(n_169), .B2(n_181), .Y(n_250) );
NAND2xp33_ASAP7_75t_L g251 ( .A(n_221), .B(n_171), .Y(n_251) );
BUFx4_ASAP7_75t_SL g252 ( .A(n_213), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_202), .B(n_161), .Y(n_253) );
INVx3_ASAP7_75t_L g254 ( .A(n_189), .Y(n_254) );
AOI22x1_ASAP7_75t_L g255 ( .A1(n_206), .A2(n_179), .B1(n_171), .B2(n_178), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_201), .B(n_157), .Y(n_256) );
INVx5_ASAP7_75t_L g257 ( .A(n_221), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_195), .B(n_157), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_189), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_219), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_195), .B(n_175), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_200), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_233), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_238), .B(n_208), .Y(n_264) );
INVx4_ASAP7_75t_L g265 ( .A(n_257), .Y(n_265) );
AOI221xp5_ASAP7_75t_L g266 ( .A1(n_243), .A2(n_211), .B1(n_229), .B2(n_228), .C(n_226), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_233), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_237), .Y(n_268) );
INVx2_ASAP7_75t_SL g269 ( .A(n_257), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_256), .B(n_225), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_237), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_257), .B(n_208), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_257), .B(n_230), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_257), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_249), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_231), .A2(n_215), .B(n_230), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_253), .B(n_205), .Y(n_277) );
AOI22xp33_ASAP7_75t_SL g278 ( .A1(n_246), .A2(n_169), .B1(n_207), .B2(n_209), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_239), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_258), .B(n_198), .Y(n_280) );
BUFx2_ASAP7_75t_L g281 ( .A(n_232), .Y(n_281) );
A2O1A1Ixp33_ASAP7_75t_L g282 ( .A1(n_240), .A2(n_166), .B(n_220), .C(n_219), .Y(n_282) );
BUFx8_ASAP7_75t_L g283 ( .A(n_246), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_261), .A2(n_220), .B1(n_222), .B2(n_216), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_258), .B(n_198), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_267), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_264), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_271), .Y(n_288) );
OAI221xp5_ASAP7_75t_L g289 ( .A1(n_266), .A2(n_250), .B1(n_236), .B2(n_235), .C(n_248), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_277), .B(n_241), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_271), .B(n_262), .Y(n_291) );
INVx5_ASAP7_75t_L g292 ( .A(n_265), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_276), .A2(n_255), .B(n_215), .Y(n_293) );
BUFx3_ASAP7_75t_L g294 ( .A(n_274), .Y(n_294) );
OAI21x1_ASAP7_75t_L g295 ( .A1(n_267), .A2(n_247), .B(n_203), .Y(n_295) );
OA21x2_ASAP7_75t_L g296 ( .A1(n_282), .A2(n_247), .B(n_172), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_267), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_284), .A2(n_234), .B1(n_259), .B2(n_254), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_279), .Y(n_299) );
OAI221xp5_ASAP7_75t_L g300 ( .A1(n_278), .A2(n_217), .B1(n_242), .B2(n_260), .C(n_173), .Y(n_300) );
AO21x2_ASAP7_75t_L g301 ( .A1(n_279), .A2(n_172), .B(n_185), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_274), .Y(n_302) );
INVx4_ASAP7_75t_L g303 ( .A(n_292), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_286), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_289), .A2(n_283), .B1(n_281), .B2(n_270), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_292), .B(n_274), .Y(n_306) );
AOI211xp5_ASAP7_75t_L g307 ( .A1(n_300), .A2(n_281), .B(n_272), .C(n_285), .Y(n_307) );
OA21x2_ASAP7_75t_L g308 ( .A1(n_295), .A2(n_279), .B(n_263), .Y(n_308) );
CKINVDCx14_ASAP7_75t_R g309 ( .A(n_292), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_286), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_288), .B(n_263), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_288), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_292), .B(n_265), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_297), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_290), .B(n_285), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_292), .Y(n_316) );
INVxp67_ASAP7_75t_L g317 ( .A(n_290), .Y(n_317) );
BUFx3_ASAP7_75t_L g318 ( .A(n_294), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_291), .B(n_268), .Y(n_319) );
NAND2xp33_ASAP7_75t_SL g320 ( .A(n_302), .B(n_265), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_287), .B(n_285), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_299), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_291), .Y(n_323) );
OR2x6_ASAP7_75t_L g324 ( .A(n_302), .B(n_273), .Y(n_324) );
BUFx2_ASAP7_75t_L g325 ( .A(n_302), .Y(n_325) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_298), .A2(n_273), .B1(n_283), .B2(n_280), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_294), .A2(n_283), .B1(n_273), .B2(n_280), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_295), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_302), .B(n_268), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_296), .Y(n_330) );
OAI21x1_ASAP7_75t_L g331 ( .A1(n_293), .A2(n_239), .B(n_245), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_319), .B(n_302), .Y(n_332) );
NAND2xp33_ASAP7_75t_R g333 ( .A(n_316), .B(n_272), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_312), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_308), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_317), .B(n_275), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_312), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_315), .B(n_272), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_303), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_308), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_323), .B(n_296), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_308), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_323), .B(n_296), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_316), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_309), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_314), .Y(n_346) );
INVx2_ASAP7_75t_SL g347 ( .A(n_316), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_321), .B(n_272), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_308), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_311), .B(n_262), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_322), .Y(n_351) );
OAI222xp33_ASAP7_75t_L g352 ( .A1(n_326), .A2(n_269), .B1(n_280), .B2(n_252), .C1(n_254), .C2(n_234), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_322), .Y(n_353) );
NOR2x1_ASAP7_75t_L g354 ( .A(n_303), .B(n_251), .Y(n_354) );
INVx4_ASAP7_75t_L g355 ( .A(n_303), .Y(n_355) );
INVx2_ASAP7_75t_SL g356 ( .A(n_313), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_325), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_328), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_304), .Y(n_359) );
OAI22xp5_ASAP7_75t_SL g360 ( .A1(n_307), .A2(n_251), .B1(n_244), .B2(n_180), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_311), .B(n_245), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_304), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_310), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_310), .B(n_301), .Y(n_364) );
INVxp67_ASAP7_75t_SL g365 ( .A(n_329), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_328), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_325), .B(n_301), .Y(n_367) );
BUFx2_ASAP7_75t_L g368 ( .A(n_318), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_329), .B(n_301), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_330), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_330), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_318), .B(n_179), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_331), .Y(n_373) );
OAI31xp33_ASAP7_75t_L g374 ( .A1(n_305), .A2(n_222), .A3(n_190), .B(n_218), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_331), .Y(n_375) );
INVx4_ASAP7_75t_L g376 ( .A(n_355), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_334), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_346), .B(n_306), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_369), .B(n_313), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_365), .B(n_324), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_346), .Y(n_381) );
NOR2xp33_ASAP7_75t_R g382 ( .A(n_333), .B(n_320), .Y(n_382) );
NAND4xp25_ASAP7_75t_SL g383 ( .A(n_374), .B(n_327), .C(n_313), .D(n_306), .Y(n_383) );
INVx2_ASAP7_75t_SL g384 ( .A(n_368), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_341), .B(n_306), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_337), .B(n_324), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_337), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_351), .B(n_324), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_345), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_343), .B(n_324), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_343), .B(n_179), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_351), .B(n_222), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_370), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_332), .B(n_171), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_335), .Y(n_395) );
BUFx2_ASAP7_75t_L g396 ( .A(n_368), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_353), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_332), .B(n_46), .Y(n_398) );
OAI222xp33_ASAP7_75t_L g399 ( .A1(n_355), .A2(n_198), .B1(n_190), .B2(n_214), .C1(n_212), .C2(n_210), .Y(n_399) );
NAND3xp33_ASAP7_75t_L g400 ( .A(n_336), .B(n_183), .C(n_215), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_371), .B(n_50), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_353), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_371), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_364), .B(n_59), .Y(n_404) );
INVx2_ASAP7_75t_SL g405 ( .A(n_339), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_359), .Y(n_406) );
OAI21xp33_ASAP7_75t_SL g407 ( .A1(n_355), .A2(n_60), .B(n_61), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_364), .B(n_64), .Y(n_408) );
NAND2xp33_ASAP7_75t_SL g409 ( .A(n_355), .B(n_215), .Y(n_409) );
AOI22x1_ASAP7_75t_L g410 ( .A1(n_339), .A2(n_210), .B1(n_218), .B2(n_214), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_359), .B(n_200), .Y(n_411) );
NOR4xp25_ASAP7_75t_SL g412 ( .A(n_357), .B(n_215), .C(n_183), .D(n_212), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_350), .B(n_223), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_362), .B(n_223), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_335), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_352), .B(n_183), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_344), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_362), .Y(n_418) );
INVxp33_ASAP7_75t_L g419 ( .A(n_382), .Y(n_419) );
AOI211xp5_ASAP7_75t_L g420 ( .A1(n_383), .A2(n_360), .B(n_356), .C(n_347), .Y(n_420) );
NAND2x1_ASAP7_75t_L g421 ( .A(n_376), .B(n_357), .Y(n_421) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_389), .A2(n_360), .B1(n_338), .B2(n_348), .C(n_354), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_377), .Y(n_423) );
NAND2xp33_ASAP7_75t_L g424 ( .A(n_405), .B(n_354), .Y(n_424) );
NAND2xp5_ASAP7_75t_SL g425 ( .A(n_376), .B(n_363), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_377), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_396), .Y(n_427) );
AOI21xp5_ASAP7_75t_L g428 ( .A1(n_409), .A2(n_349), .B(n_342), .Y(n_428) );
NAND3xp33_ASAP7_75t_SL g429 ( .A(n_400), .B(n_372), .C(n_361), .Y(n_429) );
AOI21xp33_ASAP7_75t_SL g430 ( .A1(n_407), .A2(n_363), .B(n_372), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_379), .B(n_342), .Y(n_431) );
OAI221xp5_ASAP7_75t_L g432 ( .A1(n_416), .A2(n_358), .B1(n_366), .B2(n_349), .C(n_340), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_380), .A2(n_361), .B1(n_340), .B2(n_367), .Y(n_433) );
O2A1O1Ixp33_ASAP7_75t_L g434 ( .A1(n_399), .A2(n_367), .B(n_375), .C(n_373), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_396), .Y(n_435) );
A2O1A1Ixp33_ASAP7_75t_L g436 ( .A1(n_409), .A2(n_366), .B(n_375), .C(n_373), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_384), .B(n_366), .Y(n_437) );
NOR3xp33_ASAP7_75t_L g438 ( .A(n_392), .B(n_373), .C(n_178), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_385), .B(n_176), .Y(n_439) );
OAI322xp33_ASAP7_75t_L g440 ( .A1(n_378), .A2(n_176), .A3(n_190), .B1(n_388), .B2(n_386), .C1(n_381), .C2(n_397), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_387), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_387), .Y(n_442) );
OAI31xp33_ASAP7_75t_L g443 ( .A1(n_405), .A2(n_417), .A3(n_384), .B(n_398), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_417), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_403), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_398), .A2(n_404), .B1(n_408), .B2(n_390), .Y(n_446) );
CKINVDCx16_ASAP7_75t_R g447 ( .A(n_404), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_410), .B(n_408), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_388), .B(n_386), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g450 ( .A1(n_413), .A2(n_401), .B(n_414), .C(n_411), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g451 ( .A1(n_402), .A2(n_403), .B1(n_418), .B2(n_406), .C(n_393), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_423), .Y(n_452) );
NAND2xp33_ASAP7_75t_R g453 ( .A(n_430), .B(n_412), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_444), .Y(n_454) );
XNOR2xp5_ASAP7_75t_L g455 ( .A(n_419), .B(n_394), .Y(n_455) );
HAxp5_ASAP7_75t_SL g456 ( .A(n_446), .B(n_410), .CON(n_456), .SN(n_456) );
INVx1_ASAP7_75t_SL g457 ( .A(n_427), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_426), .Y(n_458) );
NOR2x1_ASAP7_75t_L g459 ( .A(n_429), .B(n_401), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_421), .Y(n_460) );
INVx2_ASAP7_75t_SL g461 ( .A(n_425), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_422), .B(n_395), .Y(n_462) );
AND2x2_ASAP7_75t_SL g463 ( .A(n_447), .B(n_415), .Y(n_463) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_420), .B(n_443), .C(n_434), .Y(n_464) );
INVx3_ASAP7_75t_SL g465 ( .A(n_435), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_450), .B(n_391), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_428), .B(n_391), .Y(n_467) );
OAI211xp5_ASAP7_75t_SL g468 ( .A1(n_432), .A2(n_394), .B(n_434), .C(n_448), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_440), .B(n_449), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_428), .A2(n_429), .B(n_424), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_441), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_465), .Y(n_472) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_464), .A2(n_438), .B(n_436), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_452), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_463), .A2(n_431), .B1(n_433), .B2(n_437), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_458), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_460), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_462), .B(n_451), .Y(n_478) );
AOI32xp33_ASAP7_75t_L g479 ( .A1(n_459), .A2(n_439), .A3(n_451), .B1(n_442), .B2(n_445), .Y(n_479) );
INVx2_ASAP7_75t_SL g480 ( .A(n_465), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_471), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_469), .B(n_466), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_460), .B(n_463), .Y(n_483) );
XNOR2xp5_ASAP7_75t_L g484 ( .A(n_455), .B(n_454), .Y(n_484) );
INVx1_ASAP7_75t_SL g485 ( .A(n_457), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_483), .B(n_470), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_482), .B(n_469), .Y(n_487) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_480), .Y(n_488) );
INVx2_ASAP7_75t_SL g489 ( .A(n_485), .Y(n_489) );
AND2x2_ASAP7_75t_SL g490 ( .A(n_478), .B(n_456), .Y(n_490) );
XOR2x2_ASAP7_75t_L g491 ( .A(n_484), .B(n_461), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_479), .B(n_461), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_483), .A2(n_467), .B(n_468), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_475), .A2(n_453), .B1(n_474), .B2(n_476), .Y(n_494) );
OAI221xp5_ASAP7_75t_SL g495 ( .A1(n_477), .A2(n_479), .B1(n_472), .B2(n_482), .C(n_464), .Y(n_495) );
AOI221x1_ASAP7_75t_L g496 ( .A1(n_477), .A2(n_482), .B1(n_464), .B2(n_473), .C(n_478), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_481), .A2(n_464), .B1(n_482), .B2(n_469), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_488), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_487), .B(n_486), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_489), .Y(n_500) );
AO22x2_ASAP7_75t_L g501 ( .A1(n_499), .A2(n_496), .B1(n_493), .B2(n_492), .Y(n_501) );
OAI211xp5_ASAP7_75t_SL g502 ( .A1(n_500), .A2(n_497), .B(n_494), .C(n_490), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_501), .Y(n_503) );
XOR2xp5_ASAP7_75t_L g504 ( .A(n_502), .B(n_498), .Y(n_504) );
XOR2xp5_ASAP7_75t_L g505 ( .A(n_504), .B(n_491), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_505), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_506), .A2(n_503), .B(n_495), .Y(n_507) );
endmodule