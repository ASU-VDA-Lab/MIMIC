module fake_jpeg_8040_n_132 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_18),
.A2(n_0),
.B(n_1),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_5),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_15),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_30),
.B1(n_12),
.B2(n_20),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_12),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_30)
);

OAI21xp33_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_21),
.B(n_13),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_31),
.A2(n_37),
.B1(n_21),
.B2(n_13),
.Y(n_52)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_SL g39 ( 
.A(n_26),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_12),
.B(n_20),
.C(n_16),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_17),
.B(n_16),
.C(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_42),
.B(n_46),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_44),
.Y(n_65)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_24),
.Y(n_47)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_22),
.B1(n_27),
.B2(n_25),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_49),
.Y(n_66)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_22),
.B1(n_27),
.B2(n_25),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_51),
.B(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_56),
.Y(n_57)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_9),
.C(n_2),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_14),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_68),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_62),
.B(n_16),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_13),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_70),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_36),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_67),
.C(n_69),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_26),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_14),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_14),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_10),
.Y(n_84)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_80),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_48),
.B(n_51),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_79),
.B(n_60),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_46),
.B1(n_51),
.B2(n_40),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_84),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_40),
.B(n_55),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_19),
.C(n_10),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_33),
.B1(n_49),
.B2(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_82),
.Y(n_96)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_55),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_73),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_57),
.C(n_64),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_91),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_57),
.B(n_60),
.Y(n_97)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_83),
.B(n_77),
.C(n_78),
.D(n_75),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_34),
.B(n_15),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_81),
.Y(n_103)
);

AOI321xp33_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_101),
.A3(n_92),
.B1(n_88),
.B2(n_93),
.C(n_98),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_79),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_103),
.C(n_104),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_107),
.B1(n_108),
.B2(n_88),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_74),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_92),
.C(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_110),
.A2(n_101),
.B(n_106),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_111),
.B(n_114),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_113),
.C(n_44),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_89),
.C(n_82),
.Y(n_113)
);

OAI321xp33_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_82),
.A3(n_89),
.B1(n_11),
.B2(n_6),
.C(n_8),
.Y(n_114)
);

AOI321xp33_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_117),
.A3(n_118),
.B1(n_15),
.B2(n_29),
.C(n_5),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_49),
.C(n_34),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_33),
.B1(n_17),
.B2(n_11),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_17),
.B1(n_116),
.B2(n_43),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_123),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_116),
.A2(n_8),
.B(n_4),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_122),
.C(n_124),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_5),
.B1(n_6),
.B2(n_1),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_116),
.A2(n_15),
.B(n_43),
.Y(n_124)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_120),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_126),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_29),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_127),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_125),
.B(n_128),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_129),
.B(n_29),
.Y(n_132)
);


endmodule