module fake_jpeg_18227_n_336 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_30),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_7),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_27),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_36),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_29),
.B1(n_22),
.B2(n_33),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_39),
.B1(n_67),
.B2(n_22),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_60),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_66),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_32),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_75),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_29),
.B1(n_22),
.B2(n_39),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_80),
.B1(n_94),
.B2(n_38),
.Y(n_108)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_73),
.Y(n_116)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_37),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_45),
.C(n_42),
.Y(n_118)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_67),
.B1(n_39),
.B2(n_62),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_22),
.B(n_29),
.C(n_36),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_82),
.Y(n_103)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_38),
.B1(n_26),
.B2(n_18),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_27),
.B1(n_18),
.B2(n_19),
.Y(n_119)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_39),
.B1(n_38),
.B2(n_27),
.Y(n_94)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_96),
.A2(n_97),
.B1(n_57),
.B2(n_61),
.Y(n_98)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_111),
.B1(n_119),
.B2(n_74),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_66),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_110),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_108),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_47),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_60),
.B1(n_61),
.B2(n_42),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_75),
.B(n_37),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_121),
.Y(n_135)
);

XNOR2x1_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_17),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_117),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_95),
.A2(n_64),
.B1(n_18),
.B2(n_19),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_114),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_36),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_115),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_37),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_41),
.C(n_34),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_45),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_45),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_125),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_42),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_26),
.B(n_19),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_126),
.A2(n_150),
.B(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_118),
.B1(n_99),
.B2(n_115),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_128),
.A2(n_122),
.B(n_109),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_154),
.Y(n_156)
);

OAI22x1_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_88),
.B1(n_95),
.B2(n_25),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_133),
.B1(n_134),
.B2(n_155),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_131),
.A2(n_136),
.B1(n_139),
.B2(n_147),
.Y(n_160)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_74),
.B1(n_72),
.B2(n_86),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_96),
.B1(n_32),
.B2(n_24),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_41),
.B1(n_91),
.B2(n_68),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_26),
.B(n_25),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_137),
.A2(n_149),
.B(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_41),
.B1(n_91),
.B2(n_68),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_109),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_142),
.A2(n_116),
.B1(n_106),
.B2(n_123),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_23),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_148),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_73),
.B1(n_34),
.B2(n_20),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_21),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_17),
.B(n_21),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_104),
.B(n_83),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_154),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_34),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_28),
.B1(n_17),
.B2(n_34),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_156),
.B(n_161),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_162),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_100),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_120),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_165),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_164),
.A2(n_166),
.B(n_170),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_143),
.B(n_34),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_171),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_100),
.B(n_105),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_105),
.Y(n_171)
);

OAI22x1_ASAP7_75t_L g215 ( 
.A1(n_173),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_116),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_146),
.A2(n_106),
.B1(n_101),
.B2(n_28),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_176),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_17),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_185),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_130),
.B1(n_133),
.B2(n_131),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_180),
.A2(n_148),
.B1(n_150),
.B2(n_137),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_132),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_181),
.Y(n_214)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

AO22x1_ASAP7_75t_L g183 ( 
.A1(n_130),
.A2(n_106),
.B1(n_101),
.B2(n_17),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_145),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_35),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_152),
.B(n_141),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_28),
.C(n_21),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_136),
.C(n_147),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_138),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_188),
.C(n_12),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_143),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_126),
.A2(n_35),
.B(n_31),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_189),
.A2(n_35),
.B(n_31),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_192),
.B(n_0),
.C(n_1),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_194),
.A2(n_207),
.B1(n_215),
.B2(n_218),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_160),
.B1(n_168),
.B2(n_180),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_148),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_202),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_169),
.A2(n_129),
.B1(n_144),
.B2(n_155),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_204),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_164),
.A2(n_144),
.B(n_31),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_166),
.B(n_7),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_216),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_28),
.Y(n_206)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_158),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_14),
.C(n_13),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_168),
.C(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_13),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_217),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_0),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_178),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_157),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_222),
.A2(n_229),
.B(n_204),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_238),
.B1(n_192),
.B2(n_194),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_219),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_159),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_230),
.Y(n_251)
);

NOR2x1_ASAP7_75t_R g229 ( 
.A(n_205),
.B(n_215),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_179),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_235),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_190),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_167),
.C(n_170),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_177),
.Y(n_237)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_199),
.A2(n_160),
.B1(n_176),
.B2(n_167),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_195),
.B(n_157),
.C(n_183),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_183),
.C(n_178),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_210),
.B(n_158),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_241),
.B(n_242),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_193),
.B(n_196),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_189),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_221),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_209),
.C(n_216),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_250),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_253),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_232),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_255),
.Y(n_277)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_257),
.A2(n_263),
.B(n_264),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_230),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_225),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_233),
.A2(n_208),
.B1(n_191),
.B2(n_202),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_261),
.A2(n_239),
.B1(n_240),
.B2(n_231),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_197),
.C(n_206),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_265),
.C(n_221),
.Y(n_269)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_222),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_197),
.C(n_211),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_229),
.A2(n_220),
.B1(n_234),
.B2(n_224),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_9),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_267),
.A2(n_270),
.B1(n_272),
.B2(n_264),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_269),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_263),
.A2(n_244),
.B1(n_222),
.B2(n_218),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_228),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_251),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_261),
.A2(n_203),
.B1(n_228),
.B2(n_3),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_275),
.B(n_8),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_9),
.C(n_8),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_250),
.C(n_265),
.Y(n_290)
);

AOI21x1_ASAP7_75t_L g282 ( 
.A1(n_253),
.A2(n_1),
.B(n_2),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_257),
.Y(n_286)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_285),
.A2(n_298),
.B1(n_281),
.B2(n_282),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_288),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_278),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_262),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_292),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_291),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_249),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_297),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_273),
.A2(n_252),
.B1(n_248),
.B2(n_260),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_258),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_296),
.A2(n_272),
.B(n_270),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_280),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_247),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_269),
.C(n_276),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_304),
.Y(n_319)
);

INVxp33_ASAP7_75t_SL g302 ( 
.A(n_286),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_302),
.B(n_306),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_303),
.A2(n_309),
.B(n_3),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_268),
.C(n_271),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_275),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_311),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_277),
.B(n_280),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_9),
.C(n_4),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_311),
.A2(n_296),
.B1(n_292),
.B2(n_5),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_314),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_3),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_315),
.A2(n_319),
.B(n_317),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_310),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g318 ( 
.A1(n_302),
.A2(n_3),
.B(n_4),
.Y(n_318)
);

AOI21x1_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_5),
.B(n_6),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_300),
.B(n_4),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_320),
.B(n_301),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_322),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_324),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_308),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_325),
.A2(n_327),
.B(n_304),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_317),
.A2(n_299),
.B(n_307),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_328),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_330),
.B(n_329),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_326),
.C(n_5),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_6),
.B(n_331),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_6),
.Y(n_336)
);


endmodule