module real_jpeg_17511_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_74;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_1),
.A2(n_37),
.B1(n_41),
.B2(n_42),
.Y(n_36)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_2),
.Y(n_101)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_3),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_3),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_4),
.Y(n_109)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_5),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_5),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_5),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_6),
.A2(n_95),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_6),
.Y(n_142)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_7),
.B(n_109),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_7),
.B(n_79),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_7),
.B(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_8),
.A2(n_81),
.B1(n_82),
.B2(n_88),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_8),
.A2(n_81),
.B1(n_111),
.B2(n_115),
.Y(n_110)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_130),
.Y(n_10)
);

OAI21x1_ASAP7_75t_SL g11 ( 
.A1(n_12),
.A2(n_105),
.B(n_129),
.Y(n_11)
);

NOR2x1_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_49),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_13),
.B(n_49),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_26),
.B1(n_35),
.B2(n_45),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_15),
.A2(n_27),
.B1(n_110),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_22),
.A2(n_23),
.B1(n_146),
.B2(n_150),
.Y(n_145)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_27),
.A2(n_57),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_27),
.A2(n_36),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_33),
.Y(n_126)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_40),
.Y(n_116)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_44),
.Y(n_141)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g139 ( 
.A(n_46),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_90),
.B2(n_91),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_50),
.B(n_91),
.Y(n_133)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_61),
.B1(n_79),
.B2(n_80),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_57),
.B(n_58),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVxp67_ASAP7_75t_SL g89 ( 
.A(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_59),
.Y(n_58)
);

OAI32xp33_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_92),
.A3(n_94),
.B1(n_96),
.B2(n_99),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_63),
.B1(n_65),
.B2(n_67),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_60),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_61),
.A2(n_79),
.B1(n_80),
.B2(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_71),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_122),
.B(n_128),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_117),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_127),
.Y(n_128)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_164),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_134),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_143),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_153),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AO22x2_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);


endmodule