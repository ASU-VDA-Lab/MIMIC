module real_aes_5673_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_979;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_919;
wire n_857;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_958;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_356;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_680;
wire n_595;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_468;
wire n_746;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_909;
wire n_996;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_960;
wire n_504;
wire n_973;
wire n_671;
wire n_725;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_501;
wire n_488;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_756;
wire n_598;
wire n_288;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_997;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_749;
wire n_358;
wire n_385;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_1001;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_972;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_312;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_968;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_823;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_0), .A2(n_77), .B1(n_370), .B2(n_376), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g986 ( .A1(n_1), .A2(n_168), .B1(n_376), .B2(n_987), .Y(n_986) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_2), .Y(n_714) );
AND2x4_ASAP7_75t_L g725 ( .A(n_2), .B(n_272), .Y(n_725) );
AND2x4_ASAP7_75t_L g730 ( .A(n_2), .B(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_SL g748 ( .A1(n_3), .A2(n_63), .B1(n_749), .B2(n_750), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_4), .A2(n_32), .B1(n_366), .B2(n_633), .Y(n_670) );
INVx1_ASAP7_75t_L g659 ( .A(n_5), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_6), .A2(n_130), .B1(n_442), .B2(n_514), .Y(n_548) );
INVx1_ASAP7_75t_L g701 ( .A(n_7), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_8), .A2(n_241), .B1(n_404), .B2(n_405), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_9), .A2(n_112), .B1(n_384), .B2(n_628), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_10), .A2(n_121), .B1(n_722), .B2(n_726), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_11), .A2(n_253), .B1(n_477), .B2(n_568), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_12), .A2(n_57), .B1(n_384), .B2(n_628), .Y(n_671) );
INVx1_ASAP7_75t_L g998 ( .A(n_13), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_14), .A2(n_231), .B1(n_379), .B2(n_381), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_15), .A2(n_93), .B1(n_477), .B2(n_691), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_16), .A2(n_265), .B1(n_450), .B2(n_451), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_17), .A2(n_134), .B1(n_627), .B2(n_629), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_18), .B(n_340), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_19), .A2(n_34), .B1(n_441), .B2(n_442), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_20), .A2(n_28), .B1(n_396), .B2(n_451), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_21), .A2(n_170), .B1(n_404), .B2(n_405), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_22), .A2(n_96), .B1(n_384), .B2(n_386), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_23), .A2(n_109), .B1(n_379), .B2(n_563), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_24), .A2(n_140), .B1(n_411), .B2(n_412), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_25), .A2(n_186), .B1(n_370), .B2(n_633), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_26), .B(n_1000), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_27), .A2(n_67), .B1(n_323), .B2(n_465), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_29), .A2(n_215), .B1(n_314), .B2(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_30), .A2(n_51), .B1(n_472), .B2(n_552), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_31), .A2(n_139), .B1(n_398), .B2(n_467), .Y(n_678) );
INVx1_ASAP7_75t_L g966 ( .A(n_33), .Y(n_966) );
AOI211x1_ASAP7_75t_L g957 ( .A1(n_35), .A2(n_958), .B(n_960), .C(n_969), .Y(n_957) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_36), .A2(n_41), .B1(n_656), .B2(n_680), .C(n_699), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_37), .A2(n_230), .B1(n_441), .B2(n_475), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_38), .A2(n_72), .B1(n_323), .B2(n_465), .Y(n_994) );
INVx1_ASAP7_75t_L g594 ( .A(n_39), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_40), .A2(n_142), .B1(n_620), .B2(n_968), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_42), .A2(n_157), .B1(n_447), .B2(n_448), .Y(n_446) );
AOI21xp33_ASAP7_75t_L g525 ( .A1(n_43), .A2(n_396), .B(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_44), .A2(n_239), .B1(n_682), .B2(n_683), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_45), .A2(n_60), .B1(n_362), .B2(n_442), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_46), .A2(n_116), .B1(n_745), .B2(n_747), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_47), .A2(n_193), .B1(n_631), .B2(n_632), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_48), .A2(n_656), .B(n_658), .Y(n_655) );
INVx1_ASAP7_75t_L g338 ( .A(n_49), .Y(n_338) );
INVx1_ASAP7_75t_L g311 ( .A(n_50), .Y(n_311) );
INVxp67_ASAP7_75t_L g347 ( .A(n_50), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_50), .B(n_219), .Y(n_355) );
INVx1_ASAP7_75t_L g544 ( .A(n_52), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_53), .A2(n_176), .B1(n_384), .B2(n_514), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_54), .B(n_463), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_55), .A2(n_97), .B1(n_314), .B2(n_323), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_56), .A2(n_143), .B1(n_480), .B2(n_635), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_58), .A2(n_169), .B1(n_608), .B2(n_680), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_59), .A2(n_196), .B1(n_749), .B2(n_750), .Y(n_786) );
XNOR2x1_ASAP7_75t_L g602 ( .A(n_61), .B(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_61), .A2(n_264), .B1(n_756), .B2(n_777), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_62), .A2(n_90), .B1(n_407), .B2(n_408), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_64), .B(n_296), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_65), .A2(n_127), .B1(n_323), .B2(n_520), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_66), .A2(n_261), .B1(n_381), .B2(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_68), .A2(n_210), .B1(n_516), .B2(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g436 ( .A(n_69), .Y(n_436) );
INVx1_ASAP7_75t_L g423 ( .A(n_70), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_71), .A2(n_74), .B1(n_366), .B2(n_628), .Y(n_955) );
INVx1_ASAP7_75t_L g488 ( .A(n_73), .Y(n_488) );
XNOR2x1_ASAP7_75t_L g535 ( .A(n_75), .B(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_75), .A2(n_128), .B1(n_722), .B2(n_726), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_76), .A2(n_126), .B1(n_434), .B2(n_448), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_78), .A2(n_216), .B1(n_411), .B2(n_412), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_79), .A2(n_269), .B1(n_478), .B2(n_516), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_80), .A2(n_131), .B1(n_507), .B2(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g700 ( .A(n_81), .Y(n_700) );
INVx2_ASAP7_75t_L g712 ( .A(n_82), .Y(n_712) );
INVx1_ASAP7_75t_L g724 ( .A(n_83), .Y(n_724) );
AND2x4_ASAP7_75t_L g727 ( .A(n_83), .B(n_712), .Y(n_727) );
INVx1_ASAP7_75t_SL g746 ( .A(n_83), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_84), .A2(n_254), .B1(n_323), .B2(n_396), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_85), .A2(n_222), .B1(n_404), .B2(n_405), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_86), .A2(n_167), .B1(n_318), .B2(n_323), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_87), .A2(n_202), .B1(n_441), .B2(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g973 ( .A(n_88), .Y(n_973) );
XOR2xp5_ASAP7_75t_L g982 ( .A(n_89), .B(n_983), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_91), .A2(n_178), .B1(n_477), .B2(n_478), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_92), .A2(n_248), .B1(n_448), .B2(n_450), .Y(n_662) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_94), .Y(n_296) );
XNOR2x2_ASAP7_75t_SL g578 ( .A(n_95), .B(n_579), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_95), .A2(n_171), .B1(n_749), .B2(n_750), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_98), .A2(n_179), .B1(n_520), .B2(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g417 ( .A(n_99), .Y(n_417) );
INVx1_ASAP7_75t_L g774 ( .A(n_100), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_101), .A2(n_208), .B1(n_516), .B2(n_651), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_102), .A2(n_333), .B(n_337), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_103), .A2(n_278), .B1(n_745), .B2(n_747), .Y(n_785) );
INVx1_ASAP7_75t_L g974 ( .A(n_103), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_103), .A2(n_980), .B1(n_982), .B2(n_1001), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_104), .A2(n_163), .B1(n_290), .B2(n_314), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_105), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g300 ( .A(n_106), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_106), .B(n_218), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_107), .A2(n_266), .B1(n_477), .B2(n_478), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_108), .A2(n_115), .B1(n_745), .B2(n_747), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_110), .A2(n_162), .B1(n_366), .B2(n_507), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_111), .A2(n_175), .B1(n_510), .B2(n_512), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_113), .A2(n_182), .B1(n_398), .B2(n_540), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g995 ( .A1(n_114), .A2(n_996), .B(n_997), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_117), .A2(n_165), .B1(n_323), .B2(n_465), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_118), .A2(n_255), .B1(n_433), .B2(n_598), .C(n_599), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_119), .A2(n_147), .B1(n_381), .B2(n_673), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_120), .A2(n_145), .B1(n_639), .B2(n_953), .Y(n_952) );
AOI221xp5_ASAP7_75t_L g574 ( .A1(n_122), .A2(n_245), .B1(n_467), .B2(n_530), .C(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_123), .A2(n_149), .B1(n_477), .B2(n_568), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_124), .A2(n_228), .B1(n_361), .B2(n_366), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_125), .A2(n_223), .B1(n_749), .B2(n_756), .Y(n_755) );
INVxp33_ASAP7_75t_SL g780 ( .A(n_129), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_132), .A2(n_148), .B1(n_606), .B2(n_607), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_133), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g600 ( .A(n_135), .Y(n_600) );
INVx1_ASAP7_75t_L g621 ( .A(n_136), .Y(n_621) );
XNOR2x1_ASAP7_75t_L g646 ( .A(n_137), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g653 ( .A(n_138), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_141), .A2(n_177), .B1(n_729), .B2(n_732), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_144), .A2(n_257), .B1(n_414), .B2(n_415), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_146), .A2(n_250), .B1(n_404), .B2(n_405), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_150), .A2(n_271), .B1(n_407), .B2(n_408), .Y(n_665) );
XOR2x2_ASAP7_75t_L g428 ( .A(n_151), .B(n_429), .Y(n_428) );
AOI21xp33_ASAP7_75t_L g541 ( .A1(n_152), .A2(n_542), .B(n_543), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_153), .A2(n_160), .B1(n_508), .B2(n_552), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_154), .A2(n_467), .B(n_468), .Y(n_466) );
INVx1_ASAP7_75t_L g589 ( .A(n_155), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_156), .A2(n_221), .B1(n_381), .B2(n_480), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_158), .A2(n_194), .B1(n_461), .B2(n_572), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_159), .A2(n_191), .B1(n_398), .B2(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g457 ( .A(n_161), .Y(n_457) );
INVx1_ASAP7_75t_L g778 ( .A(n_164), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_166), .A2(n_200), .B1(n_398), .B2(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_172), .A2(n_204), .B1(n_637), .B2(n_638), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_173), .A2(n_185), .B1(n_411), .B2(n_412), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_174), .A2(n_258), .B1(n_407), .B2(n_408), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_180), .A2(n_189), .B1(n_314), .B2(n_542), .Y(n_993) );
XOR2xp5_ASAP7_75t_L g286 ( .A(n_181), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g517 ( .A(n_183), .B(n_518), .Y(n_517) );
INVxp67_ASAP7_75t_L g532 ( .A(n_183), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_184), .A2(n_207), .B1(n_610), .B2(n_611), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_187), .A2(n_244), .B1(n_447), .B2(n_495), .Y(n_494) );
OA22x2_ASAP7_75t_L g294 ( .A1(n_188), .A2(n_219), .B1(n_295), .B2(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g329 ( .A(n_188), .Y(n_329) );
AOI21xp33_ASAP7_75t_L g613 ( .A1(n_190), .A2(n_614), .B(n_618), .Y(n_613) );
INVx1_ASAP7_75t_L g576 ( .A(n_192), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_195), .A2(n_240), .B1(n_381), .B2(n_480), .Y(n_693) );
INVx1_ASAP7_75t_L g624 ( .A(n_197), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_198), .A2(n_268), .B1(n_729), .B2(n_732), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_199), .A2(n_203), .B1(n_404), .B2(n_405), .Y(n_452) );
INVx1_ASAP7_75t_SL g684 ( .A(n_201), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_205), .A2(n_252), .B1(n_478), .B2(n_516), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_206), .A2(n_263), .B1(n_414), .B2(n_415), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_209), .A2(n_217), .B1(n_407), .B2(n_408), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_211), .A2(n_238), .B1(n_450), .B2(n_451), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_212), .A2(n_243), .B1(n_542), .B2(n_620), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_213), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g426 ( .A(n_214), .Y(n_426) );
INVx1_ASAP7_75t_L g313 ( .A(n_218), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_218), .B(n_327), .Y(n_358) );
OAI21xp33_ASAP7_75t_L g330 ( .A1(n_219), .A2(n_237), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g824 ( .A(n_220), .Y(n_824) );
INVx1_ASAP7_75t_L g823 ( .A(n_224), .Y(n_823) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_225), .B(n_334), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_226), .A2(n_259), .B1(n_475), .B2(n_514), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_227), .A2(n_247), .B1(n_552), .B2(n_583), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_229), .A2(n_246), .B1(n_745), .B2(n_747), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_232), .A2(n_233), .B1(n_480), .B2(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g961 ( .A(n_234), .Y(n_961) );
INVx1_ASAP7_75t_L g972 ( .A(n_235), .Y(n_972) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_236), .A2(n_277), .B1(n_431), .B2(n_433), .C(n_435), .Y(n_430) );
INVx1_ASAP7_75t_L g302 ( .A(n_237), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_237), .B(n_267), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_242), .A2(n_421), .B(n_422), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_249), .A2(n_270), .B1(n_414), .B2(n_415), .Y(n_500) );
INVx1_ASAP7_75t_L g469 ( .A(n_251), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_256), .A2(n_275), .B1(n_376), .B2(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_260), .B(n_616), .Y(n_677) );
INVx1_ASAP7_75t_L g527 ( .A(n_262), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_267), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g731 ( .A(n_272), .Y(n_731) );
HB1xp67_ASAP7_75t_L g1003 ( .A(n_272), .Y(n_1003) );
INVxp33_ASAP7_75t_L g772 ( .A(n_273), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_274), .A2(n_276), .B1(n_381), .B2(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g596 ( .A(n_279), .Y(n_596) );
AOI22x1_ASAP7_75t_L g558 ( .A1(n_280), .A2(n_559), .B1(n_560), .B2(n_577), .Y(n_558) );
INVx1_ASAP7_75t_L g577 ( .A(n_280), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_706), .B(n_715), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_481), .Y(n_282) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
AOI21xp33_ASAP7_75t_L g706 ( .A1(n_284), .A2(n_482), .B(n_707), .Y(n_706) );
XNOR2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_389), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NOR2x1_ASAP7_75t_SL g287 ( .A(n_288), .B(n_359), .Y(n_287) );
NAND3xp33_ASAP7_75t_L g288 ( .A(n_289), .B(n_317), .C(n_332), .Y(n_288) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx3_ASAP7_75t_L g396 ( .A(n_292), .Y(n_396) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_292), .Y(n_467) );
BUFx3_ASAP7_75t_L g542 ( .A(n_292), .Y(n_542) );
AND2x4_ASAP7_75t_L g292 ( .A(n_293), .B(n_303), .Y(n_292) );
AND2x4_ASAP7_75t_L g320 ( .A(n_293), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g434 ( .A(n_293), .B(n_321), .Y(n_434) );
AND2x4_ASAP7_75t_L g447 ( .A(n_293), .B(n_303), .Y(n_447) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
AND2x2_ASAP7_75t_L g316 ( .A(n_294), .B(n_298), .Y(n_316) );
AND2x2_ASAP7_75t_L g345 ( .A(n_294), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g373 ( .A(n_294), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_295), .B(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp33_ASAP7_75t_L g299 ( .A(n_296), .B(n_300), .Y(n_299) );
INVx3_ASAP7_75t_L g306 ( .A(n_296), .Y(n_306) );
NAND2xp33_ASAP7_75t_L g312 ( .A(n_296), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g331 ( .A(n_296), .Y(n_331) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_296), .Y(n_343) );
AND2x4_ASAP7_75t_L g372 ( .A(n_297), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_300), .B(n_329), .Y(n_328) );
OAI21xp5_ASAP7_75t_L g346 ( .A1(n_302), .A2(n_331), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g315 ( .A(n_303), .B(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g380 ( .A(n_303), .B(n_372), .Y(n_380) );
AND2x4_ASAP7_75t_L g404 ( .A(n_303), .B(n_372), .Y(n_404) );
AND2x4_ASAP7_75t_L g450 ( .A(n_303), .B(n_316), .Y(n_450) );
AND2x4_ASAP7_75t_L g303 ( .A(n_304), .B(n_308), .Y(n_303) );
INVx2_ASAP7_75t_L g322 ( .A(n_304), .Y(n_322) );
AND2x2_ASAP7_75t_L g341 ( .A(n_304), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g364 ( .A(n_304), .B(n_365), .Y(n_364) );
AND2x4_ASAP7_75t_L g374 ( .A(n_304), .B(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_306), .B(n_311), .Y(n_310) );
INVxp67_ASAP7_75t_L g327 ( .A(n_306), .Y(n_327) );
NAND3xp33_ASAP7_75t_L g357 ( .A(n_307), .B(n_326), .C(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g321 ( .A(n_308), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g365 ( .A(n_309), .Y(n_365) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx2_ASAP7_75t_L g612 ( .A(n_314), .Y(n_612) );
BUFx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_315), .Y(n_398) );
INVx2_ASAP7_75t_L g573 ( .A(n_315), .Y(n_573) );
AND2x2_ASAP7_75t_L g336 ( .A(n_316), .B(n_321), .Y(n_336) );
AND2x4_ASAP7_75t_L g362 ( .A(n_316), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g385 ( .A(n_316), .B(n_374), .Y(n_385) );
AND2x4_ASAP7_75t_L g411 ( .A(n_316), .B(n_374), .Y(n_411) );
AND2x4_ASAP7_75t_L g412 ( .A(n_316), .B(n_368), .Y(n_412) );
AND2x2_ASAP7_75t_L g421 ( .A(n_316), .B(n_321), .Y(n_421) );
AND2x2_ASAP7_75t_L g443 ( .A(n_316), .B(n_374), .Y(n_443) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx8_ASAP7_75t_SL g419 ( .A(n_320), .Y(n_419) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_320), .Y(n_465) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_320), .Y(n_520) );
BUFx3_ASAP7_75t_L g680 ( .A(n_320), .Y(n_680) );
INVx2_ASAP7_75t_L g965 ( .A(n_320), .Y(n_965) );
AND2x4_ASAP7_75t_L g324 ( .A(n_321), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g382 ( .A(n_321), .B(n_372), .Y(n_382) );
AND2x4_ASAP7_75t_L g405 ( .A(n_321), .B(n_372), .Y(n_405) );
AND2x4_ASAP7_75t_L g448 ( .A(n_321), .B(n_325), .Y(n_448) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx3_ASAP7_75t_L g522 ( .A(n_324), .Y(n_522) );
BUFx6f_ASAP7_75t_L g608 ( .A(n_324), .Y(n_608) );
AND2x4_ASAP7_75t_L g367 ( .A(n_325), .B(n_368), .Y(n_367) );
AND2x4_ASAP7_75t_L g388 ( .A(n_325), .B(n_374), .Y(n_388) );
AND2x4_ASAP7_75t_L g408 ( .A(n_325), .B(n_368), .Y(n_408) );
AND2x4_ASAP7_75t_L g415 ( .A(n_325), .B(n_374), .Y(n_415) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_330), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
BUFx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_335), .Y(n_617) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx3_ASAP7_75t_L g432 ( .A(n_336), .Y(n_432) );
OAI21xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_339), .B(n_348), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g997 ( .A1(n_339), .A2(n_998), .B(n_999), .Y(n_997) );
INVx4_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_341), .B(n_345), .Y(n_340) );
AND2x4_ASAP7_75t_L g401 ( .A(n_341), .B(n_345), .Y(n_401) );
AND2x2_ASAP7_75t_L g451 ( .A(n_341), .B(n_345), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g353 ( .A(n_343), .Y(n_353) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_350), .B(n_469), .Y(n_468) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_351), .Y(n_528) );
INVx1_ASAP7_75t_L g683 ( .A(n_351), .Y(n_683) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx3_ASAP7_75t_L g425 ( .A(n_352), .Y(n_425) );
AO21x2_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B(n_357), .Y(n_352) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_354), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
NAND4xp25_ASAP7_75t_SL g359 ( .A(n_360), .B(n_369), .C(n_378), .D(n_383), .Y(n_359) );
BUFx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_362), .Y(n_441) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_362), .Y(n_514) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_362), .Y(n_628) );
AND2x4_ASAP7_75t_L g407 ( .A(n_363), .B(n_372), .Y(n_407) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g368 ( .A(n_364), .Y(n_368) );
INVx1_ASAP7_75t_L g375 ( .A(n_365), .Y(n_375) );
BUFx3_ASAP7_75t_L g629 ( .A(n_366), .Y(n_629) );
BUFx12f_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx6_ASAP7_75t_L g473 ( .A(n_367), .Y(n_473) );
AND2x4_ASAP7_75t_L g377 ( .A(n_368), .B(n_372), .Y(n_377) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_371), .Y(n_477) );
BUFx12f_ASAP7_75t_L g516 ( .A(n_371), .Y(n_516) );
AND2x4_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
AND2x4_ASAP7_75t_L g414 ( .A(n_372), .B(n_374), .Y(n_414) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_377), .Y(n_507) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_377), .Y(n_552) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_377), .Y(n_633) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx12f_ASAP7_75t_L g480 ( .A(n_380), .Y(n_480) );
INVx3_ASAP7_75t_L g511 ( .A(n_380), .Y(n_511) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx3_ASAP7_75t_L g512 ( .A(n_382), .Y(n_512) );
BUFx5_ASAP7_75t_L g563 ( .A(n_382), .Y(n_563) );
BUFx3_ASAP7_75t_L g637 ( .A(n_384), .Y(n_637) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx8_ASAP7_75t_L g953 ( .A(n_385), .Y(n_953) );
INVx4_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g478 ( .A(n_387), .Y(n_478) );
INVx4_ASAP7_75t_L g568 ( .A(n_387), .Y(n_568) );
INVx1_ASAP7_75t_L g639 ( .A(n_387), .Y(n_639) );
INVx1_ASAP7_75t_L g651 ( .A(n_387), .Y(n_651) );
INVx2_ASAP7_75t_L g675 ( .A(n_387), .Y(n_675) );
INVx4_ASAP7_75t_L g691 ( .A(n_387), .Y(n_691) );
INVx8_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_453), .B2(n_454), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
XNOR2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_427), .Y(n_391) );
XOR2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_426), .Y(n_392) );
NOR4xp75_ASAP7_75t_L g393 ( .A(n_394), .B(n_402), .C(n_409), .D(n_416), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_397), .Y(n_394) );
INVx2_ASAP7_75t_L g959 ( .A(n_396), .Y(n_959) );
INVx3_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g461 ( .A(n_400), .Y(n_461) );
INVx4_ASAP7_75t_L g682 ( .A(n_400), .Y(n_682) );
INVx5_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g524 ( .A(n_401), .Y(n_524) );
BUFx2_ASAP7_75t_L g540 ( .A(n_401), .Y(n_540) );
BUFx4f_ASAP7_75t_L g620 ( .A(n_401), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_406), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_410), .B(n_413), .Y(n_409) );
OAI21x1_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_418), .B(n_420), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_419), .Y(n_606) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_421), .Y(n_598) );
INVx2_ASAP7_75t_L g657 ( .A(n_421), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_424), .B(n_544), .Y(n_543) );
INVx4_ASAP7_75t_L g623 ( .A(n_424), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_424), .B(n_700), .Y(n_699) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx4_ASAP7_75t_L g437 ( .A(n_425), .Y(n_437) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND3x1_ASAP7_75t_L g429 ( .A(n_430), .B(n_438), .C(n_444), .Y(n_429) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g463 ( .A(n_432), .Y(n_463) );
INVx2_ASAP7_75t_L g530 ( .A(n_432), .Y(n_530) );
INVx2_ASAP7_75t_L g546 ( .A(n_432), .Y(n_546) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g495 ( .A(n_437), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_437), .B(n_576), .Y(n_575) );
INVx4_ASAP7_75t_L g968 ( .A(n_437), .Y(n_968) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx4f_ASAP7_75t_L g475 ( .A(n_443), .Y(n_475) );
AND4x1_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .C(n_449), .D(n_452), .Y(n_444) );
INVx2_ASAP7_75t_L g590 ( .A(n_447), .Y(n_590) );
INVx2_ASAP7_75t_L g595 ( .A(n_448), .Y(n_595) );
INVx1_ASAP7_75t_L g593 ( .A(n_450), .Y(n_593) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
XNOR2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
NOR2xp67_ASAP7_75t_L g458 ( .A(n_459), .B(n_470), .Y(n_458) );
NAND4xp25_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .C(n_464), .D(n_466), .Y(n_459) );
NAND4xp25_ASAP7_75t_SL g470 ( .A(n_471), .B(n_474), .C(n_476), .D(n_479), .Y(n_470) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx5_ASAP7_75t_L g508 ( .A(n_473), .Y(n_508) );
INVx3_ASAP7_75t_L g583 ( .A(n_473), .Y(n_583) );
INVx1_ASAP7_75t_L g987 ( .A(n_473), .Y(n_987) );
BUFx2_ASAP7_75t_SL g631 ( .A(n_477), .Y(n_631) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
XNOR2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_642), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_553), .B1(n_640), .B2(n_641), .Y(n_483) );
INVx1_ASAP7_75t_L g641 ( .A(n_484), .Y(n_641) );
XNOR2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_534), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_501), .B1(n_502), .B2(n_533), .Y(n_485) );
INVx1_ASAP7_75t_L g533 ( .A(n_486), .Y(n_533) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
XNOR2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
OR2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_496), .Y(n_489) );
NAND4xp25_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .C(n_493), .D(n_494), .Y(n_490) );
NAND4xp25_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .C(n_499), .D(n_500), .Y(n_496) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OAI22x1_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_517), .B1(n_531), .B2(n_532), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_505), .B(n_518), .Y(n_531) );
NAND4xp25_ASAP7_75t_L g505 ( .A(n_506), .B(n_509), .C(n_513), .D(n_515), .Y(n_505) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g673 ( .A(n_511), .Y(n_673) );
NAND4xp25_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .C(n_525), .D(n_529), .Y(n_518) );
INVx2_ASAP7_75t_L g654 ( .A(n_520), .Y(n_654) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g971 ( .A(n_522), .Y(n_971) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_528), .B(n_600), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_528), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g1000 ( .A(n_528), .Y(n_1000) );
INVx2_ASAP7_75t_L g962 ( .A(n_530), .Y(n_962) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NOR2x1_ASAP7_75t_L g536 ( .A(n_537), .B(n_547), .Y(n_536) );
NAND4xp25_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .C(n_541), .D(n_545), .Y(n_537) );
BUFx2_ASAP7_75t_L g610 ( .A(n_542), .Y(n_610) );
NAND4xp25_ASAP7_75t_SL g547 ( .A(n_548), .B(n_549), .C(n_550), .D(n_551), .Y(n_547) );
INVx1_ASAP7_75t_L g640 ( .A(n_553), .Y(n_640) );
XOR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_602), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_556), .B1(n_578), .B2(n_601), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND4xp75_ASAP7_75t_L g560 ( .A(n_561), .B(n_565), .C(n_569), .D(n_574), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
BUFx3_ASAP7_75t_L g635 ( .A(n_563), .Y(n_635) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g601 ( .A(n_578), .Y(n_601) );
NAND4xp75_ASAP7_75t_L g579 ( .A(n_580), .B(n_584), .C(n_587), .D(n_597), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_592), .Y(n_587) );
OAI21xp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B(n_591), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B1(n_595), .B2(n_596), .Y(n_592) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_625), .Y(n_603) );
NAND3xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_609), .C(n_613), .Y(n_604) );
BUFx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g969 ( .A1(n_612), .A2(n_970), .B1(n_972), .B2(n_973), .Y(n_969) );
INVx2_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g996 ( .A(n_617), .Y(n_996) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_621), .B1(n_622), .B2(n_624), .Y(n_618) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND4xp25_ASAP7_75t_SL g625 ( .A(n_626), .B(n_630), .C(n_634), .D(n_636), .Y(n_625) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
BUFx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_666), .B1(n_704), .B2(n_705), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_645), .Y(n_705) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND4xp75_ASAP7_75t_L g647 ( .A(n_648), .B(n_652), .C(n_660), .D(n_663), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
OA21x2_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B(n_655), .Y(n_652) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g704 ( .A(n_666), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_685), .B1(n_702), .B2(n_703), .Y(n_666) );
INVx1_ASAP7_75t_SL g702 ( .A(n_667), .Y(n_702) );
XOR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_684), .Y(n_667) );
NOR2x1_ASAP7_75t_L g668 ( .A(n_669), .B(n_676), .Y(n_668) );
NAND4xp25_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .C(n_672), .D(n_674), .Y(n_669) );
NAND4xp25_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .C(n_679), .D(n_681), .Y(n_676) );
BUFx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g703 ( .A(n_686), .Y(n_703) );
XNOR2x1_ASAP7_75t_L g686 ( .A(n_687), .B(n_701), .Y(n_686) );
NAND4xp75_ASAP7_75t_L g687 ( .A(n_688), .B(n_692), .C(n_695), .D(n_698), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
BUFx3_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_713), .C(n_714), .Y(n_709) );
AND2x2_ASAP7_75t_L g976 ( .A(n_710), .B(n_977), .Y(n_976) );
AND2x2_ASAP7_75t_L g981 ( .A(n_710), .B(n_978), .Y(n_981) );
AOI21xp5_ASAP7_75t_L g1004 ( .A1(n_710), .A2(n_714), .B(n_746), .Y(n_1004) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AO21x1_ASAP7_75t_L g1002 ( .A1(n_711), .A2(n_1003), .B(n_1004), .Y(n_1002) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g723 ( .A(n_712), .B(n_724), .Y(n_723) );
AND3x4_ASAP7_75t_L g745 ( .A(n_712), .B(n_730), .C(n_746), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_713), .B(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_714), .Y(n_978) );
OAI221xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_942), .B1(n_945), .B2(n_975), .C(n_979), .Y(n_715) );
AOI211xp5_ASAP7_75t_SL g716 ( .A1(n_717), .A2(n_733), .B(n_810), .C(n_900), .Y(n_716) );
NOR3xp33_ASAP7_75t_L g931 ( .A(n_717), .B(n_932), .C(n_933), .Y(n_931) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_718), .A2(n_842), .B1(n_848), .B2(n_867), .Y(n_841) );
AOI21xp33_ASAP7_75t_SL g884 ( .A1(n_718), .A2(n_848), .B(n_885), .Y(n_884) );
AND2x2_ASAP7_75t_L g889 ( .A(n_718), .B(n_890), .Y(n_889) );
BUFx3_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g840 ( .A(n_719), .Y(n_840) );
AND2x2_ASAP7_75t_L g887 ( .A(n_719), .B(n_768), .Y(n_887) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g847 ( .A(n_720), .Y(n_847) );
OR2x2_ASAP7_75t_L g894 ( .A(n_720), .B(n_784), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_728), .Y(n_720) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .Y(n_722) );
AND2x4_ASAP7_75t_L g729 ( .A(n_723), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g749 ( .A(n_723), .B(n_725), .Y(n_749) );
AND2x4_ASAP7_75t_L g777 ( .A(n_723), .B(n_725), .Y(n_777) );
AND2x2_ASAP7_75t_L g726 ( .A(n_725), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g750 ( .A(n_725), .B(n_727), .Y(n_750) );
AND2x4_ASAP7_75t_L g756 ( .A(n_725), .B(n_727), .Y(n_756) );
AND2x4_ASAP7_75t_L g732 ( .A(n_727), .B(n_730), .Y(n_732) );
AND2x4_ASAP7_75t_L g747 ( .A(n_727), .B(n_730), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_727), .B(n_730), .Y(n_773) );
INVx3_ASAP7_75t_L g771 ( .A(n_729), .Y(n_771) );
A2O1A1Ixp33_ASAP7_75t_SL g733 ( .A1(n_734), .A2(n_758), .B(n_781), .C(n_787), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AOI221xp5_ASAP7_75t_L g826 ( .A1(n_735), .A2(n_766), .B1(n_783), .B2(n_815), .C(n_827), .Y(n_826) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_754), .Y(n_735) );
AND2x2_ASAP7_75t_L g788 ( .A(n_736), .B(n_789), .Y(n_788) );
NOR2x1_ASAP7_75t_L g736 ( .A(n_737), .B(n_741), .Y(n_736) );
INVx2_ASAP7_75t_L g761 ( .A(n_737), .Y(n_761) );
INVx2_ASAP7_75t_L g799 ( .A(n_737), .Y(n_799) );
INVx1_ASAP7_75t_L g804 ( .A(n_737), .Y(n_804) );
AND2x2_ASAP7_75t_L g807 ( .A(n_737), .B(n_808), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_737), .B(n_814), .Y(n_813) );
BUFx6f_ASAP7_75t_L g817 ( .A(n_737), .Y(n_817) );
AND2x2_ASAP7_75t_L g850 ( .A(n_737), .B(n_765), .Y(n_850) );
AND2x2_ASAP7_75t_L g857 ( .A(n_737), .B(n_858), .Y(n_857) );
NAND2xp5_ASAP7_75t_SL g866 ( .A(n_737), .B(n_830), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_737), .B(n_878), .Y(n_877) );
NAND2xp5_ASAP7_75t_SL g907 ( .A(n_737), .B(n_865), .Y(n_907) );
NAND2xp5_ASAP7_75t_SL g910 ( .A(n_737), .B(n_911), .Y(n_910) );
AND2x2_ASAP7_75t_L g934 ( .A(n_737), .B(n_769), .Y(n_934) );
INVx4_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OR2x2_ASAP7_75t_L g837 ( .A(n_738), .B(n_763), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_738), .B(n_768), .Y(n_922) );
AND2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
AOI21xp33_ASAP7_75t_L g860 ( .A1(n_741), .A2(n_861), .B(n_862), .Y(n_860) );
INVx3_ASAP7_75t_SL g865 ( .A(n_741), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_741), .B(n_763), .Y(n_870) );
OR2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_751), .Y(n_741) );
AND2x2_ASAP7_75t_L g765 ( .A(n_742), .B(n_751), .Y(n_765) );
AND2x2_ASAP7_75t_L g814 ( .A(n_742), .B(n_789), .Y(n_814) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OR2x2_ASAP7_75t_L g792 ( .A(n_743), .B(n_751), .Y(n_792) );
AND2x2_ASAP7_75t_L g819 ( .A(n_743), .B(n_751), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_743), .B(n_754), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_743), .B(n_880), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_743), .B(n_789), .Y(n_912) );
AND2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_748), .Y(n_743) );
AND2x2_ASAP7_75t_L g802 ( .A(n_751), .B(n_763), .Y(n_802) );
INVx1_ASAP7_75t_L g859 ( .A(n_751), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_751), .B(n_789), .Y(n_861) );
AND2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx1_ASAP7_75t_SL g764 ( .A(n_754), .Y(n_764) );
INVx1_ASAP7_75t_L g789 ( .A(n_754), .Y(n_789) );
OR2x2_ASAP7_75t_L g800 ( .A(n_754), .B(n_792), .Y(n_800) );
AND2x2_ASAP7_75t_L g858 ( .A(n_754), .B(n_859), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_754), .B(n_865), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_754), .B(n_850), .Y(n_874) );
AND2x2_ASAP7_75t_L g754 ( .A(n_755), .B(n_757), .Y(n_754) );
INVx2_ASAP7_75t_L g779 ( .A(n_756), .Y(n_779) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
AOI211xp5_ASAP7_75t_SL g811 ( .A1(n_759), .A2(n_766), .B(n_812), .C(n_815), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_766), .Y(n_759) );
NAND2xp67_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_761), .B(n_856), .Y(n_862) );
AOI221xp5_ASAP7_75t_L g892 ( .A1(n_762), .A2(n_821), .B1(n_893), .B2(n_895), .C(n_897), .Y(n_892) );
O2A1O1Ixp33_ASAP7_75t_L g901 ( .A1(n_762), .A2(n_788), .B(n_889), .C(n_902), .Y(n_901) );
AND2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_765), .Y(n_762) );
AND2x4_ASAP7_75t_L g790 ( .A(n_763), .B(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g836 ( .A(n_765), .Y(n_836) );
AND2x2_ASAP7_75t_L g914 ( .A(n_765), .B(n_789), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_765), .B(n_941), .Y(n_940) );
AOI21xp5_ASAP7_75t_L g863 ( .A1(n_766), .A2(n_864), .B(n_866), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_766), .B(n_894), .Y(n_908) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
OR2x2_ASAP7_75t_L g794 ( .A(n_768), .B(n_784), .Y(n_794) );
AND2x2_ASAP7_75t_L g854 ( .A(n_768), .B(n_784), .Y(n_854) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
OR2x2_ASAP7_75t_L g805 ( .A(n_769), .B(n_784), .Y(n_805) );
INVx1_ASAP7_75t_L g808 ( .A(n_769), .Y(n_808) );
AND2x2_ASAP7_75t_L g856 ( .A(n_769), .B(n_784), .Y(n_856) );
AND2x2_ASAP7_75t_L g927 ( .A(n_769), .B(n_919), .Y(n_927) );
OR2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_775), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_770) );
OAI221xp5_ASAP7_75t_L g822 ( .A1(n_771), .A2(n_773), .B1(n_823), .B2(n_824), .C(n_825), .Y(n_822) );
INVx1_ASAP7_75t_L g944 ( .A(n_771), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_778), .B1(n_779), .B2(n_780), .Y(n_775) );
INVx3_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
OAI322xp33_ASAP7_75t_L g810 ( .A1(n_781), .A2(n_811), .A3(n_820), .B1(n_826), .B2(n_839), .C1(n_841), .C2(n_884), .Y(n_810) );
AOI221xp5_ASAP7_75t_L g904 ( .A1(n_781), .A2(n_905), .B1(n_906), .B2(n_908), .C(n_909), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g918 ( .A1(n_781), .A2(n_919), .B1(n_920), .B2(n_921), .Y(n_918) );
CKINVDCx14_ASAP7_75t_R g781 ( .A(n_782), .Y(n_781) );
CKINVDCx14_ASAP7_75t_R g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_784), .Y(n_796) );
OR2x2_ASAP7_75t_L g873 ( .A(n_784), .B(n_847), .Y(n_873) );
AND2x2_ASAP7_75t_L g881 ( .A(n_784), .B(n_846), .Y(n_881) );
AND2x2_ASAP7_75t_L g919 ( .A(n_784), .B(n_847), .Y(n_919) );
AND2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
O2A1O1Ixp33_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_790), .B(n_793), .C(n_795), .Y(n_787) );
AND2x2_ASAP7_75t_L g818 ( .A(n_789), .B(n_819), .Y(n_818) );
AND2x2_ASAP7_75t_L g878 ( .A(n_789), .B(n_859), .Y(n_878) );
NOR2x1_ASAP7_75t_R g906 ( .A(n_789), .B(n_907), .Y(n_906) );
AND2x2_ASAP7_75t_L g852 ( .A(n_790), .B(n_799), .Y(n_852) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g939 ( .A(n_792), .B(n_799), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_793), .B(n_818), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g895 ( .A(n_793), .B(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
AOI211xp5_ASAP7_75t_L g902 ( .A1(n_794), .A2(n_797), .B(n_844), .C(n_903), .Y(n_902) );
NOR2xp33_ASAP7_75t_L g941 ( .A(n_794), .B(n_804), .Y(n_941) );
OAI211xp5_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_797), .B(n_801), .C(n_806), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_796), .B(n_804), .Y(n_828) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
INVx1_ASAP7_75t_L g871 ( .A(n_799), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_799), .B(n_858), .Y(n_903) );
A2O1A1Ixp33_ASAP7_75t_L g924 ( .A1(n_799), .A2(n_887), .B(n_914), .C(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g809 ( .A(n_800), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
INVx1_ASAP7_75t_L g891 ( .A(n_802), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
INVx1_ASAP7_75t_L g890 ( .A(n_805), .Y(n_890) );
OAI221xp5_ASAP7_75t_L g935 ( .A1(n_805), .A2(n_936), .B1(n_937), .B2(n_938), .C(n_940), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_809), .Y(n_806) );
A2O1A1Ixp33_ASAP7_75t_L g868 ( .A1(n_807), .A2(n_819), .B(n_869), .C(n_872), .Y(n_868) );
INVx2_ASAP7_75t_L g833 ( .A(n_808), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_808), .B(n_840), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_809), .B(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g923 ( .A(n_814), .Y(n_923) );
AND2x2_ASAP7_75t_L g815 ( .A(n_816), .B(n_818), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_817), .B(n_854), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_819), .B(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g932 ( .A(n_819), .Y(n_932) );
AOI22xp5_ASAP7_75t_SL g916 ( .A1(n_820), .A2(n_843), .B1(n_917), .B2(n_935), .Y(n_916) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
O2A1O1Ixp33_ASAP7_75t_L g909 ( .A1(n_821), .A2(n_853), .B(n_910), .C(n_913), .Y(n_909) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_822), .B(n_840), .Y(n_839) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_822), .Y(n_844) );
OAI211xp5_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_829), .B(n_832), .C(n_838), .Y(n_827) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
OR2x2_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
AOI21xp33_ASAP7_75t_L g869 ( .A1(n_836), .A2(n_870), .B(n_871), .Y(n_869) );
INVx1_ASAP7_75t_L g899 ( .A(n_837), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_843), .B(n_845), .Y(n_842) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_SL g896 ( .A(n_845), .Y(n_896) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
A2O1A1Ixp33_ASAP7_75t_L g848 ( .A1(n_849), .A2(n_851), .B(n_853), .C(n_855), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
OAI221xp5_ASAP7_75t_L g885 ( .A1(n_851), .A2(n_886), .B1(n_888), .B2(n_891), .C(n_892), .Y(n_885) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
AOI211xp5_ASAP7_75t_SL g855 ( .A1(n_856), .A2(n_857), .B(n_860), .C(n_863), .Y(n_855) );
INVx1_ASAP7_75t_L g937 ( .A(n_856), .Y(n_937) );
NOR2xp33_ASAP7_75t_L g936 ( .A(n_857), .B(n_920), .Y(n_936) );
INVx1_ASAP7_75t_L g925 ( .A(n_861), .Y(n_925) );
INVx1_ASAP7_75t_L g915 ( .A(n_862), .Y(n_915) );
INVx1_ASAP7_75t_L g929 ( .A(n_864), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_865), .B(n_899), .Y(n_898) );
OAI21xp5_ASAP7_75t_SL g913 ( .A1(n_865), .A2(n_914), .B(n_915), .Y(n_913) );
INVx1_ASAP7_75t_L g920 ( .A(n_866), .Y(n_920) );
NAND3xp33_ASAP7_75t_L g867 ( .A(n_868), .B(n_874), .C(n_875), .Y(n_867) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g905 ( .A(n_874), .Y(n_905) );
OAI22xp33_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_879), .B1(n_881), .B2(n_882), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_893), .B(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
NAND3xp33_ASAP7_75t_L g900 ( .A(n_901), .B(n_904), .C(n_916), .Y(n_900) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
NAND5xp2_ASAP7_75t_L g917 ( .A(n_918), .B(n_924), .C(n_926), .D(n_928), .E(n_930), .Y(n_917) );
NOR2xp33_ASAP7_75t_L g921 ( .A(n_922), .B(n_923), .Y(n_921) );
INVxp67_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g942 ( .A(n_943), .Y(n_942) );
HB1xp67_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVxp67_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
HB1xp67_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
XNOR2x1_ASAP7_75t_L g949 ( .A(n_950), .B(n_974), .Y(n_949) );
NAND2x1_ASAP7_75t_L g950 ( .A(n_951), .B(n_957), .Y(n_950) );
AND4x1_ASAP7_75t_L g951 ( .A(n_952), .B(n_954), .C(n_955), .D(n_956), .Y(n_951) );
INVx2_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
OAI21xp5_ASAP7_75t_L g960 ( .A1(n_961), .A2(n_962), .B(n_963), .Y(n_960) );
INVx1_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
OAI21xp5_ASAP7_75t_SL g964 ( .A1(n_965), .A2(n_966), .B(n_967), .Y(n_964) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
CKINVDCx16_ASAP7_75t_R g975 ( .A(n_976), .Y(n_975) );
BUFx3_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
NAND4xp75_ASAP7_75t_L g984 ( .A(n_985), .B(n_989), .C(n_992), .D(n_995), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_986), .B(n_988), .Y(n_985) );
AND2x2_ASAP7_75t_L g989 ( .A(n_990), .B(n_991), .Y(n_989) );
AND2x2_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .Y(n_992) );
BUFx2_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
endmodule