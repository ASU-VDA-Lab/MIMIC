module fake_jpeg_9109_n_251 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_21),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_2),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_2),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_17),
.C(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_20),
.B1(n_34),
.B2(n_30),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_53),
.B1(n_25),
.B2(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_58),
.Y(n_81)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_57),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_34),
.B1(n_30),
.B2(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_18),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_27),
.B(n_33),
.Y(n_59)
);

OAI32xp33_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_25),
.A3(n_19),
.B1(n_28),
.B2(n_23),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_33),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_63),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_26),
.C(n_30),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_3),
.C(n_6),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_24),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_51),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_69),
.B(n_87),
.Y(n_109)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_70),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_90),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_34),
.B1(n_26),
.B2(n_31),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_94),
.B1(n_95),
.B2(n_99),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_44),
.B1(n_32),
.B2(n_31),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_77),
.B(n_8),
.CI(n_9),
.CON(n_104),
.SN(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_61),
.B1(n_67),
.B2(n_49),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_29),
.B1(n_28),
.B2(n_23),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_51),
.B1(n_62),
.B2(n_44),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_3),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_32),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_16),
.C(n_98),
.Y(n_120)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_101),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_61),
.A2(n_32),
.B1(n_4),
.B2(n_5),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_61),
.A2(n_32),
.B1(n_4),
.B2(n_5),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_60),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_52),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_100),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_46),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_104),
.B(n_106),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_105),
.A2(n_117),
.B1(n_101),
.B2(n_92),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_80),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_114),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_60),
.Y(n_114)
);

AOI32xp33_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_11),
.A3(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_124),
.B(n_109),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_96),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_119),
.B(n_125),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_77),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_81),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_16),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_79),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_87),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_126),
.B(n_122),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_127),
.B(n_88),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_68),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_132),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_131),
.B(n_137),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_68),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_81),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_146),
.B(n_153),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_108),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_143),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_100),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_82),
.B1(n_86),
.B2(n_74),
.Y(n_138)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

AO22x1_ASAP7_75t_SL g140 ( 
.A1(n_107),
.A2(n_74),
.B1(n_83),
.B2(n_88),
.Y(n_140)
);

AO22x1_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_116),
.B1(n_118),
.B2(n_127),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_129),
.B(n_142),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_110),
.B(n_88),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_145),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_115),
.B(n_104),
.C(n_73),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_107),
.A2(n_74),
.B1(n_85),
.B2(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_149),
.B1(n_111),
.B2(n_102),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_104),
.A2(n_118),
.B1(n_121),
.B2(n_117),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_89),
.B(n_121),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_154),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_156),
.A2(n_152),
.B1(n_160),
.B2(n_155),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_122),
.B(n_102),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_111),
.Y(n_166)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_161),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_168),
.A2(n_170),
.B1(n_177),
.B2(n_165),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_169),
.B(n_171),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_102),
.B(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_139),
.B(n_138),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_174),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_136),
.Y(n_175)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_133),
.Y(n_176)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_141),
.A2(n_140),
.B(n_147),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_168),
.A2(n_146),
.B1(n_150),
.B2(n_143),
.Y(n_181)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_130),
.Y(n_182)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_176),
.C(n_159),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_187),
.C(n_173),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_131),
.Y(n_185)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_186),
.A2(n_192),
.B(n_164),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_159),
.C(n_170),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_155),
.B1(n_166),
.B2(n_177),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_163),
.B1(n_157),
.B2(n_166),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_158),
.B(n_171),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_191),
.Y(n_203)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_158),
.B(n_164),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_167),
.Y(n_204)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_156),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_178),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_208),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_194),
.C(n_196),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_174),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_209),
.C(n_195),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

NOR2xp67_ASAP7_75t_SL g206 ( 
.A(n_183),
.B(n_156),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_186),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_169),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_169),
.B(n_179),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_188),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_181),
.B1(n_179),
.B2(n_202),
.Y(n_212)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_219),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_200),
.C(n_209),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_215),
.C(n_220),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_182),
.C(n_195),
.Y(n_215)
);

XOR2x2_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_197),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_221),
.A2(n_210),
.B(n_207),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_207),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_224),
.A2(n_217),
.B(n_216),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_203),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_226),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_185),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_221),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_228),
.A2(n_230),
.B1(n_231),
.B2(n_205),
.Y(n_237)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

INVxp33_ASAP7_75t_SL g233 ( 
.A(n_224),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_236),
.B(n_227),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_214),
.C(n_213),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_237),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_229),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_232),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_241),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_231),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_211),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_243),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_235),
.B(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_244),
.Y(n_247)
);

AOI321xp33_ASAP7_75t_L g248 ( 
.A1(n_246),
.A2(n_180),
.A3(n_194),
.B1(n_240),
.B2(n_245),
.C(n_233),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_248),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_249),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_247),
.Y(n_251)
);


endmodule