module real_jpeg_28934_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_337, n_11, n_14, n_336, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_336;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx11_ASAP7_75t_L g89 ( 
.A(n_0),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_0),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_L g158 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_1),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_159),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_159),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_1),
.A2(n_48),
.B1(n_50),
.B2(n_159),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_2),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_96),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_96),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_2),
.A2(n_48),
.B1(n_50),
.B2(n_96),
.Y(n_240)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_5),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_SL g173 ( 
.A1(n_5),
.A2(n_28),
.B(n_32),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_5),
.B(n_30),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_5),
.A2(n_54),
.B(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_5),
.B(n_54),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_5),
.B(n_68),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_5),
.A2(n_86),
.B1(n_89),
.B2(n_252),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_5),
.A2(n_31),
.B(n_269),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_6),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_170),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_6),
.A2(n_54),
.B1(n_55),
.B2(n_170),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_6),
.A2(n_48),
.B1(n_50),
.B2(n_170),
.Y(n_252)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_8),
.A2(n_43),
.B1(n_54),
.B2(n_55),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_8),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_9),
.A2(n_36),
.B1(n_54),
.B2(n_55),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_36),
.B1(n_48),
.B2(n_50),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_10),
.A2(n_45),
.B1(n_54),
.B2(n_55),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_45),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_10),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_11),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_47)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

OAI32xp33_ASAP7_75t_L g228 ( 
.A1(n_11),
.A2(n_50),
.A3(n_54),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_12),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_12),
.A2(n_26),
.B1(n_54),
.B2(n_55),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_12),
.A2(n_26),
.B1(n_48),
.B2(n_50),
.Y(n_121)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_14),
.A2(n_31),
.B(n_62),
.C(n_65),
.Y(n_61)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_14),
.A2(n_54),
.B1(n_55),
.B2(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_15),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_98),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g165 ( 
.A1(n_15),
.A2(n_54),
.B1(n_55),
.B2(n_98),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_15),
.A2(n_48),
.B1(n_50),
.B2(n_98),
.Y(n_184)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_16),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_17),
.A2(n_24),
.B1(n_25),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_17),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_17),
.A2(n_31),
.B1(n_32),
.B2(n_128),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_17),
.A2(n_48),
.B1(n_50),
.B2(n_128),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_17),
.A2(n_54),
.B1(n_55),
.B2(n_128),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_78),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_76),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_21),
.B(n_37),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_23),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_28),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_25),
.A2(n_34),
.B(n_168),
.C(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_30),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_27),
.A2(n_30),
.B1(n_95),
.B2(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_27),
.A2(n_30),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_27),
.A2(n_30),
.B1(n_127),
.B2(n_199),
.Y(n_213)
);

AO22x1_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_63),
.Y(n_62)
);

OAI32xp33_ASAP7_75t_L g277 ( 
.A1(n_31),
.A2(n_55),
.A3(n_63),
.B1(n_270),
.B2(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_32),
.B(n_168),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_69),
.C(n_71),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_38),
.A2(n_39),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_58),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_40),
.B(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_42),
.A2(n_73),
.B1(n_75),
.B2(n_97),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_46),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_46),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_46),
.A2(n_58),
.B1(n_137),
.B2(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_52),
.B(n_57),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_47),
.A2(n_52),
.B1(n_57),
.B2(n_107),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_47),
.A2(n_52),
.B1(n_104),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_47),
.A2(n_52),
.B1(n_123),
.B2(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_47),
.A2(n_52),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_47),
.A2(n_52),
.B1(n_226),
.B2(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_47),
.B(n_168),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_47),
.A2(n_52),
.B1(n_164),
.B2(n_295),
.Y(n_294)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_48),
.B(n_51),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_48),
.B(n_257),
.Y(n_256)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_54),
.B(n_279),
.Y(n_278)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_58),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_59),
.A2(n_60),
.B1(n_68),
.B2(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_60),
.A2(n_68),
.B1(n_113),
.B2(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_60),
.A2(n_68),
.B1(n_158),
.B2(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_60),
.A2(n_68),
.B1(n_125),
.B2(n_202),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_65),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_61),
.A2(n_65),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_61),
.A2(n_65),
.B1(n_157),
.B2(n_160),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_61),
.A2(n_65),
.B1(n_160),
.B2(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_61),
.A2(n_65),
.B1(n_182),
.B2(n_268),
.Y(n_267)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_63),
.Y(n_279)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_67),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_69),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_75),
.B1(n_94),
.B2(n_97),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_73),
.A2(n_75),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_326),
.B(n_332),
.Y(n_78)
);

OAI321xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_140),
.A3(n_149),
.B1(n_324),
.B2(n_325),
.C(n_336),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_129),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_81),
.B(n_129),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_110),
.C(n_117),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_82),
.B(n_110),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_99),
.B1(n_100),
.B2(n_109),
.Y(n_82)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_92),
.B2(n_93),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_84),
.A2(n_93),
.B(n_99),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_84),
.A2(n_85),
.B1(n_101),
.B2(n_102),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_90),
.B(n_91),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_90),
.B1(n_91),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_86),
.A2(n_90),
.B1(n_121),
.B2(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_86),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_86),
.A2(n_90),
.B1(n_246),
.B2(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_86),
.A2(n_90),
.B1(n_240),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_87),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_87),
.A2(n_88),
.B1(n_175),
.B2(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_87),
.A2(n_176),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

INVx5_ASAP7_75t_SL g241 ( 
.A(n_88),
.Y(n_241)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_90),
.Y(n_176)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_105),
.A2(n_108),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_105),
.A2(n_108),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_115),
.B(n_116),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_115),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_114),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g129 ( 
.A(n_116),
.B(n_130),
.CI(n_139),
.CON(n_129),
.SN(n_129)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_130),
.C(n_139),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_117),
.A2(n_118),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_124),
.C(n_126),
.Y(n_118)
);

FAx1_ASAP7_75t_L g307 ( 
.A(n_119),
.B(n_124),
.CI(n_126),
.CON(n_307),
.SN(n_307)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_120),
.B(n_122),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_129),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_138),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_132),
.B1(n_144),
.B2(n_147),
.Y(n_143)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_134),
.C(n_137),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_132),
.B(n_147),
.C(n_148),
.Y(n_327)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_141),
.B(n_142),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_148),
.Y(n_142)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

AOI321xp33_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_305),
.A3(n_313),
.B1(n_318),
.B2(n_323),
.C(n_337),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_204),
.C(n_216),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_186),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_152),
.B(n_186),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_171),
.C(n_178),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_153),
.B(n_302),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_166),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_161),
.B2(n_162),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_162),
.C(n_166),
.Y(n_193)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_165),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_168),
.B(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_169),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_171),
.A2(n_178),
.B1(n_179),
.B2(n_303),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_171),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_174),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_177),
.Y(n_192)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.C(n_185),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_180),
.B(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_183),
.B(n_185),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_184),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_194),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_193),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_193),
.C(n_194),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_191),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_203),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_200),
.C(n_203),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_L g319 ( 
.A1(n_205),
.A2(n_320),
.B(n_321),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_206),
.B(n_207),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_215),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_209),
.B(n_210),
.C(n_215),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_211),
.B(n_213),
.C(n_214),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_299),
.B(n_304),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_285),
.B(n_298),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_263),
.B(n_284),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_242),
.B(n_262),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_231),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_221),
.B(n_231),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_227),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_222),
.A2(n_223),
.B1(n_227),
.B2(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_238),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_236),
.C(n_238),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_237),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_239),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_249),
.B(n_261),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_244),
.B(n_248),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_254),
.B(n_260),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_251),
.B(n_253),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_264),
.B(n_265),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_276),
.B1(n_282),
.B2(n_283),
.Y(n_265)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_271),
.B1(n_274),
.B2(n_275),
.Y(n_266)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_271),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_275),
.C(n_283),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_273),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_276),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_280),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_286),
.B(n_287),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_294),
.C(n_296),
.Y(n_300)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_296),
.B2(n_297),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_293),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_294),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_300),
.B(n_301),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_310),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_310),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.C(n_309),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_308),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_307),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_314),
.A2(n_319),
.B(n_322),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_316),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);


endmodule