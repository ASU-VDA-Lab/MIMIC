module fake_netlist_1_8909_n_24 (n_3, n_1, n_2, n_0, n_24);
input n_3;
input n_1;
input n_2;
input n_0;
output n_24;
wire n_20;
wire n_5;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
wire n_6;
wire n_4;
wire n_7;
INVx3_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
NAND2xp5_ASAP7_75t_L g5 ( .A(n_2), .B(n_3), .Y(n_5) );
NAND2xp5_ASAP7_75t_L g6 ( .A(n_2), .B(n_1), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_3), .Y(n_7) );
OR2x2_ASAP7_75t_L g8 ( .A(n_3), .B(n_0), .Y(n_8) );
AOI21xp5_ASAP7_75t_L g9 ( .A1(n_6), .A2(n_0), .B(n_1), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_4), .B(n_0), .Y(n_10) );
NAND2xp5_ASAP7_75t_SL g11 ( .A(n_4), .B(n_0), .Y(n_11) );
AOI21xp5_ASAP7_75t_L g12 ( .A1(n_5), .A2(n_1), .B(n_4), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_10), .B(n_7), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_11), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_13), .B(n_9), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_16), .B(n_13), .Y(n_19) );
NAND3xp33_ASAP7_75t_SL g20 ( .A(n_19), .B(n_8), .C(n_14), .Y(n_20) );
BUFx2_ASAP7_75t_R g21 ( .A(n_18), .Y(n_21) );
AOI22xp33_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_18), .B1(n_17), .B2(n_8), .Y(n_22) );
OAI21xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_15), .B(n_7), .Y(n_23) );
AOI22xp33_ASAP7_75t_R g24 ( .A1(n_23), .A2(n_1), .B1(n_15), .B2(n_22), .Y(n_24) );
endmodule