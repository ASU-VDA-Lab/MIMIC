module fake_netlist_6_1910_n_4815 (n_992, n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_853, n_440, n_587, n_695, n_507, n_968, n_909, n_580, n_762, n_1030, n_881, n_875, n_209, n_367, n_465, n_680, n_741, n_760, n_1008, n_1027, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_828, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_1033, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_933, n_740, n_1038, n_578, n_703, n_1003, n_144, n_365, n_978, n_125, n_168, n_1061, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_820, n_1044, n_951, n_783, n_106, n_725, n_952, n_999, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_994, n_1072, n_677, n_969, n_988, n_805, n_396, n_495, n_1065, n_815, n_350, n_78, n_84, n_585, n_732, n_974, n_568, n_392, n_840, n_442, n_480, n_142, n_874, n_724, n_143, n_382, n_673, n_1020, n_180, n_1009, n_1042, n_62, n_1071, n_628, n_1067, n_883, n_557, n_823, n_349, n_643, n_233, n_617, n_698, n_898, n_1032, n_845, n_255, n_807, n_1036, n_739, n_284, n_400, n_140, n_337, n_955, n_865, n_893, n_214, n_925, n_485, n_67, n_15, n_1026, n_443, n_246, n_892, n_768, n_38, n_471, n_289, n_935, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_963, n_727, n_894, n_369, n_597, n_685, n_280, n_287, n_832, n_353, n_610, n_555, n_389, n_814, n_415, n_830, n_65, n_230, n_605, n_461, n_873, n_141, n_383, n_826, n_1024, n_669, n_200, n_447, n_176, n_872, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_1018, n_747, n_852, n_667, n_71, n_74, n_229, n_542, n_847, n_644, n_682, n_851, n_621, n_305, n_1037, n_72, n_721, n_996, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_901, n_111, n_504, n_923, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_837, n_836, n_1015, n_79, n_863, n_375, n_601, n_338, n_522, n_948, n_466, n_704, n_918, n_748, n_506, n_56, n_763, n_1057, n_360, n_945, n_977, n_603, n_1005, n_119, n_991, n_957, n_235, n_536, n_895, n_866, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_971, n_946, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_987, n_641, n_822, n_693, n_1056, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_842, n_611, n_943, n_156, n_491, n_878, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_843, n_989, n_797, n_666, n_1016, n_371, n_795, n_770, n_940, n_567, n_899, n_189, n_738, n_405, n_213, n_538, n_1035, n_294, n_302, n_499, n_380, n_838, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_844, n_448, n_886, n_953, n_20, n_1004, n_1017, n_494, n_539, n_493, n_397, n_155, n_1022, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_930, n_888, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_910, n_37, n_486, n_911, n_381, n_82, n_947, n_27, n_236, n_653, n_887, n_752, n_908, n_112, n_172, n_944, n_713, n_648, n_657, n_1049, n_576, n_1028, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_976, n_490, n_803, n_290, n_220, n_809, n_1043, n_1011, n_118, n_224, n_48, n_926, n_927, n_25, n_93, n_839, n_986, n_80, n_734, n_708, n_196, n_919, n_402, n_352, n_917, n_668, n_478, n_626, n_990, n_574, n_779, n_9, n_800, n_929, n_460, n_107, n_907, n_854, n_6, n_1058, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_870, n_366, n_904, n_777, n_407, n_913, n_450, n_103, n_808, n_867, n_272, n_526, n_921, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_937, n_390, n_473, n_293, n_1054, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_1070, n_232, n_650, n_998, n_16, n_1046, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_924, n_298, n_18, n_492, n_972, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_824, n_962, n_1000, n_279, n_686, n_796, n_1041, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_936, n_184, n_552, n_1062, n_619, n_885, n_216, n_455, n_896, n_83, n_521, n_363, n_572, n_912, n_395, n_813, n_592, n_745, n_654, n_323, n_829, n_606, n_393, n_818, n_984, n_411, n_503, n_716, n_152, n_623, n_1048, n_92, n_884, n_599, n_513, n_855, n_776, n_321, n_645, n_331, n_105, n_916, n_227, n_132, n_868, n_570, n_731, n_859, n_406, n_483, n_735, n_102, n_204, n_482, n_934, n_755, n_931, n_1021, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_958, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_942, n_792, n_880, n_476, n_981, n_714, n_2, n_291, n_219, n_543, n_889, n_357, n_150, n_264, n_263, n_985, n_589, n_860, n_481, n_788, n_819, n_939, n_997, n_821, n_325, n_938, n_1068, n_767, n_804, n_329, n_464, n_600, n_831, n_802, n_964, n_982, n_561, n_33, n_477, n_549, n_980, n_533, n_954, n_408, n_932, n_806, n_864, n_879, n_959, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_979, n_548, n_905, n_94, n_282, n_436, n_833, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_993, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_1064, n_403, n_723, n_253, n_634, n_1051, n_583, n_596, n_123, n_136, n_966, n_546, n_562, n_249, n_201, n_386, n_764, n_1039, n_556, n_159, n_1034, n_1066, n_157, n_162, n_692, n_733, n_754, n_941, n_975, n_1031, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_849, n_970, n_560, n_1014, n_753, n_642, n_995, n_276, n_569, n_441, n_221, n_811, n_882, n_1060, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_973, n_346, n_88, n_3, n_416, n_1053, n_530, n_277, n_520, n_1029, n_418, n_113, n_618, n_1055, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_861, n_674, n_857, n_871, n_967, n_775, n_922, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_1069, n_5, n_453, n_612, n_633, n_665, n_902, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_914, n_759, n_1047, n_1010, n_355, n_426, n_317, n_149, n_1040, n_915, n_632, n_702, n_431, n_90, n_347, n_812, n_24, n_459, n_54, n_1052, n_502, n_328, n_672, n_534, n_488, n_429, n_1006, n_373, n_1012, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_903, n_85, n_99, n_257, n_920, n_730, n_655, n_13, n_706, n_1045, n_786, n_670, n_203, n_286, n_254, n_207, n_834, n_242, n_835, n_928, n_19, n_47, n_690, n_29, n_850, n_75, n_401, n_324, n_743, n_766, n_816, n_335, n_430, n_1002, n_463, n_545, n_489, n_877, n_205, n_604, n_848, n_120, n_251, n_1019, n_301, n_274, n_636, n_825, n_728, n_681, n_1063, n_729, n_110, n_151, n_876, n_774, n_412, n_640, n_81, n_660, n_965, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_983, n_64, n_288, n_427, n_1059, n_479, n_496, n_598, n_422, n_696, n_906, n_688, n_722, n_961, n_862, n_135, n_165, n_351, n_869, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_890, n_637, n_295, n_385, n_701, n_817, n_950, n_629, n_388, n_190, n_858, n_262, n_484, n_613, n_736, n_187, n_897, n_900, n_846, n_501, n_841, n_956, n_960, n_531, n_827, n_1001, n_60, n_361, n_508, n_663, n_856, n_1050, n_379, n_170, n_778, n_1025, n_332, n_891, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_1013, n_1023, n_194, n_664, n_171, n_949, n_678, n_192, n_57, n_169, n_1007, n_51, n_649, n_283, n_4815);

input n_992;
input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_853;
input n_440;
input n_587;
input n_695;
input n_507;
input n_968;
input n_909;
input n_580;
input n_762;
input n_1030;
input n_881;
input n_875;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_1008;
input n_1027;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_828;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_1033;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_933;
input n_740;
input n_1038;
input n_578;
input n_703;
input n_1003;
input n_144;
input n_365;
input n_978;
input n_125;
input n_168;
input n_1061;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_820;
input n_1044;
input n_951;
input n_783;
input n_106;
input n_725;
input n_952;
input n_999;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_994;
input n_1072;
input n_677;
input n_969;
input n_988;
input n_805;
input n_396;
input n_495;
input n_1065;
input n_815;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_974;
input n_568;
input n_392;
input n_840;
input n_442;
input n_480;
input n_142;
input n_874;
input n_724;
input n_143;
input n_382;
input n_673;
input n_1020;
input n_180;
input n_1009;
input n_1042;
input n_62;
input n_1071;
input n_628;
input n_1067;
input n_883;
input n_557;
input n_823;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_898;
input n_1032;
input n_845;
input n_255;
input n_807;
input n_1036;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_955;
input n_865;
input n_893;
input n_214;
input n_925;
input n_485;
input n_67;
input n_15;
input n_1026;
input n_443;
input n_246;
input n_892;
input n_768;
input n_38;
input n_471;
input n_289;
input n_935;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_963;
input n_727;
input n_894;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_832;
input n_353;
input n_610;
input n_555;
input n_389;
input n_814;
input n_415;
input n_830;
input n_65;
input n_230;
input n_605;
input n_461;
input n_873;
input n_141;
input n_383;
input n_826;
input n_1024;
input n_669;
input n_200;
input n_447;
input n_176;
input n_872;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_1018;
input n_747;
input n_852;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_621;
input n_305;
input n_1037;
input n_72;
input n_721;
input n_996;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_901;
input n_111;
input n_504;
input n_923;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_837;
input n_836;
input n_1015;
input n_79;
input n_863;
input n_375;
input n_601;
input n_338;
input n_522;
input n_948;
input n_466;
input n_704;
input n_918;
input n_748;
input n_506;
input n_56;
input n_763;
input n_1057;
input n_360;
input n_945;
input n_977;
input n_603;
input n_1005;
input n_119;
input n_991;
input n_957;
input n_235;
input n_536;
input n_895;
input n_866;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_971;
input n_946;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_987;
input n_641;
input n_822;
input n_693;
input n_1056;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_842;
input n_611;
input n_943;
input n_156;
input n_491;
input n_878;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_843;
input n_989;
input n_797;
input n_666;
input n_1016;
input n_371;
input n_795;
input n_770;
input n_940;
input n_567;
input n_899;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_1035;
input n_294;
input n_302;
input n_499;
input n_380;
input n_838;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_844;
input n_448;
input n_886;
input n_953;
input n_20;
input n_1004;
input n_1017;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_1022;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_930;
input n_888;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_910;
input n_37;
input n_486;
input n_911;
input n_381;
input n_82;
input n_947;
input n_27;
input n_236;
input n_653;
input n_887;
input n_752;
input n_908;
input n_112;
input n_172;
input n_944;
input n_713;
input n_648;
input n_657;
input n_1049;
input n_576;
input n_1028;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_976;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_1043;
input n_1011;
input n_118;
input n_224;
input n_48;
input n_926;
input n_927;
input n_25;
input n_93;
input n_839;
input n_986;
input n_80;
input n_734;
input n_708;
input n_196;
input n_919;
input n_402;
input n_352;
input n_917;
input n_668;
input n_478;
input n_626;
input n_990;
input n_574;
input n_779;
input n_9;
input n_800;
input n_929;
input n_460;
input n_107;
input n_907;
input n_854;
input n_6;
input n_1058;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_870;
input n_366;
input n_904;
input n_777;
input n_407;
input n_913;
input n_450;
input n_103;
input n_808;
input n_867;
input n_272;
input n_526;
input n_921;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_937;
input n_390;
input n_473;
input n_293;
input n_1054;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_1070;
input n_232;
input n_650;
input n_998;
input n_16;
input n_1046;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_924;
input n_298;
input n_18;
input n_492;
input n_972;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_824;
input n_962;
input n_1000;
input n_279;
input n_686;
input n_796;
input n_1041;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_936;
input n_184;
input n_552;
input n_1062;
input n_619;
input n_885;
input n_216;
input n_455;
input n_896;
input n_83;
input n_521;
input n_363;
input n_572;
input n_912;
input n_395;
input n_813;
input n_592;
input n_745;
input n_654;
input n_323;
input n_829;
input n_606;
input n_393;
input n_818;
input n_984;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_1048;
input n_92;
input n_884;
input n_599;
input n_513;
input n_855;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_916;
input n_227;
input n_132;
input n_868;
input n_570;
input n_731;
input n_859;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_934;
input n_755;
input n_931;
input n_1021;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_958;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_942;
input n_792;
input n_880;
input n_476;
input n_981;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_889;
input n_357;
input n_150;
input n_264;
input n_263;
input n_985;
input n_589;
input n_860;
input n_481;
input n_788;
input n_819;
input n_939;
input n_997;
input n_821;
input n_325;
input n_938;
input n_1068;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_831;
input n_802;
input n_964;
input n_982;
input n_561;
input n_33;
input n_477;
input n_549;
input n_980;
input n_533;
input n_954;
input n_408;
input n_932;
input n_806;
input n_864;
input n_879;
input n_959;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_979;
input n_548;
input n_905;
input n_94;
input n_282;
input n_436;
input n_833;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_993;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_1064;
input n_403;
input n_723;
input n_253;
input n_634;
input n_1051;
input n_583;
input n_596;
input n_123;
input n_136;
input n_966;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_1039;
input n_556;
input n_159;
input n_1034;
input n_1066;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_941;
input n_975;
input n_1031;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_849;
input n_970;
input n_560;
input n_1014;
input n_753;
input n_642;
input n_995;
input n_276;
input n_569;
input n_441;
input n_221;
input n_811;
input n_882;
input n_1060;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_973;
input n_346;
input n_88;
input n_3;
input n_416;
input n_1053;
input n_530;
input n_277;
input n_520;
input n_1029;
input n_418;
input n_113;
input n_618;
input n_1055;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_861;
input n_674;
input n_857;
input n_871;
input n_967;
input n_775;
input n_922;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_1069;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_902;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_914;
input n_759;
input n_1047;
input n_1010;
input n_355;
input n_426;
input n_317;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_54;
input n_1052;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_1006;
input n_373;
input n_1012;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_903;
input n_85;
input n_99;
input n_257;
input n_920;
input n_730;
input n_655;
input n_13;
input n_706;
input n_1045;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_834;
input n_242;
input n_835;
input n_928;
input n_19;
input n_47;
input n_690;
input n_29;
input n_850;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_816;
input n_335;
input n_430;
input n_1002;
input n_463;
input n_545;
input n_489;
input n_877;
input n_205;
input n_604;
input n_848;
input n_120;
input n_251;
input n_1019;
input n_301;
input n_274;
input n_636;
input n_825;
input n_728;
input n_681;
input n_1063;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_965;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_983;
input n_64;
input n_288;
input n_427;
input n_1059;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_906;
input n_688;
input n_722;
input n_961;
input n_862;
input n_135;
input n_165;
input n_351;
input n_869;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_890;
input n_637;
input n_295;
input n_385;
input n_701;
input n_817;
input n_950;
input n_629;
input n_388;
input n_190;
input n_858;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_897;
input n_900;
input n_846;
input n_501;
input n_841;
input n_956;
input n_960;
input n_531;
input n_827;
input n_1001;
input n_60;
input n_361;
input n_508;
input n_663;
input n_856;
input n_1050;
input n_379;
input n_170;
input n_778;
input n_1025;
input n_332;
input n_891;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_1013;
input n_1023;
input n_194;
input n_664;
input n_171;
input n_949;
input n_678;
input n_192;
input n_57;
input n_169;
input n_1007;
input n_51;
input n_649;
input n_283;

output n_4815;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_4730;
wire n_4452;
wire n_3766;
wire n_1613;
wire n_4598;
wire n_1458;
wire n_2576;
wire n_1234;
wire n_3254;
wire n_3684;
wire n_4649;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_4670;
wire n_3266;
wire n_1351;
wire n_3574;
wire n_4620;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_4738;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_3783;
wire n_4177;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1581;
wire n_4504;
wire n_3844;
wire n_4388;
wire n_1237;
wire n_2534;
wire n_2353;
wire n_3301;
wire n_3089;
wire n_4395;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4517;
wire n_4168;
wire n_4372;
wire n_2451;
wire n_1738;
wire n_4490;
wire n_2243;
wire n_2324;
wire n_1854;
wire n_1575;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_1151;
wire n_4699;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_4686;
wire n_2051;
wire n_4370;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2405;
wire n_1743;
wire n_4050;
wire n_1160;
wire n_2647;
wire n_2997;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1238;
wire n_4092;
wire n_4645;
wire n_1724;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_4755;
wire n_3619;
wire n_4359;
wire n_4087;
wire n_1700;
wire n_4578;
wire n_1555;
wire n_2211;
wire n_1415;
wire n_4777;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4591;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_4702;
wire n_2291;
wire n_4754;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_2886;
wire n_2974;
wire n_1285;
wire n_1371;
wire n_3946;
wire n_1985;
wire n_4213;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_4474;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_4531;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_2247;
wire n_3106;
wire n_1711;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_4666;
wire n_2470;
wire n_2321;
wire n_4446;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_3345;
wire n_2074;
wire n_4417;
wire n_2447;
wire n_2919;
wire n_4501;
wire n_3678;
wire n_3440;
wire n_4617;
wire n_4733;
wire n_2129;
wire n_2340;
wire n_4764;
wire n_1261;
wire n_4724;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_4555;
wire n_4743;
wire n_2094;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_2356;
wire n_1143;
wire n_1511;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_4696;
wire n_4692;
wire n_1572;
wire n_4308;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_4814;
wire n_1902;
wire n_1842;
wire n_2739;
wire n_2044;
wire n_1954;
wire n_2510;
wire n_1620;
wire n_1541;
wire n_2480;
wire n_1300;
wire n_3023;
wire n_1735;
wire n_3232;
wire n_2791;
wire n_1313;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_3877;
wire n_3316;
wire n_4325;
wire n_4602;
wire n_2212;
wire n_3929;
wire n_3048;
wire n_3063;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_1455;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_4767;
wire n_2703;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_4722;
wire n_4606;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_4187;
wire n_1971;
wire n_1781;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_1471;
wire n_1094;
wire n_3737;
wire n_3624;
wire n_3077;
wire n_3979;
wire n_2873;
wire n_1345;
wire n_3452;
wire n_3655;
wire n_1820;
wire n_4556;
wire n_3107;
wire n_4563;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_4687;
wire n_3948;
wire n_2836;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_4619;
wire n_2378;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_4414;
wire n_1280;
wire n_3765;
wire n_2655;
wire n_4600;
wire n_4125;
wire n_2625;
wire n_1400;
wire n_3296;
wire n_4646;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_1088;
wire n_4262;
wire n_4392;
wire n_1894;
wire n_2996;
wire n_1231;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_4071;
wire n_4255;
wire n_4403;
wire n_4729;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_1967;
wire n_1193;
wire n_3999;
wire n_3928;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_4751;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_4605;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_4549;
wire n_4575;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_3943;
wire n_4320;
wire n_4305;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_4349;
wire n_4102;
wire n_4297;
wire n_2113;
wire n_1641;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_4662;
wire n_1843;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_4227;
wire n_2778;
wire n_2850;
wire n_4314;
wire n_2080;
wire n_1909;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_1441;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_3910;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4415;
wire n_4296;
wire n_2633;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2059;
wire n_4507;
wire n_2198;
wire n_3319;
wire n_3728;
wire n_2669;
wire n_2925;
wire n_4094;
wire n_4499;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_4677;
wire n_3272;
wire n_4765;
wire n_3193;
wire n_2522;
wire n_3949;
wire n_4364;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_4354;
wire n_2616;
wire n_3912;
wire n_4732;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_4393;
wire n_1162;
wire n_1530;
wire n_3798;
wire n_3488;
wire n_2811;
wire n_1543;
wire n_1302;
wire n_1599;
wire n_3732;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_2832;
wire n_4581;
wire n_4226;
wire n_1762;
wire n_4641;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_4377;
wire n_3446;
wire n_4158;
wire n_4366;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_4795;
wire n_3630;
wire n_4698;
wire n_3518;
wire n_4445;
wire n_3824;
wire n_4792;
wire n_4810;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_2692;
wire n_1680;
wire n_3842;
wire n_3248;
wire n_2031;
wire n_4544;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_4477;
wire n_3888;
wire n_4511;
wire n_2908;
wire n_3168;
wire n_4468;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4130;
wire n_4161;
wire n_4337;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_3403;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3092;
wire n_3055;
wire n_3492;
wire n_3895;
wire n_3966;
wire n_4369;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_4454;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_4742;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_4520;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_4502;
wire n_4503;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_3746;
wire n_4375;
wire n_1111;
wire n_2971;
wire n_1713;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4277;
wire n_4526;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1950;
wire n_1726;
wire n_1912;
wire n_1563;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_4441;
wire n_4613;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_4478;
wire n_1167;
wire n_2818;
wire n_1359;
wire n_2428;
wire n_3581;
wire n_4717;
wire n_3794;
wire n_3247;
wire n_3069;
wire n_3921;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_2664;
wire n_2641;
wire n_1664;
wire n_1722;
wire n_4585;
wire n_4731;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_4773;
wire n_3933;
wire n_2749;
wire n_2008;
wire n_3298;
wire n_2192;
wire n_3346;
wire n_2254;
wire n_2345;
wire n_3281;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_4467;
wire n_2311;
wire n_1386;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_1747;
wire n_3691;
wire n_4427;
wire n_3861;
wire n_2624;
wire n_4066;
wire n_4485;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_4681;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4220;
wire n_4523;
wire n_4752;
wire n_1214;
wire n_2347;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_3917;
wire n_1654;
wire n_4371;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_4552;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_4043;
wire n_4673;
wire n_4313;
wire n_4353;
wire n_2916;
wire n_3415;
wire n_4292;
wire n_4607;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_4381;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_3434;
wire n_4510;
wire n_1515;
wire n_4473;
wire n_4356;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_4169;
wire n_4055;
wire n_2377;
wire n_2178;
wire n_3271;
wire n_4362;
wire n_4248;
wire n_2812;
wire n_4518;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_3009;
wire n_1709;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_4361;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_1630;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_4589;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_4367;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_2271;
wire n_3192;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_4560;
wire n_4737;
wire n_4685;
wire n_4394;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_4675;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_2431;
wire n_3073;
wire n_4018;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_2943;
wire n_1294;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_1634;
wire n_2078;
wire n_3252;
wire n_2932;
wire n_3253;
wire n_3337;
wire n_3431;
wire n_1465;
wire n_1767;
wire n_1779;
wire n_3450;
wire n_4002;
wire n_3209;
wire n_2622;
wire n_1858;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_3021;
wire n_1712;
wire n_4603;
wire n_1391;
wire n_4663;
wire n_2750;
wire n_2558;
wire n_2893;
wire n_1523;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_4697;
wire n_2954;
wire n_3477;
wire n_4289;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4288;
wire n_2684;
wire n_2712;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_4653;
wire n_1487;
wire n_4435;
wire n_2691;
wire n_3421;
wire n_2913;
wire n_3614;
wire n_4471;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_4802;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_4728;
wire n_4385;
wire n_1952;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_1932;
wire n_1101;
wire n_2535;
wire n_3442;
wire n_1880;
wire n_3366;
wire n_2631;
wire n_4191;
wire n_4636;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_4701;
wire n_4651;
wire n_1451;
wire n_3941;
wire n_2767;
wire n_3793;
wire n_1839;
wire n_2341;
wire n_4576;
wire n_3727;
wire n_1765;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_1514;
wire n_1863;
wire n_4615;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1139;
wire n_1714;
wire n_3922;
wire n_3179;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_2897;
wire n_2537;
wire n_4389;
wire n_3970;
wire n_4483;
wire n_4345;
wire n_2554;
wire n_4661;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_2747;
wire n_1513;
wire n_3924;
wire n_3171;
wire n_1913;
wire n_4621;
wire n_4216;
wire n_3608;
wire n_4540;
wire n_4664;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_3053;
wire n_1808;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_2339;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_4785;
wire n_3470;
wire n_4683;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_4713;
wire n_4098;
wire n_4021;
wire n_4476;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_4688;
wire n_3166;
wire n_4753;
wire n_2316;
wire n_1771;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_3435;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_4022;
wire n_2239;
wire n_3082;
wire n_1707;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_4775;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_4674;
wire n_2191;
wire n_2717;
wire n_1723;
wire n_4481;
wire n_1246;
wire n_4528;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_4475;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_2335;
wire n_1529;
wire n_2473;
wire n_4443;
wire n_3887;
wire n_4634;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_2667;
wire n_4123;
wire n_1431;
wire n_1615;
wire n_4114;
wire n_3312;
wire n_1474;
wire n_1571;
wire n_3835;
wire n_4587;
wire n_4286;
wire n_3119;
wire n_1809;
wire n_4280;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_4379;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_4718;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_4525;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_4218;
wire n_4440;
wire n_4402;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_2848;
wire n_1849;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_4541;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4551;
wire n_4264;
wire n_4484;
wire n_2857;
wire n_3693;
wire n_4497;
wire n_3788;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_4459;
wire n_1299;
wire n_4545;
wire n_4708;
wire n_2896;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_4627;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_4464;
wire n_2403;
wire n_3342;
wire n_4624;
wire n_2837;
wire n_4175;
wire n_4700;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_4659;
wire n_4771;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3867;
wire n_3341;
wire n_4455;
wire n_4453;
wire n_1073;
wire n_1195;
wire n_3559;
wire n_4514;
wire n_3025;
wire n_2137;
wire n_3191;
wire n_1626;
wire n_4005;
wire n_2482;
wire n_1507;
wire n_3810;
wire n_3546;
wire n_4798;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4564;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_3987;
wire n_1857;
wire n_4806;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_2424;
wire n_2296;
wire n_1604;
wire n_3201;
wire n_3633;
wire n_4487;
wire n_3447;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_1774;
wire n_3103;
wire n_2354;
wire n_1201;
wire n_2682;
wire n_3032;
wire n_1475;
wire n_1398;
wire n_3638;
wire n_4573;
wire n_4592;
wire n_2589;
wire n_4535;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_3393;
wire n_2442;
wire n_1207;
wire n_3627;
wire n_3451;
wire n_3480;
wire n_1368;
wire n_1791;
wire n_1418;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_3087;
wire n_3072;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_4695;
wire n_2545;
wire n_3577;
wire n_3540;
wire n_4401;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_4368;
wire n_1478;
wire n_4796;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_2966;
wire n_2294;
wire n_2581;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_3591;
wire n_3641;
wire n_3777;
wire n_1314;
wire n_2218;
wire n_2788;
wire n_1837;
wire n_4533;
wire n_4756;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_4419;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_1410;
wire n_4746;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1564;
wire n_1736;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_4658;
wire n_2331;
wire n_1372;
wire n_2860;
wire n_2292;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_2416;
wire n_1427;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_3909;
wire n_3944;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2323;
wire n_1220;
wire n_1893;
wire n_2784;
wire n_2301;
wire n_2209;
wire n_3582;
wire n_4665;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_4431;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_4387;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_4654;
wire n_4633;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_3481;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_4584;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_4276;
wire n_2990;
wire n_3847;
wire n_1775;
wire n_1286;
wire n_1773;
wire n_2115;
wire n_4430;
wire n_2410;
wire n_2552;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_1093;
wire n_4428;
wire n_4597;
wire n_1783;
wire n_1533;
wire n_2929;
wire n_3364;
wire n_2780;
wire n_3226;
wire n_3323;
wire n_1597;
wire n_4020;
wire n_4176;
wire n_4489;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_4404;
wire n_1153;
wire n_3407;
wire n_1618;
wire n_1531;
wire n_4618;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4204;
wire n_4261;
wire n_1745;
wire n_4679;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_4496;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_4805;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_4513;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_3646;
wire n_2801;
wire n_2920;
wire n_4015;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_1374;
wire n_2556;
wire n_4706;
wire n_2648;
wire n_4747;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_4570;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_3188;
wire n_1459;
wire n_1892;
wire n_1614;
wire n_3742;
wire n_4410;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4034;
wire n_1617;
wire n_4056;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_4622;
wire n_4721;
wire n_4807;
wire n_3093;
wire n_3175;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_2732;
wire n_4693;
wire n_2928;
wire n_4206;
wire n_4448;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_3284;
wire n_1281;
wire n_1267;
wire n_1881;
wire n_1806;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_2720;
wire n_1520;
wire n_3126;
wire n_2159;
wire n_2289;
wire n_1390;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_3663;
wire n_4132;
wire n_4386;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_3360;
wire n_2087;
wire n_1855;
wire n_3051;
wire n_1636;
wire n_1437;
wire n_4609;
wire n_4438;
wire n_2135;
wire n_3956;
wire n_4707;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4676;
wire n_4001;
wire n_1687;
wire n_2328;
wire n_1439;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_2627;
wire n_4355;
wire n_3234;
wire n_2276;
wire n_4422;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_3016;
wire n_2993;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_4647;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_1129;
wire n_3870;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1995;
wire n_2181;
wire n_1594;
wire n_3751;
wire n_3625;
wire n_2911;
wire n_1869;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_4655;
wire n_1429;
wire n_4632;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_4470;
wire n_3466;
wire n_4801;
wire n_3554;
wire n_1593;
wire n_4546;
wire n_4813;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_4583;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_2942;
wire n_1635;
wire n_4014;
wire n_1079;
wire n_4704;
wire n_4714;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_4357;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_4509;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_2327;
wire n_4374;
wire n_2201;
wire n_3919;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_4668;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4635;
wire n_2984;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_3276;
wire n_2597;
wire n_2375;
wire n_3194;
wire n_3250;
wire n_1934;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_4582;
wire n_1728;
wire n_3973;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_3886;
wire n_2924;
wire n_4761;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_4420;
wire n_4710;
wire n_1510;
wire n_3637;
wire n_4574;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_2598;
wire n_1916;
wire n_1683;
wire n_1270;
wire n_2549;
wire n_4690;
wire n_1187;
wire n_4405;
wire n_4304;
wire n_4234;
wire n_4413;
wire n_1403;
wire n_1669;
wire n_4558;
wire n_1852;
wire n_4488;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_4759;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_2052;
wire n_1847;
wire n_3634;
wire n_2302;
wire n_4211;
wire n_4667;
wire n_4182;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_1397;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_1409;
wire n_4230;
wire n_4656;
wire n_1841;
wire n_4660;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_4637;
wire n_4274;
wire n_2423;
wire n_3277;
wire n_4797;
wire n_3108;
wire n_2548;
wire n_2785;
wire n_1657;
wire n_4189;
wire n_4270;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1108;
wire n_3730;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_4397;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_4155;
wire n_2740;
wire n_4238;
wire n_3011;
wire n_1601;
wire n_1960;
wire n_4808;
wire n_2694;
wire n_2061;
wire n_4611;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_3042;
wire n_1356;
wire n_1589;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_4610;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_4472;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_2716;
wire n_3249;
wire n_1320;
wire n_3657;
wire n_3081;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_4725;
wire n_4590;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_3137;
wire n_3382;
wire n_1535;
wire n_4406;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_4380;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_4398;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_2472;
wire n_3529;
wire n_2171;
wire n_1213;
wire n_1891;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_4614;
wire n_3536;
wire n_4109;
wire n_4192;
wire n_1443;
wire n_2392;
wire n_1272;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_4565;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4195;
wire n_4159;
wire n_4567;
wire n_3784;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_4554;
wire n_3594;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_4586;
wire n_4778;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_2050;
wire n_2373;
wire n_1472;
wire n_4626;
wire n_4595;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4144;
wire n_2964;
wire n_1870;
wire n_4174;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_4734;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3475;
wire n_3501;
wire n_4442;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_4434;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_4680;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_2257;
wire n_3692;
wire n_4515;
wire n_4689;
wire n_4616;
wire n_2017;
wire n_1682;
wire n_4516;
wire n_4258;
wire n_2699;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_3029;
wire n_2200;
wire n_1828;
wire n_4547;
wire n_3597;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_4548;
wire n_4643;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_2376;
wire n_1405;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_3878;
wire n_4601;
wire n_2766;
wire n_2670;
wire n_1332;
wire n_2700;
wire n_4323;
wire n_2346;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_4623;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_4553;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_3439;
wire n_1407;
wire n_3588;
wire n_2768;
wire n_1795;
wire n_4135;
wire n_2871;
wire n_4279;
wire n_2688;
wire n_3858;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_4183;
wire n_1489;
wire n_4321;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_3292;
wire n_1271;
wire n_1496;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_4644;
wire n_4790;
wire n_2258;
wire n_1485;
wire n_1544;
wire n_1640;
wire n_4040;
wire n_4561;
wire n_4461;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4209;
wire n_4111;
wire n_2390;
wire n_4007;
wire n_3712;
wire n_4608;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_4716;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_3381;
wire n_1548;
wire n_3562;
wire n_3044;
wire n_4757;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_3007;
wire n_2809;
wire n_2172;
wire n_3528;
wire n_4682;
wire n_3489;
wire n_4571;
wire n_4343;
wire n_2835;
wire n_4715;
wire n_4530;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_3074;
wire n_1086;
wire n_3102;
wire n_1948;
wire n_4694;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_4672;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_2154;
wire n_2962;
wire n_3377;
wire n_4604;
wire n_2939;
wire n_4782;
wire n_3305;
wire n_1484;
wire n_2992;
wire n_1906;
wire n_1321;
wire n_1241;
wire n_2533;
wire n_3157;
wire n_1672;
wire n_3530;
wire n_4185;
wire n_3221;
wire n_3752;
wire n_3267;
wire n_1758;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_4378;
wire n_4407;
wire n_1914;
wire n_1318;
wire n_1235;
wire n_3457;
wire n_2759;
wire n_1229;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_3762;
wire n_3469;
wire n_3932;
wire n_2266;
wire n_2960;
wire n_3958;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_4519;
wire n_2388;
wire n_3984;
wire n_4774;
wire n_2056;
wire n_4205;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_4358;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_4524;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_4469;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_1931;
wire n_2083;
wire n_1269;
wire n_2834;
wire n_4572;
wire n_3207;
wire n_2668;
wire n_4424;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_4776;
wire n_1941;
wire n_1375;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_4726;
wire n_1794;
wire n_3506;
wire n_1962;
wire n_1236;
wire n_1650;
wire n_2398;
wire n_1559;
wire n_1928;
wire n_1725;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_4736;
wire n_4317;
wire n_4493;
wire n_4723;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_3124;
wire n_1741;
wire n_1325;
wire n_1746;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_3524;
wire n_4315;
wire n_2671;
wire n_2888;
wire n_2761;
wire n_2923;
wire n_2793;
wire n_2715;
wire n_2885;
wire n_1804;
wire n_3711;
wire n_3776;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_4650;
wire n_4788;
wire n_2062;
wire n_4539;
wire n_2041;
wire n_2975;
wire n_4421;
wire n_1477;
wire n_4719;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_4793;
wire n_2874;
wire n_1200;
wire n_4498;
wire n_2070;
wire n_2588;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_1154;
wire n_4492;
wire n_3308;
wire n_1113;
wire n_2833;
wire n_1600;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_4799;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_4423;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_4789;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_4376;
wire n_1800;
wire n_2241;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_4203;
wire n_3808;
wire n_3190;
wire n_1742;
wire n_4505;
wire n_4657;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_4365;
wire n_1826;
wire n_2951;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_4512;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1929;
wire n_2369;
wire n_1378;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_4542;
wire n_3199;
wire n_2931;
wire n_4462;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_1953;
wire n_4450;
wire n_4536;
wire n_4741;
wire n_4543;
wire n_3343;
wire n_3303;
wire n_4157;
wire n_2752;
wire n_4173;
wire n_3135;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_4630;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_4550;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_2140;
wire n_4652;
wire n_3503;
wire n_3160;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_2358;
wire n_1401;
wire n_1255;
wire n_3658;
wire n_1516;
wire n_4534;
wire n_1536;
wire n_3846;
wire n_2163;
wire n_2186;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_1132;
wire n_4748;
wire n_1074;
wire n_1394;
wire n_4439;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_4783;
wire n_3874;
wire n_2814;
wire n_2528;
wire n_1379;
wire n_4639;
wire n_2969;
wire n_2787;
wire n_1097;
wire n_1338;
wire n_2395;
wire n_3027;
wire n_3231;
wire n_1554;
wire n_4083;
wire n_4494;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_4786;
wire n_4295;
wire n_1120;
wire n_1583;
wire n_4480;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_4579;
wire n_2020;
wire n_1643;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_4225;
wire n_4811;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_3432;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_3583;
wire n_2883;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_2385;
wire n_1283;
wire n_4112;
wire n_4009;
wire n_1785;
wire n_1114;
wire n_1147;
wire n_1848;
wire n_3268;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3701;
wire n_3154;
wire n_4027;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_3473;
wire n_4557;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_4432;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_4352;
wire n_4391;
wire n_4416;
wire n_2702;
wire n_3241;
wire n_4593;
wire n_2906;
wire n_1303;
wire n_2769;
wire n_4342;
wire n_4465;
wire n_3622;
wire n_4568;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_4495;
wire n_1173;
wire n_1924;
wire n_1721;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4436;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_2180;
wire n_1689;
wire n_4569;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_4559;
wire n_1347;
wire n_4106;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4373;
wire n_1245;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_4711;
wire n_2952;
wire n_3068;
wire n_3853;
wire n_4740;
wire n_2117;
wire n_2234;
wire n_4631;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_3811;
wire n_4720;
wire n_3494;
wire n_1656;
wire n_1460;
wire n_2112;
wire n_2255;
wire n_1737;
wire n_2430;
wire n_1464;
wire n_3584;
wire n_3486;
wire n_1414;
wire n_4678;
wire n_4086;
wire n_2721;
wire n_2649;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_3836;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_4068;
wire n_2032;
wire n_4625;
wire n_4812;
wire n_4409;
wire n_2744;
wire n_4363;
wire n_4309;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_4521;
wire n_2444;
wire n_2437;
wire n_1215;
wire n_2743;
wire n_3962;
wire n_4629;
wire n_4638;
wire n_1973;
wire n_4766;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_1500;
wire n_1537;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_3404;
wire n_1122;
wire n_1253;
wire n_2242;
wire n_1266;
wire n_3362;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4744;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_4142;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_1584;
wire n_2425;
wire n_3461;
wire n_3408;
wire n_1582;
wire n_3680;
wire n_4265;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_4532;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_4383;
wire n_4491;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_2666;
wire n_4105;
wire n_1851;
wire n_1585;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_4244;
wire n_4486;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_1156;
wire n_1362;
wire n_4259;
wire n_3123;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_4612;
wire n_3038;
wire n_2033;
wire n_3086;
wire n_4104;
wire n_2531;
wire n_1789;
wire n_1770;
wire n_4787;
wire n_3285;
wire n_4208;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_4529;
wire n_3361;
wire n_3596;
wire n_3478;
wire n_4537;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_4346;
wire n_4351;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_4316;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_4779;
wire n_4640;
wire n_3521;
wire n_3233;
wire n_4599;
wire n_2800;
wire n_1710;
wire n_2161;
wire n_3496;
wire n_4437;
wire n_1301;
wire n_2805;
wire n_4769;
wire n_3310;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4390;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_4628;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_4784;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_4396;
wire n_4508;
wire n_1763;
wire n_4594;
wire n_1998;
wire n_3066;
wire n_4727;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_3989;
wire n_2303;
wire n_2478;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_4451;
wire n_1606;
wire n_4332;
wire n_4108;
wire n_1133;
wire n_4460;
wire n_3374;
wire n_1194;
wire n_4429;
wire n_4506;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_4538;
wire n_2640;
wire n_3695;
wire n_4642;
wire n_4051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_4293;
wire n_3552;
wire n_3206;
wire n_1305;
wire n_2578;
wire n_2363;
wire n_4562;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_3383;
wire n_3709;
wire n_4684;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_3187;
wire n_2540;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_4580;
wire n_3330;
wire n_1479;
wire n_4768;
wire n_2217;
wire n_2197;
wire n_1675;
wire n_4758;
wire n_4781;
wire n_2065;
wire n_2879;
wire n_3717;
wire n_4522;
wire n_4148;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_4341;
wire n_1884;
wire n_2040;
wire n_4057;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_1170;
wire n_2221;
wire n_1629;
wire n_4263;
wire n_2055;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_4447;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_1578;
wire n_1861;
wire n_3110;
wire n_3017;
wire n_1632;
wire n_1890;
wire n_3955;
wire n_2477;
wire n_1805;
wire n_1888;
wire n_2280;
wire n_1557;
wire n_3903;
wire n_3945;
wire n_1311;
wire n_1833;
wire n_4780;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_1612;
wire n_2162;
wire n_3908;
wire n_2333;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_4803;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_4463;
wire n_1417;
wire n_2185;
wire n_2086;
wire n_1242;
wire n_2927;
wire n_3673;
wire n_4750;
wire n_3833;
wire n_1836;
wire n_4281;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_4648;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_3333;
wire n_2899;
wire n_3274;
wire n_4129;
wire n_3186;
wire n_1322;
wire n_4457;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_4804;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_4794;
wire n_4500;
wire n_2105;
wire n_3079;
wire n_4360;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1423;
wire n_1935;
wire n_4039;
wire n_4745;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4566;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_4275;
wire n_4482;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_4426;
wire n_2912;
wire n_4703;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_4425;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_4449;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_4762;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_4030;
wire n_3113;
wire n_1240;
wire n_4809;

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_818),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_749),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_353),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_20),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_328),
.Y(n_1077)
);

CKINVDCx14_ASAP7_75t_R g1078 ( 
.A(n_661),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_241),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_126),
.Y(n_1080)
);

BUFx10_ASAP7_75t_L g1081 ( 
.A(n_656),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_666),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_689),
.Y(n_1083)
);

INVx2_ASAP7_75t_SL g1084 ( 
.A(n_62),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_797),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_984),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_934),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_565),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_383),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_614),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_913),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_242),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_916),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_816),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_245),
.Y(n_1095)
);

BUFx10_ASAP7_75t_L g1096 ( 
.A(n_1066),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_240),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_780),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_1052),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_908),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_836),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_300),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_142),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_901),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_502),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_709),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_374),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_54),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_897),
.Y(n_1109)
);

CKINVDCx20_ASAP7_75t_R g1110 ( 
.A(n_964),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_677),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_310),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_557),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_984),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_78),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_843),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_216),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_829),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_28),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_630),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_373),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_403),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_278),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_1071),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_1062),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_297),
.Y(n_1127)
);

BUFx10_ASAP7_75t_L g1128 ( 
.A(n_0),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_643),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_636),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_101),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_309),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_160),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_628),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_461),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_995),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_570),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_391),
.Y(n_1138)
);

INVx1_ASAP7_75t_SL g1139 ( 
.A(n_875),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_297),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_154),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_819),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_227),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_405),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_229),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_758),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_923),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_425),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_413),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_925),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_154),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_398),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_192),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_240),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_844),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_957),
.Y(n_1156)
);

CKINVDCx16_ASAP7_75t_R g1157 ( 
.A(n_116),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_805),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_1039),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_419),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1011),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1005),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_380),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_939),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_930),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_736),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_211),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_851),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_719),
.Y(n_1169)
);

CKINVDCx20_ASAP7_75t_R g1170 ( 
.A(n_827),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_65),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_629),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_483),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_236),
.Y(n_1174)
);

BUFx10_ASAP7_75t_L g1175 ( 
.A(n_267),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_782),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_573),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_927),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_361),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_816),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_348),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_823),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_941),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_535),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1065),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_798),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_330),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_581),
.Y(n_1188)
);

CKINVDCx16_ASAP7_75t_R g1189 ( 
.A(n_588),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_520),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_247),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_918),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_656),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_367),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_895),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_864),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_519),
.Y(n_1197)
);

CKINVDCx20_ASAP7_75t_R g1198 ( 
.A(n_677),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_551),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_903),
.Y(n_1200)
);

INVx1_ASAP7_75t_SL g1201 ( 
.A(n_1025),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_486),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1003),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_461),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_778),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1027),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_857),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_920),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_614),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_348),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_805),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_969),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_456),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_327),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_234),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_578),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_443),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_793),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_413),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_716),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_637),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_765),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_994),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_810),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_884),
.Y(n_1225)
);

BUFx10_ASAP7_75t_L g1226 ( 
.A(n_455),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_980),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1064),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_868),
.Y(n_1229)
);

HB1xp67_ASAP7_75t_L g1230 ( 
.A(n_616),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_428),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_519),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_38),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_822),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_842),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_197),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_769),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_902),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_798),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_670),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_447),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_839),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_494),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_184),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_186),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_170),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_722),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_893),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_570),
.Y(n_1249)
);

CKINVDCx16_ASAP7_75t_R g1250 ( 
.A(n_534),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_649),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_292),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_657),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_43),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_455),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_508),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_364),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_18),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_380),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_837),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_529),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_537),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_579),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_444),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_454),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_176),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_959),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_910),
.Y(n_1268)
);

BUFx10_ASAP7_75t_L g1269 ( 
.A(n_1025),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_99),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_701),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_384),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_837),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_433),
.Y(n_1274)
);

INVxp67_ASAP7_75t_L g1275 ( 
.A(n_533),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_527),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_965),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_946),
.Y(n_1278)
);

CKINVDCx14_ASAP7_75t_R g1279 ( 
.A(n_410),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_869),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_342),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_51),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_808),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_925),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_890),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_378),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_887),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_878),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_734),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_898),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_820),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_64),
.Y(n_1292)
);

INVx2_ASAP7_75t_SL g1293 ( 
.A(n_917),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_793),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_655),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_921),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_752),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_596),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_23),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_144),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_849),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_139),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_881),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_97),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_454),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1063),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_506),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_212),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_595),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_617),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_326),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_612),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_549),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_130),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_667),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_667),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_72),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_905),
.Y(n_1318)
);

BUFx10_ASAP7_75t_L g1319 ( 
.A(n_563),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_232),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_486),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_703),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_675),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_202),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_598),
.Y(n_1325)
);

CKINVDCx16_ASAP7_75t_R g1326 ( 
.A(n_533),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_549),
.Y(n_1327)
);

BUFx10_ASAP7_75t_L g1328 ( 
.A(n_958),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_836),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_838),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_775),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_121),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_870),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_287),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_888),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_992),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1046),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_886),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_777),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_121),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_658),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_702),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_415),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_227),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_871),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_610),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_933),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_942),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_573),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_791),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_548),
.Y(n_1351)
);

BUFx2_ASAP7_75t_R g1352 ( 
.A(n_506),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_219),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_865),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_835),
.Y(n_1355)
);

INVxp67_ASAP7_75t_SL g1356 ( 
.A(n_159),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_699),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_36),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_114),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_69),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_2),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_170),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_391),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_838),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_502),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_0),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_604),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_954),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_15),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_35),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_42),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_474),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_662),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_457),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_631),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_536),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1044),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1001),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_661),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_571),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_382),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_410),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_862),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_314),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_289),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_940),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_663),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_216),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_317),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_546),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_515),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_125),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_810),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_886),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_534),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_751),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_174),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_145),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_119),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_895),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_582),
.Y(n_1401)
);

BUFx5_ASAP7_75t_L g1402 ( 
.A(n_587),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1067),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_293),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_865),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_564),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_163),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_912),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_891),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_937),
.Y(n_1410)
);

BUFx10_ASAP7_75t_L g1411 ( 
.A(n_503),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_927),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_971),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_83),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_914),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_777),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_114),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_911),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_128),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_772),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_358),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_176),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_965),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_472),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_936),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_107),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_546),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_618),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_974),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1013),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_341),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_482),
.Y(n_1432)
);

INVx2_ASAP7_75t_SL g1433 ( 
.A(n_128),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_234),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_68),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_295),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_741),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_158),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_403),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_912),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_324),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_872),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_786),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_173),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_560),
.Y(n_1445)
);

BUFx6f_ASAP7_75t_L g1446 ( 
.A(n_212),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_390),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_443),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_982),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_58),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_640),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_152),
.Y(n_1452)
);

BUFx2_ASAP7_75t_L g1453 ( 
.A(n_509),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_13),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_134),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_264),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_460),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_802),
.Y(n_1458)
);

CKINVDCx16_ASAP7_75t_R g1459 ( 
.A(n_765),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_346),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_867),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_808),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_719),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_919),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_852),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_977),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_330),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_482),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_977),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_663),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_599),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_780),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_904),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_853),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_846),
.Y(n_1475)
);

CKINVDCx12_ASAP7_75t_R g1476 ( 
.A(n_967),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_126),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_855),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_820),
.Y(n_1479)
);

CKINVDCx16_ASAP7_75t_R g1480 ( 
.A(n_55),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_944),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_527),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_948),
.Y(n_1483)
);

CKINVDCx16_ASAP7_75t_R g1484 ( 
.A(n_1024),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_290),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_196),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_142),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_163),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_840),
.Y(n_1489)
);

BUFx10_ASAP7_75t_L g1490 ( 
.A(n_845),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_253),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_463),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_894),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_856),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_446),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_978),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_817),
.Y(n_1497)
);

CKINVDCx16_ASAP7_75t_R g1498 ( 
.A(n_951),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_877),
.Y(n_1499)
);

INVxp67_ASAP7_75t_L g1500 ( 
.A(n_359),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_270),
.Y(n_1501)
);

BUFx5_ASAP7_75t_L g1502 ( 
.A(n_1050),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_947),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_833),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_161),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_872),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_720),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_896),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_498),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_572),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_985),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_340),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_498),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_148),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_686),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_864),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_441),
.Y(n_1517)
);

BUFx10_ASAP7_75t_L g1518 ( 
.A(n_556),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_476),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_396),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_432),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_852),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_744),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_664),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_335),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_462),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_919),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_913),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_162),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_730),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_876),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_494),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_516),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_904),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_964),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_52),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_92),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_333),
.Y(n_1538)
);

CKINVDCx20_ASAP7_75t_R g1539 ( 
.A(n_595),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_553),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_177),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_448),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_473),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_826),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_358),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_541),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_185),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_950),
.Y(n_1548)
);

INVx1_ASAP7_75t_SL g1549 ( 
.A(n_683),
.Y(n_1549)
);

CKINVDCx20_ASAP7_75t_R g1550 ( 
.A(n_487),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_409),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_522),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_695),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_702),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1042),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_900),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_237),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_394),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_67),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_938),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_860),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_929),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_335),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_188),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_571),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_321),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_300),
.Y(n_1567)
);

INVxp67_ASAP7_75t_SL g1568 ( 
.A(n_876),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_434),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_307),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_440),
.Y(n_1571)
);

INVx1_ASAP7_75t_SL g1572 ( 
.A(n_1001),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_100),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_971),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_368),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_849),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1054),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_603),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_48),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_966),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_505),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_888),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_38),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_998),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_844),
.Y(n_1585)
);

BUFx10_ASAP7_75t_L g1586 ( 
.A(n_310),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_665),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_210),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_959),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_186),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_911),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_232),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_604),
.Y(n_1593)
);

CKINVDCx20_ASAP7_75t_R g1594 ( 
.A(n_13),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_202),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_349),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_935),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_850),
.Y(n_1598)
);

CKINVDCx20_ASAP7_75t_R g1599 ( 
.A(n_1022),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_630),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_572),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_383),
.Y(n_1602)
);

CKINVDCx20_ASAP7_75t_R g1603 ( 
.A(n_708),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_692),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1023),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_643),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_381),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_376),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_968),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_106),
.Y(n_1610)
);

INVx1_ASAP7_75t_SL g1611 ( 
.A(n_932),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_699),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_444),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_963),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_272),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1028),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_428),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_85),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_93),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_897),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_250),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_744),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_205),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_201),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_675),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_857),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_221),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_458),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_230),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_650),
.Y(n_1630)
);

CKINVDCx20_ASAP7_75t_R g1631 ( 
.A(n_821),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_859),
.Y(n_1632)
);

INVx2_ASAP7_75t_SL g1633 ( 
.A(n_664),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_222),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_961),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_809),
.Y(n_1636)
);

BUFx10_ASAP7_75t_L g1637 ( 
.A(n_674),
.Y(n_1637)
);

CKINVDCx16_ASAP7_75t_R g1638 ( 
.A(n_797),
.Y(n_1638)
);

INVx2_ASAP7_75t_SL g1639 ( 
.A(n_1014),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_242),
.Y(n_1640)
);

BUFx10_ASAP7_75t_L g1641 ( 
.A(n_160),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_260),
.Y(n_1642)
);

CKINVDCx20_ASAP7_75t_R g1643 ( 
.A(n_531),
.Y(n_1643)
);

CKINVDCx20_ASAP7_75t_R g1644 ( 
.A(n_552),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_543),
.Y(n_1645)
);

CKINVDCx20_ASAP7_75t_R g1646 ( 
.A(n_928),
.Y(n_1646)
);

CKINVDCx20_ASAP7_75t_R g1647 ( 
.A(n_874),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_943),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_401),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_991),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_869),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_430),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_563),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_204),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_878),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_689),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1057),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_818),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_811),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_246),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_253),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_465),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_505),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_949),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_298),
.Y(n_1665)
);

CKINVDCx20_ASAP7_75t_R g1666 ( 
.A(n_809),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_826),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_962),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_825),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_557),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_794),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_824),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_564),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_439),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_425),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_205),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_511),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_8),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_605),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_522),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_628),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_866),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_129),
.Y(n_1683)
);

CKINVDCx20_ASAP7_75t_R g1684 ( 
.A(n_774),
.Y(n_1684)
);

BUFx3_ASAP7_75t_L g1685 ( 
.A(n_636),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_887),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_423),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_626),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_92),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_247),
.Y(n_1690)
);

CKINVDCx14_ASAP7_75t_R g1691 ( 
.A(n_1021),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_306),
.Y(n_1692)
);

BUFx10_ASAP7_75t_L g1693 ( 
.A(n_159),
.Y(n_1693)
);

CKINVDCx20_ASAP7_75t_R g1694 ( 
.A(n_196),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_764),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_634),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_681),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_779),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_651),
.Y(n_1699)
);

INVx1_ASAP7_75t_SL g1700 ( 
.A(n_262),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_69),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_926),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_464),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_558),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_594),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_576),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_499),
.Y(n_1707)
);

CKINVDCx16_ASAP7_75t_R g1708 ( 
.A(n_1003),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_956),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_562),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_386),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_292),
.Y(n_1712)
);

CKINVDCx20_ASAP7_75t_R g1713 ( 
.A(n_713),
.Y(n_1713)
);

BUFx10_ASAP7_75t_L g1714 ( 
.A(n_357),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_331),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_238),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_997),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_882),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_263),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1056),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_470),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1017),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_736),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_998),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_885),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_989),
.Y(n_1726)
);

CKINVDCx20_ASAP7_75t_R g1727 ( 
.A(n_46),
.Y(n_1727)
);

BUFx3_ASAP7_75t_L g1728 ( 
.A(n_1041),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_453),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_225),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_91),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_985),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_655),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_285),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1014),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_700),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_867),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_213),
.Y(n_1738)
);

CKINVDCx16_ASAP7_75t_R g1739 ( 
.A(n_324),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_239),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_999),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_265),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_858),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_182),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_879),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_415),
.Y(n_1746)
);

CKINVDCx20_ASAP7_75t_R g1747 ( 
.A(n_396),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_795),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_945),
.Y(n_1749)
);

BUFx3_ASAP7_75t_L g1750 ( 
.A(n_331),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_513),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_850),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_378),
.Y(n_1753)
);

CKINVDCx16_ASAP7_75t_R g1754 ( 
.A(n_278),
.Y(n_1754)
);

BUFx3_ASAP7_75t_L g1755 ( 
.A(n_841),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_907),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_674),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_994),
.Y(n_1758)
);

BUFx3_ASAP7_75t_L g1759 ( 
.A(n_366),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_730),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_624),
.Y(n_1761)
);

INVx2_ASAP7_75t_SL g1762 ( 
.A(n_909),
.Y(n_1762)
);

INVx2_ASAP7_75t_SL g1763 ( 
.A(n_583),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_62),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_123),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_394),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_922),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_704),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_565),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_880),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_83),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_540),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_828),
.Y(n_1773)
);

CKINVDCx20_ASAP7_75t_R g1774 ( 
.A(n_917),
.Y(n_1774)
);

INVx2_ASAP7_75t_SL g1775 ( 
.A(n_6),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_620),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_187),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_21),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_10),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_566),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_579),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_830),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_847),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_464),
.Y(n_1784)
);

INVxp67_ASAP7_75t_SL g1785 ( 
.A(n_715),
.Y(n_1785)
);

INVx2_ASAP7_75t_SL g1786 ( 
.A(n_963),
.Y(n_1786)
);

CKINVDCx20_ASAP7_75t_R g1787 ( 
.A(n_693),
.Y(n_1787)
);

BUFx6f_ASAP7_75t_L g1788 ( 
.A(n_831),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_993),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_569),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_832),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_615),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_757),
.Y(n_1793)
);

CKINVDCx16_ASAP7_75t_R g1794 ( 
.A(n_899),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_824),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_955),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_41),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_993),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_108),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_853),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_883),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_860),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_308),
.Y(n_1803)
);

BUFx3_ASAP7_75t_L g1804 ( 
.A(n_848),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_537),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_400),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_275),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_463),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_766),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_1011),
.Y(n_1810)
);

CKINVDCx20_ASAP7_75t_R g1811 ( 
.A(n_442),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_523),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_181),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1033),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_758),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_901),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_791),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_940),
.Y(n_1818)
);

INVx1_ASAP7_75t_SL g1819 ( 
.A(n_787),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_58),
.Y(n_1820)
);

CKINVDCx14_ASAP7_75t_R g1821 ( 
.A(n_265),
.Y(n_1821)
);

INVx1_ASAP7_75t_SL g1822 ( 
.A(n_72),
.Y(n_1822)
);

INVx2_ASAP7_75t_SL g1823 ( 
.A(n_117),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_283),
.Y(n_1824)
);

CKINVDCx20_ASAP7_75t_R g1825 ( 
.A(n_952),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_392),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_779),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_67),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_756),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_376),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_712),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_287),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_109),
.Y(n_1833)
);

BUFx6f_ASAP7_75t_L g1834 ( 
.A(n_286),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_720),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_559),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_757),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_617),
.Y(n_1838)
);

BUFx2_ASAP7_75t_L g1839 ( 
.A(n_518),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_514),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_727),
.Y(n_1841)
);

CKINVDCx20_ASAP7_75t_R g1842 ( 
.A(n_1028),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_550),
.Y(n_1843)
);

HB1xp67_ASAP7_75t_L g1844 ( 
.A(n_889),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_282),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_304),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_594),
.Y(n_1847)
);

CKINVDCx20_ASAP7_75t_R g1848 ( 
.A(n_755),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_327),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_949),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_447),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_907),
.Y(n_1852)
);

BUFx3_ASAP7_75t_L g1853 ( 
.A(n_577),
.Y(n_1853)
);

BUFx3_ASAP7_75t_L g1854 ( 
.A(n_210),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_735),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_931),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_529),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_108),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_892),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_510),
.Y(n_1860)
);

BUFx10_ASAP7_75t_L g1861 ( 
.A(n_924),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_359),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_762),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_9),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_560),
.Y(n_1865)
);

BUFx3_ASAP7_75t_L g1866 ( 
.A(n_937),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_708),
.Y(n_1867)
);

BUFx6f_ASAP7_75t_L g1868 ( 
.A(n_155),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_183),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_475),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_236),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_416),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_63),
.Y(n_1873)
);

INVx1_ASAP7_75t_SL g1874 ( 
.A(n_395),
.Y(n_1874)
);

CKINVDCx20_ASAP7_75t_R g1875 ( 
.A(n_446),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_861),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_148),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_421),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_1020),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_282),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_492),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_194),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_485),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1047),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_642),
.Y(n_1885)
);

INVx2_ASAP7_75t_SL g1886 ( 
.A(n_942),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_87),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_588),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_344),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_741),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_559),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_495),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_513),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_11),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_133),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_367),
.Y(n_1896)
);

INVx1_ASAP7_75t_SL g1897 ( 
.A(n_147),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_641),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_266),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_873),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_321),
.Y(n_1901)
);

BUFx5_ASAP7_75t_L g1902 ( 
.A(n_329),
.Y(n_1902)
);

CKINVDCx20_ASAP7_75t_R g1903 ( 
.A(n_197),
.Y(n_1903)
);

CKINVDCx20_ASAP7_75t_R g1904 ( 
.A(n_440),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_373),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_686),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_155),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_915),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_906),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_854),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1037),
.Y(n_1911)
);

BUFx2_ASAP7_75t_L g1912 ( 
.A(n_672),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_39),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_960),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_504),
.Y(n_1915)
);

BUFx3_ASAP7_75t_L g1916 ( 
.A(n_900),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_863),
.Y(n_1917)
);

BUFx2_ASAP7_75t_L g1918 ( 
.A(n_497),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_788),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_866),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_903),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_953),
.Y(n_1922)
);

INVx1_ASAP7_75t_SL g1923 ( 
.A(n_397),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_10),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_319),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_996),
.Y(n_1926)
);

BUFx6f_ASAP7_75t_L g1927 ( 
.A(n_181),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_834),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_1049),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_445),
.Y(n_1930)
);

CKINVDCx12_ASAP7_75t_R g1931 ( 
.A(n_27),
.Y(n_1931)
);

BUFx5_ASAP7_75t_L g1932 ( 
.A(n_540),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_716),
.Y(n_1933)
);

CKINVDCx20_ASAP7_75t_R g1934 ( 
.A(n_1078),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_1099),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1402),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1402),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1402),
.Y(n_1938)
);

INVxp67_ASAP7_75t_SL g1939 ( 
.A(n_1728),
.Y(n_1939)
);

INVxp67_ASAP7_75t_SL g1940 ( 
.A(n_1728),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1402),
.Y(n_1941)
);

INVxp33_ASAP7_75t_L g1942 ( 
.A(n_1162),
.Y(n_1942)
);

INVxp67_ASAP7_75t_SL g1943 ( 
.A(n_1230),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1402),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1402),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1125),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1402),
.Y(n_1947)
);

CKINVDCx20_ASAP7_75t_R g1948 ( 
.A(n_1078),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1902),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1932),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1902),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1159),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_1306),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1902),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1902),
.Y(n_1955)
);

INVx1_ASAP7_75t_SL g1956 ( 
.A(n_1369),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1902),
.Y(n_1957)
);

INVxp33_ASAP7_75t_SL g1958 ( 
.A(n_1253),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1902),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1902),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1932),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1932),
.Y(n_1962)
);

CKINVDCx16_ASAP7_75t_R g1963 ( 
.A(n_1157),
.Y(n_1963)
);

CKINVDCx20_ASAP7_75t_R g1964 ( 
.A(n_1279),
.Y(n_1964)
);

BUFx3_ASAP7_75t_L g1965 ( 
.A(n_1096),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1476),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1337),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1932),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1932),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1932),
.Y(n_1970)
);

CKINVDCx16_ASAP7_75t_R g1971 ( 
.A(n_1189),
.Y(n_1971)
);

BUFx2_ASAP7_75t_SL g1972 ( 
.A(n_1096),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1932),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1403),
.Y(n_1974)
);

CKINVDCx20_ASAP7_75t_R g1975 ( 
.A(n_1279),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1927),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1104),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1577),
.Y(n_1978)
);

INVxp67_ASAP7_75t_SL g1979 ( 
.A(n_1355),
.Y(n_1979)
);

BUFx2_ASAP7_75t_SL g1980 ( 
.A(n_1096),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1104),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1105),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1105),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1181),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1181),
.Y(n_1985)
);

CKINVDCx20_ASAP7_75t_R g1986 ( 
.A(n_1691),
.Y(n_1986)
);

INVxp67_ASAP7_75t_SL g1987 ( 
.A(n_1508),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1196),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1196),
.Y(n_1989)
);

INVx3_ASAP7_75t_L g1990 ( 
.A(n_1094),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1094),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1206),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1206),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1212),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1657),
.Y(n_1995)
);

INVxp67_ASAP7_75t_L g1996 ( 
.A(n_1382),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1212),
.Y(n_1997)
);

INVxp67_ASAP7_75t_SL g1998 ( 
.A(n_1840),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1214),
.Y(n_1999)
);

INVxp67_ASAP7_75t_L g2000 ( 
.A(n_1453),
.Y(n_2000)
);

BUFx3_ASAP7_75t_L g2001 ( 
.A(n_1214),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1931),
.Y(n_2002)
);

INVxp33_ASAP7_75t_L g2003 ( 
.A(n_1844),
.Y(n_2003)
);

INVxp33_ASAP7_75t_L g2004 ( 
.A(n_1483),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1216),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1216),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1258),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1927),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1258),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1270),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1270),
.Y(n_2011)
);

CKINVDCx16_ASAP7_75t_R g2012 ( 
.A(n_1250),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1578),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1578),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1720),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1596),
.Y(n_2016)
);

HB1xp67_ASAP7_75t_L g2017 ( 
.A(n_1326),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1596),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1685),
.Y(n_2019)
);

INVxp67_ASAP7_75t_SL g2020 ( 
.A(n_1094),
.Y(n_2020)
);

CKINVDCx5p33_ASAP7_75t_R g2021 ( 
.A(n_1884),
.Y(n_2021)
);

CKINVDCx20_ASAP7_75t_R g2022 ( 
.A(n_1691),
.Y(n_2022)
);

CKINVDCx20_ASAP7_75t_R g2023 ( 
.A(n_1821),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1685),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1750),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1750),
.Y(n_2026)
);

CKINVDCx16_ASAP7_75t_R g2027 ( 
.A(n_1459),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1755),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1755),
.Y(n_2029)
);

INVxp67_ASAP7_75t_SL g2030 ( 
.A(n_1094),
.Y(n_2030)
);

INVxp33_ASAP7_75t_SL g2031 ( 
.A(n_1556),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1759),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1927),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1927),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1108),
.Y(n_2035)
);

CKINVDCx5p33_ASAP7_75t_R g2036 ( 
.A(n_1929),
.Y(n_2036)
);

CKINVDCx5p33_ASAP7_75t_R g2037 ( 
.A(n_1480),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1759),
.Y(n_2038)
);

INVxp67_ASAP7_75t_SL g2039 ( 
.A(n_1108),
.Y(n_2039)
);

INVxp67_ASAP7_75t_L g2040 ( 
.A(n_1634),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1804),
.Y(n_2041)
);

CKINVDCx16_ASAP7_75t_R g2042 ( 
.A(n_1484),
.Y(n_2042)
);

INVxp33_ASAP7_75t_SL g2043 ( 
.A(n_1839),
.Y(n_2043)
);

BUFx3_ASAP7_75t_L g2044 ( 
.A(n_1804),
.Y(n_2044)
);

INVxp67_ASAP7_75t_SL g2045 ( 
.A(n_1108),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_1498),
.Y(n_2046)
);

CKINVDCx20_ASAP7_75t_R g2047 ( 
.A(n_1821),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1853),
.Y(n_2048)
);

CKINVDCx16_ASAP7_75t_R g2049 ( 
.A(n_1638),
.Y(n_2049)
);

INVxp33_ASAP7_75t_SL g2050 ( 
.A(n_1912),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1853),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1854),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_1708),
.Y(n_2053)
);

INVxp33_ASAP7_75t_L g2054 ( 
.A(n_1918),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1854),
.Y(n_2055)
);

BUFx10_ASAP7_75t_L g2056 ( 
.A(n_1073),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_1739),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1108),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1866),
.Y(n_2059)
);

HB1xp67_ASAP7_75t_L g2060 ( 
.A(n_1754),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1866),
.Y(n_2061)
);

CKINVDCx16_ASAP7_75t_R g2062 ( 
.A(n_1794),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1916),
.Y(n_2063)
);

INVxp67_ASAP7_75t_L g2064 ( 
.A(n_1281),
.Y(n_2064)
);

CKINVDCx20_ASAP7_75t_R g2065 ( 
.A(n_1083),
.Y(n_2065)
);

INVxp67_ASAP7_75t_SL g2066 ( 
.A(n_1148),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1916),
.Y(n_2067)
);

INVxp33_ASAP7_75t_SL g2068 ( 
.A(n_1074),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_1077),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1148),
.Y(n_2070)
);

INVxp33_ASAP7_75t_L g2071 ( 
.A(n_1075),
.Y(n_2071)
);

BUFx3_ASAP7_75t_L g2072 ( 
.A(n_1081),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1148),
.Y(n_2073)
);

NOR2xp33_ASAP7_75t_L g2074 ( 
.A(n_1126),
.B(n_2),
.Y(n_2074)
);

CKINVDCx16_ASAP7_75t_R g2075 ( 
.A(n_1081),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1148),
.Y(n_2076)
);

INVx1_ASAP7_75t_SL g2077 ( 
.A(n_1076),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1173),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1173),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1173),
.Y(n_2080)
);

CKINVDCx5p33_ASAP7_75t_R g2081 ( 
.A(n_1919),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1173),
.Y(n_2082)
);

INVxp67_ASAP7_75t_SL g2083 ( 
.A(n_1274),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1274),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_1274),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1274),
.Y(n_2086)
);

BUFx2_ASAP7_75t_L g2087 ( 
.A(n_1082),
.Y(n_2087)
);

CKINVDCx20_ASAP7_75t_R g2088 ( 
.A(n_1083),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1289),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1289),
.Y(n_2090)
);

CKINVDCx5p33_ASAP7_75t_R g2091 ( 
.A(n_1924),
.Y(n_2091)
);

HB1xp67_ASAP7_75t_L g2092 ( 
.A(n_1925),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1289),
.Y(n_2093)
);

CKINVDCx20_ASAP7_75t_R g2094 ( 
.A(n_1110),
.Y(n_2094)
);

CKINVDCx16_ASAP7_75t_R g2095 ( 
.A(n_1081),
.Y(n_2095)
);

INVxp67_ASAP7_75t_L g2096 ( 
.A(n_1128),
.Y(n_2096)
);

CKINVDCx20_ASAP7_75t_R g2097 ( 
.A(n_1110),
.Y(n_2097)
);

INVxp67_ASAP7_75t_SL g2098 ( 
.A(n_1289),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1311),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1311),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1311),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_1933),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1311),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1368),
.Y(n_2104)
);

CKINVDCx20_ASAP7_75t_R g2105 ( 
.A(n_1111),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1368),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1368),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1368),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1376),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1376),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1376),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1376),
.Y(n_2112)
);

CKINVDCx5p33_ASAP7_75t_R g2113 ( 
.A(n_1910),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1387),
.Y(n_2114)
);

INVxp67_ASAP7_75t_SL g2115 ( 
.A(n_1387),
.Y(n_2115)
);

HB1xp67_ASAP7_75t_L g2116 ( 
.A(n_1913),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1387),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1387),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1410),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1410),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1410),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1410),
.Y(n_2122)
);

HB1xp67_ASAP7_75t_L g2123 ( 
.A(n_1915),
.Y(n_2123)
);

INVxp67_ASAP7_75t_SL g2124 ( 
.A(n_1412),
.Y(n_2124)
);

CKINVDCx20_ASAP7_75t_R g2125 ( 
.A(n_1111),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1412),
.Y(n_2126)
);

INVxp67_ASAP7_75t_L g2127 ( 
.A(n_1128),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1412),
.Y(n_2128)
);

INVx1_ASAP7_75t_SL g2129 ( 
.A(n_1100),
.Y(n_2129)
);

INVxp67_ASAP7_75t_L g2130 ( 
.A(n_1281),
.Y(n_2130)
);

BUFx6f_ASAP7_75t_L g2131 ( 
.A(n_1976),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1935),
.B(n_1185),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2020),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1991),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_2008),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_2033),
.Y(n_2136)
);

OAI21x1_ASAP7_75t_L g2137 ( 
.A1(n_1950),
.A2(n_1377),
.B(n_1228),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2030),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2034),
.Y(n_2139)
);

NOR2xp33_ASAP7_75t_L g2140 ( 
.A(n_2068),
.B(n_1555),
.Y(n_2140)
);

BUFx2_ASAP7_75t_L g2141 ( 
.A(n_2037),
.Y(n_2141)
);

BUFx2_ASAP7_75t_L g2142 ( 
.A(n_2046),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2035),
.Y(n_2143)
);

AND2x4_ASAP7_75t_L g2144 ( 
.A(n_1965),
.B(n_2072),
.Y(n_2144)
);

AOI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_2031),
.A2(n_2043),
.B1(n_2050),
.B2(n_1958),
.Y(n_2145)
);

NAND2xp33_ASAP7_75t_L g2146 ( 
.A(n_2069),
.B(n_1412),
.Y(n_2146)
);

BUFx6f_ASAP7_75t_L g2147 ( 
.A(n_2058),
.Y(n_2147)
);

BUFx6f_ASAP7_75t_L g2148 ( 
.A(n_2085),
.Y(n_2148)
);

INVx5_ASAP7_75t_L g2149 ( 
.A(n_2056),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_L g2150 ( 
.A(n_2081),
.B(n_1911),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2039),
.Y(n_2151)
);

INVx3_ASAP7_75t_L g2152 ( 
.A(n_2001),
.Y(n_2152)
);

AND2x6_ASAP7_75t_L g2153 ( 
.A(n_1977),
.B(n_1139),
.Y(n_2153)
);

OA21x2_ASAP7_75t_L g2154 ( 
.A1(n_1936),
.A2(n_1087),
.B(n_1079),
.Y(n_2154)
);

BUFx2_ASAP7_75t_L g2155 ( 
.A(n_2053),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1946),
.B(n_1502),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_2099),
.Y(n_2157)
);

OR2x6_ASAP7_75t_L g2158 ( 
.A(n_1972),
.B(n_1293),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_2114),
.Y(n_2159)
);

OA21x2_ASAP7_75t_L g2160 ( 
.A1(n_1937),
.A2(n_1087),
.B(n_1079),
.Y(n_2160)
);

INVx3_ASAP7_75t_L g2161 ( 
.A(n_2044),
.Y(n_2161)
);

NAND2xp33_ASAP7_75t_L g2162 ( 
.A(n_2091),
.B(n_1444),
.Y(n_2162)
);

AOI22xp33_ASAP7_75t_SL g2163 ( 
.A1(n_1980),
.A2(n_1137),
.B1(n_1170),
.B2(n_1154),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2118),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2045),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1990),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2066),
.Y(n_2167)
);

NOR2xp33_ASAP7_75t_L g2168 ( 
.A(n_2102),
.B(n_1293),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1952),
.B(n_1502),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2083),
.Y(n_2170)
);

HB1xp67_ASAP7_75t_L g2171 ( 
.A(n_2057),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1990),
.Y(n_2172)
);

BUFx2_ASAP7_75t_L g2173 ( 
.A(n_1934),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_2113),
.B(n_1416),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2098),
.Y(n_2175)
);

OA21x2_ASAP7_75t_L g2176 ( 
.A1(n_1938),
.A2(n_1944),
.B(n_1941),
.Y(n_2176)
);

CKINVDCx14_ASAP7_75t_R g2177 ( 
.A(n_1948),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2092),
.B(n_2116),
.Y(n_2178)
);

BUFx6f_ASAP7_75t_L g2179 ( 
.A(n_2070),
.Y(n_2179)
);

INVx5_ASAP7_75t_L g2180 ( 
.A(n_2056),
.Y(n_2180)
);

OAI21x1_ASAP7_75t_L g2181 ( 
.A1(n_1969),
.A2(n_1970),
.B(n_1947),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1953),
.B(n_1502),
.Y(n_2182)
);

AOI22xp5_ASAP7_75t_L g2183 ( 
.A1(n_1964),
.A2(n_1568),
.B1(n_1785),
.B2(n_1356),
.Y(n_2183)
);

BUFx8_ASAP7_75t_SL g2184 ( 
.A(n_2065),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2073),
.Y(n_2185)
);

AND2x4_ASAP7_75t_L g2186 ( 
.A(n_2087),
.B(n_1084),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2115),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2124),
.Y(n_2188)
);

AND2x6_ASAP7_75t_L g2189 ( 
.A(n_1981),
.B(n_1201),
.Y(n_2189)
);

BUFx12f_ASAP7_75t_L g2190 ( 
.A(n_1967),
.Y(n_2190)
);

INVx2_ASAP7_75t_SL g2191 ( 
.A(n_2123),
.Y(n_2191)
);

BUFx6f_ASAP7_75t_L g2192 ( 
.A(n_2076),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_2078),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_1939),
.B(n_1128),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2079),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_2080),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2082),
.Y(n_2197)
);

AND2x4_ASAP7_75t_L g2198 ( 
.A(n_1943),
.B(n_1433),
.Y(n_2198)
);

INVxp67_ASAP7_75t_L g2199 ( 
.A(n_2017),
.Y(n_2199)
);

AND2x4_ASAP7_75t_L g2200 ( 
.A(n_1979),
.B(n_1633),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_1940),
.B(n_1175),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2084),
.Y(n_2202)
);

INVx3_ASAP7_75t_L g2203 ( 
.A(n_2086),
.Y(n_2203)
);

OAI22xp5_ASAP7_75t_SL g2204 ( 
.A1(n_1975),
.A2(n_1154),
.B1(n_1170),
.B2(n_1137),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1974),
.B(n_1502),
.Y(n_2205)
);

INVx6_ASAP7_75t_L g2206 ( 
.A(n_2075),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2077),
.B(n_1175),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2089),
.Y(n_2208)
);

BUFx6f_ASAP7_75t_L g2209 ( 
.A(n_2090),
.Y(n_2209)
);

INVx3_ASAP7_75t_L g2210 ( 
.A(n_2093),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2100),
.Y(n_2211)
);

BUFx6f_ASAP7_75t_L g2212 ( 
.A(n_2101),
.Y(n_2212)
);

INVx6_ASAP7_75t_L g2213 ( 
.A(n_2095),
.Y(n_2213)
);

HB1xp67_ASAP7_75t_L g2214 ( 
.A(n_2077),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2103),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_1987),
.B(n_1639),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2104),
.Y(n_2217)
);

NAND2xp33_ASAP7_75t_L g2218 ( 
.A(n_1956),
.B(n_1444),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2106),
.Y(n_2219)
);

CKINVDCx6p67_ASAP7_75t_R g2220 ( 
.A(n_1986),
.Y(n_2220)
);

OA21x2_ASAP7_75t_L g2221 ( 
.A1(n_1945),
.A2(n_1144),
.B(n_1122),
.Y(n_2221)
);

AOI22xp5_ASAP7_75t_L g2222 ( 
.A1(n_2022),
.A2(n_1085),
.B1(n_1089),
.B2(n_1088),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2107),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2108),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2109),
.Y(n_2225)
);

CKINVDCx6p67_ASAP7_75t_R g2226 ( 
.A(n_2023),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2110),
.Y(n_2227)
);

INVx2_ASAP7_75t_SL g2228 ( 
.A(n_1966),
.Y(n_2228)
);

INVx4_ASAP7_75t_L g2229 ( 
.A(n_1978),
.Y(n_2229)
);

AND2x4_ASAP7_75t_L g2230 ( 
.A(n_1998),
.B(n_1762),
.Y(n_2230)
);

AND2x4_ASAP7_75t_L g2231 ( 
.A(n_1996),
.B(n_1763),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2129),
.B(n_1175),
.Y(n_2232)
);

AOI22x1_ASAP7_75t_SL g2233 ( 
.A1(n_2088),
.A2(n_1178),
.B1(n_1180),
.B2(n_1176),
.Y(n_2233)
);

BUFx6f_ASAP7_75t_L g2234 ( 
.A(n_2111),
.Y(n_2234)
);

BUFx6f_ASAP7_75t_L g2235 ( 
.A(n_2112),
.Y(n_2235)
);

AND2x4_ASAP7_75t_L g2236 ( 
.A(n_2000),
.B(n_1775),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_2117),
.Y(n_2237)
);

OA21x2_ASAP7_75t_L g2238 ( 
.A1(n_1949),
.A2(n_1144),
.B(n_1122),
.Y(n_2238)
);

AND2x4_ASAP7_75t_L g2239 ( 
.A(n_2002),
.B(n_1786),
.Y(n_2239)
);

OAI22xp5_ASAP7_75t_L g2240 ( 
.A1(n_1956),
.A2(n_1086),
.B1(n_1500),
.B2(n_1275),
.Y(n_2240)
);

BUFx3_ASAP7_75t_L g2241 ( 
.A(n_1982),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2129),
.B(n_1226),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_1995),
.B(n_2015),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2021),
.B(n_1502),
.Y(n_2244)
);

BUFx6f_ASAP7_75t_L g2245 ( 
.A(n_2119),
.Y(n_2245)
);

INVx2_ASAP7_75t_SL g2246 ( 
.A(n_2036),
.Y(n_2246)
);

INVx3_ASAP7_75t_L g2247 ( 
.A(n_2120),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_1983),
.B(n_1502),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2121),
.Y(n_2249)
);

INVx3_ASAP7_75t_L g2250 ( 
.A(n_2122),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2126),
.Y(n_2251)
);

BUFx6f_ASAP7_75t_L g2252 ( 
.A(n_2128),
.Y(n_2252)
);

OA21x2_ASAP7_75t_L g2253 ( 
.A1(n_1951),
.A2(n_1210),
.B(n_1194),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1984),
.Y(n_2254)
);

AOI22xp5_ASAP7_75t_L g2255 ( 
.A1(n_2047),
.A2(n_1090),
.B1(n_1093),
.B2(n_1091),
.Y(n_2255)
);

AND2x4_ASAP7_75t_L g2256 ( 
.A(n_2040),
.B(n_1823),
.Y(n_2256)
);

BUFx6f_ASAP7_75t_L g2257 ( 
.A(n_1954),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1955),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_1957),
.Y(n_2259)
);

BUFx6f_ASAP7_75t_L g2260 ( 
.A(n_1959),
.Y(n_2260)
);

AND2x4_ASAP7_75t_L g2261 ( 
.A(n_2040),
.B(n_1886),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1960),
.Y(n_2262)
);

INVx4_ASAP7_75t_L g2263 ( 
.A(n_1963),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1985),
.Y(n_2264)
);

BUFx6f_ASAP7_75t_L g2265 ( 
.A(n_1961),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1988),
.Y(n_2266)
);

BUFx6f_ASAP7_75t_L g2267 ( 
.A(n_1962),
.Y(n_2267)
);

AND2x4_ASAP7_75t_L g2268 ( 
.A(n_2096),
.B(n_1416),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_1968),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_1989),
.B(n_1502),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_1971),
.B(n_1444),
.Y(n_2271)
);

CKINVDCx5p33_ASAP7_75t_R g2272 ( 
.A(n_2012),
.Y(n_2272)
);

BUFx6f_ASAP7_75t_L g2273 ( 
.A(n_1973),
.Y(n_2273)
);

OAI22xp5_ASAP7_75t_L g2274 ( 
.A1(n_2004),
.A2(n_1097),
.B1(n_1098),
.B2(n_1095),
.Y(n_2274)
);

INVx4_ASAP7_75t_L g2275 ( 
.A(n_2027),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1992),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1993),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1994),
.Y(n_2278)
);

AOI22xp5_ASAP7_75t_L g2279 ( 
.A1(n_2042),
.A2(n_1103),
.B1(n_1106),
.B2(n_1102),
.Y(n_2279)
);

BUFx6f_ASAP7_75t_L g2280 ( 
.A(n_1997),
.Y(n_2280)
);

OAI22xp5_ASAP7_75t_SL g2281 ( 
.A1(n_2094),
.A2(n_1178),
.B1(n_1180),
.B2(n_1176),
.Y(n_2281)
);

CKINVDCx11_ASAP7_75t_R g2282 ( 
.A(n_2097),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2054),
.B(n_1942),
.Y(n_2283)
);

AND2x4_ASAP7_75t_L g2284 ( 
.A(n_2127),
.B(n_1080),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2003),
.B(n_1226),
.Y(n_2285)
);

AND2x6_ASAP7_75t_L g2286 ( 
.A(n_1999),
.B(n_1277),
.Y(n_2286)
);

OAI21x1_ASAP7_75t_L g2287 ( 
.A1(n_2005),
.A2(n_1210),
.B(n_1194),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2006),
.B(n_1444),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2007),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_2049),
.B(n_1446),
.Y(n_2290)
);

AOI22xp5_ASAP7_75t_L g2291 ( 
.A1(n_2062),
.A2(n_1112),
.B1(n_1113),
.B2(n_1109),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2009),
.Y(n_2292)
);

INVx3_ASAP7_75t_L g2293 ( 
.A(n_2010),
.Y(n_2293)
);

BUFx6f_ASAP7_75t_L g2294 ( 
.A(n_2011),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2013),
.B(n_1446),
.Y(n_2295)
);

BUFx6f_ASAP7_75t_L g2296 ( 
.A(n_2014),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2016),
.Y(n_2297)
);

INVx5_ASAP7_75t_L g2298 ( 
.A(n_2071),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2018),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2019),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2024),
.Y(n_2301)
);

OA21x2_ASAP7_75t_L g2302 ( 
.A1(n_2025),
.A2(n_1255),
.B(n_1222),
.Y(n_2302)
);

OAI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2060),
.A2(n_1116),
.B1(n_1117),
.B2(n_1114),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_2026),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2028),
.B(n_1446),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2029),
.Y(n_2306)
);

OA21x2_ASAP7_75t_L g2307 ( 
.A1(n_2032),
.A2(n_1255),
.B(n_1222),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2038),
.B(n_2041),
.Y(n_2308)
);

BUFx6f_ASAP7_75t_L g2309 ( 
.A(n_2048),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2051),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2052),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2055),
.Y(n_2312)
);

AND2x4_ASAP7_75t_L g2313 ( 
.A(n_2059),
.B(n_1092),
.Y(n_2313)
);

BUFx6f_ASAP7_75t_L g2314 ( 
.A(n_2061),
.Y(n_2314)
);

BUFx2_ASAP7_75t_L g2315 ( 
.A(n_2105),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2063),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_SL g2317 ( 
.A(n_2074),
.B(n_1446),
.Y(n_2317)
);

CKINVDCx5p33_ASAP7_75t_R g2318 ( 
.A(n_2125),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_2067),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2064),
.Y(n_2320)
);

OA21x2_ASAP7_75t_L g2321 ( 
.A1(n_2064),
.A2(n_1301),
.B(n_1271),
.Y(n_2321)
);

INVx3_ASAP7_75t_L g2322 ( 
.A(n_2130),
.Y(n_2322)
);

AND2x6_ASAP7_75t_L g2323 ( 
.A(n_2130),
.B(n_1321),
.Y(n_2323)
);

BUFx6f_ASAP7_75t_L g2324 ( 
.A(n_1976),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2020),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2020),
.Y(n_2326)
);

BUFx6f_ASAP7_75t_L g2327 ( 
.A(n_1976),
.Y(n_2327)
);

BUFx2_ASAP7_75t_L g2328 ( 
.A(n_2037),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_1976),
.Y(n_2329)
);

OA21x2_ASAP7_75t_L g2330 ( 
.A1(n_1936),
.A2(n_1301),
.B(n_1271),
.Y(n_2330)
);

INVx3_ASAP7_75t_L g2331 ( 
.A(n_2001),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_1935),
.B(n_1452),
.Y(n_2332)
);

INVx3_ASAP7_75t_L g2333 ( 
.A(n_2001),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_1976),
.Y(n_2334)
);

BUFx6f_ASAP7_75t_L g2335 ( 
.A(n_1976),
.Y(n_2335)
);

AOI22xp5_ASAP7_75t_SL g2336 ( 
.A1(n_1934),
.A2(n_1198),
.B1(n_1204),
.B2(n_1193),
.Y(n_2336)
);

OAI22xp5_ASAP7_75t_SL g2337 ( 
.A1(n_1934),
.A2(n_1198),
.B1(n_1204),
.B2(n_1193),
.Y(n_2337)
);

BUFx6f_ASAP7_75t_L g2338 ( 
.A(n_1976),
.Y(n_2338)
);

BUFx12f_ASAP7_75t_L g2339 ( 
.A(n_2037),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_1976),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2020),
.Y(n_2341)
);

NOR2x1_ASAP7_75t_L g2342 ( 
.A(n_1965),
.B(n_1101),
.Y(n_2342)
);

AOI22x1_ASAP7_75t_SL g2343 ( 
.A1(n_2065),
.A2(n_1219),
.B1(n_1245),
.B2(n_1217),
.Y(n_2343)
);

BUFx6f_ASAP7_75t_L g2344 ( 
.A(n_1976),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_1935),
.B(n_1452),
.Y(n_2345)
);

CKINVDCx5p33_ASAP7_75t_R g2346 ( 
.A(n_1935),
.Y(n_2346)
);

INVx3_ASAP7_75t_L g2347 ( 
.A(n_2001),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2020),
.Y(n_2348)
);

INVx3_ASAP7_75t_L g2349 ( 
.A(n_2001),
.Y(n_2349)
);

BUFx6f_ASAP7_75t_L g2350 ( 
.A(n_1976),
.Y(n_2350)
);

INVx3_ASAP7_75t_L g2351 ( 
.A(n_2001),
.Y(n_2351)
);

BUFx2_ASAP7_75t_L g2352 ( 
.A(n_2037),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_1976),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_1935),
.B(n_1452),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_1976),
.Y(n_2355)
);

AOI22x1_ASAP7_75t_SL g2356 ( 
.A1(n_2065),
.A2(n_1219),
.B1(n_1245),
.B2(n_1217),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_1935),
.B(n_1452),
.Y(n_2357)
);

BUFx6f_ASAP7_75t_L g2358 ( 
.A(n_1976),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2020),
.Y(n_2359)
);

OAI21x1_ASAP7_75t_L g2360 ( 
.A1(n_1950),
.A2(n_1381),
.B(n_1344),
.Y(n_2360)
);

BUFx6f_ASAP7_75t_L g2361 ( 
.A(n_1976),
.Y(n_2361)
);

AND2x4_ASAP7_75t_L g2362 ( 
.A(n_1965),
.B(n_1107),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_1976),
.Y(n_2363)
);

BUFx2_ASAP7_75t_L g2364 ( 
.A(n_2037),
.Y(n_2364)
);

AND2x6_ASAP7_75t_L g2365 ( 
.A(n_1965),
.B(n_1325),
.Y(n_2365)
);

AOI22xp5_ASAP7_75t_L g2366 ( 
.A1(n_2031),
.A2(n_1118),
.B1(n_1120),
.B2(n_1119),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_1976),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2020),
.Y(n_2368)
);

BUFx8_ASAP7_75t_L g2369 ( 
.A(n_2087),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2020),
.Y(n_2370)
);

INVx3_ASAP7_75t_L g2371 ( 
.A(n_2001),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2020),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_1976),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2020),
.Y(n_2374)
);

BUFx8_ASAP7_75t_L g2375 ( 
.A(n_2087),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2020),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_SL g2377 ( 
.A(n_1963),
.B(n_1517),
.Y(n_2377)
);

AOI22xp5_ASAP7_75t_SL g2378 ( 
.A1(n_1934),
.A2(n_1260),
.B1(n_1261),
.B2(n_1246),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_1976),
.Y(n_2379)
);

OAI22xp5_ASAP7_75t_L g2380 ( 
.A1(n_2031),
.A2(n_1124),
.B1(n_1127),
.B2(n_1123),
.Y(n_2380)
);

BUFx6f_ASAP7_75t_L g2381 ( 
.A(n_1976),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2020),
.Y(n_2382)
);

AND2x4_ASAP7_75t_L g2383 ( 
.A(n_1965),
.B(n_1115),
.Y(n_2383)
);

OA21x2_ASAP7_75t_L g2384 ( 
.A1(n_1936),
.A2(n_1381),
.B(n_1344),
.Y(n_2384)
);

AND2x4_ASAP7_75t_L g2385 ( 
.A(n_1965),
.B(n_1121),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2020),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2020),
.Y(n_2387)
);

AOI22xp5_ASAP7_75t_L g2388 ( 
.A1(n_2031),
.A2(n_1130),
.B1(n_1132),
.B2(n_1131),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2020),
.Y(n_2389)
);

AND2x4_ASAP7_75t_L g2390 ( 
.A(n_1965),
.B(n_1129),
.Y(n_2390)
);

BUFx6f_ASAP7_75t_L g2391 ( 
.A(n_1976),
.Y(n_2391)
);

NOR2xp33_ASAP7_75t_L g2392 ( 
.A(n_2068),
.B(n_1517),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2020),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2020),
.Y(n_2394)
);

INVx3_ASAP7_75t_L g2395 ( 
.A(n_2001),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_2092),
.B(n_1226),
.Y(n_2396)
);

AND2x4_ASAP7_75t_L g2397 ( 
.A(n_1965),
.B(n_1134),
.Y(n_2397)
);

AOI22xp5_ASAP7_75t_L g2398 ( 
.A1(n_2031),
.A2(n_1135),
.B1(n_1138),
.B2(n_1133),
.Y(n_2398)
);

HB1xp67_ASAP7_75t_L g2399 ( 
.A(n_2037),
.Y(n_2399)
);

BUFx6f_ASAP7_75t_L g2400 ( 
.A(n_1976),
.Y(n_2400)
);

AND2x4_ASAP7_75t_L g2401 ( 
.A(n_1965),
.B(n_1136),
.Y(n_2401)
);

BUFx6f_ASAP7_75t_L g2402 ( 
.A(n_1976),
.Y(n_2402)
);

BUFx3_ASAP7_75t_L g2403 ( 
.A(n_2001),
.Y(n_2403)
);

HB1xp67_ASAP7_75t_L g2404 ( 
.A(n_2037),
.Y(n_2404)
);

AND2x4_ASAP7_75t_L g2405 ( 
.A(n_1965),
.B(n_1140),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_1935),
.B(n_1517),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_1935),
.B(n_1517),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_1976),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2092),
.B(n_1269),
.Y(n_2409)
);

HB1xp67_ASAP7_75t_L g2410 ( 
.A(n_2037),
.Y(n_2410)
);

INVxp67_ASAP7_75t_L g2411 ( 
.A(n_1972),
.Y(n_2411)
);

BUFx8_ASAP7_75t_SL g2412 ( 
.A(n_2065),
.Y(n_2412)
);

CKINVDCx5p33_ASAP7_75t_R g2413 ( 
.A(n_1935),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2020),
.Y(n_2414)
);

INVx2_ASAP7_75t_SL g2415 ( 
.A(n_2056),
.Y(n_2415)
);

OAI22xp5_ASAP7_75t_SL g2416 ( 
.A1(n_1934),
.A2(n_1260),
.B1(n_1261),
.B2(n_1246),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2092),
.B(n_1269),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_1976),
.Y(n_2418)
);

BUFx3_ASAP7_75t_L g2419 ( 
.A(n_2001),
.Y(n_2419)
);

BUFx3_ASAP7_75t_L g2420 ( 
.A(n_2001),
.Y(n_2420)
);

AND2x4_ASAP7_75t_L g2421 ( 
.A(n_1965),
.B(n_1142),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_1976),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_L g2423 ( 
.A(n_2068),
.B(n_1525),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_1976),
.Y(n_2424)
);

OAI21x1_ASAP7_75t_L g2425 ( 
.A1(n_1950),
.A2(n_1413),
.B(n_1397),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2020),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_SL g2427 ( 
.A(n_1963),
.B(n_1525),
.Y(n_2427)
);

AND2x6_ASAP7_75t_L g2428 ( 
.A(n_1965),
.B(n_1354),
.Y(n_2428)
);

INVx2_ASAP7_75t_SL g2429 ( 
.A(n_2056),
.Y(n_2429)
);

BUFx6f_ASAP7_75t_L g2430 ( 
.A(n_1976),
.Y(n_2430)
);

BUFx2_ASAP7_75t_L g2431 ( 
.A(n_2037),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2020),
.Y(n_2432)
);

OAI22x1_ASAP7_75t_SL g2433 ( 
.A1(n_2065),
.A2(n_1284),
.B1(n_1288),
.B2(n_1273),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_1976),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2020),
.Y(n_2435)
);

BUFx6f_ASAP7_75t_L g2436 ( 
.A(n_1976),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_1976),
.Y(n_2437)
);

INVxp67_ASAP7_75t_L g2438 ( 
.A(n_1972),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_1935),
.B(n_1525),
.Y(n_2439)
);

BUFx6f_ASAP7_75t_L g2440 ( 
.A(n_1976),
.Y(n_2440)
);

AOI22xp5_ASAP7_75t_SL g2441 ( 
.A1(n_1934),
.A2(n_1284),
.B1(n_1288),
.B2(n_1273),
.Y(n_2441)
);

OAI21x1_ASAP7_75t_L g2442 ( 
.A1(n_1950),
.A2(n_1413),
.B(n_1397),
.Y(n_2442)
);

INVx6_ASAP7_75t_L g2443 ( 
.A(n_2056),
.Y(n_2443)
);

INVx4_ASAP7_75t_L g2444 ( 
.A(n_1935),
.Y(n_2444)
);

AND2x2_ASAP7_75t_L g2445 ( 
.A(n_2092),
.B(n_1269),
.Y(n_2445)
);

AND2x6_ASAP7_75t_L g2446 ( 
.A(n_1965),
.B(n_1364),
.Y(n_2446)
);

BUFx6f_ASAP7_75t_L g2447 ( 
.A(n_1976),
.Y(n_2447)
);

BUFx6f_ASAP7_75t_L g2448 ( 
.A(n_1976),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2020),
.Y(n_2449)
);

OAI22x1_ASAP7_75t_L g2450 ( 
.A1(n_1956),
.A2(n_1428),
.B1(n_1458),
.B2(n_1419),
.Y(n_2450)
);

BUFx3_ASAP7_75t_L g2451 ( 
.A(n_2001),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2092),
.B(n_1319),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_1976),
.Y(n_2453)
);

INVx4_ASAP7_75t_L g2454 ( 
.A(n_1935),
.Y(n_2454)
);

BUFx3_ASAP7_75t_L g2455 ( 
.A(n_2001),
.Y(n_2455)
);

AND2x4_ASAP7_75t_L g2456 ( 
.A(n_1965),
.B(n_1145),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2020),
.Y(n_2457)
);

OA21x2_ASAP7_75t_L g2458 ( 
.A1(n_1936),
.A2(n_1442),
.B(n_1431),
.Y(n_2458)
);

OAI21x1_ASAP7_75t_L g2459 ( 
.A1(n_1950),
.A2(n_1442),
.B(n_1431),
.Y(n_2459)
);

BUFx6f_ASAP7_75t_L g2460 ( 
.A(n_1976),
.Y(n_2460)
);

BUFx2_ASAP7_75t_L g2461 ( 
.A(n_2037),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2020),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_1935),
.B(n_1525),
.Y(n_2463)
);

AOI22xp5_ASAP7_75t_L g2464 ( 
.A1(n_2031),
.A2(n_1143),
.B1(n_1146),
.B2(n_1141),
.Y(n_2464)
);

INVx3_ASAP7_75t_L g2465 ( 
.A(n_2001),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_1976),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_1935),
.B(n_1551),
.Y(n_2467)
);

NOR2x1_ASAP7_75t_L g2468 ( 
.A(n_1965),
.B(n_1151),
.Y(n_2468)
);

AND2x4_ASAP7_75t_L g2469 ( 
.A(n_1965),
.B(n_1156),
.Y(n_2469)
);

INVx3_ASAP7_75t_L g2470 ( 
.A(n_2001),
.Y(n_2470)
);

OAI22x1_ASAP7_75t_L g2471 ( 
.A1(n_1956),
.A2(n_1497),
.B1(n_1501),
.B2(n_1467),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_1935),
.B(n_1551),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_2131),
.Y(n_2473)
);

INVxp67_ASAP7_75t_SL g2474 ( 
.A(n_2152),
.Y(n_2474)
);

NOR2xp33_ASAP7_75t_R g2475 ( 
.A(n_2177),
.B(n_2346),
.Y(n_2475)
);

CKINVDCx5p33_ASAP7_75t_R g2476 ( 
.A(n_2413),
.Y(n_2476)
);

CKINVDCx5p33_ASAP7_75t_R g2477 ( 
.A(n_2184),
.Y(n_2477)
);

CKINVDCx5p33_ASAP7_75t_R g2478 ( 
.A(n_2412),
.Y(n_2478)
);

CKINVDCx5p33_ASAP7_75t_R g2479 ( 
.A(n_2190),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_2282),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2254),
.Y(n_2481)
);

BUFx6f_ASAP7_75t_L g2482 ( 
.A(n_2287),
.Y(n_2482)
);

CKINVDCx20_ASAP7_75t_R g2483 ( 
.A(n_2318),
.Y(n_2483)
);

CKINVDCx5p33_ASAP7_75t_R g2484 ( 
.A(n_2214),
.Y(n_2484)
);

CKINVDCx20_ASAP7_75t_R g2485 ( 
.A(n_2220),
.Y(n_2485)
);

CKINVDCx5p33_ASAP7_75t_R g2486 ( 
.A(n_2339),
.Y(n_2486)
);

CKINVDCx5p33_ASAP7_75t_R g2487 ( 
.A(n_2272),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_2229),
.Y(n_2488)
);

BUFx2_ASAP7_75t_L g2489 ( 
.A(n_2283),
.Y(n_2489)
);

CKINVDCx5p33_ASAP7_75t_R g2490 ( 
.A(n_2444),
.Y(n_2490)
);

NOR2xp33_ASAP7_75t_R g2491 ( 
.A(n_2146),
.B(n_2162),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2264),
.Y(n_2492)
);

CKINVDCx5p33_ASAP7_75t_R g2493 ( 
.A(n_2454),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2131),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2147),
.Y(n_2495)
);

CKINVDCx5p33_ASAP7_75t_R g2496 ( 
.A(n_2226),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2266),
.Y(n_2497)
);

CKINVDCx5p33_ASAP7_75t_R g2498 ( 
.A(n_2246),
.Y(n_2498)
);

CKINVDCx5p33_ASAP7_75t_R g2499 ( 
.A(n_2243),
.Y(n_2499)
);

AND2x4_ASAP7_75t_L g2500 ( 
.A(n_2362),
.B(n_1160),
.Y(n_2500)
);

CKINVDCx5p33_ASAP7_75t_R g2501 ( 
.A(n_2141),
.Y(n_2501)
);

INVxp33_ASAP7_75t_SL g2502 ( 
.A(n_2204),
.Y(n_2502)
);

NOR2xp33_ASAP7_75t_R g2503 ( 
.A(n_2415),
.B(n_1147),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2332),
.B(n_2345),
.Y(n_2504)
);

CKINVDCx5p33_ASAP7_75t_R g2505 ( 
.A(n_2142),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_2155),
.Y(n_2506)
);

CKINVDCx5p33_ASAP7_75t_R g2507 ( 
.A(n_2328),
.Y(n_2507)
);

CKINVDCx5p33_ASAP7_75t_R g2508 ( 
.A(n_2352),
.Y(n_2508)
);

CKINVDCx5p33_ASAP7_75t_R g2509 ( 
.A(n_2364),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_2207),
.B(n_1319),
.Y(n_2510)
);

INVxp67_ASAP7_75t_SL g2511 ( 
.A(n_2161),
.Y(n_2511)
);

CKINVDCx5p33_ASAP7_75t_R g2512 ( 
.A(n_2431),
.Y(n_2512)
);

CKINVDCx5p33_ASAP7_75t_R g2513 ( 
.A(n_2461),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2276),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2354),
.B(n_1551),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2277),
.Y(n_2516)
);

CKINVDCx5p33_ASAP7_75t_R g2517 ( 
.A(n_2443),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2278),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2289),
.Y(n_2519)
);

CKINVDCx5p33_ASAP7_75t_R g2520 ( 
.A(n_2149),
.Y(n_2520)
);

OA21x2_ASAP7_75t_L g2521 ( 
.A1(n_2360),
.A2(n_1506),
.B(n_1460),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2292),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2297),
.Y(n_2523)
);

CKINVDCx5p33_ASAP7_75t_R g2524 ( 
.A(n_2149),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2147),
.Y(n_2525)
);

CKINVDCx20_ASAP7_75t_R g2526 ( 
.A(n_2315),
.Y(n_2526)
);

BUFx3_ASAP7_75t_L g2527 ( 
.A(n_2403),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2357),
.B(n_1551),
.Y(n_2528)
);

CKINVDCx5p33_ASAP7_75t_R g2529 ( 
.A(n_2180),
.Y(n_2529)
);

CKINVDCx5p33_ASAP7_75t_R g2530 ( 
.A(n_2180),
.Y(n_2530)
);

CKINVDCx5p33_ASAP7_75t_R g2531 ( 
.A(n_2369),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2148),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2148),
.Y(n_2533)
);

CKINVDCx5p33_ASAP7_75t_R g2534 ( 
.A(n_2375),
.Y(n_2534)
);

NAND2xp33_ASAP7_75t_R g2535 ( 
.A(n_2178),
.B(n_1149),
.Y(n_2535)
);

BUFx3_ASAP7_75t_L g2536 ( 
.A(n_2419),
.Y(n_2536)
);

CKINVDCx20_ASAP7_75t_R g2537 ( 
.A(n_2173),
.Y(n_2537)
);

CKINVDCx5p33_ASAP7_75t_R g2538 ( 
.A(n_2206),
.Y(n_2538)
);

CKINVDCx5p33_ASAP7_75t_R g2539 ( 
.A(n_2213),
.Y(n_2539)
);

CKINVDCx5p33_ASAP7_75t_R g2540 ( 
.A(n_2171),
.Y(n_2540)
);

CKINVDCx5p33_ASAP7_75t_R g2541 ( 
.A(n_2399),
.Y(n_2541)
);

CKINVDCx5p33_ASAP7_75t_R g2542 ( 
.A(n_2404),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2299),
.Y(n_2543)
);

INVx3_ASAP7_75t_L g2544 ( 
.A(n_2324),
.Y(n_2544)
);

BUFx10_ASAP7_75t_L g2545 ( 
.A(n_2429),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2324),
.Y(n_2546)
);

CKINVDCx5p33_ASAP7_75t_R g2547 ( 
.A(n_2410),
.Y(n_2547)
);

CKINVDCx20_ASAP7_75t_R g2548 ( 
.A(n_2263),
.Y(n_2548)
);

XOR2x2_ASAP7_75t_L g2549 ( 
.A(n_2336),
.B(n_1503),
.Y(n_2549)
);

CKINVDCx5p33_ASAP7_75t_R g2550 ( 
.A(n_2411),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2300),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2327),
.Y(n_2552)
);

NOR2xp33_ASAP7_75t_R g2553 ( 
.A(n_2191),
.B(n_1150),
.Y(n_2553)
);

CKINVDCx5p33_ASAP7_75t_R g2554 ( 
.A(n_2438),
.Y(n_2554)
);

CKINVDCx5p33_ASAP7_75t_R g2555 ( 
.A(n_2420),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2232),
.B(n_1319),
.Y(n_2556)
);

CKINVDCx5p33_ASAP7_75t_R g2557 ( 
.A(n_2451),
.Y(n_2557)
);

HB1xp67_ASAP7_75t_L g2558 ( 
.A(n_2298),
.Y(n_2558)
);

BUFx3_ASAP7_75t_L g2559 ( 
.A(n_2455),
.Y(n_2559)
);

CKINVDCx20_ASAP7_75t_R g2560 ( 
.A(n_2275),
.Y(n_2560)
);

CKINVDCx5p33_ASAP7_75t_R g2561 ( 
.A(n_2158),
.Y(n_2561)
);

BUFx6f_ASAP7_75t_L g2562 ( 
.A(n_2425),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2327),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2301),
.Y(n_2564)
);

CKINVDCx5p33_ASAP7_75t_R g2565 ( 
.A(n_2150),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2306),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2311),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2312),
.Y(n_2568)
);

CKINVDCx5p33_ASAP7_75t_R g2569 ( 
.A(n_2298),
.Y(n_2569)
);

CKINVDCx5p33_ASAP7_75t_R g2570 ( 
.A(n_2406),
.Y(n_2570)
);

CKINVDCx5p33_ASAP7_75t_R g2571 ( 
.A(n_2407),
.Y(n_2571)
);

CKINVDCx5p33_ASAP7_75t_R g2572 ( 
.A(n_2439),
.Y(n_2572)
);

CKINVDCx20_ASAP7_75t_R g2573 ( 
.A(n_2145),
.Y(n_2573)
);

CKINVDCx5p33_ASAP7_75t_R g2574 ( 
.A(n_2463),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2257),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2335),
.Y(n_2576)
);

HB1xp67_ASAP7_75t_L g2577 ( 
.A(n_2242),
.Y(n_2577)
);

CKINVDCx5p33_ASAP7_75t_R g2578 ( 
.A(n_2467),
.Y(n_2578)
);

CKINVDCx5p33_ASAP7_75t_R g2579 ( 
.A(n_2472),
.Y(n_2579)
);

CKINVDCx5p33_ASAP7_75t_R g2580 ( 
.A(n_2156),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2257),
.Y(n_2581)
);

CKINVDCx5p33_ASAP7_75t_R g2582 ( 
.A(n_2169),
.Y(n_2582)
);

CKINVDCx5p33_ASAP7_75t_R g2583 ( 
.A(n_2182),
.Y(n_2583)
);

NOR2xp67_ASAP7_75t_L g2584 ( 
.A(n_2322),
.B(n_1036),
.Y(n_2584)
);

CKINVDCx5p33_ASAP7_75t_R g2585 ( 
.A(n_2205),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2335),
.Y(n_2586)
);

CKINVDCx5p33_ASAP7_75t_R g2587 ( 
.A(n_2244),
.Y(n_2587)
);

CKINVDCx5p33_ASAP7_75t_R g2588 ( 
.A(n_2144),
.Y(n_2588)
);

CKINVDCx5p33_ASAP7_75t_R g2589 ( 
.A(n_2140),
.Y(n_2589)
);

CKINVDCx5p33_ASAP7_75t_R g2590 ( 
.A(n_2331),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2338),
.Y(n_2591)
);

AND2x2_ASAP7_75t_L g2592 ( 
.A(n_2285),
.B(n_2396),
.Y(n_2592)
);

CKINVDCx5p33_ASAP7_75t_R g2593 ( 
.A(n_2333),
.Y(n_2593)
);

BUFx10_ASAP7_75t_L g2594 ( 
.A(n_2168),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2409),
.B(n_1328),
.Y(n_2595)
);

CKINVDCx5p33_ASAP7_75t_R g2596 ( 
.A(n_2347),
.Y(n_2596)
);

INVx3_ASAP7_75t_L g2597 ( 
.A(n_2338),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2260),
.Y(n_2598)
);

CKINVDCx5p33_ASAP7_75t_R g2599 ( 
.A(n_2349),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2344),
.Y(n_2600)
);

NOR2xp33_ASAP7_75t_L g2601 ( 
.A(n_2132),
.B(n_1152),
.Y(n_2601)
);

CKINVDCx5p33_ASAP7_75t_R g2602 ( 
.A(n_2351),
.Y(n_2602)
);

CKINVDCx20_ASAP7_75t_R g2603 ( 
.A(n_2281),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2260),
.Y(n_2604)
);

HB1xp67_ASAP7_75t_L g2605 ( 
.A(n_2371),
.Y(n_2605)
);

CKINVDCx5p33_ASAP7_75t_R g2606 ( 
.A(n_2395),
.Y(n_2606)
);

CKINVDCx5p33_ASAP7_75t_R g2607 ( 
.A(n_2465),
.Y(n_2607)
);

AOI22xp5_ASAP7_75t_L g2608 ( 
.A1(n_2183),
.A2(n_1549),
.B1(n_1565),
.B2(n_1532),
.Y(n_2608)
);

CKINVDCx5p33_ASAP7_75t_R g2609 ( 
.A(n_2470),
.Y(n_2609)
);

OAI22xp33_ASAP7_75t_L g2610 ( 
.A1(n_2366),
.A2(n_1611),
.B1(n_1621),
.B2(n_1572),
.Y(n_2610)
);

CKINVDCx5p33_ASAP7_75t_R g2611 ( 
.A(n_2392),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2265),
.Y(n_2612)
);

BUFx2_ASAP7_75t_L g2613 ( 
.A(n_2323),
.Y(n_2613)
);

INVxp67_ASAP7_75t_SL g2614 ( 
.A(n_2265),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2344),
.Y(n_2615)
);

CKINVDCx5p33_ASAP7_75t_R g2616 ( 
.A(n_2423),
.Y(n_2616)
);

CKINVDCx5p33_ASAP7_75t_R g2617 ( 
.A(n_2380),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2267),
.Y(n_2618)
);

AND2x4_ASAP7_75t_L g2619 ( 
.A(n_2383),
.B(n_1163),
.Y(n_2619)
);

BUFx6f_ASAP7_75t_L g2620 ( 
.A(n_2442),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2350),
.Y(n_2621)
);

CKINVDCx20_ASAP7_75t_R g2622 ( 
.A(n_2222),
.Y(n_2622)
);

CKINVDCx5p33_ASAP7_75t_R g2623 ( 
.A(n_2174),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2133),
.B(n_1588),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2267),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2350),
.Y(n_2626)
);

CKINVDCx5p33_ASAP7_75t_R g2627 ( 
.A(n_2337),
.Y(n_2627)
);

CKINVDCx5p33_ASAP7_75t_R g2628 ( 
.A(n_2416),
.Y(n_2628)
);

CKINVDCx5p33_ASAP7_75t_R g2629 ( 
.A(n_2255),
.Y(n_2629)
);

CKINVDCx20_ASAP7_75t_R g2630 ( 
.A(n_2199),
.Y(n_2630)
);

BUFx3_ASAP7_75t_L g2631 ( 
.A(n_2241),
.Y(n_2631)
);

CKINVDCx5p33_ASAP7_75t_R g2632 ( 
.A(n_2303),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2273),
.Y(n_2633)
);

HB1xp67_ASAP7_75t_L g2634 ( 
.A(n_2417),
.Y(n_2634)
);

CKINVDCx16_ASAP7_75t_R g2635 ( 
.A(n_2233),
.Y(n_2635)
);

HB1xp67_ASAP7_75t_L g2636 ( 
.A(n_2445),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2358),
.Y(n_2637)
);

NAND2xp33_ASAP7_75t_SL g2638 ( 
.A(n_2450),
.B(n_1299),
.Y(n_2638)
);

BUFx2_ASAP7_75t_L g2639 ( 
.A(n_2323),
.Y(n_2639)
);

CKINVDCx5p33_ASAP7_75t_R g2640 ( 
.A(n_2433),
.Y(n_2640)
);

NOR2xp33_ASAP7_75t_R g2641 ( 
.A(n_2138),
.B(n_1153),
.Y(n_2641)
);

CKINVDCx5p33_ASAP7_75t_R g2642 ( 
.A(n_2279),
.Y(n_2642)
);

CKINVDCx20_ASAP7_75t_R g2643 ( 
.A(n_2291),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2273),
.Y(n_2644)
);

CKINVDCx5p33_ASAP7_75t_R g2645 ( 
.A(n_2343),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2280),
.Y(n_2646)
);

CKINVDCx20_ASAP7_75t_R g2647 ( 
.A(n_2378),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2280),
.Y(n_2648)
);

CKINVDCx5p33_ASAP7_75t_R g2649 ( 
.A(n_2356),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2294),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_2365),
.Y(n_2651)
);

CKINVDCx5p33_ASAP7_75t_R g2652 ( 
.A(n_2365),
.Y(n_2652)
);

CKINVDCx16_ASAP7_75t_R g2653 ( 
.A(n_2452),
.Y(n_2653)
);

CKINVDCx5p33_ASAP7_75t_R g2654 ( 
.A(n_2428),
.Y(n_2654)
);

BUFx8_ASAP7_75t_SL g2655 ( 
.A(n_2284),
.Y(n_2655)
);

CKINVDCx5p33_ASAP7_75t_R g2656 ( 
.A(n_2428),
.Y(n_2656)
);

CKINVDCx5p33_ASAP7_75t_R g2657 ( 
.A(n_2446),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2294),
.Y(n_2658)
);

CKINVDCx5p33_ASAP7_75t_R g2659 ( 
.A(n_2446),
.Y(n_2659)
);

CKINVDCx5p33_ASAP7_75t_R g2660 ( 
.A(n_2388),
.Y(n_2660)
);

NOR2xp67_ASAP7_75t_L g2661 ( 
.A(n_2293),
.B(n_1038),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2358),
.Y(n_2662)
);

CKINVDCx5p33_ASAP7_75t_R g2663 ( 
.A(n_2398),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2296),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2361),
.Y(n_2665)
);

CKINVDCx5p33_ASAP7_75t_R g2666 ( 
.A(n_2464),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2151),
.B(n_1588),
.Y(n_2667)
);

CKINVDCx5p33_ASAP7_75t_R g2668 ( 
.A(n_2274),
.Y(n_2668)
);

AND3x2_ASAP7_75t_L g2669 ( 
.A(n_2194),
.B(n_1506),
.C(n_1460),
.Y(n_2669)
);

CKINVDCx5p33_ASAP7_75t_R g2670 ( 
.A(n_2441),
.Y(n_2670)
);

HB1xp67_ASAP7_75t_L g2671 ( 
.A(n_2320),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2296),
.Y(n_2672)
);

HB1xp67_ASAP7_75t_L g2673 ( 
.A(n_2228),
.Y(n_2673)
);

CKINVDCx20_ASAP7_75t_R g2674 ( 
.A(n_2271),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2361),
.Y(n_2675)
);

BUFx10_ASAP7_75t_L g2676 ( 
.A(n_2231),
.Y(n_2676)
);

HB1xp67_ASAP7_75t_L g2677 ( 
.A(n_2201),
.Y(n_2677)
);

BUFx3_ASAP7_75t_L g2678 ( 
.A(n_2308),
.Y(n_2678)
);

CKINVDCx20_ASAP7_75t_R g2679 ( 
.A(n_2290),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2379),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2309),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2379),
.Y(n_2682)
);

INVx3_ASAP7_75t_L g2683 ( 
.A(n_2381),
.Y(n_2683)
);

NOR2xp33_ASAP7_75t_R g2684 ( 
.A(n_2165),
.B(n_1155),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2309),
.Y(n_2685)
);

NOR2xp33_ASAP7_75t_R g2686 ( 
.A(n_2167),
.B(n_1158),
.Y(n_2686)
);

BUFx10_ASAP7_75t_L g2687 ( 
.A(n_2236),
.Y(n_2687)
);

CKINVDCx5p33_ASAP7_75t_R g2688 ( 
.A(n_2163),
.Y(n_2688)
);

CKINVDCx5p33_ASAP7_75t_R g2689 ( 
.A(n_2186),
.Y(n_2689)
);

CKINVDCx5p33_ASAP7_75t_R g2690 ( 
.A(n_2170),
.Y(n_2690)
);

BUFx6f_ASAP7_75t_SL g2691 ( 
.A(n_2153),
.Y(n_2691)
);

CKINVDCx5p33_ASAP7_75t_R g2692 ( 
.A(n_2175),
.Y(n_2692)
);

INVx3_ASAP7_75t_L g2693 ( 
.A(n_2381),
.Y(n_2693)
);

NOR2xp33_ASAP7_75t_R g2694 ( 
.A(n_2187),
.B(n_1161),
.Y(n_2694)
);

BUFx6f_ASAP7_75t_L g2695 ( 
.A(n_2459),
.Y(n_2695)
);

CKINVDCx5p33_ASAP7_75t_R g2696 ( 
.A(n_2188),
.Y(n_2696)
);

BUFx2_ASAP7_75t_L g2697 ( 
.A(n_2153),
.Y(n_2697)
);

CKINVDCx5p33_ASAP7_75t_R g2698 ( 
.A(n_2325),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2314),
.Y(n_2699)
);

CKINVDCx5p33_ASAP7_75t_R g2700 ( 
.A(n_2326),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2314),
.Y(n_2701)
);

CKINVDCx5p33_ASAP7_75t_R g2702 ( 
.A(n_2341),
.Y(n_2702)
);

CKINVDCx5p33_ASAP7_75t_R g2703 ( 
.A(n_2348),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2304),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2310),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2316),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2319),
.Y(n_2707)
);

CKINVDCx16_ASAP7_75t_R g2708 ( 
.A(n_2239),
.Y(n_2708)
);

BUFx2_ASAP7_75t_L g2709 ( 
.A(n_2189),
.Y(n_2709)
);

CKINVDCx5p33_ASAP7_75t_R g2710 ( 
.A(n_2359),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2154),
.Y(n_2711)
);

CKINVDCx5p33_ASAP7_75t_R g2712 ( 
.A(n_2368),
.Y(n_2712)
);

INVx3_ASAP7_75t_L g2713 ( 
.A(n_2391),
.Y(n_2713)
);

OAI22xp5_ASAP7_75t_SL g2714 ( 
.A1(n_2471),
.A2(n_1302),
.B1(n_1330),
.B2(n_1299),
.Y(n_2714)
);

NOR2xp33_ASAP7_75t_L g2715 ( 
.A(n_2370),
.B(n_1164),
.Y(n_2715)
);

CKINVDCx20_ASAP7_75t_R g2716 ( 
.A(n_2377),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2372),
.B(n_1588),
.Y(n_2717)
);

BUFx2_ASAP7_75t_L g2718 ( 
.A(n_2189),
.Y(n_2718)
);

CKINVDCx5p33_ASAP7_75t_R g2719 ( 
.A(n_2374),
.Y(n_2719)
);

CKINVDCx20_ASAP7_75t_R g2720 ( 
.A(n_2427),
.Y(n_2720)
);

CKINVDCx5p33_ASAP7_75t_R g2721 ( 
.A(n_2376),
.Y(n_2721)
);

CKINVDCx5p33_ASAP7_75t_R g2722 ( 
.A(n_2382),
.Y(n_2722)
);

CKINVDCx20_ASAP7_75t_R g2723 ( 
.A(n_2317),
.Y(n_2723)
);

CKINVDCx5p33_ASAP7_75t_R g2724 ( 
.A(n_2386),
.Y(n_2724)
);

CKINVDCx20_ASAP7_75t_R g2725 ( 
.A(n_2387),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2391),
.Y(n_2726)
);

HB1xp67_ASAP7_75t_L g2727 ( 
.A(n_2385),
.Y(n_2727)
);

CKINVDCx20_ASAP7_75t_R g2728 ( 
.A(n_2389),
.Y(n_2728)
);

CKINVDCx20_ASAP7_75t_R g2729 ( 
.A(n_2393),
.Y(n_2729)
);

NOR2xp67_ASAP7_75t_L g2730 ( 
.A(n_2203),
.B(n_1040),
.Y(n_2730)
);

NOR2xp67_ASAP7_75t_L g2731 ( 
.A(n_2210),
.B(n_1043),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_SL g2732 ( 
.A(n_2198),
.B(n_1328),
.Y(n_2732)
);

BUFx16f_ASAP7_75t_R g2733 ( 
.A(n_2268),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2160),
.Y(n_2734)
);

CKINVDCx5p33_ASAP7_75t_R g2735 ( 
.A(n_2394),
.Y(n_2735)
);

CKINVDCx5p33_ASAP7_75t_R g2736 ( 
.A(n_2414),
.Y(n_2736)
);

NOR2xp33_ASAP7_75t_L g2737 ( 
.A(n_2426),
.B(n_1165),
.Y(n_2737)
);

CKINVDCx5p33_ASAP7_75t_R g2738 ( 
.A(n_2432),
.Y(n_2738)
);

HB1xp67_ASAP7_75t_L g2739 ( 
.A(n_2390),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2200),
.B(n_1328),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2221),
.Y(n_2741)
);

CKINVDCx5p33_ASAP7_75t_R g2742 ( 
.A(n_2435),
.Y(n_2742)
);

CKINVDCx5p33_ASAP7_75t_R g2743 ( 
.A(n_2449),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2400),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2238),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_2457),
.Y(n_2746)
);

INVx3_ASAP7_75t_L g2747 ( 
.A(n_2400),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2253),
.Y(n_2748)
);

CKINVDCx5p33_ASAP7_75t_R g2749 ( 
.A(n_2462),
.Y(n_2749)
);

HB1xp67_ASAP7_75t_L g2750 ( 
.A(n_2397),
.Y(n_2750)
);

NOR2xp33_ASAP7_75t_R g2751 ( 
.A(n_2218),
.B(n_1166),
.Y(n_2751)
);

CKINVDCx5p33_ASAP7_75t_R g2752 ( 
.A(n_2216),
.Y(n_2752)
);

CKINVDCx5p33_ASAP7_75t_R g2753 ( 
.A(n_2230),
.Y(n_2753)
);

HB1xp67_ASAP7_75t_L g2754 ( 
.A(n_2401),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2330),
.Y(n_2755)
);

CKINVDCx5p33_ASAP7_75t_R g2756 ( 
.A(n_2286),
.Y(n_2756)
);

INVx3_ASAP7_75t_L g2757 ( 
.A(n_2402),
.Y(n_2757)
);

CKINVDCx5p33_ASAP7_75t_R g2758 ( 
.A(n_2286),
.Y(n_2758)
);

CKINVDCx5p33_ASAP7_75t_R g2759 ( 
.A(n_2405),
.Y(n_2759)
);

CKINVDCx5p33_ASAP7_75t_R g2760 ( 
.A(n_2421),
.Y(n_2760)
);

CKINVDCx5p33_ASAP7_75t_R g2761 ( 
.A(n_2456),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2384),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2402),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2430),
.Y(n_2764)
);

CKINVDCx5p33_ASAP7_75t_R g2765 ( 
.A(n_2469),
.Y(n_2765)
);

CKINVDCx5p33_ASAP7_75t_R g2766 ( 
.A(n_2256),
.Y(n_2766)
);

CKINVDCx5p33_ASAP7_75t_R g2767 ( 
.A(n_2261),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2458),
.Y(n_2768)
);

AND2x2_ASAP7_75t_L g2769 ( 
.A(n_2342),
.B(n_1411),
.Y(n_2769)
);

CKINVDCx5p33_ASAP7_75t_R g2770 ( 
.A(n_2240),
.Y(n_2770)
);

INVxp67_ASAP7_75t_L g2771 ( 
.A(n_2468),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2258),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2430),
.Y(n_2773)
);

NOR2xp33_ASAP7_75t_L g2774 ( 
.A(n_2195),
.B(n_1169),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2436),
.Y(n_2775)
);

CKINVDCx5p33_ASAP7_75t_R g2776 ( 
.A(n_2436),
.Y(n_2776)
);

CKINVDCx5p33_ASAP7_75t_R g2777 ( 
.A(n_2440),
.Y(n_2777)
);

CKINVDCx5p33_ASAP7_75t_R g2778 ( 
.A(n_2440),
.Y(n_2778)
);

CKINVDCx5p33_ASAP7_75t_R g2779 ( 
.A(n_2447),
.Y(n_2779)
);

CKINVDCx20_ASAP7_75t_R g2780 ( 
.A(n_2248),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2772),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2481),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_2580),
.B(n_2259),
.Y(n_2783)
);

OR2x2_ASAP7_75t_L g2784 ( 
.A(n_2577),
.B(n_2321),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_SL g2785 ( 
.A(n_2570),
.B(n_2447),
.Y(n_2785)
);

INVx3_ASAP7_75t_L g2786 ( 
.A(n_2631),
.Y(n_2786)
);

AO21x2_ASAP7_75t_L g2787 ( 
.A1(n_2504),
.A2(n_2137),
.B(n_2270),
.Y(n_2787)
);

BUFx3_ASAP7_75t_L g2788 ( 
.A(n_2527),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_SL g2789 ( 
.A(n_2517),
.B(n_1352),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2492),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_2582),
.B(n_2262),
.Y(n_2791)
);

AND2x2_ASAP7_75t_L g2792 ( 
.A(n_2510),
.B(n_2313),
.Y(n_2792)
);

AOI22xp33_ASAP7_75t_L g2793 ( 
.A1(n_2711),
.A2(n_2176),
.B1(n_2269),
.B2(n_2181),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2704),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2497),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2705),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_SL g2797 ( 
.A(n_2571),
.B(n_2448),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2583),
.B(n_2302),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_SL g2799 ( 
.A(n_2572),
.B(n_2448),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2585),
.B(n_2307),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_SL g2801 ( 
.A(n_2574),
.B(n_2460),
.Y(n_2801)
);

INVx2_ASAP7_75t_SL g2802 ( 
.A(n_2484),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2514),
.Y(n_2803)
);

INVx4_ASAP7_75t_L g2804 ( 
.A(n_2776),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_2706),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2707),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2516),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2518),
.Y(n_2808)
);

BUFx2_ASAP7_75t_L g2809 ( 
.A(n_2526),
.Y(n_2809)
);

INVx2_ASAP7_75t_SL g2810 ( 
.A(n_2676),
.Y(n_2810)
);

INVx2_ASAP7_75t_SL g2811 ( 
.A(n_2676),
.Y(n_2811)
);

AND2x6_ASAP7_75t_L g2812 ( 
.A(n_2734),
.B(n_1524),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2519),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2522),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2523),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2543),
.Y(n_2816)
);

AND2x2_ASAP7_75t_L g2817 ( 
.A(n_2556),
.B(n_2288),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2587),
.B(n_2460),
.Y(n_2818)
);

BUFx2_ASAP7_75t_L g2819 ( 
.A(n_2613),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2551),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2564),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2566),
.Y(n_2822)
);

AND2x4_ASAP7_75t_L g2823 ( 
.A(n_2536),
.B(n_2197),
.Y(n_2823)
);

AOI22xp33_ASAP7_75t_L g2824 ( 
.A1(n_2741),
.A2(n_2748),
.B1(n_2755),
.B2(n_2745),
.Y(n_2824)
);

INVx3_ASAP7_75t_L g2825 ( 
.A(n_2777),
.Y(n_2825)
);

AND2x4_ASAP7_75t_L g2826 ( 
.A(n_2559),
.B(n_2202),
.Y(n_2826)
);

BUFx2_ASAP7_75t_L g2827 ( 
.A(n_2639),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2567),
.Y(n_2828)
);

NOR2xp33_ASAP7_75t_L g2829 ( 
.A(n_2589),
.B(n_1700),
.Y(n_2829)
);

BUFx3_ASAP7_75t_L g2830 ( 
.A(n_2778),
.Y(n_2830)
);

BUFx6f_ASAP7_75t_L g2831 ( 
.A(n_2544),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_R g2832 ( 
.A(n_2477),
.B(n_1172),
.Y(n_2832)
);

BUFx3_ASAP7_75t_L g2833 ( 
.A(n_2779),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_SL g2834 ( 
.A(n_2578),
.B(n_2179),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2568),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2592),
.B(n_2295),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2544),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2579),
.B(n_2134),
.Y(n_2838)
);

AND2x4_ASAP7_75t_SL g2839 ( 
.A(n_2545),
.B(n_1411),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2678),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2671),
.Y(n_2841)
);

NOR2xp33_ASAP7_75t_L g2842 ( 
.A(n_2565),
.B(n_1803),
.Y(n_2842)
);

AOI22xp5_ASAP7_75t_L g2843 ( 
.A1(n_2668),
.A2(n_2217),
.B1(n_2219),
.B2(n_2215),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2601),
.B(n_2135),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_SL g2845 ( 
.A(n_2623),
.B(n_2179),
.Y(n_2845)
);

INVx1_ASAP7_75t_SL g2846 ( 
.A(n_2630),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_2595),
.B(n_2305),
.Y(n_2847)
);

NOR2xp33_ASAP7_75t_L g2848 ( 
.A(n_2611),
.B(n_1819),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2762),
.Y(n_2849)
);

CKINVDCx5p33_ASAP7_75t_R g2850 ( 
.A(n_2476),
.Y(n_2850)
);

AO22x2_ASAP7_75t_L g2851 ( 
.A1(n_2549),
.A2(n_1874),
.B1(n_1897),
.B2(n_1822),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2597),
.Y(n_2852)
);

INVx4_ASAP7_75t_L g2853 ( 
.A(n_2538),
.Y(n_2853)
);

AND2x4_ASAP7_75t_L g2854 ( 
.A(n_2646),
.B(n_2224),
.Y(n_2854)
);

AND2x4_ASAP7_75t_L g2855 ( 
.A(n_2648),
.B(n_2225),
.Y(n_2855)
);

CKINVDCx5p33_ASAP7_75t_R g2856 ( 
.A(n_2475),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2768),
.Y(n_2857)
);

AND2x6_ASAP7_75t_L g2858 ( 
.A(n_2482),
.B(n_1524),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2597),
.Y(n_2859)
);

INVx3_ASAP7_75t_L g2860 ( 
.A(n_2473),
.Y(n_2860)
);

AOI22xp33_ASAP7_75t_L g2861 ( 
.A1(n_2482),
.A2(n_1595),
.B1(n_1652),
.B2(n_1588),
.Y(n_2861)
);

NOR2xp33_ASAP7_75t_L g2862 ( 
.A(n_2616),
.B(n_1923),
.Y(n_2862)
);

BUFx3_ASAP7_75t_L g2863 ( 
.A(n_2483),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2515),
.B(n_2136),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2494),
.Y(n_2865)
);

INVx3_ASAP7_75t_L g2866 ( 
.A(n_2495),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2683),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_SL g2868 ( 
.A(n_2653),
.B(n_2192),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2525),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_2528),
.B(n_2139),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2683),
.Y(n_2871)
);

HB1xp67_ASAP7_75t_L g2872 ( 
.A(n_2489),
.Y(n_2872)
);

AND2x4_ASAP7_75t_L g2873 ( 
.A(n_2650),
.B(n_2227),
.Y(n_2873)
);

BUFx3_ASAP7_75t_L g2874 ( 
.A(n_2539),
.Y(n_2874)
);

INVx2_ASAP7_75t_SL g2875 ( 
.A(n_2687),
.Y(n_2875)
);

BUFx3_ASAP7_75t_L g2876 ( 
.A(n_2555),
.Y(n_2876)
);

AOI22xp5_ASAP7_75t_L g2877 ( 
.A1(n_2780),
.A2(n_2251),
.B1(n_2196),
.B2(n_2208),
.Y(n_2877)
);

INVx2_ASAP7_75t_L g2878 ( 
.A(n_2693),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2532),
.Y(n_2879)
);

INVx2_ASAP7_75t_SL g2880 ( 
.A(n_2687),
.Y(n_2880)
);

INVx3_ASAP7_75t_L g2881 ( 
.A(n_2533),
.Y(n_2881)
);

NAND3xp33_ASAP7_75t_L g2882 ( 
.A(n_2677),
.B(n_1182),
.C(n_1179),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_SL g2883 ( 
.A(n_2690),
.B(n_2192),
.Y(n_2883)
);

NOR2xp33_ASAP7_75t_L g2884 ( 
.A(n_2692),
.B(n_1183),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2546),
.Y(n_2885)
);

OR2x6_ASAP7_75t_L g2886 ( 
.A(n_2697),
.B(n_1574),
.Y(n_2886)
);

AND2x2_ASAP7_75t_SL g2887 ( 
.A(n_2709),
.B(n_2718),
.Y(n_2887)
);

INVxp67_ASAP7_75t_L g2888 ( 
.A(n_2535),
.Y(n_2888)
);

INVx4_ASAP7_75t_L g2889 ( 
.A(n_2557),
.Y(n_2889)
);

BUFx3_ASAP7_75t_L g2890 ( 
.A(n_2537),
.Y(n_2890)
);

AND2x6_ASAP7_75t_L g2891 ( 
.A(n_2482),
.B(n_1574),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2614),
.B(n_2143),
.Y(n_2892)
);

AND2x6_ASAP7_75t_L g2893 ( 
.A(n_2562),
.B(n_1576),
.Y(n_2893)
);

OR2x2_ASAP7_75t_SL g2894 ( 
.A(n_2708),
.B(n_1576),
.Y(n_2894)
);

AOI22xp5_ASAP7_75t_L g2895 ( 
.A1(n_2723),
.A2(n_2211),
.B1(n_2223),
.B2(n_2185),
.Y(n_2895)
);

AOI22xp5_ASAP7_75t_L g2896 ( 
.A1(n_2660),
.A2(n_2249),
.B1(n_2237),
.B2(n_2172),
.Y(n_2896)
);

AND2x6_ASAP7_75t_L g2897 ( 
.A(n_2562),
.B(n_1604),
.Y(n_2897)
);

HB1xp67_ASAP7_75t_L g2898 ( 
.A(n_2634),
.Y(n_2898)
);

NAND3xp33_ASAP7_75t_L g2899 ( 
.A(n_2696),
.B(n_1187),
.C(n_1186),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2552),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2563),
.Y(n_2901)
);

AND2x2_ASAP7_75t_L g2902 ( 
.A(n_2636),
.B(n_1411),
.Y(n_2902)
);

AND2x2_ASAP7_75t_L g2903 ( 
.A(n_2740),
.B(n_1490),
.Y(n_2903)
);

OAI21xp33_ASAP7_75t_L g2904 ( 
.A1(n_2641),
.A2(n_2686),
.B(n_2684),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2698),
.B(n_2157),
.Y(n_2905)
);

BUFx6f_ASAP7_75t_L g2906 ( 
.A(n_2693),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2576),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2713),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2586),
.Y(n_2909)
);

AND2x4_ASAP7_75t_L g2910 ( 
.A(n_2658),
.B(n_2166),
.Y(n_2910)
);

AND2x2_ASAP7_75t_L g2911 ( 
.A(n_2700),
.B(n_1490),
.Y(n_2911)
);

NOR2xp33_ASAP7_75t_L g2912 ( 
.A(n_2702),
.B(n_1188),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2591),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2600),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2615),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_SL g2916 ( 
.A(n_2703),
.B(n_2193),
.Y(n_2916)
);

NOR2xp33_ASAP7_75t_L g2917 ( 
.A(n_2710),
.B(n_1191),
.Y(n_2917)
);

BUFx6f_ASAP7_75t_L g2918 ( 
.A(n_2713),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2712),
.B(n_2159),
.Y(n_2919)
);

NOR2xp33_ASAP7_75t_L g2920 ( 
.A(n_2719),
.B(n_1192),
.Y(n_2920)
);

AOI22xp33_ASAP7_75t_L g2921 ( 
.A1(n_2521),
.A2(n_1652),
.B1(n_1659),
.B2(n_1595),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2747),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2747),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2621),
.Y(n_2924)
);

BUFx3_ASAP7_75t_L g2925 ( 
.A(n_2590),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2626),
.Y(n_2926)
);

AND2x4_ASAP7_75t_L g2927 ( 
.A(n_2664),
.B(n_2164),
.Y(n_2927)
);

BUFx10_ASAP7_75t_L g2928 ( 
.A(n_2478),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2637),
.Y(n_2929)
);

OR2x2_ASAP7_75t_L g2930 ( 
.A(n_2673),
.B(n_1197),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2721),
.B(n_2329),
.Y(n_2931)
);

BUFx3_ASAP7_75t_L g2932 ( 
.A(n_2593),
.Y(n_2932)
);

INVx3_ASAP7_75t_L g2933 ( 
.A(n_2662),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2665),
.Y(n_2934)
);

BUFx10_ASAP7_75t_L g2935 ( 
.A(n_2531),
.Y(n_2935)
);

BUFx3_ASAP7_75t_L g2936 ( 
.A(n_2596),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2675),
.Y(n_2937)
);

BUFx3_ASAP7_75t_L g2938 ( 
.A(n_2599),
.Y(n_2938)
);

AOI22xp5_ASAP7_75t_L g2939 ( 
.A1(n_2663),
.A2(n_2340),
.B1(n_2353),
.B2(n_2334),
.Y(n_2939)
);

INVx3_ASAP7_75t_L g2940 ( 
.A(n_2680),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2757),
.Y(n_2941)
);

CKINVDCx5p33_ASAP7_75t_R g2942 ( 
.A(n_2488),
.Y(n_2942)
);

INVx5_ASAP7_75t_L g2943 ( 
.A(n_2655),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2682),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2722),
.B(n_2355),
.Y(n_2945)
);

AND2x2_ASAP7_75t_L g2946 ( 
.A(n_2724),
.B(n_1490),
.Y(n_2946)
);

AND2x2_ASAP7_75t_L g2947 ( 
.A(n_2735),
.B(n_2736),
.Y(n_2947)
);

BUFx6f_ASAP7_75t_L g2948 ( 
.A(n_2757),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2726),
.Y(n_2949)
);

AND2x6_ASAP7_75t_L g2950 ( 
.A(n_2562),
.B(n_1604),
.Y(n_2950)
);

AOI22xp33_ASAP7_75t_L g2951 ( 
.A1(n_2521),
.A2(n_1652),
.B1(n_1659),
.B2(n_1595),
.Y(n_2951)
);

CKINVDCx5p33_ASAP7_75t_R g2952 ( 
.A(n_2490),
.Y(n_2952)
);

AND2x6_ASAP7_75t_L g2953 ( 
.A(n_2620),
.B(n_1625),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2738),
.B(n_1518),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2744),
.Y(n_2955)
);

AOI22xp33_ASAP7_75t_L g2956 ( 
.A1(n_2620),
.A2(n_1652),
.B1(n_1659),
.B2(n_1595),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2763),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2764),
.Y(n_2958)
);

AND2x4_ASAP7_75t_L g2959 ( 
.A(n_2672),
.B(n_2363),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2773),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2775),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2681),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2620),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2742),
.B(n_2367),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2695),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2685),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2699),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2701),
.Y(n_2968)
);

INVx2_ASAP7_75t_SL g2969 ( 
.A(n_2766),
.Y(n_2969)
);

INVx3_ASAP7_75t_L g2970 ( 
.A(n_2602),
.Y(n_2970)
);

BUFx4f_ASAP7_75t_L g2971 ( 
.A(n_2769),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2743),
.B(n_2373),
.Y(n_2972)
);

NOR2xp33_ASAP7_75t_L g2973 ( 
.A(n_2746),
.B(n_1199),
.Y(n_2973)
);

INVx1_ASAP7_75t_SL g2974 ( 
.A(n_2725),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2624),
.Y(n_2975)
);

AND2x2_ASAP7_75t_L g2976 ( 
.A(n_2749),
.B(n_1518),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_2695),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2667),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2717),
.Y(n_2979)
);

BUFx3_ASAP7_75t_L g2980 ( 
.A(n_2606),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2695),
.Y(n_2981)
);

BUFx3_ASAP7_75t_L g2982 ( 
.A(n_2607),
.Y(n_2982)
);

AND2x2_ASAP7_75t_L g2983 ( 
.A(n_2594),
.B(n_1518),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2575),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2605),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2715),
.B(n_2408),
.Y(n_2986)
);

BUFx6f_ASAP7_75t_L g2987 ( 
.A(n_2500),
.Y(n_2987)
);

AND2x4_ASAP7_75t_L g2988 ( 
.A(n_2474),
.B(n_2418),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2727),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2737),
.B(n_2422),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_2581),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2739),
.Y(n_2992)
);

BUFx3_ASAP7_75t_L g2993 ( 
.A(n_2609),
.Y(n_2993)
);

NAND3xp33_ASAP7_75t_L g2994 ( 
.A(n_2774),
.B(n_1202),
.C(n_1200),
.Y(n_2994)
);

BUFx3_ASAP7_75t_L g2995 ( 
.A(n_2548),
.Y(n_2995)
);

BUFx6f_ASAP7_75t_L g2996 ( 
.A(n_2500),
.Y(n_2996)
);

INVxp67_ASAP7_75t_L g2997 ( 
.A(n_2750),
.Y(n_2997)
);

BUFx3_ASAP7_75t_L g2998 ( 
.A(n_2560),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2511),
.B(n_2424),
.Y(n_2999)
);

AOI22xp33_ASAP7_75t_L g3000 ( 
.A1(n_2610),
.A2(n_1726),
.B1(n_1761),
.B2(n_1659),
.Y(n_3000)
);

INVxp67_ASAP7_75t_SL g3001 ( 
.A(n_2598),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2604),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2754),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2619),
.Y(n_3004)
);

NOR2xp33_ASAP7_75t_L g3005 ( 
.A(n_2594),
.B(n_1205),
.Y(n_3005)
);

INVx3_ASAP7_75t_L g3006 ( 
.A(n_2545),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2612),
.B(n_2434),
.Y(n_3007)
);

BUFx2_ASAP7_75t_L g3008 ( 
.A(n_2728),
.Y(n_3008)
);

INVx8_ASAP7_75t_L g3009 ( 
.A(n_2691),
.Y(n_3009)
);

AND2x2_ASAP7_75t_L g3010 ( 
.A(n_2752),
.B(n_1586),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_SL g3011 ( 
.A(n_2753),
.B(n_2193),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2619),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2618),
.Y(n_3013)
);

AND2x6_ASAP7_75t_L g3014 ( 
.A(n_2625),
.B(n_1625),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2633),
.Y(n_3015)
);

NOR2xp33_ASAP7_75t_L g3016 ( 
.A(n_2550),
.B(n_1208),
.Y(n_3016)
);

INVx4_ASAP7_75t_L g3017 ( 
.A(n_2487),
.Y(n_3017)
);

AND2x6_ASAP7_75t_L g3018 ( 
.A(n_2644),
.B(n_1640),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2729),
.Y(n_3019)
);

AND2x4_ASAP7_75t_L g3020 ( 
.A(n_2558),
.B(n_2669),
.Y(n_3020)
);

NAND2x1_ASAP7_75t_L g3021 ( 
.A(n_2730),
.B(n_2437),
.Y(n_3021)
);

NAND3xp33_ASAP7_75t_L g3022 ( 
.A(n_2629),
.B(n_1211),
.C(n_1209),
.Y(n_3022)
);

INVx3_ASAP7_75t_L g3023 ( 
.A(n_2689),
.Y(n_3023)
);

AND2x2_ASAP7_75t_L g3024 ( 
.A(n_2498),
.B(n_1586),
.Y(n_3024)
);

AND2x4_ASAP7_75t_L g3025 ( 
.A(n_2588),
.B(n_2453),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2584),
.Y(n_3026)
);

HB1xp67_ASAP7_75t_L g3027 ( 
.A(n_2767),
.Y(n_3027)
);

HB1xp67_ASAP7_75t_L g3028 ( 
.A(n_2759),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2836),
.B(n_2817),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_SL g3030 ( 
.A(n_2971),
.B(n_2499),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_2813),
.Y(n_3031)
);

BUFx6f_ASAP7_75t_L g3032 ( 
.A(n_2987),
.Y(n_3032)
);

NAND3xp33_ASAP7_75t_L g3033 ( 
.A(n_2842),
.B(n_2688),
.C(n_2770),
.Y(n_3033)
);

AND2x4_ASAP7_75t_L g3034 ( 
.A(n_2830),
.B(n_2485),
.Y(n_3034)
);

O2A1O1Ixp33_ASAP7_75t_L g3035 ( 
.A1(n_2784),
.A2(n_2732),
.B(n_2771),
.C(n_2502),
.Y(n_3035)
);

AOI21xp5_ASAP7_75t_L g3036 ( 
.A1(n_2798),
.A2(n_2731),
.B(n_2661),
.Y(n_3036)
);

INVx3_ASAP7_75t_L g3037 ( 
.A(n_2833),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2847),
.B(n_2493),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_SL g3039 ( 
.A(n_2904),
.B(n_2501),
.Y(n_3039)
);

AOI22xp33_ASAP7_75t_L g3040 ( 
.A1(n_2975),
.A2(n_2638),
.B1(n_2632),
.B2(n_2666),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2821),
.Y(n_3041)
);

OR2x2_ASAP7_75t_L g3042 ( 
.A(n_2974),
.B(n_2505),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_SL g3043 ( 
.A(n_2947),
.B(n_2506),
.Y(n_3043)
);

NOR2xp33_ASAP7_75t_L g3044 ( 
.A(n_2829),
.B(n_2642),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2782),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2835),
.Y(n_3046)
);

NAND3xp33_ASAP7_75t_L g3047 ( 
.A(n_2848),
.B(n_2608),
.C(n_2554),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2790),
.Y(n_3048)
);

OR2x6_ASAP7_75t_L g3049 ( 
.A(n_3009),
.B(n_2714),
.Y(n_3049)
);

A2O1A1Ixp33_ASAP7_75t_L g3050 ( 
.A1(n_2862),
.A2(n_2617),
.B(n_2679),
.C(n_2674),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2783),
.B(n_2694),
.Y(n_3051)
);

AOI22xp5_ASAP7_75t_L g3052 ( 
.A1(n_2888),
.A2(n_2716),
.B1(n_2720),
.B2(n_2622),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2795),
.Y(n_3053)
);

INVx3_ASAP7_75t_L g3054 ( 
.A(n_2831),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_L g3055 ( 
.A(n_2791),
.B(n_2553),
.Y(n_3055)
);

INVx2_ASAP7_75t_L g3056 ( 
.A(n_2849),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2803),
.Y(n_3057)
);

NOR2xp33_ASAP7_75t_L g3058 ( 
.A(n_2884),
.B(n_2507),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_2978),
.B(n_2491),
.Y(n_3059)
);

NOR2xp33_ASAP7_75t_L g3060 ( 
.A(n_2912),
.B(n_2508),
.Y(n_3060)
);

INVx2_ASAP7_75t_L g3061 ( 
.A(n_2857),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_2807),
.Y(n_3062)
);

NOR3xp33_ASAP7_75t_L g3063 ( 
.A(n_2917),
.B(n_2758),
.C(n_2756),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2808),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2814),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2815),
.Y(n_3066)
);

INVx2_ASAP7_75t_SL g3067 ( 
.A(n_2872),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_2816),
.Y(n_3068)
);

INVxp67_ASAP7_75t_L g3069 ( 
.A(n_2911),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_SL g3070 ( 
.A(n_2942),
.B(n_2509),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_SL g3071 ( 
.A(n_2952),
.B(n_2512),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_SL g3072 ( 
.A(n_2987),
.B(n_2513),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2979),
.B(n_2751),
.Y(n_3073)
);

OAI22xp5_ASAP7_75t_L g3074 ( 
.A1(n_2824),
.A2(n_2643),
.B1(n_2541),
.B2(n_2542),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2844),
.B(n_2986),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2820),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_2990),
.B(n_2503),
.Y(n_3077)
);

AND2x6_ASAP7_75t_SL g3078 ( 
.A(n_3019),
.B(n_3005),
.Y(n_3078)
);

AOI21xp5_ASAP7_75t_L g3079 ( 
.A1(n_2800),
.A2(n_2761),
.B(n_2760),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_SL g3080 ( 
.A(n_2996),
.B(n_2825),
.Y(n_3080)
);

NOR2xp33_ASAP7_75t_L g3081 ( 
.A(n_2920),
.B(n_2540),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2838),
.B(n_2765),
.Y(n_3082)
);

NOR2xp33_ASAP7_75t_L g3083 ( 
.A(n_2973),
.B(n_2547),
.Y(n_3083)
);

INVx2_ASAP7_75t_SL g3084 ( 
.A(n_2898),
.Y(n_3084)
);

INVx2_ASAP7_75t_SL g3085 ( 
.A(n_3025),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2822),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2828),
.Y(n_3087)
);

INVx2_ASAP7_75t_L g3088 ( 
.A(n_2781),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2946),
.B(n_2651),
.Y(n_3089)
);

INVx2_ASAP7_75t_SL g3090 ( 
.A(n_2886),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2794),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2818),
.B(n_2905),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2796),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2919),
.B(n_2652),
.Y(n_3094)
);

OAI22xp5_ASAP7_75t_L g3095 ( 
.A1(n_3026),
.A2(n_2656),
.B1(n_2657),
.B2(n_2654),
.Y(n_3095)
);

CKINVDCx5p33_ASAP7_75t_R g3096 ( 
.A(n_2850),
.Y(n_3096)
);

NAND2xp5_ASAP7_75t_SL g3097 ( 
.A(n_2996),
.B(n_2659),
.Y(n_3097)
);

BUFx3_ASAP7_75t_L g3098 ( 
.A(n_2874),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2931),
.B(n_2520),
.Y(n_3099)
);

INVx8_ASAP7_75t_L g3100 ( 
.A(n_3009),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_2945),
.B(n_2524),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2964),
.B(n_2529),
.Y(n_3102)
);

NAND3xp33_ASAP7_75t_L g3103 ( 
.A(n_3016),
.B(n_2670),
.C(n_2628),
.Y(n_3103)
);

INVx2_ASAP7_75t_SL g3104 ( 
.A(n_2886),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2972),
.B(n_2530),
.Y(n_3105)
);

AND2x2_ASAP7_75t_L g3106 ( 
.A(n_2954),
.B(n_2569),
.Y(n_3106)
);

A2O1A1Ixp33_ASAP7_75t_L g3107 ( 
.A1(n_2792),
.A2(n_2627),
.B(n_2573),
.C(n_1168),
.Y(n_3107)
);

AOI22xp5_ASAP7_75t_L g3108 ( 
.A1(n_2812),
.A2(n_2691),
.B1(n_2561),
.B2(n_2647),
.Y(n_3108)
);

OAI22xp33_ASAP7_75t_L g3109 ( 
.A1(n_2841),
.A2(n_2496),
.B1(n_2479),
.B2(n_2486),
.Y(n_3109)
);

BUFx3_ASAP7_75t_L g3110 ( 
.A(n_2788),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_2963),
.B(n_2466),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2965),
.B(n_2247),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2805),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_SL g3114 ( 
.A(n_2970),
.B(n_2480),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_SL g3115 ( 
.A(n_2802),
.B(n_2733),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_SL g3116 ( 
.A(n_2976),
.B(n_2209),
.Y(n_3116)
);

HB1xp67_ASAP7_75t_L g3117 ( 
.A(n_2989),
.Y(n_3117)
);

AOI22xp5_ASAP7_75t_L g3118 ( 
.A1(n_2812),
.A2(n_2858),
.B1(n_2891),
.B2(n_2893),
.Y(n_3118)
);

AOI22xp33_ASAP7_75t_L g3119 ( 
.A1(n_2812),
.A2(n_2603),
.B1(n_1761),
.B2(n_1788),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2977),
.B(n_2250),
.Y(n_3120)
);

O2A1O1Ixp33_ASAP7_75t_L g3121 ( 
.A1(n_3000),
.A2(n_1669),
.B(n_1701),
.C(n_1640),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2981),
.B(n_2209),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_SL g3123 ( 
.A(n_2804),
.B(n_2212),
.Y(n_3123)
);

NOR2xp33_ASAP7_75t_L g3124 ( 
.A(n_2997),
.B(n_2983),
.Y(n_3124)
);

INVx2_ASAP7_75t_L g3125 ( 
.A(n_2806),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2927),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_3007),
.Y(n_3127)
);

A2O1A1Ixp33_ASAP7_75t_L g3128 ( 
.A1(n_2882),
.A2(n_1171),
.B(n_1174),
.C(n_1167),
.Y(n_3128)
);

AOI22xp33_ASAP7_75t_L g3129 ( 
.A1(n_2858),
.A2(n_1761),
.B1(n_1788),
.B2(n_1726),
.Y(n_3129)
);

INVx1_ASAP7_75t_SL g3130 ( 
.A(n_2846),
.Y(n_3130)
);

INVx2_ASAP7_75t_SL g3131 ( 
.A(n_2831),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_SL g3132 ( 
.A(n_2889),
.B(n_2840),
.Y(n_3132)
);

AOI22xp33_ASAP7_75t_L g3133 ( 
.A1(n_2858),
.A2(n_1761),
.B1(n_1788),
.B2(n_1726),
.Y(n_3133)
);

INVx2_ASAP7_75t_L g3134 ( 
.A(n_2959),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_2988),
.B(n_2212),
.Y(n_3135)
);

BUFx6f_ASAP7_75t_L g3136 ( 
.A(n_2906),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2910),
.Y(n_3137)
);

INVxp67_ASAP7_75t_SL g3138 ( 
.A(n_2786),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_SL g3139 ( 
.A(n_3024),
.B(n_3006),
.Y(n_3139)
);

AOI22xp5_ASAP7_75t_L g3140 ( 
.A1(n_2891),
.A2(n_2235),
.B1(n_2245),
.B2(n_2234),
.Y(n_3140)
);

OR2x2_ASAP7_75t_L g3141 ( 
.A(n_3008),
.B(n_2635),
.Y(n_3141)
);

AOI22xp33_ASAP7_75t_L g3142 ( 
.A1(n_2891),
.A2(n_2897),
.B1(n_2950),
.B2(n_2893),
.Y(n_3142)
);

OR2x2_ASAP7_75t_L g3143 ( 
.A(n_2809),
.B(n_2640),
.Y(n_3143)
);

NOR2xp67_ASAP7_75t_L g3144 ( 
.A(n_2853),
.B(n_3017),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2893),
.B(n_2234),
.Y(n_3145)
);

NOR3xp33_ASAP7_75t_L g3146 ( 
.A(n_3022),
.B(n_2649),
.C(n_2645),
.Y(n_3146)
);

NOR2xp33_ASAP7_75t_L g3147 ( 
.A(n_2930),
.B(n_1302),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_SL g3148 ( 
.A(n_2925),
.B(n_2235),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_2949),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_2955),
.Y(n_3150)
);

NOR2xp33_ASAP7_75t_L g3151 ( 
.A(n_2992),
.B(n_1330),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2962),
.Y(n_3152)
);

CKINVDCx20_ASAP7_75t_R g3153 ( 
.A(n_2856),
.Y(n_3153)
);

AOI22xp33_ASAP7_75t_L g3154 ( 
.A1(n_2897),
.A2(n_1788),
.B1(n_1834),
.B2(n_1726),
.Y(n_3154)
);

AND2x4_ASAP7_75t_L g3155 ( 
.A(n_2890),
.B(n_2823),
.Y(n_3155)
);

AND2x2_ASAP7_75t_L g3156 ( 
.A(n_2902),
.B(n_1586),
.Y(n_3156)
);

AND2x2_ASAP7_75t_L g3157 ( 
.A(n_2903),
.B(n_1637),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_2897),
.B(n_2245),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_2966),
.Y(n_3159)
);

OAI21xp5_ASAP7_75t_L g3160 ( 
.A1(n_2793),
.A2(n_1184),
.B(n_1177),
.Y(n_3160)
);

AOI22xp5_ASAP7_75t_L g3161 ( 
.A1(n_2950),
.A2(n_2953),
.B1(n_2843),
.B2(n_3004),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2950),
.B(n_2252),
.Y(n_3162)
);

INVxp67_ASAP7_75t_SL g3163 ( 
.A(n_2906),
.Y(n_3163)
);

AOI21xp5_ASAP7_75t_L g3164 ( 
.A1(n_2864),
.A2(n_2252),
.B(n_1195),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_SL g3165 ( 
.A(n_2932),
.B(n_2534),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2953),
.B(n_1834),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2960),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_2984),
.Y(n_3168)
);

AND2x4_ASAP7_75t_SL g3169 ( 
.A(n_2928),
.B(n_3023),
.Y(n_3169)
);

INVx2_ASAP7_75t_L g3170 ( 
.A(n_2991),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_2953),
.B(n_1834),
.Y(n_3171)
);

NOR2xp33_ASAP7_75t_L g3172 ( 
.A(n_3003),
.B(n_1391),
.Y(n_3172)
);

OAI22xp5_ASAP7_75t_L g3173 ( 
.A1(n_2921),
.A2(n_1400),
.B1(n_1401),
.B2(n_1391),
.Y(n_3173)
);

INVx4_ASAP7_75t_L g3174 ( 
.A(n_2876),
.Y(n_3174)
);

O2A1O1Ixp33_ASAP7_75t_L g3175 ( 
.A1(n_2845),
.A2(n_1701),
.B(n_1856),
.C(n_1669),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2967),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2999),
.B(n_1834),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_SL g3178 ( 
.A(n_2936),
.B(n_1400),
.Y(n_3178)
);

OR2x6_ASAP7_75t_L g3179 ( 
.A(n_2969),
.B(n_1856),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_L g3180 ( 
.A(n_2899),
.B(n_1401),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2968),
.Y(n_3181)
);

INVx3_ASAP7_75t_L g3182 ( 
.A(n_2918),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_3013),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2951),
.B(n_1868),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_3001),
.B(n_1868),
.Y(n_3185)
);

INVx2_ASAP7_75t_SL g3186 ( 
.A(n_2918),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_3015),
.Y(n_3187)
);

NOR2xp33_ASAP7_75t_SL g3188 ( 
.A(n_2789),
.B(n_2943),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2870),
.B(n_1868),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_3002),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_L g3191 ( 
.A(n_2834),
.B(n_1868),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_SL g3192 ( 
.A(n_2938),
.B(n_1432),
.Y(n_3192)
);

INVx3_ASAP7_75t_L g3193 ( 
.A(n_2948),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_2892),
.B(n_1213),
.Y(n_3194)
);

AOI22xp33_ASAP7_75t_L g3195 ( 
.A1(n_2994),
.A2(n_1451),
.B1(n_1461),
.B2(n_1432),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_2785),
.B(n_1218),
.Y(n_3196)
);

INVx3_ASAP7_75t_L g3197 ( 
.A(n_2948),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2797),
.B(n_1220),
.Y(n_3198)
);

NOR3xp33_ASAP7_75t_L g3199 ( 
.A(n_2868),
.B(n_1225),
.C(n_1223),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2799),
.B(n_1227),
.Y(n_3200)
);

INVxp33_ASAP7_75t_L g3201 ( 
.A(n_3010),
.Y(n_3201)
);

INVxp33_ASAP7_75t_L g3202 ( 
.A(n_3027),
.Y(n_3202)
);

NAND2xp33_ASAP7_75t_L g3203 ( 
.A(n_3014),
.B(n_1229),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_2837),
.Y(n_3204)
);

INVx2_ASAP7_75t_L g3205 ( 
.A(n_2852),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_2801),
.B(n_1231),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_3012),
.B(n_1233),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_2980),
.B(n_1637),
.Y(n_3208)
);

OAI22xp33_ASAP7_75t_L g3209 ( 
.A1(n_2982),
.A2(n_1461),
.B1(n_1523),
.B2(n_1451),
.Y(n_3209)
);

NOR2xp33_ASAP7_75t_SL g3210 ( 
.A(n_2943),
.B(n_1523),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_SL g3211 ( 
.A(n_2993),
.B(n_1539),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2854),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2855),
.Y(n_3213)
);

OAI22xp5_ASAP7_75t_L g3214 ( 
.A1(n_2861),
.A2(n_1550),
.B1(n_1594),
.B2(n_1539),
.Y(n_3214)
);

OAI22xp33_ASAP7_75t_L g3215 ( 
.A1(n_2877),
.A2(n_1594),
.B1(n_1599),
.B2(n_1550),
.Y(n_3215)
);

OAI22xp5_ASAP7_75t_SL g3216 ( 
.A1(n_2887),
.A2(n_1603),
.B1(n_1631),
.B2(n_1599),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_2939),
.B(n_1234),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_SL g3218 ( 
.A(n_2985),
.B(n_2896),
.Y(n_3218)
);

INVx8_ASAP7_75t_L g3219 ( 
.A(n_3014),
.Y(n_3219)
);

INVx3_ASAP7_75t_L g3220 ( 
.A(n_2826),
.Y(n_3220)
);

NAND2xp33_ASAP7_75t_L g3221 ( 
.A(n_3014),
.B(n_3018),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_2859),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2787),
.B(n_1236),
.Y(n_3223)
);

BUFx3_ASAP7_75t_L g3224 ( 
.A(n_2863),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_2956),
.B(n_1237),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2873),
.Y(n_3226)
);

NAND3xp33_ASAP7_75t_L g3227 ( 
.A(n_2895),
.B(n_2916),
.C(n_2883),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2865),
.Y(n_3228)
);

AND2x2_ASAP7_75t_SL g3229 ( 
.A(n_2839),
.B(n_1859),
.Y(n_3229)
);

NOR2xp33_ASAP7_75t_L g3230 ( 
.A(n_2819),
.B(n_1603),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_2867),
.Y(n_3231)
);

AND2x2_ASAP7_75t_L g3232 ( 
.A(n_3044),
.B(n_2827),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_SL g3233 ( 
.A(n_3038),
.B(n_3028),
.Y(n_3233)
);

NOR2xp33_ASAP7_75t_L g3234 ( 
.A(n_3092),
.B(n_2995),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_3075),
.B(n_2871),
.Y(n_3235)
);

AOI21xp33_ASAP7_75t_L g3236 ( 
.A1(n_3081),
.A2(n_2851),
.B(n_2811),
.Y(n_3236)
);

NOR2xp33_ASAP7_75t_L g3237 ( 
.A(n_3083),
.B(n_3051),
.Y(n_3237)
);

OAI22xp5_ASAP7_75t_L g3238 ( 
.A1(n_3029),
.A2(n_2894),
.B1(n_2875),
.B2(n_2880),
.Y(n_3238)
);

NOR2xp33_ASAP7_75t_SL g3239 ( 
.A(n_3096),
.B(n_2935),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3056),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_3077),
.B(n_2878),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_3127),
.B(n_2908),
.Y(n_3242)
);

AND2x2_ASAP7_75t_L g3243 ( 
.A(n_3058),
.B(n_2998),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_3055),
.B(n_2922),
.Y(n_3244)
);

BUFx6f_ASAP7_75t_L g3245 ( 
.A(n_3136),
.Y(n_3245)
);

AND2x2_ASAP7_75t_L g3246 ( 
.A(n_3060),
.B(n_2810),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_3059),
.B(n_3061),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_3073),
.B(n_2923),
.Y(n_3248)
);

AOI21xp5_ASAP7_75t_L g3249 ( 
.A1(n_3036),
.A2(n_3021),
.B(n_3011),
.Y(n_3249)
);

INVx2_ASAP7_75t_L g3250 ( 
.A(n_3062),
.Y(n_3250)
);

OAI21xp5_ASAP7_75t_L g3251 ( 
.A1(n_3223),
.A2(n_2879),
.B(n_2869),
.Y(n_3251)
);

NOR2xp33_ASAP7_75t_L g3252 ( 
.A(n_3033),
.B(n_2885),
.Y(n_3252)
);

INVx3_ASAP7_75t_L g3253 ( 
.A(n_3098),
.Y(n_3253)
);

AOI21xp5_ASAP7_75t_L g3254 ( 
.A1(n_3135),
.A2(n_2941),
.B(n_2901),
.Y(n_3254)
);

AND2x4_ASAP7_75t_L g3255 ( 
.A(n_3110),
.B(n_3020),
.Y(n_3255)
);

AOI21xp5_ASAP7_75t_L g3256 ( 
.A1(n_3221),
.A2(n_2907),
.B(n_2900),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_3045),
.B(n_2909),
.Y(n_3257)
);

BUFx2_ASAP7_75t_L g3258 ( 
.A(n_3067),
.Y(n_3258)
);

A2O1A1Ixp33_ASAP7_75t_L g3259 ( 
.A1(n_3035),
.A2(n_2914),
.B(n_2915),
.C(n_2913),
.Y(n_3259)
);

AOI21xp5_ASAP7_75t_L g3260 ( 
.A1(n_3111),
.A2(n_2926),
.B(n_2924),
.Y(n_3260)
);

NOR2xp33_ASAP7_75t_L g3261 ( 
.A(n_3094),
.B(n_2929),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_SL g3262 ( 
.A(n_3082),
.B(n_2860),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_3048),
.B(n_2934),
.Y(n_3263)
);

AOI21xp5_ASAP7_75t_L g3264 ( 
.A1(n_3177),
.A2(n_2944),
.B(n_2937),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_L g3265 ( 
.A(n_3053),
.B(n_2957),
.Y(n_3265)
);

AOI21xp5_ASAP7_75t_L g3266 ( 
.A1(n_3122),
.A2(n_2961),
.B(n_2958),
.Y(n_3266)
);

AOI21xp5_ASAP7_75t_L g3267 ( 
.A1(n_3218),
.A2(n_2881),
.B(n_2866),
.Y(n_3267)
);

OAI22xp5_ASAP7_75t_L g3268 ( 
.A1(n_3040),
.A2(n_2940),
.B1(n_2933),
.B2(n_1643),
.Y(n_3268)
);

NAND2x1_ASAP7_75t_L g3269 ( 
.A(n_3136),
.B(n_3204),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_3068),
.Y(n_3270)
);

NAND3xp33_ASAP7_75t_L g3271 ( 
.A(n_3180),
.B(n_1241),
.C(n_1240),
.Y(n_3271)
);

AOI21xp5_ASAP7_75t_L g3272 ( 
.A1(n_3112),
.A2(n_1203),
.B(n_1190),
.Y(n_3272)
);

OAI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_3184),
.A2(n_3018),
.B(n_1215),
.Y(n_3273)
);

AOI21xp5_ASAP7_75t_L g3274 ( 
.A1(n_3120),
.A2(n_1221),
.B(n_1207),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_3057),
.B(n_3018),
.Y(n_3275)
);

NAND3xp33_ASAP7_75t_L g3276 ( 
.A(n_3047),
.B(n_1247),
.C(n_1244),
.Y(n_3276)
);

INVx2_ASAP7_75t_L g3277 ( 
.A(n_3086),
.Y(n_3277)
);

AOI21xp5_ASAP7_75t_L g3278 ( 
.A1(n_3138),
.A2(n_1232),
.B(n_1224),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_3064),
.B(n_2832),
.Y(n_3279)
);

NOR2x1_ASAP7_75t_R g3280 ( 
.A(n_3174),
.B(n_1248),
.Y(n_3280)
);

AOI21xp5_ASAP7_75t_L g3281 ( 
.A1(n_3194),
.A2(n_1238),
.B(n_1235),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_L g3282 ( 
.A(n_3065),
.B(n_1249),
.Y(n_3282)
);

OAI21xp5_ASAP7_75t_L g3283 ( 
.A1(n_3189),
.A2(n_1242),
.B(n_1239),
.Y(n_3283)
);

AOI21xp5_ASAP7_75t_L g3284 ( 
.A1(n_3079),
.A2(n_1256),
.B(n_1243),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_3066),
.B(n_1251),
.Y(n_3285)
);

AOI21xp5_ASAP7_75t_L g3286 ( 
.A1(n_3099),
.A2(n_1263),
.B(n_1262),
.Y(n_3286)
);

AOI22xp5_ASAP7_75t_L g3287 ( 
.A1(n_3227),
.A2(n_1643),
.B1(n_1644),
.B2(n_1631),
.Y(n_3287)
);

AOI21xp5_ASAP7_75t_L g3288 ( 
.A1(n_3101),
.A2(n_1268),
.B(n_1267),
.Y(n_3288)
);

A2O1A1Ixp33_ASAP7_75t_L g3289 ( 
.A1(n_3147),
.A2(n_1282),
.B(n_1285),
.C(n_1278),
.Y(n_3289)
);

NOR2xp33_ASAP7_75t_L g3290 ( 
.A(n_3074),
.B(n_1644),
.Y(n_3290)
);

NOR2xp33_ASAP7_75t_L g3291 ( 
.A(n_3201),
.B(n_1646),
.Y(n_3291)
);

A2O1A1Ixp33_ASAP7_75t_L g3292 ( 
.A1(n_3161),
.A2(n_3124),
.B(n_3119),
.C(n_3087),
.Y(n_3292)
);

INVx3_ASAP7_75t_L g3293 ( 
.A(n_3032),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3076),
.B(n_3031),
.Y(n_3294)
);

AOI33xp33_ASAP7_75t_L g3295 ( 
.A1(n_3195),
.A2(n_1292),
.A3(n_1287),
.B1(n_1307),
.B2(n_1290),
.B3(n_1286),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_3041),
.B(n_1252),
.Y(n_3296)
);

AOI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_3102),
.A2(n_1313),
.B(n_1310),
.Y(n_3297)
);

A2O1A1Ixp33_ASAP7_75t_L g3298 ( 
.A1(n_3160),
.A2(n_1316),
.B(n_1317),
.C(n_1314),
.Y(n_3298)
);

AOI21xp5_ASAP7_75t_L g3299 ( 
.A1(n_3105),
.A2(n_3132),
.B(n_3116),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_SL g3300 ( 
.A(n_3144),
.B(n_3037),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_SL g3301 ( 
.A(n_3069),
.B(n_1646),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_3046),
.B(n_1254),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_3093),
.B(n_1257),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_SL g3304 ( 
.A(n_3084),
.B(n_1647),
.Y(n_3304)
);

AOI21xp5_ASAP7_75t_L g3305 ( 
.A1(n_3145),
.A2(n_1324),
.B(n_1318),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_3088),
.B(n_1259),
.Y(n_3306)
);

AOI21xp5_ASAP7_75t_L g3307 ( 
.A1(n_3158),
.A2(n_1339),
.B(n_1333),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_3091),
.B(n_1264),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3113),
.B(n_1265),
.Y(n_3309)
);

INVx3_ASAP7_75t_L g3310 ( 
.A(n_3032),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3125),
.B(n_1266),
.Y(n_3311)
);

NOR2xp33_ASAP7_75t_L g3312 ( 
.A(n_3050),
.B(n_1647),
.Y(n_3312)
);

AOI21xp5_ASAP7_75t_L g3313 ( 
.A1(n_3162),
.A2(n_1359),
.B(n_1343),
.Y(n_3313)
);

AOI21xp5_ASAP7_75t_L g3314 ( 
.A1(n_3142),
.A2(n_3185),
.B(n_3207),
.Y(n_3314)
);

AOI21xp5_ASAP7_75t_L g3315 ( 
.A1(n_3080),
.A2(n_3118),
.B(n_3139),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3152),
.B(n_1272),
.Y(n_3316)
);

BUFx3_ASAP7_75t_L g3317 ( 
.A(n_3100),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_SL g3318 ( 
.A(n_3103),
.B(n_1666),
.Y(n_3318)
);

NOR2x1_ASAP7_75t_L g3319 ( 
.A(n_3153),
.B(n_1666),
.Y(n_3319)
);

HB1xp67_ASAP7_75t_L g3320 ( 
.A(n_3117),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_3159),
.B(n_1276),
.Y(n_3321)
);

AOI21xp33_ASAP7_75t_L g3322 ( 
.A1(n_3215),
.A2(n_1694),
.B(n_1684),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_3176),
.B(n_1280),
.Y(n_3323)
);

NOR2xp33_ASAP7_75t_L g3324 ( 
.A(n_3230),
.B(n_1684),
.Y(n_3324)
);

AO21x1_ASAP7_75t_L g3325 ( 
.A1(n_3166),
.A2(n_1363),
.B(n_1361),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3181),
.Y(n_3326)
);

AOI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_3171),
.A2(n_1373),
.B(n_1370),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3183),
.B(n_1283),
.Y(n_3328)
);

INVx3_ASAP7_75t_L g3329 ( 
.A(n_3155),
.Y(n_3329)
);

AOI21xp5_ASAP7_75t_L g3330 ( 
.A1(n_3196),
.A2(n_1379),
.B(n_1375),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_SL g3331 ( 
.A(n_3085),
.B(n_1694),
.Y(n_3331)
);

NOR3xp33_ASAP7_75t_L g3332 ( 
.A(n_3173),
.B(n_3192),
.C(n_3178),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_3187),
.B(n_1291),
.Y(n_3333)
);

OAI21xp5_ASAP7_75t_L g3334 ( 
.A1(n_3217),
.A2(n_1384),
.B(n_1383),
.Y(n_3334)
);

AOI21x1_ASAP7_75t_L g3335 ( 
.A1(n_3191),
.A2(n_1388),
.B(n_1386),
.Y(n_3335)
);

AOI222xp33_ASAP7_75t_L g3336 ( 
.A1(n_3216),
.A2(n_1848),
.B1(n_1713),
.B2(n_1747),
.C1(n_1787),
.C2(n_1774),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_3156),
.B(n_1294),
.Y(n_3337)
);

OAI321xp33_ASAP7_75t_L g3338 ( 
.A1(n_3214),
.A2(n_1406),
.A3(n_1399),
.B1(n_1409),
.B2(n_1404),
.C(n_1393),
.Y(n_3338)
);

AOI21xp5_ASAP7_75t_L g3339 ( 
.A1(n_3198),
.A2(n_1418),
.B(n_1415),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3228),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_3157),
.B(n_3168),
.Y(n_3341)
);

O2A1O1Ixp33_ASAP7_75t_L g3342 ( 
.A1(n_3107),
.A2(n_1429),
.B(n_1435),
.C(n_1424),
.Y(n_3342)
);

NOR2xp33_ASAP7_75t_SL g3343 ( 
.A(n_3188),
.B(n_1713),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_3170),
.B(n_1295),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_3190),
.B(n_1296),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_3149),
.B(n_1297),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3150),
.Y(n_3347)
);

NOR2xp33_ASAP7_75t_L g3348 ( 
.A(n_3130),
.B(n_1727),
.Y(n_3348)
);

AOI21xp5_ASAP7_75t_L g3349 ( 
.A1(n_3200),
.A2(n_1440),
.B(n_1439),
.Y(n_3349)
);

INVx3_ASAP7_75t_L g3350 ( 
.A(n_3136),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_3167),
.B(n_1298),
.Y(n_3351)
);

NOR2xp33_ASAP7_75t_L g3352 ( 
.A(n_3202),
.B(n_1727),
.Y(n_3352)
);

AOI21xp5_ASAP7_75t_L g3353 ( 
.A1(n_3206),
.A2(n_1445),
.B(n_1443),
.Y(n_3353)
);

INVx4_ASAP7_75t_L g3354 ( 
.A(n_3100),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3205),
.B(n_1300),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3222),
.B(n_1303),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3231),
.Y(n_3357)
);

NOR2xp33_ASAP7_75t_L g3358 ( 
.A(n_3151),
.B(n_1747),
.Y(n_3358)
);

O2A1O1Ixp33_ASAP7_75t_L g3359 ( 
.A1(n_3128),
.A2(n_1463),
.B(n_1466),
.C(n_1462),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3137),
.Y(n_3360)
);

INVx2_ASAP7_75t_L g3361 ( 
.A(n_3126),
.Y(n_3361)
);

INVx2_ASAP7_75t_L g3362 ( 
.A(n_3134),
.Y(n_3362)
);

AND2x4_ASAP7_75t_L g3363 ( 
.A(n_3224),
.B(n_1471),
.Y(n_3363)
);

INVx4_ASAP7_75t_L g3364 ( 
.A(n_3169),
.Y(n_3364)
);

NOR2xp67_ASAP7_75t_SL g3365 ( 
.A(n_3220),
.B(n_1859),
.Y(n_3365)
);

AOI21xp5_ASAP7_75t_L g3366 ( 
.A1(n_3039),
.A2(n_1477),
.B(n_1475),
.Y(n_3366)
);

AOI21xp5_ASAP7_75t_L g3367 ( 
.A1(n_3163),
.A2(n_1485),
.B(n_1481),
.Y(n_3367)
);

BUFx6f_ASAP7_75t_L g3368 ( 
.A(n_3219),
.Y(n_3368)
);

AOI21xp5_ASAP7_75t_L g3369 ( 
.A1(n_3219),
.A2(n_1494),
.B(n_1486),
.Y(n_3369)
);

AOI22xp33_ASAP7_75t_L g3370 ( 
.A1(n_3199),
.A2(n_1787),
.B1(n_1811),
.B2(n_1774),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3089),
.B(n_1304),
.Y(n_3371)
);

BUFx6f_ASAP7_75t_L g3372 ( 
.A(n_3131),
.Y(n_3372)
);

AOI21xp5_ASAP7_75t_L g3373 ( 
.A1(n_3123),
.A2(n_1505),
.B(n_1495),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_3054),
.Y(n_3374)
);

AOI21xp5_ASAP7_75t_L g3375 ( 
.A1(n_3030),
.A2(n_1514),
.B(n_1513),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_3164),
.B(n_1305),
.Y(n_3376)
);

OAI21xp5_ASAP7_75t_L g3377 ( 
.A1(n_3225),
.A2(n_1520),
.B(n_1515),
.Y(n_3377)
);

O2A1O1Ixp33_ASAP7_75t_L g3378 ( 
.A1(n_3175),
.A2(n_1534),
.B(n_1536),
.C(n_1533),
.Y(n_3378)
);

AOI21xp5_ASAP7_75t_L g3379 ( 
.A1(n_3097),
.A2(n_1538),
.B(n_1537),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_3182),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3212),
.Y(n_3381)
);

AND2x4_ASAP7_75t_L g3382 ( 
.A(n_3090),
.B(n_3104),
.Y(n_3382)
);

INVx2_ASAP7_75t_L g3383 ( 
.A(n_3193),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3326),
.Y(n_3384)
);

OAI22xp5_ASAP7_75t_L g3385 ( 
.A1(n_3237),
.A2(n_3292),
.B1(n_3247),
.B2(n_3234),
.Y(n_3385)
);

BUFx2_ASAP7_75t_L g3386 ( 
.A(n_3258),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_SL g3387 ( 
.A(n_3343),
.B(n_3210),
.Y(n_3387)
);

INVx4_ASAP7_75t_L g3388 ( 
.A(n_3253),
.Y(n_3388)
);

AOI21xp5_ASAP7_75t_L g3389 ( 
.A1(n_3249),
.A2(n_3203),
.B(n_3072),
.Y(n_3389)
);

NOR2xp33_ASAP7_75t_R g3390 ( 
.A(n_3239),
.B(n_3078),
.Y(n_3390)
);

INVx3_ASAP7_75t_L g3391 ( 
.A(n_3364),
.Y(n_3391)
);

AOI22xp5_ASAP7_75t_L g3392 ( 
.A1(n_3358),
.A2(n_3052),
.B1(n_3043),
.B2(n_3063),
.Y(n_3392)
);

CKINVDCx5p33_ASAP7_75t_R g3393 ( 
.A(n_3243),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3340),
.Y(n_3394)
);

BUFx6f_ASAP7_75t_L g3395 ( 
.A(n_3245),
.Y(n_3395)
);

INVx3_ASAP7_75t_L g3396 ( 
.A(n_3354),
.Y(n_3396)
);

OAI21x1_ASAP7_75t_L g3397 ( 
.A1(n_3256),
.A2(n_3140),
.B(n_3133),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_SL g3398 ( 
.A(n_3232),
.B(n_3209),
.Y(n_3398)
);

AOI21xp5_ASAP7_75t_L g3399 ( 
.A1(n_3251),
.A2(n_3148),
.B(n_3129),
.Y(n_3399)
);

AOI22xp5_ASAP7_75t_L g3400 ( 
.A1(n_3324),
.A2(n_3290),
.B1(n_3312),
.B2(n_3332),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_3261),
.B(n_3172),
.Y(n_3401)
);

AOI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_3314),
.A2(n_3154),
.B(n_3213),
.Y(n_3402)
);

NOR2xp33_ASAP7_75t_L g3403 ( 
.A(n_3322),
.B(n_3211),
.Y(n_3403)
);

A2O1A1Ixp33_ASAP7_75t_L g3404 ( 
.A1(n_3334),
.A2(n_3121),
.B(n_3106),
.C(n_3208),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3294),
.Y(n_3405)
);

BUFx12f_ASAP7_75t_L g3406 ( 
.A(n_3255),
.Y(n_3406)
);

AOI21xp5_ASAP7_75t_L g3407 ( 
.A1(n_3235),
.A2(n_3226),
.B(n_3095),
.Y(n_3407)
);

BUFx12f_ASAP7_75t_L g3408 ( 
.A(n_3372),
.Y(n_3408)
);

AND3x4_ASAP7_75t_L g3409 ( 
.A(n_3319),
.B(n_3146),
.C(n_3034),
.Y(n_3409)
);

AOI21xp5_ASAP7_75t_L g3410 ( 
.A1(n_3299),
.A2(n_3114),
.B(n_3186),
.Y(n_3410)
);

A2O1A1Ixp33_ASAP7_75t_L g3411 ( 
.A1(n_3377),
.A2(n_3252),
.B(n_3315),
.C(n_3271),
.Y(n_3411)
);

AOI21xp5_ASAP7_75t_L g3412 ( 
.A1(n_3273),
.A2(n_3115),
.B(n_3197),
.Y(n_3412)
);

AOI21xp5_ASAP7_75t_L g3413 ( 
.A1(n_3244),
.A2(n_3229),
.B(n_3071),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_3341),
.B(n_3246),
.Y(n_3414)
);

INVx2_ASAP7_75t_SL g3415 ( 
.A(n_3372),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3240),
.Y(n_3416)
);

BUFx12f_ASAP7_75t_L g3417 ( 
.A(n_3372),
.Y(n_3417)
);

OAI21x1_ASAP7_75t_L g3418 ( 
.A1(n_3264),
.A2(n_3165),
.B(n_1872),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3250),
.Y(n_3419)
);

NOR2xp33_ASAP7_75t_L g3420 ( 
.A(n_3348),
.B(n_3042),
.Y(n_3420)
);

O2A1O1Ixp5_ASAP7_75t_L g3421 ( 
.A1(n_3283),
.A2(n_3070),
.B(n_1872),
.C(n_1542),
.Y(n_3421)
);

INVx1_ASAP7_75t_SL g3422 ( 
.A(n_3320),
.Y(n_3422)
);

AOI22xp33_ASAP7_75t_L g3423 ( 
.A1(n_3336),
.A2(n_3179),
.B1(n_3049),
.B2(n_3108),
.Y(n_3423)
);

AOI22xp5_ASAP7_75t_L g3424 ( 
.A1(n_3318),
.A2(n_3109),
.B1(n_3143),
.B2(n_3141),
.Y(n_3424)
);

BUFx2_ASAP7_75t_L g3425 ( 
.A(n_3245),
.Y(n_3425)
);

CKINVDCx5p33_ASAP7_75t_R g3426 ( 
.A(n_3317),
.Y(n_3426)
);

O2A1O1Ixp5_ASAP7_75t_L g3427 ( 
.A1(n_3365),
.A2(n_1543),
.B(n_1544),
.C(n_1540),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_3241),
.B(n_3179),
.Y(n_3428)
);

BUFx6f_ASAP7_75t_L g3429 ( 
.A(n_3245),
.Y(n_3429)
);

AND2x2_ASAP7_75t_L g3430 ( 
.A(n_3291),
.B(n_3049),
.Y(n_3430)
);

BUFx2_ASAP7_75t_L g3431 ( 
.A(n_3293),
.Y(n_3431)
);

OAI22x1_ASAP7_75t_L g3432 ( 
.A1(n_3287),
.A2(n_1309),
.B1(n_1312),
.B2(n_1308),
.Y(n_3432)
);

AO32x1_ASAP7_75t_L g3433 ( 
.A1(n_3238),
.A2(n_1566),
.A3(n_1569),
.B1(n_1562),
.B2(n_1560),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3270),
.Y(n_3434)
);

BUFx6f_ASAP7_75t_L g3435 ( 
.A(n_3368),
.Y(n_3435)
);

OAI22xp5_ASAP7_75t_L g3436 ( 
.A1(n_3248),
.A2(n_3279),
.B1(n_3277),
.B2(n_3242),
.Y(n_3436)
);

BUFx3_ASAP7_75t_L g3437 ( 
.A(n_3329),
.Y(n_3437)
);

CKINVDCx6p67_ASAP7_75t_R g3438 ( 
.A(n_3368),
.Y(n_3438)
);

INVx5_ASAP7_75t_L g3439 ( 
.A(n_3368),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3257),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_3295),
.B(n_1571),
.Y(n_3441)
);

AOI21xp5_ASAP7_75t_L g3442 ( 
.A1(n_3262),
.A2(n_1581),
.B(n_1580),
.Y(n_3442)
);

AND2x4_ASAP7_75t_L g3443 ( 
.A(n_3382),
.B(n_1584),
.Y(n_3443)
);

O2A1O1Ixp33_ASAP7_75t_L g3444 ( 
.A1(n_3289),
.A2(n_1590),
.B(n_1598),
.C(n_1587),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_3337),
.B(n_1605),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_L g3446 ( 
.A(n_3352),
.B(n_1811),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3347),
.Y(n_3447)
);

AOI21xp5_ASAP7_75t_L g3448 ( 
.A1(n_3267),
.A2(n_1610),
.B(n_1606),
.Y(n_3448)
);

INVx2_ASAP7_75t_L g3449 ( 
.A(n_3357),
.Y(n_3449)
);

INVx1_ASAP7_75t_SL g3450 ( 
.A(n_3382),
.Y(n_3450)
);

AOI21xp5_ASAP7_75t_L g3451 ( 
.A1(n_3275),
.A2(n_1620),
.B(n_1615),
.Y(n_3451)
);

AND2x2_ASAP7_75t_L g3452 ( 
.A(n_3371),
.B(n_1637),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_3282),
.B(n_1624),
.Y(n_3453)
);

AOI22xp5_ASAP7_75t_L g3454 ( 
.A1(n_3233),
.A2(n_1842),
.B1(n_1848),
.B2(n_1825),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_SL g3455 ( 
.A(n_3236),
.B(n_1825),
.Y(n_3455)
);

NOR3xp33_ASAP7_75t_L g3456 ( 
.A(n_3338),
.B(n_3276),
.C(n_3304),
.Y(n_3456)
);

AOI21xp5_ASAP7_75t_L g3457 ( 
.A1(n_3260),
.A2(n_1635),
.B(n_1629),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_SL g3458 ( 
.A(n_3268),
.B(n_1842),
.Y(n_3458)
);

INVxp67_ASAP7_75t_SL g3459 ( 
.A(n_3310),
.Y(n_3459)
);

BUFx4f_ASAP7_75t_L g3460 ( 
.A(n_3363),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_3263),
.Y(n_3461)
);

INVx2_ASAP7_75t_L g3462 ( 
.A(n_3265),
.Y(n_3462)
);

AO22x1_ASAP7_75t_L g3463 ( 
.A1(n_3381),
.A2(n_1320),
.B1(n_1322),
.B2(n_1315),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3360),
.Y(n_3464)
);

AOI21xp5_ASAP7_75t_L g3465 ( 
.A1(n_3254),
.A2(n_1653),
.B(n_1645),
.Y(n_3465)
);

INVxp67_ASAP7_75t_SL g3466 ( 
.A(n_3350),
.Y(n_3466)
);

O2A1O1Ixp33_ASAP7_75t_L g3467 ( 
.A1(n_3342),
.A2(n_1655),
.B(n_1668),
.C(n_1661),
.Y(n_3467)
);

AOI21xp5_ASAP7_75t_L g3468 ( 
.A1(n_3266),
.A2(n_1672),
.B(n_1671),
.Y(n_3468)
);

CKINVDCx20_ASAP7_75t_R g3469 ( 
.A(n_3300),
.Y(n_3469)
);

AOI21xp5_ASAP7_75t_L g3470 ( 
.A1(n_3259),
.A2(n_1678),
.B(n_1676),
.Y(n_3470)
);

NOR2xp33_ASAP7_75t_L g3471 ( 
.A(n_3331),
.B(n_1875),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3361),
.Y(n_3472)
);

NOR2xp33_ASAP7_75t_L g3473 ( 
.A(n_3301),
.B(n_1875),
.Y(n_3473)
);

O2A1O1Ixp33_ASAP7_75t_L g3474 ( 
.A1(n_3298),
.A2(n_1680),
.B(n_1689),
.C(n_1686),
.Y(n_3474)
);

AOI22xp33_ASAP7_75t_L g3475 ( 
.A1(n_3362),
.A2(n_1904),
.B1(n_1903),
.B2(n_1693),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3285),
.B(n_1695),
.Y(n_3476)
);

NOR2xp33_ASAP7_75t_L g3477 ( 
.A(n_3370),
.B(n_1903),
.Y(n_3477)
);

OAI22xp5_ASAP7_75t_L g3478 ( 
.A1(n_3316),
.A2(n_1904),
.B1(n_1327),
.B2(n_1329),
.Y(n_3478)
);

AOI22xp33_ASAP7_75t_L g3479 ( 
.A1(n_3321),
.A2(n_1693),
.B1(n_1714),
.B2(n_1641),
.Y(n_3479)
);

AOI21xp5_ASAP7_75t_L g3480 ( 
.A1(n_3376),
.A2(n_1704),
.B(n_1702),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3323),
.B(n_1707),
.Y(n_3481)
);

AOI22xp33_ASAP7_75t_L g3482 ( 
.A1(n_3328),
.A2(n_1693),
.B1(n_1714),
.B2(n_1641),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_3333),
.B(n_1710),
.Y(n_3483)
);

NOR2xp33_ASAP7_75t_R g3484 ( 
.A(n_3335),
.B(n_1045),
.Y(n_3484)
);

AND2x2_ASAP7_75t_L g3485 ( 
.A(n_3383),
.B(n_1641),
.Y(n_3485)
);

AOI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_3296),
.A2(n_3306),
.B(n_3302),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3303),
.B(n_3308),
.Y(n_3487)
);

AND3x1_ASAP7_75t_SL g3488 ( 
.A(n_3280),
.B(n_1930),
.C(n_1922),
.Y(n_3488)
);

BUFx6f_ASAP7_75t_L g3489 ( 
.A(n_3374),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_SL g3490 ( 
.A(n_3380),
.B(n_1714),
.Y(n_3490)
);

CKINVDCx16_ASAP7_75t_R g3491 ( 
.A(n_3309),
.Y(n_3491)
);

AOI22x1_ASAP7_75t_L g3492 ( 
.A1(n_3284),
.A2(n_1331),
.B1(n_1332),
.B2(n_1323),
.Y(n_3492)
);

AND2x2_ASAP7_75t_L g3493 ( 
.A(n_3311),
.B(n_1861),
.Y(n_3493)
);

CKINVDCx6p67_ASAP7_75t_R g3494 ( 
.A(n_3344),
.Y(n_3494)
);

INVx2_ASAP7_75t_L g3495 ( 
.A(n_3269),
.Y(n_3495)
);

NOR2xp33_ASAP7_75t_L g3496 ( 
.A(n_3345),
.B(n_3351),
.Y(n_3496)
);

AOI22xp33_ASAP7_75t_L g3497 ( 
.A1(n_3346),
.A2(n_1861),
.B1(n_1717),
.B2(n_1718),
.Y(n_3497)
);

NAND3xp33_ASAP7_75t_L g3498 ( 
.A(n_3286),
.B(n_1335),
.C(n_1334),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3281),
.B(n_1711),
.Y(n_3499)
);

INVx2_ASAP7_75t_L g3500 ( 
.A(n_3355),
.Y(n_3500)
);

OAI22xp5_ASAP7_75t_L g3501 ( 
.A1(n_3356),
.A2(n_1338),
.B1(n_1340),
.B2(n_1336),
.Y(n_3501)
);

O2A1O1Ixp33_ASAP7_75t_L g3502 ( 
.A1(n_3288),
.A2(n_1731),
.B(n_1733),
.C(n_1723),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3278),
.Y(n_3503)
);

AOI22xp33_ASAP7_75t_SL g3504 ( 
.A1(n_3297),
.A2(n_1861),
.B1(n_1342),
.B2(n_1345),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3272),
.Y(n_3505)
);

AOI21xp5_ASAP7_75t_L g3506 ( 
.A1(n_3330),
.A2(n_1744),
.B(n_1737),
.Y(n_3506)
);

BUFx6f_ASAP7_75t_L g3507 ( 
.A(n_3369),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3339),
.B(n_1745),
.Y(n_3508)
);

AOI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_3349),
.A2(n_1749),
.B(n_1748),
.Y(n_3509)
);

INVxp67_ASAP7_75t_SL g3510 ( 
.A(n_3378),
.Y(n_3510)
);

NOR3xp33_ASAP7_75t_SL g3511 ( 
.A(n_3366),
.B(n_1346),
.C(n_1341),
.Y(n_3511)
);

OR2x2_ASAP7_75t_L g3512 ( 
.A(n_3353),
.B(n_1347),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3274),
.Y(n_3513)
);

OAI22xp33_ASAP7_75t_L g3514 ( 
.A1(n_3367),
.A2(n_3375),
.B1(n_3379),
.B2(n_3373),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3359),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_L g3516 ( 
.A(n_3305),
.B(n_1757),
.Y(n_3516)
);

AO32x1_ASAP7_75t_L g3517 ( 
.A1(n_3325),
.A2(n_1769),
.A3(n_1771),
.B1(n_1768),
.B2(n_1764),
.Y(n_3517)
);

AND2x2_ASAP7_75t_SL g3518 ( 
.A(n_3307),
.B(n_1778),
.Y(n_3518)
);

BUFx2_ASAP7_75t_L g3519 ( 
.A(n_3313),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3327),
.B(n_1781),
.Y(n_3520)
);

OAI21xp5_ASAP7_75t_L g3521 ( 
.A1(n_3314),
.A2(n_1798),
.B(n_1783),
.Y(n_3521)
);

NOR2xp33_ASAP7_75t_L g3522 ( 
.A(n_3237),
.B(n_1348),
.Y(n_3522)
);

OR2x6_ASAP7_75t_L g3523 ( 
.A(n_3364),
.B(n_1801),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3384),
.Y(n_3524)
);

NOR2x1_ASAP7_75t_SL g3525 ( 
.A(n_3385),
.B(n_1812),
.Y(n_3525)
);

OAI21x1_ASAP7_75t_L g3526 ( 
.A1(n_3389),
.A2(n_1817),
.B(n_1815),
.Y(n_3526)
);

NAND3xp33_ASAP7_75t_L g3527 ( 
.A(n_3400),
.B(n_1350),
.C(n_1349),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_3447),
.Y(n_3528)
);

OAI21x1_ASAP7_75t_L g3529 ( 
.A1(n_3402),
.A2(n_1826),
.B(n_1824),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3394),
.Y(n_3530)
);

OAI22xp5_ASAP7_75t_L g3531 ( 
.A1(n_3401),
.A2(n_1353),
.B1(n_1357),
.B2(n_1351),
.Y(n_3531)
);

CKINVDCx5p33_ASAP7_75t_R g3532 ( 
.A(n_3393),
.Y(n_3532)
);

NOR2xp33_ASAP7_75t_R g3533 ( 
.A(n_3426),
.B(n_1048),
.Y(n_3533)
);

OAI21xp5_ASAP7_75t_SL g3534 ( 
.A1(n_3477),
.A2(n_1828),
.B(n_1827),
.Y(n_3534)
);

INVx2_ASAP7_75t_L g3535 ( 
.A(n_3449),
.Y(n_3535)
);

AO31x2_ASAP7_75t_L g3536 ( 
.A1(n_3411),
.A2(n_1830),
.A3(n_1835),
.B(n_1829),
.Y(n_3536)
);

A2O1A1Ixp33_ASAP7_75t_L g3537 ( 
.A1(n_3522),
.A2(n_1851),
.B(n_1855),
.C(n_1847),
.Y(n_3537)
);

AOI221xp5_ASAP7_75t_SL g3538 ( 
.A1(n_3403),
.A2(n_1867),
.B1(n_1870),
.B2(n_1865),
.C(n_1862),
.Y(n_3538)
);

OAI21xp5_ASAP7_75t_L g3539 ( 
.A1(n_3496),
.A2(n_1883),
.B(n_1876),
.Y(n_3539)
);

AO31x2_ASAP7_75t_L g3540 ( 
.A1(n_3470),
.A2(n_1887),
.A3(n_1889),
.B(n_1885),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3440),
.B(n_1358),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3464),
.Y(n_3542)
);

OA21x2_ASAP7_75t_L g3543 ( 
.A1(n_3521),
.A2(n_1900),
.B(n_1894),
.Y(n_3543)
);

O2A1O1Ixp33_ASAP7_75t_L g3544 ( 
.A1(n_3458),
.A2(n_1917),
.B(n_1914),
.C(n_1362),
.Y(n_3544)
);

OR2x2_ASAP7_75t_L g3545 ( 
.A(n_3414),
.B(n_1360),
.Y(n_3545)
);

INVx2_ASAP7_75t_L g3546 ( 
.A(n_3419),
.Y(n_3546)
);

NAND3xp33_ASAP7_75t_L g3547 ( 
.A(n_3456),
.B(n_1366),
.C(n_1365),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3416),
.Y(n_3548)
);

AND2x2_ASAP7_75t_L g3549 ( 
.A(n_3452),
.B(n_1367),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3461),
.B(n_1371),
.Y(n_3550)
);

AO21x1_ASAP7_75t_L g3551 ( 
.A1(n_3399),
.A2(n_1),
.B(n_3),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_3462),
.B(n_1372),
.Y(n_3552)
);

AOI22xp5_ASAP7_75t_L g3553 ( 
.A1(n_3446),
.A2(n_1378),
.B1(n_1380),
.B2(n_1374),
.Y(n_3553)
);

O2A1O1Ixp5_ASAP7_75t_SL g3554 ( 
.A1(n_3455),
.A2(n_3505),
.B(n_3436),
.C(n_3503),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3405),
.B(n_1385),
.Y(n_3555)
);

OAI21x1_ASAP7_75t_L g3556 ( 
.A1(n_3418),
.A2(n_1053),
.B(n_1051),
.Y(n_3556)
);

INVx4_ASAP7_75t_L g3557 ( 
.A(n_3439),
.Y(n_3557)
);

OAI21xp5_ASAP7_75t_L g3558 ( 
.A1(n_3486),
.A2(n_1390),
.B(n_1389),
.Y(n_3558)
);

NAND3xp33_ASAP7_75t_L g3559 ( 
.A(n_3404),
.B(n_3420),
.C(n_3504),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_3434),
.Y(n_3560)
);

OAI21xp5_ASAP7_75t_L g3561 ( 
.A1(n_3487),
.A2(n_1896),
.B(n_1895),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3500),
.B(n_1392),
.Y(n_3562)
);

O2A1O1Ixp33_ASAP7_75t_SL g3563 ( 
.A1(n_3514),
.A2(n_5),
.B(n_3),
.C(n_4),
.Y(n_3563)
);

CKINVDCx20_ASAP7_75t_R g3564 ( 
.A(n_3469),
.Y(n_3564)
);

AND2x4_ASAP7_75t_L g3565 ( 
.A(n_3439),
.B(n_3437),
.Y(n_3565)
);

AND2x2_ASAP7_75t_L g3566 ( 
.A(n_3493),
.B(n_3491),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3472),
.Y(n_3567)
);

OAI21x1_ASAP7_75t_L g3568 ( 
.A1(n_3410),
.A2(n_1058),
.B(n_1055),
.Y(n_3568)
);

AOI21x1_ASAP7_75t_L g3569 ( 
.A1(n_3412),
.A2(n_1060),
.B(n_1059),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_SL g3570 ( 
.A(n_3392),
.B(n_1908),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3473),
.B(n_1394),
.Y(n_3571)
);

OAI21x1_ASAP7_75t_L g3572 ( 
.A1(n_3397),
.A2(n_1068),
.B(n_1061),
.Y(n_3572)
);

AO31x2_ASAP7_75t_L g3573 ( 
.A1(n_3465),
.A2(n_1070),
.A3(n_1072),
.B(n_1069),
.Y(n_3573)
);

NOR4xp25_ASAP7_75t_L g3574 ( 
.A(n_3467),
.B(n_14),
.C(n_22),
.D(n_4),
.Y(n_3574)
);

BUFx2_ASAP7_75t_L g3575 ( 
.A(n_3386),
.Y(n_3575)
);

BUFx8_ASAP7_75t_SL g3576 ( 
.A(n_3408),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3398),
.B(n_1395),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_SL g3578 ( 
.A(n_3413),
.B(n_3424),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3428),
.B(n_1396),
.Y(n_3579)
);

BUFx6f_ASAP7_75t_L g3580 ( 
.A(n_3417),
.Y(n_3580)
);

HB1xp67_ASAP7_75t_L g3581 ( 
.A(n_3422),
.Y(n_3581)
);

OAI21x1_ASAP7_75t_L g3582 ( 
.A1(n_3448),
.A2(n_5),
.B(n_6),
.Y(n_3582)
);

OR2x2_ASAP7_75t_L g3583 ( 
.A(n_3445),
.B(n_1398),
.Y(n_3583)
);

A2O1A1Ixp33_ASAP7_75t_L g3584 ( 
.A1(n_3407),
.A2(n_1407),
.B(n_1408),
.C(n_1405),
.Y(n_3584)
);

OAI21x1_ASAP7_75t_L g3585 ( 
.A1(n_3457),
.A2(n_7),
.B(n_8),
.Y(n_3585)
);

OAI21xp5_ASAP7_75t_L g3586 ( 
.A1(n_3421),
.A2(n_1920),
.B(n_1909),
.Y(n_3586)
);

AOI21xp5_ASAP7_75t_L g3587 ( 
.A1(n_3513),
.A2(n_1417),
.B(n_1414),
.Y(n_3587)
);

AOI21xp5_ASAP7_75t_L g3588 ( 
.A1(n_3519),
.A2(n_1421),
.B(n_1420),
.Y(n_3588)
);

OAI22x1_ASAP7_75t_L g3589 ( 
.A1(n_3454),
.A2(n_1423),
.B1(n_1425),
.B2(n_1422),
.Y(n_3589)
);

AO31x2_ASAP7_75t_L g3590 ( 
.A1(n_3468),
.A2(n_11),
.A3(n_7),
.B(n_9),
.Y(n_3590)
);

OAI21x1_ASAP7_75t_L g3591 ( 
.A1(n_3451),
.A2(n_12),
.B(n_14),
.Y(n_3591)
);

CKINVDCx16_ASAP7_75t_R g3592 ( 
.A(n_3390),
.Y(n_3592)
);

BUFx8_ASAP7_75t_L g3593 ( 
.A(n_3435),
.Y(n_3593)
);

OAI21xp5_ASAP7_75t_L g3594 ( 
.A1(n_3510),
.A2(n_1901),
.B(n_1899),
.Y(n_3594)
);

INVx2_ASAP7_75t_L g3595 ( 
.A(n_3489),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_3489),
.Y(n_3596)
);

OAI21x1_ASAP7_75t_L g3597 ( 
.A1(n_3427),
.A2(n_12),
.B(n_15),
.Y(n_3597)
);

OAI21xp5_ASAP7_75t_L g3598 ( 
.A1(n_3453),
.A2(n_3481),
.B(n_3476),
.Y(n_3598)
);

OA21x2_ASAP7_75t_L g3599 ( 
.A1(n_3515),
.A2(n_1427),
.B(n_1426),
.Y(n_3599)
);

OAI21x1_ASAP7_75t_L g3600 ( 
.A1(n_3480),
.A2(n_16),
.B(n_17),
.Y(n_3600)
);

NAND3x1_ASAP7_75t_L g3601 ( 
.A(n_3430),
.B(n_16),
.C(n_17),
.Y(n_3601)
);

INVx1_ASAP7_75t_SL g3602 ( 
.A(n_3450),
.Y(n_3602)
);

AOI21xp5_ASAP7_75t_L g3603 ( 
.A1(n_3483),
.A2(n_1434),
.B(n_1430),
.Y(n_3603)
);

NOR2x1_ASAP7_75t_L g3604 ( 
.A(n_3391),
.B(n_1436),
.Y(n_3604)
);

OAI22x1_ASAP7_75t_L g3605 ( 
.A1(n_3387),
.A2(n_1438),
.B1(n_1441),
.B2(n_1437),
.Y(n_3605)
);

OAI21x1_ASAP7_75t_L g3606 ( 
.A1(n_3495),
.A2(n_18),
.B(n_19),
.Y(n_3606)
);

AOI21xp5_ASAP7_75t_L g3607 ( 
.A1(n_3507),
.A2(n_1448),
.B(n_1447),
.Y(n_3607)
);

AOI211x1_ASAP7_75t_L g3608 ( 
.A1(n_3463),
.A2(n_1450),
.B(n_1454),
.C(n_1449),
.Y(n_3608)
);

O2A1O1Ixp5_ASAP7_75t_L g3609 ( 
.A1(n_3441),
.A2(n_1456),
.B(n_1457),
.C(n_1455),
.Y(n_3609)
);

O2A1O1Ixp33_ASAP7_75t_L g3610 ( 
.A1(n_3512),
.A2(n_1465),
.B(n_1468),
.C(n_1464),
.Y(n_3610)
);

O2A1O1Ixp5_ASAP7_75t_L g3611 ( 
.A1(n_3490),
.A2(n_1470),
.B(n_1472),
.C(n_1469),
.Y(n_3611)
);

AOI221xp5_ASAP7_75t_L g3612 ( 
.A1(n_3478),
.A2(n_1478),
.B1(n_1479),
.B2(n_1474),
.C(n_1473),
.Y(n_3612)
);

OAI21xp5_ASAP7_75t_L g3613 ( 
.A1(n_3498),
.A2(n_1905),
.B(n_1898),
.Y(n_3613)
);

OAI22xp33_ASAP7_75t_L g3614 ( 
.A1(n_3494),
.A2(n_1487),
.B1(n_1488),
.B2(n_1482),
.Y(n_3614)
);

O2A1O1Ixp33_ASAP7_75t_SL g3615 ( 
.A1(n_3499),
.A2(n_3508),
.B(n_3516),
.C(n_3520),
.Y(n_3615)
);

AOI21xp5_ASAP7_75t_L g3616 ( 
.A1(n_3507),
.A2(n_1491),
.B(n_1489),
.Y(n_3616)
);

OAI21x1_ASAP7_75t_L g3617 ( 
.A1(n_3442),
.A2(n_19),
.B(n_20),
.Y(n_3617)
);

INVx3_ASAP7_75t_L g3618 ( 
.A(n_3388),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3471),
.B(n_1492),
.Y(n_3619)
);

OR2x2_ASAP7_75t_L g3620 ( 
.A(n_3423),
.B(n_1493),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3475),
.B(n_1496),
.Y(n_3621)
);

INVx3_ASAP7_75t_L g3622 ( 
.A(n_3406),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3474),
.Y(n_3623)
);

AOI21xp5_ASAP7_75t_L g3624 ( 
.A1(n_3518),
.A2(n_1504),
.B(n_1499),
.Y(n_3624)
);

AOI221x1_ASAP7_75t_L g3625 ( 
.A1(n_3432),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.C(n_24),
.Y(n_3625)
);

BUFx3_ASAP7_75t_L g3626 ( 
.A(n_3435),
.Y(n_3626)
);

OAI21xp5_ASAP7_75t_L g3627 ( 
.A1(n_3501),
.A2(n_3482),
.B(n_3479),
.Y(n_3627)
);

A2O1A1Ixp33_ASAP7_75t_L g3628 ( 
.A1(n_3511),
.A2(n_1509),
.B(n_1510),
.C(n_1507),
.Y(n_3628)
);

AO31x2_ASAP7_75t_L g3629 ( 
.A1(n_3506),
.A2(n_26),
.A3(n_24),
.B(n_25),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3444),
.Y(n_3630)
);

OAI21x1_ASAP7_75t_L g3631 ( 
.A1(n_3509),
.A2(n_25),
.B(n_26),
.Y(n_3631)
);

OAI21xp5_ASAP7_75t_L g3632 ( 
.A1(n_3497),
.A2(n_1512),
.B(n_1511),
.Y(n_3632)
);

AOI21xp5_ASAP7_75t_L g3633 ( 
.A1(n_3517),
.A2(n_1519),
.B(n_1516),
.Y(n_3633)
);

AOI21x1_ASAP7_75t_L g3634 ( 
.A1(n_3425),
.A2(n_27),
.B(n_28),
.Y(n_3634)
);

OAI21x1_ASAP7_75t_L g3635 ( 
.A1(n_3556),
.A2(n_3502),
.B(n_3492),
.Y(n_3635)
);

OAI21x1_ASAP7_75t_L g3636 ( 
.A1(n_3572),
.A2(n_3396),
.B(n_3466),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3524),
.Y(n_3637)
);

OR2x2_ASAP7_75t_L g3638 ( 
.A(n_3581),
.B(n_3443),
.Y(n_3638)
);

INVx8_ASAP7_75t_L g3639 ( 
.A(n_3576),
.Y(n_3639)
);

AOI222xp33_ASAP7_75t_L g3640 ( 
.A1(n_3539),
.A2(n_1527),
.B1(n_1559),
.B2(n_1597),
.C1(n_1579),
.C2(n_1546),
.Y(n_3640)
);

AO21x2_ASAP7_75t_L g3641 ( 
.A1(n_3578),
.A2(n_3484),
.B(n_3485),
.Y(n_3641)
);

OA21x2_ASAP7_75t_L g3642 ( 
.A1(n_3538),
.A2(n_3459),
.B(n_3517),
.Y(n_3642)
);

AND2x2_ASAP7_75t_L g3643 ( 
.A(n_3566),
.B(n_3528),
.Y(n_3643)
);

AOI22xp33_ASAP7_75t_L g3644 ( 
.A1(n_3559),
.A2(n_3409),
.B1(n_3523),
.B2(n_3460),
.Y(n_3644)
);

AO21x1_ASAP7_75t_L g3645 ( 
.A1(n_3570),
.A2(n_3433),
.B(n_3488),
.Y(n_3645)
);

INVx2_ASAP7_75t_L g3646 ( 
.A(n_3535),
.Y(n_3646)
);

OAI21xp5_ASAP7_75t_L g3647 ( 
.A1(n_3547),
.A2(n_3523),
.B(n_3431),
.Y(n_3647)
);

OAI21x1_ASAP7_75t_L g3648 ( 
.A1(n_3526),
.A2(n_3433),
.B(n_3438),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_3546),
.Y(n_3649)
);

AOI21xp5_ASAP7_75t_L g3650 ( 
.A1(n_3615),
.A2(n_3439),
.B(n_3415),
.Y(n_3650)
);

OA21x2_ASAP7_75t_L g3651 ( 
.A1(n_3529),
.A2(n_1522),
.B(n_1521),
.Y(n_3651)
);

OA21x2_ASAP7_75t_L g3652 ( 
.A1(n_3551),
.A2(n_3597),
.B(n_3585),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3530),
.Y(n_3653)
);

OAI21xp5_ASAP7_75t_L g3654 ( 
.A1(n_3598),
.A2(n_1528),
.B(n_1526),
.Y(n_3654)
);

INVx5_ASAP7_75t_L g3655 ( 
.A(n_3557),
.Y(n_3655)
);

AND2x2_ASAP7_75t_L g3656 ( 
.A(n_3560),
.B(n_3395),
.Y(n_3656)
);

AOI22x1_ASAP7_75t_L g3657 ( 
.A1(n_3589),
.A2(n_1530),
.B1(n_1531),
.B2(n_1529),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3567),
.Y(n_3658)
);

OAI211xp5_ASAP7_75t_SL g3659 ( 
.A1(n_3534),
.A2(n_1541),
.B(n_1545),
.C(n_1535),
.Y(n_3659)
);

AOI22xp33_ASAP7_75t_L g3660 ( 
.A1(n_3627),
.A2(n_1548),
.B1(n_1552),
.B2(n_1547),
.Y(n_3660)
);

NOR2x1_ASAP7_75t_R g3661 ( 
.A(n_3532),
.B(n_3395),
.Y(n_3661)
);

OAI21x1_ASAP7_75t_L g3662 ( 
.A1(n_3568),
.A2(n_3429),
.B(n_29),
.Y(n_3662)
);

NAND2xp33_ASAP7_75t_L g3663 ( 
.A(n_3601),
.B(n_3429),
.Y(n_3663)
);

CKINVDCx6p67_ASAP7_75t_R g3664 ( 
.A(n_3592),
.Y(n_3664)
);

AOI22xp33_ASAP7_75t_L g3665 ( 
.A1(n_3527),
.A2(n_1554),
.B1(n_1557),
.B2(n_1553),
.Y(n_3665)
);

XOR2xp5_ASAP7_75t_L g3666 ( 
.A(n_3564),
.B(n_1558),
.Y(n_3666)
);

BUFx3_ASAP7_75t_L g3667 ( 
.A(n_3593),
.Y(n_3667)
);

BUFx2_ASAP7_75t_L g3668 ( 
.A(n_3575),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_3542),
.Y(n_3669)
);

NOR2xp33_ASAP7_75t_L g3670 ( 
.A(n_3602),
.B(n_1561),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3548),
.Y(n_3671)
);

AND2x2_ASAP7_75t_L g3672 ( 
.A(n_3599),
.B(n_29),
.Y(n_3672)
);

AO32x2_ASAP7_75t_L g3673 ( 
.A1(n_3531),
.A2(n_3574),
.A3(n_3625),
.B1(n_3554),
.B2(n_3563),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_SL g3674 ( 
.A(n_3594),
.B(n_1563),
.Y(n_3674)
);

OAI22xp5_ASAP7_75t_L g3675 ( 
.A1(n_3620),
.A2(n_1567),
.B1(n_1570),
.B2(n_1564),
.Y(n_3675)
);

AO21x2_ASAP7_75t_L g3676 ( 
.A1(n_3525),
.A2(n_1575),
.B(n_1573),
.Y(n_3676)
);

OAI22xp33_ASAP7_75t_L g3677 ( 
.A1(n_3571),
.A2(n_1882),
.B1(n_1888),
.B2(n_1881),
.Y(n_3677)
);

AO31x2_ASAP7_75t_L g3678 ( 
.A1(n_3584),
.A2(n_32),
.A3(n_30),
.B(n_31),
.Y(n_3678)
);

OAI21x1_ASAP7_75t_L g3679 ( 
.A1(n_3569),
.A2(n_30),
.B(n_31),
.Y(n_3679)
);

OAI21x1_ASAP7_75t_L g3680 ( 
.A1(n_3582),
.A2(n_32),
.B(n_33),
.Y(n_3680)
);

AND2x2_ASAP7_75t_L g3681 ( 
.A(n_3605),
.B(n_33),
.Y(n_3681)
);

AO31x2_ASAP7_75t_L g3682 ( 
.A1(n_3633),
.A2(n_36),
.A3(n_34),
.B(n_35),
.Y(n_3682)
);

OAI22xp33_ASAP7_75t_L g3683 ( 
.A1(n_3619),
.A2(n_1926),
.B1(n_1928),
.B2(n_1921),
.Y(n_3683)
);

OAI22xp33_ASAP7_75t_L g3684 ( 
.A1(n_3577),
.A2(n_1583),
.B1(n_1585),
.B2(n_1582),
.Y(n_3684)
);

OAI21x1_ASAP7_75t_L g3685 ( 
.A1(n_3631),
.A2(n_34),
.B(n_37),
.Y(n_3685)
);

OAI21x1_ASAP7_75t_L g3686 ( 
.A1(n_3617),
.A2(n_37),
.B(n_39),
.Y(n_3686)
);

AND2x2_ASAP7_75t_L g3687 ( 
.A(n_3595),
.B(n_40),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3536),
.Y(n_3688)
);

AO21x2_ASAP7_75t_L g3689 ( 
.A1(n_3558),
.A2(n_1591),
.B(n_1589),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3536),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3590),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3590),
.Y(n_3692)
);

AOI22xp33_ASAP7_75t_SL g3693 ( 
.A1(n_3561),
.A2(n_3621),
.B1(n_3543),
.B2(n_3630),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3629),
.Y(n_3694)
);

AO21x2_ASAP7_75t_L g3695 ( 
.A1(n_3587),
.A2(n_1593),
.B(n_1592),
.Y(n_3695)
);

BUFx3_ASAP7_75t_L g3696 ( 
.A(n_3626),
.Y(n_3696)
);

NOR2xp33_ASAP7_75t_L g3697 ( 
.A(n_3614),
.B(n_1600),
.Y(n_3697)
);

INVx1_ASAP7_75t_SL g3698 ( 
.A(n_3596),
.Y(n_3698)
);

INVx2_ASAP7_75t_L g3699 ( 
.A(n_3606),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3545),
.B(n_1891),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3541),
.B(n_1892),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3600),
.Y(n_3702)
);

INVx4_ASAP7_75t_L g3703 ( 
.A(n_3580),
.Y(n_3703)
);

OAI21x1_ASAP7_75t_SL g3704 ( 
.A1(n_3634),
.A2(n_40),
.B(n_41),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3629),
.Y(n_3705)
);

OAI21xp5_ASAP7_75t_L g3706 ( 
.A1(n_3609),
.A2(n_1602),
.B(n_1601),
.Y(n_3706)
);

OAI21x1_ASAP7_75t_L g3707 ( 
.A1(n_3591),
.A2(n_42),
.B(n_43),
.Y(n_3707)
);

AOI21xp5_ASAP7_75t_L g3708 ( 
.A1(n_3623),
.A2(n_1608),
.B(n_1607),
.Y(n_3708)
);

BUFx2_ASAP7_75t_L g3709 ( 
.A(n_3565),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3540),
.Y(n_3710)
);

OR2x2_ASAP7_75t_L g3711 ( 
.A(n_3691),
.B(n_3540),
.Y(n_3711)
);

AOI21xp5_ASAP7_75t_L g3712 ( 
.A1(n_3689),
.A2(n_3610),
.B(n_3544),
.Y(n_3712)
);

AO21x2_ASAP7_75t_L g3713 ( 
.A1(n_3710),
.A2(n_3586),
.B(n_3588),
.Y(n_3713)
);

CKINVDCx5p33_ASAP7_75t_R g3714 ( 
.A(n_3664),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3643),
.B(n_3555),
.Y(n_3715)
);

AND2x4_ASAP7_75t_L g3716 ( 
.A(n_3668),
.B(n_3622),
.Y(n_3716)
);

INVxp67_ASAP7_75t_SL g3717 ( 
.A(n_3692),
.Y(n_3717)
);

OA21x2_ASAP7_75t_L g3718 ( 
.A1(n_3679),
.A2(n_3537),
.B(n_3607),
.Y(n_3718)
);

OA21x2_ASAP7_75t_L g3719 ( 
.A1(n_3680),
.A2(n_3616),
.B(n_3611),
.Y(n_3719)
);

INVx2_ASAP7_75t_L g3720 ( 
.A(n_3649),
.Y(n_3720)
);

OR2x2_ASAP7_75t_L g3721 ( 
.A(n_3637),
.B(n_3579),
.Y(n_3721)
);

OAI21x1_ASAP7_75t_L g3722 ( 
.A1(n_3662),
.A2(n_3604),
.B(n_3613),
.Y(n_3722)
);

OR2x6_ASAP7_75t_L g3723 ( 
.A(n_3639),
.B(n_3580),
.Y(n_3723)
);

O2A1O1Ixp33_ASAP7_75t_L g3724 ( 
.A1(n_3674),
.A2(n_3628),
.B(n_3632),
.C(n_3624),
.Y(n_3724)
);

BUFx2_ASAP7_75t_L g3725 ( 
.A(n_3709),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3653),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3658),
.B(n_3550),
.Y(n_3727)
);

AND2x4_ASAP7_75t_L g3728 ( 
.A(n_3656),
.B(n_3618),
.Y(n_3728)
);

OAI21x1_ASAP7_75t_L g3729 ( 
.A1(n_3635),
.A2(n_3702),
.B(n_3648),
.Y(n_3729)
);

OR2x2_ASAP7_75t_L g3730 ( 
.A(n_3694),
.B(n_3573),
.Y(n_3730)
);

INVx2_ASAP7_75t_L g3731 ( 
.A(n_3669),
.Y(n_3731)
);

OAI21xp5_ASAP7_75t_L g3732 ( 
.A1(n_3693),
.A2(n_3553),
.B(n_3603),
.Y(n_3732)
);

CKINVDCx11_ASAP7_75t_R g3733 ( 
.A(n_3639),
.Y(n_3733)
);

INVx1_ASAP7_75t_SL g3734 ( 
.A(n_3638),
.Y(n_3734)
);

AO31x2_ASAP7_75t_L g3735 ( 
.A1(n_3705),
.A2(n_3552),
.A3(n_3562),
.B(n_3573),
.Y(n_3735)
);

BUFx2_ASAP7_75t_L g3736 ( 
.A(n_3696),
.Y(n_3736)
);

AO31x2_ASAP7_75t_L g3737 ( 
.A1(n_3688),
.A2(n_3608),
.A3(n_46),
.B(n_44),
.Y(n_3737)
);

INVx2_ASAP7_75t_SL g3738 ( 
.A(n_3667),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_3646),
.B(n_3549),
.Y(n_3739)
);

BUFx6f_ASAP7_75t_L g3740 ( 
.A(n_3703),
.Y(n_3740)
);

AOI21xp5_ASAP7_75t_L g3741 ( 
.A1(n_3641),
.A2(n_3583),
.B(n_3612),
.Y(n_3741)
);

AOI21xp5_ASAP7_75t_L g3742 ( 
.A1(n_3650),
.A2(n_3654),
.B(n_3651),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_3671),
.Y(n_3743)
);

NAND2x1p5_ASAP7_75t_L g3744 ( 
.A(n_3655),
.B(n_3533),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3690),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_3698),
.B(n_1609),
.Y(n_3746)
);

OA21x2_ASAP7_75t_L g3747 ( 
.A1(n_3685),
.A2(n_3707),
.B(n_3686),
.Y(n_3747)
);

OR2x2_ASAP7_75t_L g3748 ( 
.A(n_3699),
.B(n_44),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3678),
.Y(n_3749)
);

OA21x2_ASAP7_75t_L g3750 ( 
.A1(n_3636),
.A2(n_1613),
.B(n_1612),
.Y(n_3750)
);

BUFx2_ASAP7_75t_SL g3751 ( 
.A(n_3655),
.Y(n_3751)
);

BUFx2_ASAP7_75t_L g3752 ( 
.A(n_3661),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3678),
.Y(n_3753)
);

OAI21x1_ASAP7_75t_SL g3754 ( 
.A1(n_3645),
.A2(n_45),
.B(n_47),
.Y(n_3754)
);

OAI21x1_ASAP7_75t_L g3755 ( 
.A1(n_3652),
.A2(n_45),
.B(n_47),
.Y(n_3755)
);

AOI21xp5_ASAP7_75t_L g3756 ( 
.A1(n_3695),
.A2(n_1616),
.B(n_1614),
.Y(n_3756)
);

AOI21xp5_ASAP7_75t_L g3757 ( 
.A1(n_3652),
.A2(n_1618),
.B(n_1617),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_3687),
.Y(n_3758)
);

HB1xp67_ASAP7_75t_L g3759 ( 
.A(n_3642),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3672),
.Y(n_3760)
);

OA21x2_ASAP7_75t_L g3761 ( 
.A1(n_3704),
.A2(n_1622),
.B(n_1619),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_3681),
.B(n_1623),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_3644),
.B(n_1626),
.Y(n_3763)
);

AO21x2_ASAP7_75t_L g3764 ( 
.A1(n_3706),
.A2(n_3708),
.B(n_3647),
.Y(n_3764)
);

INVx4_ASAP7_75t_L g3765 ( 
.A(n_3655),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3682),
.Y(n_3766)
);

OA21x2_ASAP7_75t_L g3767 ( 
.A1(n_3657),
.A2(n_1628),
.B(n_1627),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3726),
.Y(n_3768)
);

OR2x6_ASAP7_75t_L g3769 ( 
.A(n_3751),
.B(n_3700),
.Y(n_3769)
);

INVx3_ASAP7_75t_L g3770 ( 
.A(n_3728),
.Y(n_3770)
);

OAI21xp5_ASAP7_75t_L g3771 ( 
.A1(n_3741),
.A2(n_3697),
.B(n_3660),
.Y(n_3771)
);

INVx2_ASAP7_75t_L g3772 ( 
.A(n_3731),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3743),
.Y(n_3773)
);

OAI21x1_ASAP7_75t_L g3774 ( 
.A1(n_3729),
.A2(n_3701),
.B(n_3673),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3745),
.Y(n_3775)
);

OA21x2_ASAP7_75t_L g3776 ( 
.A1(n_3742),
.A2(n_3665),
.B(n_3670),
.Y(n_3776)
);

OAI21x1_ASAP7_75t_L g3777 ( 
.A1(n_3755),
.A2(n_3673),
.B(n_3682),
.Y(n_3777)
);

INVx2_ASAP7_75t_L g3778 ( 
.A(n_3720),
.Y(n_3778)
);

HB1xp67_ASAP7_75t_L g3779 ( 
.A(n_3760),
.Y(n_3779)
);

HB1xp67_ASAP7_75t_L g3780 ( 
.A(n_3734),
.Y(n_3780)
);

AOI21x1_ASAP7_75t_L g3781 ( 
.A1(n_3759),
.A2(n_3675),
.B(n_3666),
.Y(n_3781)
);

AO21x2_ASAP7_75t_L g3782 ( 
.A1(n_3766),
.A2(n_3676),
.B(n_3677),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3717),
.Y(n_3783)
);

HB1xp67_ASAP7_75t_L g3784 ( 
.A(n_3749),
.Y(n_3784)
);

OR2x2_ASAP7_75t_L g3785 ( 
.A(n_3711),
.B(n_3684),
.Y(n_3785)
);

AO21x2_ASAP7_75t_L g3786 ( 
.A1(n_3754),
.A2(n_3683),
.B(n_3663),
.Y(n_3786)
);

OR2x2_ASAP7_75t_L g3787 ( 
.A(n_3711),
.B(n_48),
.Y(n_3787)
);

AND2x2_ASAP7_75t_L g3788 ( 
.A(n_3725),
.B(n_49),
.Y(n_3788)
);

BUFx6f_ASAP7_75t_L g3789 ( 
.A(n_3733),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3753),
.Y(n_3790)
);

AOI21xp5_ASAP7_75t_L g3791 ( 
.A1(n_3712),
.A2(n_3659),
.B(n_3640),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3730),
.Y(n_3792)
);

OAI21x1_ASAP7_75t_L g3793 ( 
.A1(n_3730),
.A2(n_49),
.B(n_50),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3721),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3748),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3727),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3735),
.Y(n_3797)
);

BUFx2_ASAP7_75t_L g3798 ( 
.A(n_3765),
.Y(n_3798)
);

NAND2x1_ASAP7_75t_L g3799 ( 
.A(n_3736),
.B(n_50),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3735),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3739),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3758),
.Y(n_3802)
);

BUFx2_ASAP7_75t_L g3803 ( 
.A(n_3716),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3747),
.Y(n_3804)
);

AND2x2_ASAP7_75t_L g3805 ( 
.A(n_3752),
.B(n_51),
.Y(n_3805)
);

OAI21xp5_ASAP7_75t_L g3806 ( 
.A1(n_3732),
.A2(n_1632),
.B(n_1630),
.Y(n_3806)
);

INVxp67_ASAP7_75t_L g3807 ( 
.A(n_3715),
.Y(n_3807)
);

INVxp67_ASAP7_75t_L g3808 ( 
.A(n_3746),
.Y(n_3808)
);

INVx2_ASAP7_75t_L g3809 ( 
.A(n_3713),
.Y(n_3809)
);

AND2x2_ASAP7_75t_L g3810 ( 
.A(n_3738),
.B(n_52),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3737),
.Y(n_3811)
);

BUFx6f_ASAP7_75t_L g3812 ( 
.A(n_3740),
.Y(n_3812)
);

INVx2_ASAP7_75t_L g3813 ( 
.A(n_3750),
.Y(n_3813)
);

OR2x2_ASAP7_75t_L g3814 ( 
.A(n_3762),
.B(n_53),
.Y(n_3814)
);

INVxp67_ASAP7_75t_R g3815 ( 
.A(n_3722),
.Y(n_3815)
);

AND2x2_ASAP7_75t_L g3816 ( 
.A(n_3714),
.B(n_53),
.Y(n_3816)
);

INVx2_ASAP7_75t_L g3817 ( 
.A(n_3737),
.Y(n_3817)
);

HB1xp67_ASAP7_75t_L g3818 ( 
.A(n_3764),
.Y(n_3818)
);

AND2x2_ASAP7_75t_L g3819 ( 
.A(n_3723),
.B(n_54),
.Y(n_3819)
);

AND2x2_ASAP7_75t_L g3820 ( 
.A(n_3723),
.B(n_55),
.Y(n_3820)
);

OA21x2_ASAP7_75t_L g3821 ( 
.A1(n_3757),
.A2(n_1642),
.B(n_1636),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3761),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3719),
.Y(n_3823)
);

AND2x2_ASAP7_75t_L g3824 ( 
.A(n_3740),
.B(n_3744),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3718),
.Y(n_3825)
);

NOR2x1_ASAP7_75t_L g3826 ( 
.A(n_3767),
.B(n_56),
.Y(n_3826)
);

AOI22xp33_ASAP7_75t_SL g3827 ( 
.A1(n_3771),
.A2(n_3763),
.B1(n_3756),
.B2(n_3724),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3768),
.Y(n_3828)
);

BUFx3_ASAP7_75t_L g3829 ( 
.A(n_3789),
.Y(n_3829)
);

OAI33xp33_ASAP7_75t_L g3830 ( 
.A1(n_3787),
.A2(n_1651),
.A3(n_1649),
.B1(n_1654),
.B2(n_1650),
.B3(n_1648),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_3796),
.B(n_1656),
.Y(n_3831)
);

AO22x1_ASAP7_75t_L g3832 ( 
.A1(n_3789),
.A2(n_1660),
.B1(n_1662),
.B2(n_1658),
.Y(n_3832)
);

OAI21xp33_ASAP7_75t_SL g3833 ( 
.A1(n_3774),
.A2(n_56),
.B(n_57),
.Y(n_3833)
);

BUFx2_ASAP7_75t_L g3834 ( 
.A(n_3803),
.Y(n_3834)
);

BUFx3_ASAP7_75t_L g3835 ( 
.A(n_3812),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_3801),
.B(n_1663),
.Y(n_3836)
);

AOI22xp5_ASAP7_75t_L g3837 ( 
.A1(n_3776),
.A2(n_1665),
.B1(n_1667),
.B2(n_1664),
.Y(n_3837)
);

AOI221xp5_ASAP7_75t_L g3838 ( 
.A1(n_3806),
.A2(n_1674),
.B1(n_1675),
.B2(n_1673),
.C(n_1670),
.Y(n_3838)
);

OAI21x1_ASAP7_75t_L g3839 ( 
.A1(n_3809),
.A2(n_3777),
.B(n_3823),
.Y(n_3839)
);

INVxp67_ASAP7_75t_L g3840 ( 
.A(n_3780),
.Y(n_3840)
);

AND2x2_ASAP7_75t_L g3841 ( 
.A(n_3803),
.B(n_57),
.Y(n_3841)
);

AOI22xp33_ASAP7_75t_SL g3842 ( 
.A1(n_3776),
.A2(n_1679),
.B1(n_1681),
.B2(n_1677),
.Y(n_3842)
);

OAI22xp33_ASAP7_75t_L g3843 ( 
.A1(n_3791),
.A2(n_1683),
.B1(n_1687),
.B2(n_1682),
.Y(n_3843)
);

AOI22xp5_ASAP7_75t_L g3844 ( 
.A1(n_3786),
.A2(n_1690),
.B1(n_1692),
.B2(n_1688),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3772),
.Y(n_3845)
);

OAI22xp5_ASAP7_75t_L g3846 ( 
.A1(n_3769),
.A2(n_1697),
.B1(n_1698),
.B2(n_1696),
.Y(n_3846)
);

INVxp67_ASAP7_75t_L g3847 ( 
.A(n_3779),
.Y(n_3847)
);

AOI22xp33_ASAP7_75t_L g3848 ( 
.A1(n_3821),
.A2(n_1860),
.B1(n_1863),
.B2(n_1858),
.Y(n_3848)
);

AOI222xp33_ASAP7_75t_L g3849 ( 
.A1(n_3808),
.A2(n_1706),
.B1(n_1703),
.B2(n_1709),
.C1(n_1705),
.C2(n_1699),
.Y(n_3849)
);

AND2x2_ASAP7_75t_L g3850 ( 
.A(n_3794),
.B(n_59),
.Y(n_3850)
);

AOI22xp33_ASAP7_75t_SL g3851 ( 
.A1(n_3821),
.A2(n_1715),
.B1(n_1716),
.B2(n_1712),
.Y(n_3851)
);

AOI22xp33_ASAP7_75t_SL g3852 ( 
.A1(n_3822),
.A2(n_1721),
.B1(n_1722),
.B2(n_1719),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_L g3853 ( 
.A(n_3807),
.B(n_1724),
.Y(n_3853)
);

AOI22xp33_ASAP7_75t_L g3854 ( 
.A1(n_3826),
.A2(n_1729),
.B1(n_1730),
.B2(n_1725),
.Y(n_3854)
);

OR2x6_ASAP7_75t_L g3855 ( 
.A(n_3769),
.B(n_59),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3775),
.Y(n_3856)
);

AND2x2_ASAP7_75t_L g3857 ( 
.A(n_3770),
.B(n_60),
.Y(n_3857)
);

OAI21xp5_ASAP7_75t_L g3858 ( 
.A1(n_3781),
.A2(n_1734),
.B(n_1732),
.Y(n_3858)
);

OAI211xp5_ASAP7_75t_L g3859 ( 
.A1(n_3781),
.A2(n_1751),
.B(n_1767),
.C(n_1735),
.Y(n_3859)
);

INVx2_ASAP7_75t_L g3860 ( 
.A(n_3773),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3828),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3856),
.Y(n_3862)
);

AND2x2_ASAP7_75t_L g3863 ( 
.A(n_3834),
.B(n_3798),
.Y(n_3863)
);

AOI22xp33_ASAP7_75t_L g3864 ( 
.A1(n_3827),
.A2(n_3813),
.B1(n_3818),
.B2(n_3782),
.Y(n_3864)
);

OR2x2_ASAP7_75t_L g3865 ( 
.A(n_3840),
.B(n_3792),
.Y(n_3865)
);

INVxp67_ASAP7_75t_SL g3866 ( 
.A(n_3847),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3860),
.Y(n_3867)
);

AND2x4_ASAP7_75t_L g3868 ( 
.A(n_3845),
.B(n_3798),
.Y(n_3868)
);

AND2x2_ASAP7_75t_SL g3869 ( 
.A(n_3837),
.B(n_3824),
.Y(n_3869)
);

BUFx2_ASAP7_75t_L g3870 ( 
.A(n_3855),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3839),
.Y(n_3871)
);

INVx2_ASAP7_75t_L g3872 ( 
.A(n_3850),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3841),
.B(n_3795),
.Y(n_3873)
);

AND2x2_ASAP7_75t_L g3874 ( 
.A(n_3835),
.B(n_3802),
.Y(n_3874)
);

AND2x2_ASAP7_75t_L g3875 ( 
.A(n_3829),
.B(n_3815),
.Y(n_3875)
);

AND2x2_ASAP7_75t_L g3876 ( 
.A(n_3855),
.B(n_3778),
.Y(n_3876)
);

AND2x4_ASAP7_75t_L g3877 ( 
.A(n_3857),
.B(n_3790),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3836),
.Y(n_3878)
);

AND2x2_ASAP7_75t_L g3879 ( 
.A(n_3853),
.B(n_3783),
.Y(n_3879)
);

INVx2_ASAP7_75t_L g3880 ( 
.A(n_3831),
.Y(n_3880)
);

AND2x4_ASAP7_75t_L g3881 ( 
.A(n_3844),
.B(n_3784),
.Y(n_3881)
);

BUFx2_ASAP7_75t_L g3882 ( 
.A(n_3833),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3842),
.B(n_3785),
.Y(n_3883)
);

AND2x4_ASAP7_75t_L g3884 ( 
.A(n_3858),
.B(n_3811),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3846),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3859),
.Y(n_3886)
);

INVx2_ASAP7_75t_SL g3887 ( 
.A(n_3832),
.Y(n_3887)
);

INVx2_ASAP7_75t_L g3888 ( 
.A(n_3830),
.Y(n_3888)
);

INVx3_ASAP7_75t_L g3889 ( 
.A(n_3843),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3854),
.Y(n_3890)
);

INVx2_ASAP7_75t_L g3891 ( 
.A(n_3851),
.Y(n_3891)
);

AOI22xp33_ASAP7_75t_L g3892 ( 
.A1(n_3838),
.A2(n_3817),
.B1(n_3805),
.B2(n_3814),
.Y(n_3892)
);

INVx1_ASAP7_75t_L g3893 ( 
.A(n_3848),
.Y(n_3893)
);

NAND3xp33_ASAP7_75t_L g3894 ( 
.A(n_3864),
.B(n_3893),
.C(n_3889),
.Y(n_3894)
);

INVx2_ASAP7_75t_L g3895 ( 
.A(n_3868),
.Y(n_3895)
);

AND2x2_ASAP7_75t_L g3896 ( 
.A(n_3875),
.B(n_3788),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3862),
.Y(n_3897)
);

AND2x2_ASAP7_75t_L g3898 ( 
.A(n_3863),
.B(n_3812),
.Y(n_3898)
);

HB1xp67_ASAP7_75t_L g3899 ( 
.A(n_3882),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3862),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3861),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_3868),
.Y(n_3902)
);

AND2x4_ASAP7_75t_SL g3903 ( 
.A(n_3876),
.B(n_3819),
.Y(n_3903)
);

NAND2x1p5_ASAP7_75t_L g3904 ( 
.A(n_3870),
.B(n_3799),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3865),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3867),
.Y(n_3906)
);

HB1xp67_ASAP7_75t_L g3907 ( 
.A(n_3866),
.Y(n_3907)
);

OR2x2_ASAP7_75t_L g3908 ( 
.A(n_3873),
.B(n_3872),
.Y(n_3908)
);

AND2x2_ASAP7_75t_L g3909 ( 
.A(n_3879),
.B(n_3820),
.Y(n_3909)
);

HB1xp67_ASAP7_75t_L g3910 ( 
.A(n_3880),
.Y(n_3910)
);

OAI22xp5_ASAP7_75t_L g3911 ( 
.A1(n_3869),
.A2(n_3852),
.B1(n_3825),
.B2(n_3797),
.Y(n_3911)
);

INVx3_ASAP7_75t_SL g3912 ( 
.A(n_3887),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_L g3913 ( 
.A(n_3878),
.B(n_3793),
.Y(n_3913)
);

OAI22xp5_ASAP7_75t_L g3914 ( 
.A1(n_3884),
.A2(n_3800),
.B1(n_3804),
.B2(n_3816),
.Y(n_3914)
);

INVxp67_ASAP7_75t_L g3915 ( 
.A(n_3886),
.Y(n_3915)
);

AND2x2_ASAP7_75t_L g3916 ( 
.A(n_3877),
.B(n_3810),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_L g3917 ( 
.A(n_3881),
.B(n_3849),
.Y(n_3917)
);

AND2x2_ASAP7_75t_L g3918 ( 
.A(n_3877),
.B(n_60),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3871),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3874),
.Y(n_3920)
);

OR2x2_ASAP7_75t_L g3921 ( 
.A(n_3881),
.B(n_61),
.Y(n_3921)
);

AND2x4_ASAP7_75t_SL g3922 ( 
.A(n_3889),
.B(n_3884),
.Y(n_3922)
);

INVxp33_ASAP7_75t_SL g3923 ( 
.A(n_3883),
.Y(n_3923)
);

OR2x2_ASAP7_75t_L g3924 ( 
.A(n_3885),
.B(n_61),
.Y(n_3924)
);

AND2x2_ASAP7_75t_L g3925 ( 
.A(n_3892),
.B(n_3891),
.Y(n_3925)
);

AND2x2_ASAP7_75t_L g3926 ( 
.A(n_3890),
.B(n_63),
.Y(n_3926)
);

OR2x2_ASAP7_75t_L g3927 ( 
.A(n_3888),
.B(n_64),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3866),
.B(n_1736),
.Y(n_3928)
);

OAI22xp33_ASAP7_75t_L g3929 ( 
.A1(n_3899),
.A2(n_1740),
.B1(n_1741),
.B2(n_1738),
.Y(n_3929)
);

OAI221xp5_ASAP7_75t_L g3930 ( 
.A1(n_3911),
.A2(n_1746),
.B1(n_1752),
.B2(n_1743),
.C(n_1742),
.Y(n_3930)
);

AND2x2_ASAP7_75t_L g3931 ( 
.A(n_3912),
.B(n_3922),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_SL g3932 ( 
.A(n_3923),
.B(n_1753),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3897),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_3903),
.Y(n_3934)
);

NAND5xp2_ASAP7_75t_L g3935 ( 
.A(n_3904),
.B(n_68),
.C(n_65),
.D(n_66),
.E(n_70),
.Y(n_3935)
);

OR2x2_ASAP7_75t_L g3936 ( 
.A(n_3907),
.B(n_66),
.Y(n_3936)
);

AO21x2_ASAP7_75t_L g3937 ( 
.A1(n_3894),
.A2(n_3919),
.B(n_3928),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3897),
.Y(n_3938)
);

INVx1_ASAP7_75t_SL g3939 ( 
.A(n_3921),
.Y(n_3939)
);

AND2x2_ASAP7_75t_L g3940 ( 
.A(n_3920),
.B(n_70),
.Y(n_3940)
);

NAND3xp33_ASAP7_75t_L g3941 ( 
.A(n_3917),
.B(n_1879),
.C(n_1758),
.Y(n_3941)
);

INVx2_ASAP7_75t_L g3942 ( 
.A(n_3898),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3900),
.Y(n_3943)
);

INVx1_ASAP7_75t_SL g3944 ( 
.A(n_3924),
.Y(n_3944)
);

AOI22xp33_ASAP7_75t_L g3945 ( 
.A1(n_3925),
.A2(n_1760),
.B1(n_1765),
.B2(n_1756),
.Y(n_3945)
);

AND2x2_ASAP7_75t_L g3946 ( 
.A(n_3895),
.B(n_71),
.Y(n_3946)
);

OAI33xp33_ASAP7_75t_L g3947 ( 
.A1(n_3915),
.A2(n_1773),
.A3(n_1770),
.B1(n_1776),
.B2(n_1772),
.B3(n_1766),
.Y(n_3947)
);

OR2x2_ASAP7_75t_L g3948 ( 
.A(n_3908),
.B(n_71),
.Y(n_3948)
);

AND2x2_ASAP7_75t_L g3949 ( 
.A(n_3902),
.B(n_73),
.Y(n_3949)
);

BUFx2_ASAP7_75t_L g3950 ( 
.A(n_3910),
.Y(n_3950)
);

OR2x2_ASAP7_75t_L g3951 ( 
.A(n_3905),
.B(n_73),
.Y(n_3951)
);

OAI21xp5_ASAP7_75t_SL g3952 ( 
.A1(n_3914),
.A2(n_76),
.B(n_75),
.Y(n_3952)
);

OR2x2_ASAP7_75t_L g3953 ( 
.A(n_3913),
.B(n_74),
.Y(n_3953)
);

OAI22xp33_ASAP7_75t_L g3954 ( 
.A1(n_3901),
.A2(n_1779),
.B1(n_1780),
.B2(n_1777),
.Y(n_3954)
);

AND2x2_ASAP7_75t_L g3955 ( 
.A(n_3916),
.B(n_74),
.Y(n_3955)
);

OAI211xp5_ASAP7_75t_SL g3956 ( 
.A1(n_3927),
.A2(n_1784),
.B(n_1789),
.C(n_1782),
.Y(n_3956)
);

OR2x2_ASAP7_75t_L g3957 ( 
.A(n_3906),
.B(n_75),
.Y(n_3957)
);

AND2x2_ASAP7_75t_L g3958 ( 
.A(n_3896),
.B(n_76),
.Y(n_3958)
);

INVxp67_ASAP7_75t_SL g3959 ( 
.A(n_3906),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_L g3960 ( 
.A(n_3918),
.B(n_1790),
.Y(n_3960)
);

AND2x2_ASAP7_75t_L g3961 ( 
.A(n_3909),
.B(n_77),
.Y(n_3961)
);

BUFx2_ASAP7_75t_L g3962 ( 
.A(n_3931),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3933),
.Y(n_3963)
);

INVx2_ASAP7_75t_SL g3964 ( 
.A(n_3950),
.Y(n_3964)
);

NAND3xp33_ASAP7_75t_SL g3965 ( 
.A(n_3952),
.B(n_3926),
.C(n_3919),
.Y(n_3965)
);

INVx3_ASAP7_75t_L g3966 ( 
.A(n_3942),
.Y(n_3966)
);

NAND4xp75_ASAP7_75t_L g3967 ( 
.A(n_3932),
.B(n_3937),
.C(n_3961),
.D(n_3958),
.Y(n_3967)
);

AND2x4_ASAP7_75t_L g3968 ( 
.A(n_3934),
.B(n_77),
.Y(n_3968)
);

AND2x2_ASAP7_75t_L g3969 ( 
.A(n_3939),
.B(n_3944),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_L g3970 ( 
.A(n_3929),
.B(n_1791),
.Y(n_3970)
);

NAND4xp25_ASAP7_75t_L g3971 ( 
.A(n_3935),
.B(n_3941),
.C(n_3945),
.D(n_3930),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3933),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3955),
.B(n_78),
.Y(n_3973)
);

INVx1_ASAP7_75t_SL g3974 ( 
.A(n_3936),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3938),
.Y(n_3975)
);

AND2x4_ASAP7_75t_L g3976 ( 
.A(n_3959),
.B(n_79),
.Y(n_3976)
);

INVx4_ASAP7_75t_L g3977 ( 
.A(n_3946),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3948),
.B(n_1792),
.Y(n_3978)
);

OR2x2_ASAP7_75t_L g3979 ( 
.A(n_3953),
.B(n_79),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3949),
.B(n_3940),
.Y(n_3980)
);

NAND2xp5_ASAP7_75t_L g3981 ( 
.A(n_3951),
.B(n_1793),
.Y(n_3981)
);

INVx2_ASAP7_75t_L g3982 ( 
.A(n_3943),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3957),
.B(n_1795),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_L g3984 ( 
.A(n_3960),
.B(n_1796),
.Y(n_3984)
);

OR2x2_ASAP7_75t_L g3985 ( 
.A(n_3943),
.B(n_3954),
.Y(n_3985)
);

AOI22xp5_ASAP7_75t_L g3986 ( 
.A1(n_3947),
.A2(n_1799),
.B1(n_1800),
.B2(n_1797),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3956),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_3939),
.B(n_1802),
.Y(n_3988)
);

HB1xp67_ASAP7_75t_L g3989 ( 
.A(n_3950),
.Y(n_3989)
);

HB1xp67_ASAP7_75t_L g3990 ( 
.A(n_3950),
.Y(n_3990)
);

INVx2_ASAP7_75t_SL g3991 ( 
.A(n_3931),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_SL g3992 ( 
.A(n_3931),
.B(n_1805),
.Y(n_3992)
);

AND2x4_ASAP7_75t_L g3993 ( 
.A(n_3931),
.B(n_80),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_3933),
.Y(n_3994)
);

AND2x2_ASAP7_75t_L g3995 ( 
.A(n_3931),
.B(n_80),
.Y(n_3995)
);

OR2x2_ASAP7_75t_L g3996 ( 
.A(n_3939),
.B(n_81),
.Y(n_3996)
);

AND2x2_ASAP7_75t_L g3997 ( 
.A(n_3931),
.B(n_81),
.Y(n_3997)
);

INVx2_ASAP7_75t_L g3998 ( 
.A(n_3931),
.Y(n_3998)
);

OR2x2_ASAP7_75t_L g3999 ( 
.A(n_3939),
.B(n_82),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3933),
.Y(n_4000)
);

AND2x2_ASAP7_75t_L g4001 ( 
.A(n_3931),
.B(n_82),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3939),
.B(n_1806),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3933),
.Y(n_4003)
);

AND2x2_ASAP7_75t_L g4004 ( 
.A(n_3931),
.B(n_84),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3933),
.Y(n_4005)
);

NAND3xp33_ASAP7_75t_L g4006 ( 
.A(n_3952),
.B(n_1808),
.C(n_1807),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_L g4007 ( 
.A(n_3964),
.B(n_3989),
.Y(n_4007)
);

AND2x2_ASAP7_75t_L g4008 ( 
.A(n_3962),
.B(n_84),
.Y(n_4008)
);

AND2x2_ASAP7_75t_L g4009 ( 
.A(n_3962),
.B(n_85),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3990),
.Y(n_4010)
);

OR2x2_ASAP7_75t_L g4011 ( 
.A(n_3974),
.B(n_86),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3969),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3963),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3972),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_3994),
.Y(n_4015)
);

AND2x2_ASAP7_75t_SL g4016 ( 
.A(n_3977),
.B(n_86),
.Y(n_4016)
);

HB1xp67_ASAP7_75t_L g4017 ( 
.A(n_3976),
.Y(n_4017)
);

OR2x2_ASAP7_75t_L g4018 ( 
.A(n_3985),
.B(n_87),
.Y(n_4018)
);

AOI21xp33_ASAP7_75t_L g4019 ( 
.A1(n_3991),
.A2(n_1845),
.B(n_1831),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_4000),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_4003),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_4005),
.Y(n_4022)
);

OR2x2_ASAP7_75t_L g4023 ( 
.A(n_3966),
.B(n_88),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3982),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_L g4025 ( 
.A(n_3980),
.B(n_1809),
.Y(n_4025)
);

INVx2_ASAP7_75t_L g4026 ( 
.A(n_3993),
.Y(n_4026)
);

OR2x2_ASAP7_75t_L g4027 ( 
.A(n_3965),
.B(n_88),
.Y(n_4027)
);

INVx1_ASAP7_75t_SL g4028 ( 
.A(n_3996),
.Y(n_4028)
);

AND2x2_ASAP7_75t_L g4029 ( 
.A(n_3998),
.B(n_89),
.Y(n_4029)
);

NAND2x2_ASAP7_75t_L g4030 ( 
.A(n_3999),
.B(n_89),
.Y(n_4030)
);

OR2x2_ASAP7_75t_L g4031 ( 
.A(n_3979),
.B(n_90),
.Y(n_4031)
);

HB1xp67_ASAP7_75t_L g4032 ( 
.A(n_3976),
.Y(n_4032)
);

BUFx2_ASAP7_75t_L g4033 ( 
.A(n_3995),
.Y(n_4033)
);

OR2x2_ASAP7_75t_L g4034 ( 
.A(n_3967),
.B(n_90),
.Y(n_4034)
);

INVx3_ASAP7_75t_L g4035 ( 
.A(n_3968),
.Y(n_4035)
);

XOR2xp5_ASAP7_75t_L g4036 ( 
.A(n_3971),
.B(n_4006),
.Y(n_4036)
);

NOR2xp33_ASAP7_75t_L g4037 ( 
.A(n_3992),
.B(n_1810),
.Y(n_4037)
);

INVxp67_ASAP7_75t_L g4038 ( 
.A(n_3997),
.Y(n_4038)
);

AND2x2_ASAP7_75t_L g4039 ( 
.A(n_4001),
.B(n_91),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_4004),
.B(n_1813),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_3975),
.Y(n_4041)
);

AND2x2_ASAP7_75t_L g4042 ( 
.A(n_3973),
.B(n_93),
.Y(n_4042)
);

AND2x4_ASAP7_75t_L g4043 ( 
.A(n_3987),
.B(n_94),
.Y(n_4043)
);

AOI211x1_ASAP7_75t_SL g4044 ( 
.A1(n_3988),
.A2(n_96),
.B(n_94),
.C(n_95),
.Y(n_4044)
);

AND2x2_ASAP7_75t_L g4045 ( 
.A(n_4002),
.B(n_95),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3983),
.Y(n_4046)
);

AND2x2_ASAP7_75t_L g4047 ( 
.A(n_3978),
.B(n_96),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_3981),
.Y(n_4048)
);

AND2x2_ASAP7_75t_L g4049 ( 
.A(n_3984),
.B(n_97),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_L g4050 ( 
.A(n_3970),
.B(n_1814),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_3986),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3989),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_L g4053 ( 
.A(n_3964),
.B(n_1816),
.Y(n_4053)
);

AND2x4_ASAP7_75t_L g4054 ( 
.A(n_3962),
.B(n_98),
.Y(n_4054)
);

INVx2_ASAP7_75t_L g4055 ( 
.A(n_3962),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3989),
.Y(n_4056)
);

OR2x2_ASAP7_75t_L g4057 ( 
.A(n_3974),
.B(n_98),
.Y(n_4057)
);

INVx2_ASAP7_75t_SL g4058 ( 
.A(n_3962),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3989),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_3964),
.B(n_1818),
.Y(n_4060)
);

AND2x2_ASAP7_75t_L g4061 ( 
.A(n_3962),
.B(n_99),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_L g4062 ( 
.A(n_3964),
.B(n_1820),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_L g4063 ( 
.A(n_3964),
.B(n_1832),
.Y(n_4063)
);

AND2x2_ASAP7_75t_L g4064 ( 
.A(n_3962),
.B(n_100),
.Y(n_4064)
);

AND2x2_ASAP7_75t_L g4065 ( 
.A(n_3962),
.B(n_101),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_3989),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3964),
.B(n_1833),
.Y(n_4067)
);

INVx2_ASAP7_75t_SL g4068 ( 
.A(n_3962),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_3989),
.Y(n_4069)
);

OR2x2_ASAP7_75t_L g4070 ( 
.A(n_3974),
.B(n_102),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_L g4071 ( 
.A(n_3964),
.B(n_1836),
.Y(n_4071)
);

INVx2_ASAP7_75t_L g4072 ( 
.A(n_4058),
.Y(n_4072)
);

INVx1_ASAP7_75t_SL g4073 ( 
.A(n_4016),
.Y(n_4073)
);

INVx2_ASAP7_75t_L g4074 ( 
.A(n_4068),
.Y(n_4074)
);

CKINVDCx14_ASAP7_75t_R g4075 ( 
.A(n_4033),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_4017),
.Y(n_4076)
);

AND2x4_ASAP7_75t_SL g4077 ( 
.A(n_4035),
.B(n_4026),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_4032),
.Y(n_4078)
);

OAI31xp33_ASAP7_75t_L g4079 ( 
.A1(n_4034),
.A2(n_104),
.A3(n_102),
.B(n_103),
.Y(n_4079)
);

INVx1_ASAP7_75t_SL g4080 ( 
.A(n_4008),
.Y(n_4080)
);

OAI21xp5_ASAP7_75t_L g4081 ( 
.A1(n_4036),
.A2(n_1838),
.B(n_1837),
.Y(n_4081)
);

OAI22xp5_ASAP7_75t_L g4082 ( 
.A1(n_4055),
.A2(n_1843),
.B1(n_1846),
.B2(n_1841),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_L g4083 ( 
.A(n_4009),
.B(n_1849),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_4010),
.Y(n_4084)
);

INVxp33_ASAP7_75t_L g4085 ( 
.A(n_4007),
.Y(n_4085)
);

AOI32xp33_ASAP7_75t_L g4086 ( 
.A1(n_4012),
.A2(n_1857),
.A3(n_1864),
.B1(n_1852),
.B2(n_1850),
.Y(n_4086)
);

OR2x2_ASAP7_75t_L g4087 ( 
.A(n_4018),
.B(n_103),
.Y(n_4087)
);

INVx1_ASAP7_75t_SL g4088 ( 
.A(n_4061),
.Y(n_4088)
);

INVx2_ASAP7_75t_L g4089 ( 
.A(n_4054),
.Y(n_4089)
);

OAI221xp5_ASAP7_75t_L g4090 ( 
.A1(n_4027),
.A2(n_1890),
.B1(n_1873),
.B2(n_1877),
.C(n_1871),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_4052),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_L g4092 ( 
.A(n_4064),
.B(n_1869),
.Y(n_4092)
);

NAND2x1p5_ASAP7_75t_L g4093 ( 
.A(n_4054),
.B(n_104),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_4056),
.Y(n_4094)
);

OAI211xp5_ASAP7_75t_L g4095 ( 
.A1(n_4059),
.A2(n_1880),
.B(n_1893),
.C(n_1878),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_4066),
.Y(n_4096)
);

AOI32xp33_ASAP7_75t_L g4097 ( 
.A1(n_4069),
.A2(n_1907),
.A3(n_1906),
.B1(n_107),
.B2(n_105),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_4065),
.Y(n_4098)
);

INVxp67_ASAP7_75t_L g4099 ( 
.A(n_4011),
.Y(n_4099)
);

O2A1O1Ixp33_ASAP7_75t_L g4100 ( 
.A1(n_4051),
.A2(n_109),
.B(n_105),
.C(n_106),
.Y(n_4100)
);

NOR2x1_ASAP7_75t_L g4101 ( 
.A(n_4057),
.B(n_110),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_L g4102 ( 
.A(n_4028),
.B(n_110),
.Y(n_4102)
);

INVx1_ASAP7_75t_SL g4103 ( 
.A(n_4070),
.Y(n_4103)
);

NOR2x1_ASAP7_75t_L g4104 ( 
.A(n_4023),
.B(n_111),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_4031),
.Y(n_4105)
);

INVx2_ASAP7_75t_L g4106 ( 
.A(n_4043),
.Y(n_4106)
);

AND2x2_ASAP7_75t_L g4107 ( 
.A(n_4038),
.B(n_1032),
.Y(n_4107)
);

OAI32xp33_ASAP7_75t_L g4108 ( 
.A1(n_4044),
.A2(n_4030),
.A3(n_4041),
.B1(n_4015),
.B2(n_4020),
.Y(n_4108)
);

OAI21xp5_ASAP7_75t_L g4109 ( 
.A1(n_4048),
.A2(n_111),
.B(n_112),
.Y(n_4109)
);

INVxp67_ASAP7_75t_SL g4110 ( 
.A(n_4040),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_L g4111 ( 
.A(n_4029),
.B(n_112),
.Y(n_4111)
);

OAI21xp33_ASAP7_75t_L g4112 ( 
.A1(n_4046),
.A2(n_113),
.B(n_115),
.Y(n_4112)
);

AOI22xp5_ASAP7_75t_L g4113 ( 
.A1(n_4025),
.A2(n_4043),
.B1(n_4024),
.B2(n_4039),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_4013),
.Y(n_4114)
);

INVx2_ASAP7_75t_SL g4115 ( 
.A(n_4042),
.Y(n_4115)
);

AND2x2_ASAP7_75t_L g4116 ( 
.A(n_4049),
.B(n_1034),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_L g4117 ( 
.A(n_4047),
.B(n_113),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_4014),
.Y(n_4118)
);

INVx2_ASAP7_75t_L g4119 ( 
.A(n_4021),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_4022),
.Y(n_4120)
);

OAI21xp5_ASAP7_75t_L g4121 ( 
.A1(n_4050),
.A2(n_115),
.B(n_116),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_4045),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_4053),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_4060),
.Y(n_4124)
);

OR2x2_ASAP7_75t_L g4125 ( 
.A(n_4062),
.B(n_117),
.Y(n_4125)
);

OAI21xp33_ASAP7_75t_L g4126 ( 
.A1(n_4063),
.A2(n_118),
.B(n_119),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_4067),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_4071),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_4037),
.Y(n_4129)
);

OAI21xp5_ASAP7_75t_L g4130 ( 
.A1(n_4019),
.A2(n_118),
.B(n_120),
.Y(n_4130)
);

AOI221xp5_ASAP7_75t_L g4131 ( 
.A1(n_4010),
.A2(n_123),
.B1(n_120),
.B2(n_122),
.C(n_124),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_4017),
.Y(n_4132)
);

OAI221xp5_ASAP7_75t_L g4133 ( 
.A1(n_4034),
.A2(n_125),
.B1(n_122),
.B2(n_124),
.C(n_127),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_4017),
.Y(n_4134)
);

INVx1_ASAP7_75t_L g4135 ( 
.A(n_4017),
.Y(n_4135)
);

OAI32xp33_ASAP7_75t_L g4136 ( 
.A1(n_4034),
.A2(n_130),
.A3(n_127),
.B1(n_129),
.B2(n_131),
.Y(n_4136)
);

AND2x2_ASAP7_75t_L g4137 ( 
.A(n_4033),
.B(n_1032),
.Y(n_4137)
);

INVx2_ASAP7_75t_L g4138 ( 
.A(n_4058),
.Y(n_4138)
);

O2A1O1Ixp33_ASAP7_75t_L g4139 ( 
.A1(n_4034),
.A2(n_133),
.B(n_131),
.C(n_132),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_4017),
.Y(n_4140)
);

OAI21xp5_ASAP7_75t_L g4141 ( 
.A1(n_4034),
.A2(n_132),
.B(n_134),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_4017),
.Y(n_4142)
);

AOI21xp5_ASAP7_75t_L g4143 ( 
.A1(n_4036),
.A2(n_135),
.B(n_136),
.Y(n_4143)
);

AOI22xp5_ASAP7_75t_L g4144 ( 
.A1(n_4036),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_4017),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_4017),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_4017),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_4017),
.Y(n_4148)
);

AOI32xp33_ASAP7_75t_L g4149 ( 
.A1(n_4034),
.A2(n_139),
.A3(n_137),
.B1(n_138),
.B2(n_140),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_4017),
.Y(n_4150)
);

INVx2_ASAP7_75t_L g4151 ( 
.A(n_4058),
.Y(n_4151)
);

AND2x4_ASAP7_75t_L g4152 ( 
.A(n_4058),
.B(n_140),
.Y(n_4152)
);

NAND3xp33_ASAP7_75t_SL g4153 ( 
.A(n_4034),
.B(n_138),
.C(n_141),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_4017),
.Y(n_4154)
);

HB1xp67_ASAP7_75t_L g4155 ( 
.A(n_4058),
.Y(n_4155)
);

INVx2_ASAP7_75t_L g4156 ( 
.A(n_4058),
.Y(n_4156)
);

NOR2xp33_ASAP7_75t_L g4157 ( 
.A(n_4035),
.B(n_1024),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_4017),
.Y(n_4158)
);

OAI22xp5_ASAP7_75t_L g4159 ( 
.A1(n_4075),
.A2(n_144),
.B1(n_141),
.B2(n_143),
.Y(n_4159)
);

AND2x2_ASAP7_75t_L g4160 ( 
.A(n_4073),
.B(n_143),
.Y(n_4160)
);

INVxp67_ASAP7_75t_L g4161 ( 
.A(n_4155),
.Y(n_4161)
);

OAI211xp5_ASAP7_75t_SL g4162 ( 
.A1(n_4099),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_4077),
.B(n_146),
.Y(n_4163)
);

BUFx2_ASAP7_75t_L g4164 ( 
.A(n_4152),
.Y(n_4164)
);

OAI322xp33_ASAP7_75t_L g4165 ( 
.A1(n_4084),
.A2(n_156),
.A3(n_153),
.B1(n_151),
.B2(n_149),
.C1(n_150),
.C2(n_152),
.Y(n_4165)
);

INVx2_ASAP7_75t_L g4166 ( 
.A(n_4093),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_4076),
.Y(n_4167)
);

INVxp67_ASAP7_75t_SL g4168 ( 
.A(n_4101),
.Y(n_4168)
);

OR2x2_ASAP7_75t_L g4169 ( 
.A(n_4080),
.B(n_149),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_4078),
.Y(n_4170)
);

NOR2xp33_ASAP7_75t_L g4171 ( 
.A(n_4085),
.B(n_150),
.Y(n_4171)
);

AOI21xp5_ASAP7_75t_L g4172 ( 
.A1(n_4139),
.A2(n_151),
.B(n_153),
.Y(n_4172)
);

AOI21xp33_ASAP7_75t_SL g4173 ( 
.A1(n_4115),
.A2(n_156),
.B(n_157),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4132),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_4088),
.B(n_157),
.Y(n_4175)
);

OAI21xp5_ASAP7_75t_SL g4176 ( 
.A1(n_4113),
.A2(n_1023),
.B(n_1022),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_4134),
.Y(n_4177)
);

OAI21xp5_ASAP7_75t_L g4178 ( 
.A1(n_4143),
.A2(n_158),
.B(n_161),
.Y(n_4178)
);

HB1xp67_ASAP7_75t_L g4179 ( 
.A(n_4152),
.Y(n_4179)
);

HB1xp67_ASAP7_75t_L g4180 ( 
.A(n_4104),
.Y(n_4180)
);

AOI22xp5_ASAP7_75t_L g4181 ( 
.A1(n_4153),
.A2(n_165),
.B1(n_162),
.B2(n_164),
.Y(n_4181)
);

INVx1_ASAP7_75t_SL g4182 ( 
.A(n_4137),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_L g4183 ( 
.A(n_4106),
.B(n_164),
.Y(n_4183)
);

AOI32xp33_ASAP7_75t_L g4184 ( 
.A1(n_4072),
.A2(n_4138),
.A3(n_4156),
.B1(n_4151),
.B2(n_4074),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_4135),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_4140),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_4142),
.Y(n_4187)
);

AOI22xp5_ASAP7_75t_SL g4188 ( 
.A1(n_4158),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_4188)
);

AND2x2_ASAP7_75t_L g4189 ( 
.A(n_4089),
.B(n_166),
.Y(n_4189)
);

AOI21xp5_ASAP7_75t_L g4190 ( 
.A1(n_4141),
.A2(n_167),
.B(n_168),
.Y(n_4190)
);

NOR2xp33_ASAP7_75t_L g4191 ( 
.A(n_4103),
.B(n_168),
.Y(n_4191)
);

AOI22x1_ASAP7_75t_L g4192 ( 
.A1(n_4098),
.A2(n_172),
.B1(n_169),
.B2(n_171),
.Y(n_4192)
);

OR2x2_ASAP7_75t_L g4193 ( 
.A(n_4145),
.B(n_169),
.Y(n_4193)
);

OAI22xp5_ASAP7_75t_L g4194 ( 
.A1(n_4144),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_4194)
);

OAI21xp33_ASAP7_75t_SL g4195 ( 
.A1(n_4146),
.A2(n_174),
.B(n_175),
.Y(n_4195)
);

OAI21x1_ASAP7_75t_SL g4196 ( 
.A1(n_4147),
.A2(n_175),
.B(n_177),
.Y(n_4196)
);

OAI22xp33_ASAP7_75t_L g4197 ( 
.A1(n_4133),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_4197)
);

NOR2xp33_ASAP7_75t_L g4198 ( 
.A(n_4108),
.B(n_178),
.Y(n_4198)
);

OR2x2_ASAP7_75t_L g4199 ( 
.A(n_4148),
.B(n_179),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4150),
.Y(n_4200)
);

AND2x2_ASAP7_75t_L g4201 ( 
.A(n_4154),
.B(n_180),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_L g4202 ( 
.A(n_4149),
.B(n_182),
.Y(n_4202)
);

NAND2xp5_ASAP7_75t_L g4203 ( 
.A(n_4122),
.B(n_183),
.Y(n_4203)
);

INVx2_ASAP7_75t_L g4204 ( 
.A(n_4116),
.Y(n_4204)
);

O2A1O1Ixp33_ASAP7_75t_SL g4205 ( 
.A1(n_4136),
.A2(n_187),
.B(n_184),
.C(n_185),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_4107),
.Y(n_4206)
);

OAI221xp5_ASAP7_75t_L g4207 ( 
.A1(n_4079),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.C(n_191),
.Y(n_4207)
);

NOR2xp33_ASAP7_75t_L g4208 ( 
.A(n_4105),
.B(n_189),
.Y(n_4208)
);

NOR2xp33_ASAP7_75t_L g4209 ( 
.A(n_4102),
.B(n_190),
.Y(n_4209)
);

OAI321xp33_ASAP7_75t_L g4210 ( 
.A1(n_4091),
.A2(n_193),
.A3(n_195),
.B1(n_191),
.B2(n_192),
.C(n_194),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_4087),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_4111),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_4117),
.Y(n_4213)
);

INVx2_ASAP7_75t_SL g4214 ( 
.A(n_4094),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_4096),
.Y(n_4215)
);

OAI21xp33_ASAP7_75t_L g4216 ( 
.A1(n_4110),
.A2(n_193),
.B(n_195),
.Y(n_4216)
);

AOI21xp33_ASAP7_75t_L g4217 ( 
.A1(n_4123),
.A2(n_1021),
.B(n_1020),
.Y(n_4217)
);

OAI21xp33_ASAP7_75t_L g4218 ( 
.A1(n_4124),
.A2(n_198),
.B(n_199),
.Y(n_4218)
);

INVx2_ASAP7_75t_SL g4219 ( 
.A(n_4119),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4157),
.Y(n_4220)
);

NAND2xp5_ASAP7_75t_L g4221 ( 
.A(n_4097),
.B(n_198),
.Y(n_4221)
);

OAI321xp33_ASAP7_75t_L g4222 ( 
.A1(n_4114),
.A2(n_4120),
.A3(n_4118),
.B1(n_4109),
.B2(n_4127),
.C(n_4131),
.Y(n_4222)
);

AND2x4_ASAP7_75t_L g4223 ( 
.A(n_4128),
.B(n_199),
.Y(n_4223)
);

OR2x2_ASAP7_75t_L g4224 ( 
.A(n_4129),
.B(n_4083),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_4125),
.Y(n_4225)
);

OR2x2_ASAP7_75t_L g4226 ( 
.A(n_4092),
.B(n_200),
.Y(n_4226)
);

INVx2_ASAP7_75t_L g4227 ( 
.A(n_4090),
.Y(n_4227)
);

AOI21xp33_ASAP7_75t_L g4228 ( 
.A1(n_4095),
.A2(n_1030),
.B(n_1029),
.Y(n_4228)
);

AND2x2_ASAP7_75t_L g4229 ( 
.A(n_4121),
.B(n_200),
.Y(n_4229)
);

AND2x2_ASAP7_75t_L g4230 ( 
.A(n_4130),
.B(n_201),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4112),
.Y(n_4231)
);

NOR2xp33_ASAP7_75t_SL g4232 ( 
.A(n_4126),
.B(n_203),
.Y(n_4232)
);

AOI222xp33_ASAP7_75t_L g4233 ( 
.A1(n_4081),
.A2(n_233),
.B1(n_214),
.B2(n_245),
.C1(n_223),
.C2(n_203),
.Y(n_4233)
);

OAI22xp33_ASAP7_75t_SL g4234 ( 
.A1(n_4082),
.A2(n_1035),
.B1(n_1034),
.B2(n_207),
.Y(n_4234)
);

INVx1_ASAP7_75t_SL g4235 ( 
.A(n_4100),
.Y(n_4235)
);

AND2x2_ASAP7_75t_L g4236 ( 
.A(n_4086),
.B(n_204),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_4155),
.Y(n_4237)
);

XOR2x2_ASAP7_75t_L g4238 ( 
.A(n_4101),
.B(n_206),
.Y(n_4238)
);

A2O1A1Ixp33_ASAP7_75t_L g4239 ( 
.A1(n_4139),
.A2(n_208),
.B(n_206),
.C(n_207),
.Y(n_4239)
);

INVx2_ASAP7_75t_SL g4240 ( 
.A(n_4155),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_4155),
.Y(n_4241)
);

AOI22xp33_ASAP7_75t_SL g4242 ( 
.A1(n_4075),
.A2(n_211),
.B1(n_208),
.B2(n_209),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_4155),
.Y(n_4243)
);

OAI221xp5_ASAP7_75t_L g4244 ( 
.A1(n_4073),
.A2(n_214),
.B1(n_209),
.B2(n_213),
.C(n_215),
.Y(n_4244)
);

INVx2_ASAP7_75t_SL g4245 ( 
.A(n_4155),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_4155),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4155),
.Y(n_4247)
);

INVx1_ASAP7_75t_L g4248 ( 
.A(n_4155),
.Y(n_4248)
);

OAI211xp5_ASAP7_75t_L g4249 ( 
.A1(n_4075),
.A2(n_218),
.B(n_215),
.C(n_217),
.Y(n_4249)
);

AOI21xp5_ASAP7_75t_L g4250 ( 
.A1(n_4073),
.A2(n_217),
.B(n_218),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_4073),
.B(n_219),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_4155),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_SL g4253 ( 
.A(n_4073),
.B(n_220),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_4155),
.Y(n_4254)
);

AND2x2_ASAP7_75t_L g4255 ( 
.A(n_4075),
.B(n_220),
.Y(n_4255)
);

OAI22xp33_ASAP7_75t_L g4256 ( 
.A1(n_4085),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_4073),
.B(n_224),
.Y(n_4257)
);

OAI32xp33_ASAP7_75t_L g4258 ( 
.A1(n_4073),
.A2(n_226),
.A3(n_229),
.B1(n_225),
.B2(n_228),
.Y(n_4258)
);

OAI21xp5_ASAP7_75t_L g4259 ( 
.A1(n_4139),
.A2(n_224),
.B(n_226),
.Y(n_4259)
);

INVx2_ASAP7_75t_L g4260 ( 
.A(n_4093),
.Y(n_4260)
);

AOI21xp5_ASAP7_75t_L g4261 ( 
.A1(n_4073),
.A2(n_228),
.B(n_230),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4155),
.Y(n_4262)
);

AOI221xp5_ASAP7_75t_L g4263 ( 
.A1(n_4108),
.A2(n_255),
.B1(n_263),
.B2(n_244),
.C(n_231),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_4155),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_L g4265 ( 
.A(n_4073),
.B(n_231),
.Y(n_4265)
);

NAND4xp25_ASAP7_75t_L g4266 ( 
.A(n_4080),
.B(n_237),
.C(n_233),
.D(n_235),
.Y(n_4266)
);

AOI21xp33_ASAP7_75t_SL g4267 ( 
.A1(n_4155),
.A2(n_235),
.B(n_238),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4155),
.Y(n_4268)
);

OAI322xp33_ASAP7_75t_L g4269 ( 
.A1(n_4075),
.A2(n_248),
.A3(n_246),
.B1(n_243),
.B2(n_239),
.C1(n_241),
.C2(n_244),
.Y(n_4269)
);

OAI21xp5_ASAP7_75t_L g4270 ( 
.A1(n_4139),
.A2(n_243),
.B(n_248),
.Y(n_4270)
);

NOR2xp33_ASAP7_75t_L g4271 ( 
.A(n_4073),
.B(n_249),
.Y(n_4271)
);

AND2x2_ASAP7_75t_L g4272 ( 
.A(n_4075),
.B(n_249),
.Y(n_4272)
);

INVxp67_ASAP7_75t_L g4273 ( 
.A(n_4155),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_4073),
.B(n_250),
.Y(n_4274)
);

INVxp67_ASAP7_75t_L g4275 ( 
.A(n_4155),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_L g4276 ( 
.A(n_4073),
.B(n_251),
.Y(n_4276)
);

AOI21xp33_ASAP7_75t_SL g4277 ( 
.A1(n_4155),
.A2(n_251),
.B(n_252),
.Y(n_4277)
);

INVx2_ASAP7_75t_L g4278 ( 
.A(n_4093),
.Y(n_4278)
);

NAND3xp33_ASAP7_75t_L g4279 ( 
.A(n_4075),
.B(n_252),
.C(n_254),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_4155),
.Y(n_4280)
);

OR2x2_ASAP7_75t_L g4281 ( 
.A(n_4073),
.B(n_254),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4155),
.Y(n_4282)
);

NOR2xp33_ASAP7_75t_L g4283 ( 
.A(n_4073),
.B(n_255),
.Y(n_4283)
);

A2O1A1Ixp33_ASAP7_75t_L g4284 ( 
.A1(n_4139),
.A2(n_258),
.B(n_256),
.C(n_257),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4155),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_L g4286 ( 
.A(n_4073),
.B(n_256),
.Y(n_4286)
);

INVxp67_ASAP7_75t_SL g4287 ( 
.A(n_4155),
.Y(n_4287)
);

INVx2_ASAP7_75t_L g4288 ( 
.A(n_4093),
.Y(n_4288)
);

INVx2_ASAP7_75t_SL g4289 ( 
.A(n_4155),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_L g4290 ( 
.A(n_4073),
.B(n_257),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4155),
.Y(n_4291)
);

INVxp67_ASAP7_75t_L g4292 ( 
.A(n_4155),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4155),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_4155),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_4073),
.B(n_258),
.Y(n_4295)
);

AOI21xp5_ASAP7_75t_SL g4296 ( 
.A1(n_4139),
.A2(n_259),
.B(n_260),
.Y(n_4296)
);

AOI22xp33_ASAP7_75t_L g4297 ( 
.A1(n_4075),
.A2(n_262),
.B1(n_259),
.B2(n_261),
.Y(n_4297)
);

INVx2_ASAP7_75t_L g4298 ( 
.A(n_4093),
.Y(n_4298)
);

OR2x6_ASAP7_75t_L g4299 ( 
.A(n_4093),
.B(n_264),
.Y(n_4299)
);

OAI22xp33_ASAP7_75t_L g4300 ( 
.A1(n_4085),
.A2(n_267),
.B1(n_261),
.B2(n_266),
.Y(n_4300)
);

AND2x2_ASAP7_75t_L g4301 ( 
.A(n_4075),
.B(n_268),
.Y(n_4301)
);

INVx2_ASAP7_75t_L g4302 ( 
.A(n_4093),
.Y(n_4302)
);

NAND2xp5_ASAP7_75t_SL g4303 ( 
.A(n_4073),
.B(n_268),
.Y(n_4303)
);

NOR3xp33_ASAP7_75t_L g4304 ( 
.A(n_4073),
.B(n_269),
.C(n_270),
.Y(n_4304)
);

OAI321xp33_ASAP7_75t_L g4305 ( 
.A1(n_4076),
.A2(n_272),
.A3(n_274),
.B1(n_269),
.B2(n_271),
.C(n_273),
.Y(n_4305)
);

AO22x1_ASAP7_75t_L g4306 ( 
.A1(n_4101),
.A2(n_274),
.B1(n_271),
.B2(n_273),
.Y(n_4306)
);

INVxp67_ASAP7_75t_L g4307 ( 
.A(n_4155),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_SL g4308 ( 
.A(n_4073),
.B(n_275),
.Y(n_4308)
);

AOI22xp5_ASAP7_75t_L g4309 ( 
.A1(n_4198),
.A2(n_1029),
.B1(n_1030),
.B2(n_1027),
.Y(n_4309)
);

OAI31xp33_ASAP7_75t_L g4310 ( 
.A1(n_4249),
.A2(n_279),
.A3(n_276),
.B(n_277),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4179),
.Y(n_4311)
);

AOI22xp33_ASAP7_75t_L g4312 ( 
.A1(n_4263),
.A2(n_279),
.B1(n_276),
.B2(n_277),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4164),
.Y(n_4313)
);

AOI322xp5_ASAP7_75t_L g4314 ( 
.A1(n_4235),
.A2(n_286),
.A3(n_285),
.B1(n_283),
.B2(n_280),
.C1(n_281),
.C2(n_284),
.Y(n_4314)
);

AND2x2_ASAP7_75t_L g4315 ( 
.A(n_4255),
.B(n_280),
.Y(n_4315)
);

AND2x2_ASAP7_75t_L g4316 ( 
.A(n_4272),
.B(n_281),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4180),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4287),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_L g4319 ( 
.A(n_4301),
.B(n_284),
.Y(n_4319)
);

AOI22xp5_ASAP7_75t_L g4320 ( 
.A1(n_4240),
.A2(n_1015),
.B1(n_1016),
.B2(n_1013),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_4245),
.B(n_288),
.Y(n_4321)
);

AOI22xp5_ASAP7_75t_L g4322 ( 
.A1(n_4289),
.A2(n_1016),
.B1(n_1017),
.B2(n_1015),
.Y(n_4322)
);

OAI221xp5_ASAP7_75t_SL g4323 ( 
.A1(n_4184),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.C(n_291),
.Y(n_4323)
);

O2A1O1Ixp33_ASAP7_75t_SL g4324 ( 
.A1(n_4239),
.A2(n_294),
.B(n_291),
.C(n_293),
.Y(n_4324)
);

AOI22xp33_ASAP7_75t_SL g4325 ( 
.A1(n_4168),
.A2(n_4237),
.B1(n_4243),
.B2(n_4241),
.Y(n_4325)
);

OAI22xp5_ASAP7_75t_L g4326 ( 
.A1(n_4161),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_4306),
.B(n_296),
.Y(n_4327)
);

INVxp67_ASAP7_75t_L g4328 ( 
.A(n_4299),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4160),
.Y(n_4329)
);

AND2x2_ASAP7_75t_L g4330 ( 
.A(n_4166),
.B(n_298),
.Y(n_4330)
);

AO221x1_ASAP7_75t_L g4331 ( 
.A1(n_4273),
.A2(n_302),
.B1(n_299),
.B2(n_301),
.C(n_303),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_4281),
.Y(n_4332)
);

OAI211xp5_ASAP7_75t_L g4333 ( 
.A1(n_4296),
.A2(n_4292),
.B(n_4275),
.C(n_4307),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_L g4334 ( 
.A(n_4242),
.B(n_299),
.Y(n_4334)
);

OAI32xp33_ASAP7_75t_L g4335 ( 
.A1(n_4195),
.A2(n_318),
.A3(n_329),
.B1(n_309),
.B2(n_301),
.Y(n_4335)
);

OAI221xp5_ASAP7_75t_L g4336 ( 
.A1(n_4259),
.A2(n_1012),
.B1(n_1018),
.B2(n_1010),
.C(n_1009),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_4246),
.Y(n_4337)
);

OAI21xp5_ASAP7_75t_SL g4338 ( 
.A1(n_4182),
.A2(n_302),
.B(n_303),
.Y(n_4338)
);

AND2x2_ASAP7_75t_L g4339 ( 
.A(n_4260),
.B(n_304),
.Y(n_4339)
);

AOI21xp5_ASAP7_75t_L g4340 ( 
.A1(n_4222),
.A2(n_305),
.B(n_306),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_4247),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_4248),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_4252),
.B(n_305),
.Y(n_4343)
);

AOI22xp5_ASAP7_75t_L g4344 ( 
.A1(n_4254),
.A2(n_1031),
.B1(n_1033),
.B2(n_1026),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_4262),
.Y(n_4345)
);

AND2x2_ASAP7_75t_L g4346 ( 
.A(n_4278),
.B(n_4288),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4264),
.Y(n_4347)
);

AND2x2_ASAP7_75t_L g4348 ( 
.A(n_4298),
.B(n_307),
.Y(n_4348)
);

INVxp67_ASAP7_75t_L g4349 ( 
.A(n_4299),
.Y(n_4349)
);

OAI211xp5_ASAP7_75t_SL g4350 ( 
.A1(n_4225),
.A2(n_4211),
.B(n_4212),
.C(n_4213),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4268),
.Y(n_4351)
);

AOI32xp33_ASAP7_75t_L g4352 ( 
.A1(n_4304),
.A2(n_312),
.A3(n_308),
.B1(n_311),
.B2(n_313),
.Y(n_4352)
);

AOI22xp33_ASAP7_75t_L g4353 ( 
.A1(n_4280),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.Y(n_4353)
);

AOI32xp33_ASAP7_75t_L g4354 ( 
.A1(n_4282),
.A2(n_316),
.A3(n_314),
.B1(n_315),
.B2(n_317),
.Y(n_4354)
);

INVx1_ASAP7_75t_SL g4355 ( 
.A(n_4238),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4285),
.Y(n_4356)
);

OR2x6_ASAP7_75t_L g4357 ( 
.A(n_4163),
.B(n_315),
.Y(n_4357)
);

NAND2xp5_ASAP7_75t_L g4358 ( 
.A(n_4291),
.B(n_316),
.Y(n_4358)
);

OAI21xp33_ASAP7_75t_L g4359 ( 
.A1(n_4293),
.A2(n_318),
.B(n_319),
.Y(n_4359)
);

INVx2_ASAP7_75t_L g4360 ( 
.A(n_4302),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_L g4361 ( 
.A(n_4294),
.B(n_320),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_4189),
.Y(n_4362)
);

INVx1_ASAP7_75t_SL g4363 ( 
.A(n_4188),
.Y(n_4363)
);

AOI22xp5_ASAP7_75t_L g4364 ( 
.A1(n_4232),
.A2(n_1010),
.B1(n_1012),
.B2(n_1009),
.Y(n_4364)
);

OAI321xp33_ASAP7_75t_L g4365 ( 
.A1(n_4167),
.A2(n_323),
.A3(n_326),
.B1(n_320),
.B2(n_322),
.C(n_325),
.Y(n_4365)
);

AND2x2_ASAP7_75t_L g4366 ( 
.A(n_4204),
.B(n_322),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_L g4367 ( 
.A(n_4267),
.B(n_323),
.Y(n_4367)
);

NOR2xp33_ASAP7_75t_L g4368 ( 
.A(n_4253),
.B(n_325),
.Y(n_4368)
);

OAI22xp5_ASAP7_75t_L g4369 ( 
.A1(n_4181),
.A2(n_333),
.B1(n_328),
.B2(n_332),
.Y(n_4369)
);

INVxp67_ASAP7_75t_SL g4370 ( 
.A(n_4303),
.Y(n_4370)
);

OAI22xp33_ASAP7_75t_L g4371 ( 
.A1(n_4266),
.A2(n_4202),
.B1(n_4305),
.B2(n_4221),
.Y(n_4371)
);

AOI22xp5_ASAP7_75t_L g4372 ( 
.A1(n_4231),
.A2(n_999),
.B1(n_1000),
.B2(n_997),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_L g4373 ( 
.A(n_4277),
.B(n_4271),
.Y(n_4373)
);

AOI211xp5_ASAP7_75t_L g4374 ( 
.A1(n_4269),
.A2(n_342),
.B(n_351),
.C(n_332),
.Y(n_4374)
);

OR2x2_ASAP7_75t_L g4375 ( 
.A(n_4169),
.B(n_334),
.Y(n_4375)
);

AND2x2_ASAP7_75t_L g4376 ( 
.A(n_4206),
.B(n_334),
.Y(n_4376)
);

AOI221xp5_ASAP7_75t_L g4377 ( 
.A1(n_4205),
.A2(n_1006),
.B1(n_1007),
.B2(n_1005),
.C(n_1004),
.Y(n_4377)
);

INVxp67_ASAP7_75t_L g4378 ( 
.A(n_4283),
.Y(n_4378)
);

O2A1O1Ixp5_ASAP7_75t_L g4379 ( 
.A1(n_4170),
.A2(n_338),
.B(n_336),
.C(n_337),
.Y(n_4379)
);

INVx2_ASAP7_75t_L g4380 ( 
.A(n_4223),
.Y(n_4380)
);

AOI21xp33_ASAP7_75t_L g4381 ( 
.A1(n_4220),
.A2(n_336),
.B(n_337),
.Y(n_4381)
);

AND2x2_ASAP7_75t_L g4382 ( 
.A(n_4201),
.B(n_338),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_4251),
.Y(n_4383)
);

OAI21xp33_ASAP7_75t_SL g4384 ( 
.A1(n_4214),
.A2(n_339),
.B(n_340),
.Y(n_4384)
);

AOI21xp33_ASAP7_75t_L g4385 ( 
.A1(n_4227),
.A2(n_339),
.B(n_341),
.Y(n_4385)
);

INVxp67_ASAP7_75t_SL g4386 ( 
.A(n_4308),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4257),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_L g4388 ( 
.A(n_4173),
.B(n_343),
.Y(n_4388)
);

AOI22xp5_ASAP7_75t_L g4389 ( 
.A1(n_4279),
.A2(n_1035),
.B1(n_1031),
.B2(n_345),
.Y(n_4389)
);

AOI21xp33_ASAP7_75t_SL g4390 ( 
.A1(n_4171),
.A2(n_1026),
.B(n_343),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4265),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4274),
.Y(n_4392)
);

OAI22xp5_ASAP7_75t_L g4393 ( 
.A1(n_4297),
.A2(n_346),
.B1(n_344),
.B2(n_345),
.Y(n_4393)
);

INVx2_ASAP7_75t_L g4394 ( 
.A(n_4223),
.Y(n_4394)
);

OAI221xp5_ASAP7_75t_L g4395 ( 
.A1(n_4270),
.A2(n_996),
.B1(n_1000),
.B2(n_995),
.C(n_992),
.Y(n_4395)
);

OAI21xp33_ASAP7_75t_SL g4396 ( 
.A1(n_4219),
.A2(n_347),
.B(n_349),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4276),
.Y(n_4397)
);

OAI221xp5_ASAP7_75t_L g4398 ( 
.A1(n_4176),
.A2(n_1007),
.B1(n_1008),
.B2(n_1006),
.C(n_1004),
.Y(n_4398)
);

INVx2_ASAP7_75t_L g4399 ( 
.A(n_4193),
.Y(n_4399)
);

NAND2xp5_ASAP7_75t_L g4400 ( 
.A(n_4250),
.B(n_347),
.Y(n_4400)
);

AOI222xp33_ASAP7_75t_L g4401 ( 
.A1(n_4178),
.A2(n_352),
.B1(n_354),
.B2(n_350),
.C1(n_351),
.C2(n_353),
.Y(n_4401)
);

NOR2xp33_ASAP7_75t_L g4402 ( 
.A(n_4286),
.B(n_350),
.Y(n_4402)
);

OAI21xp5_ASAP7_75t_L g4403 ( 
.A1(n_4172),
.A2(n_355),
.B(n_354),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_L g4404 ( 
.A(n_4261),
.B(n_352),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4290),
.Y(n_4405)
);

AOI22xp5_ASAP7_75t_L g4406 ( 
.A1(n_4191),
.A2(n_982),
.B1(n_983),
.B2(n_981),
.Y(n_4406)
);

AND2x2_ASAP7_75t_L g4407 ( 
.A(n_4174),
.B(n_355),
.Y(n_4407)
);

NAND2xp5_ASAP7_75t_L g4408 ( 
.A(n_4177),
.B(n_356),
.Y(n_4408)
);

INVxp67_ASAP7_75t_L g4409 ( 
.A(n_4196),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4295),
.Y(n_4410)
);

INVx1_ASAP7_75t_SL g4411 ( 
.A(n_4199),
.Y(n_4411)
);

AOI22xp5_ASAP7_75t_L g4412 ( 
.A1(n_4185),
.A2(n_986),
.B1(n_987),
.B2(n_983),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4183),
.Y(n_4413)
);

BUFx3_ASAP7_75t_L g4414 ( 
.A(n_4186),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_L g4415 ( 
.A(n_4187),
.B(n_356),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4175),
.Y(n_4416)
);

INVx2_ASAP7_75t_SL g4417 ( 
.A(n_4200),
.Y(n_4417)
);

OAI21xp5_ASAP7_75t_SL g4418 ( 
.A1(n_4233),
.A2(n_357),
.B(n_360),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_L g4419 ( 
.A(n_4159),
.B(n_360),
.Y(n_4419)
);

AND2x2_ASAP7_75t_SL g4420 ( 
.A(n_4224),
.B(n_361),
.Y(n_4420)
);

AOI221xp5_ASAP7_75t_L g4421 ( 
.A1(n_4210),
.A2(n_991),
.B1(n_1002),
.B2(n_990),
.C(n_989),
.Y(n_4421)
);

OAI22xp5_ASAP7_75t_L g4422 ( 
.A1(n_4284),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_4422)
);

INVx2_ASAP7_75t_L g4423 ( 
.A(n_4192),
.Y(n_4423)
);

NAND2xp5_ASAP7_75t_L g4424 ( 
.A(n_4229),
.B(n_362),
.Y(n_4424)
);

INVxp67_ASAP7_75t_SL g4425 ( 
.A(n_4256),
.Y(n_4425)
);

OAI21xp5_ASAP7_75t_L g4426 ( 
.A1(n_4190),
.A2(n_366),
.B(n_365),
.Y(n_4426)
);

OAI21xp5_ASAP7_75t_L g4427 ( 
.A1(n_4244),
.A2(n_368),
.B(n_365),
.Y(n_4427)
);

OAI221xp5_ASAP7_75t_SL g4428 ( 
.A1(n_4333),
.A2(n_4215),
.B1(n_4207),
.B2(n_4216),
.C(n_4197),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_L g4429 ( 
.A(n_4363),
.B(n_4208),
.Y(n_4429)
);

NAND2xp33_ASAP7_75t_L g4430 ( 
.A(n_4318),
.B(n_4218),
.Y(n_4430)
);

OAI21xp5_ASAP7_75t_SL g4431 ( 
.A1(n_4325),
.A2(n_4228),
.B(n_4162),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_L g4432 ( 
.A(n_4313),
.B(n_4236),
.Y(n_4432)
);

OAI221xp5_ASAP7_75t_L g4433 ( 
.A1(n_4340),
.A2(n_4203),
.B1(n_4194),
.B2(n_4217),
.C(n_4209),
.Y(n_4433)
);

NOR3xp33_ASAP7_75t_L g4434 ( 
.A(n_4350),
.B(n_4234),
.C(n_4230),
.Y(n_4434)
);

OAI21xp5_ASAP7_75t_SL g4435 ( 
.A1(n_4418),
.A2(n_4300),
.B(n_4226),
.Y(n_4435)
);

NAND4xp25_ASAP7_75t_L g4436 ( 
.A(n_4355),
.B(n_4346),
.C(n_4311),
.D(n_4329),
.Y(n_4436)
);

NOR3xp33_ASAP7_75t_L g4437 ( 
.A(n_4328),
.B(n_4165),
.C(n_4258),
.Y(n_4437)
);

OAI32xp33_ASAP7_75t_L g4438 ( 
.A1(n_4423),
.A2(n_370),
.A3(n_372),
.B1(n_369),
.B2(n_371),
.Y(n_4438)
);

AOI221x1_ASAP7_75t_L g4439 ( 
.A1(n_4317),
.A2(n_370),
.B1(n_363),
.B2(n_369),
.C(n_371),
.Y(n_4439)
);

O2A1O1Ixp33_ASAP7_75t_L g4440 ( 
.A1(n_4323),
.A2(n_375),
.B(n_372),
.C(n_374),
.Y(n_4440)
);

AO21x1_ASAP7_75t_L g4441 ( 
.A1(n_4327),
.A2(n_1018),
.B(n_980),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_SL g4442 ( 
.A(n_4377),
.B(n_375),
.Y(n_4442)
);

A2O1A1Ixp33_ASAP7_75t_L g4443 ( 
.A1(n_4310),
.A2(n_388),
.B(n_399),
.C(n_377),
.Y(n_4443)
);

AOI21xp5_ASAP7_75t_L g4444 ( 
.A1(n_4400),
.A2(n_377),
.B(n_379),
.Y(n_4444)
);

NAND3x1_ASAP7_75t_L g4445 ( 
.A(n_4309),
.B(n_4367),
.C(n_4379),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_4315),
.Y(n_4446)
);

NAND3xp33_ASAP7_75t_L g4447 ( 
.A(n_4374),
.B(n_379),
.C(n_381),
.Y(n_4447)
);

AOI32xp33_ASAP7_75t_L g4448 ( 
.A1(n_4371),
.A2(n_385),
.A3(n_382),
.B1(n_384),
.B2(n_386),
.Y(n_4448)
);

AOI21xp33_ASAP7_75t_L g4449 ( 
.A1(n_4349),
.A2(n_385),
.B(n_387),
.Y(n_4449)
);

NAND3x1_ASAP7_75t_L g4450 ( 
.A(n_4388),
.B(n_387),
.C(n_388),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_4316),
.Y(n_4451)
);

AOI222xp33_ASAP7_75t_L g4452 ( 
.A1(n_4425),
.A2(n_392),
.B1(n_395),
.B2(n_389),
.C1(n_390),
.C2(n_393),
.Y(n_4452)
);

AOI211xp5_ASAP7_75t_L g4453 ( 
.A1(n_4409),
.A2(n_979),
.B(n_981),
.C(n_978),
.Y(n_4453)
);

XNOR2xp5_ASAP7_75t_L g4454 ( 
.A(n_4364),
.B(n_389),
.Y(n_4454)
);

OAI21xp33_ASAP7_75t_L g4455 ( 
.A1(n_4373),
.A2(n_393),
.B(n_397),
.Y(n_4455)
);

NAND2xp5_ASAP7_75t_L g4456 ( 
.A(n_4420),
.B(n_398),
.Y(n_4456)
);

NOR2xp33_ASAP7_75t_L g4457 ( 
.A(n_4380),
.B(n_399),
.Y(n_4457)
);

OAI211xp5_ASAP7_75t_L g4458 ( 
.A1(n_4421),
.A2(n_4396),
.B(n_4384),
.C(n_4312),
.Y(n_4458)
);

INVx2_ASAP7_75t_L g4459 ( 
.A(n_4394),
.Y(n_4459)
);

OR2x2_ASAP7_75t_L g4460 ( 
.A(n_4360),
.B(n_400),
.Y(n_4460)
);

OAI21xp33_ASAP7_75t_L g4461 ( 
.A1(n_4370),
.A2(n_401),
.B(n_402),
.Y(n_4461)
);

OAI211xp5_ASAP7_75t_L g4462 ( 
.A1(n_4386),
.A2(n_405),
.B(n_402),
.C(n_404),
.Y(n_4462)
);

AOI222xp33_ASAP7_75t_L g4463 ( 
.A1(n_4337),
.A2(n_407),
.B1(n_409),
.B2(n_404),
.C1(n_406),
.C2(n_408),
.Y(n_4463)
);

AOI311xp33_ASAP7_75t_L g4464 ( 
.A1(n_4341),
.A2(n_408),
.A3(n_406),
.B(n_407),
.C(n_411),
.Y(n_4464)
);

OAI21xp33_ASAP7_75t_L g4465 ( 
.A1(n_4378),
.A2(n_411),
.B(n_412),
.Y(n_4465)
);

AOI311xp33_ASAP7_75t_L g4466 ( 
.A1(n_4342),
.A2(n_416),
.A3(n_412),
.B(n_414),
.C(n_417),
.Y(n_4466)
);

AOI221xp5_ASAP7_75t_L g4467 ( 
.A1(n_4345),
.A2(n_418),
.B1(n_414),
.B2(n_417),
.C(n_419),
.Y(n_4467)
);

OAI21xp5_ASAP7_75t_SL g4468 ( 
.A1(n_4338),
.A2(n_418),
.B(n_420),
.Y(n_4468)
);

AOI221xp5_ASAP7_75t_L g4469 ( 
.A1(n_4347),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.C(n_423),
.Y(n_4469)
);

OAI21xp33_ASAP7_75t_SL g4470 ( 
.A1(n_4411),
.A2(n_422),
.B(n_424),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_L g4471 ( 
.A(n_4331),
.B(n_424),
.Y(n_4471)
);

AOI211xp5_ASAP7_75t_L g4472 ( 
.A1(n_4335),
.A2(n_972),
.B(n_973),
.C(n_970),
.Y(n_4472)
);

OAI22xp33_ASAP7_75t_L g4473 ( 
.A1(n_4334),
.A2(n_429),
.B1(n_426),
.B2(n_427),
.Y(n_4473)
);

AOI221xp5_ASAP7_75t_L g4474 ( 
.A1(n_4351),
.A2(n_429),
.B1(n_426),
.B2(n_427),
.C(n_430),
.Y(n_4474)
);

AOI221xp5_ASAP7_75t_L g4475 ( 
.A1(n_4356),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.C(n_434),
.Y(n_4475)
);

NAND2xp5_ASAP7_75t_SL g4476 ( 
.A(n_4352),
.B(n_431),
.Y(n_4476)
);

NAND4xp25_ASAP7_75t_L g4477 ( 
.A(n_4362),
.B(n_437),
.C(n_435),
.D(n_436),
.Y(n_4477)
);

OAI21xp33_ASAP7_75t_L g4478 ( 
.A1(n_4332),
.A2(n_4414),
.B(n_4387),
.Y(n_4478)
);

OAI211xp5_ASAP7_75t_L g4479 ( 
.A1(n_4314),
.A2(n_437),
.B(n_435),
.C(n_436),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_4319),
.Y(n_4480)
);

NAND2xp5_ASAP7_75t_L g4481 ( 
.A(n_4382),
.B(n_438),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_L g4482 ( 
.A(n_4330),
.B(n_438),
.Y(n_4482)
);

AOI222xp33_ASAP7_75t_L g4483 ( 
.A1(n_4427),
.A2(n_442),
.B1(n_448),
.B2(n_439),
.C1(n_441),
.C2(n_445),
.Y(n_4483)
);

AOI311xp33_ASAP7_75t_L g4484 ( 
.A1(n_4383),
.A2(n_451),
.A3(n_449),
.B(n_450),
.C(n_452),
.Y(n_4484)
);

INVx2_ASAP7_75t_SL g4485 ( 
.A(n_4339),
.Y(n_4485)
);

AOI22xp33_ASAP7_75t_SL g4486 ( 
.A1(n_4417),
.A2(n_451),
.B1(n_449),
.B2(n_450),
.Y(n_4486)
);

OAI211xp5_ASAP7_75t_L g4487 ( 
.A1(n_4401),
.A2(n_456),
.B(n_452),
.C(n_453),
.Y(n_4487)
);

OAI221xp5_ASAP7_75t_SL g4488 ( 
.A1(n_4391),
.A2(n_987),
.B1(n_988),
.B2(n_986),
.C(n_979),
.Y(n_4488)
);

AOI222xp33_ASAP7_75t_L g4489 ( 
.A1(n_4403),
.A2(n_459),
.B1(n_462),
.B2(n_457),
.C1(n_458),
.C2(n_460),
.Y(n_4489)
);

NOR3xp33_ASAP7_75t_L g4490 ( 
.A(n_4392),
.B(n_459),
.C(n_465),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_4348),
.Y(n_4491)
);

AOI22xp33_ASAP7_75t_L g4492 ( 
.A1(n_4397),
.A2(n_468),
.B1(n_466),
.B2(n_467),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_4366),
.Y(n_4493)
);

AOI21xp5_ASAP7_75t_L g4494 ( 
.A1(n_4404),
.A2(n_466),
.B(n_467),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_4321),
.Y(n_4495)
);

AOI22xp5_ASAP7_75t_L g4496 ( 
.A1(n_4405),
.A2(n_470),
.B1(n_468),
.B2(n_469),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_4375),
.Y(n_4497)
);

OAI22xp33_ASAP7_75t_L g4498 ( 
.A1(n_4389),
.A2(n_472),
.B1(n_469),
.B2(n_471),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_4376),
.B(n_4354),
.Y(n_4499)
);

AOI21xp5_ASAP7_75t_L g4500 ( 
.A1(n_4324),
.A2(n_471),
.B(n_473),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4407),
.Y(n_4501)
);

AOI21xp33_ASAP7_75t_SL g4502 ( 
.A1(n_4422),
.A2(n_476),
.B(n_475),
.Y(n_4502)
);

NAND2xp5_ASAP7_75t_SL g4503 ( 
.A(n_4390),
.B(n_474),
.Y(n_4503)
);

OAI22xp33_ASAP7_75t_L g4504 ( 
.A1(n_4365),
.A2(n_479),
.B1(n_477),
.B2(n_478),
.Y(n_4504)
);

OAI21xp33_ASAP7_75t_SL g4505 ( 
.A1(n_4410),
.A2(n_477),
.B(n_478),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4357),
.Y(n_4506)
);

OAI21x1_ASAP7_75t_L g4507 ( 
.A1(n_4399),
.A2(n_1019),
.B(n_1008),
.Y(n_4507)
);

A2O1A1Ixp33_ASAP7_75t_L g4508 ( 
.A1(n_4426),
.A2(n_489),
.B(n_499),
.C(n_479),
.Y(n_4508)
);

NOR3xp33_ASAP7_75t_L g4509 ( 
.A(n_4416),
.B(n_480),
.C(n_481),
.Y(n_4509)
);

NAND3xp33_ASAP7_75t_L g4510 ( 
.A(n_4343),
.B(n_480),
.C(n_481),
.Y(n_4510)
);

AND2x2_ASAP7_75t_L g4511 ( 
.A(n_4357),
.B(n_483),
.Y(n_4511)
);

AOI221xp5_ASAP7_75t_L g4512 ( 
.A1(n_4385),
.A2(n_487),
.B1(n_484),
.B2(n_485),
.C(n_488),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_4358),
.Y(n_4513)
);

AOI21xp5_ASAP7_75t_L g4514 ( 
.A1(n_4424),
.A2(n_484),
.B(n_488),
.Y(n_4514)
);

O2A1O1Ixp5_ASAP7_75t_L g4515 ( 
.A1(n_4413),
.A2(n_491),
.B(n_489),
.C(n_490),
.Y(n_4515)
);

AOI221xp5_ASAP7_75t_L g4516 ( 
.A1(n_4336),
.A2(n_492),
.B1(n_490),
.B2(n_491),
.C(n_493),
.Y(n_4516)
);

INVx1_ASAP7_75t_SL g4517 ( 
.A(n_4419),
.Y(n_4517)
);

NAND4xp75_ASAP7_75t_L g4518 ( 
.A(n_4361),
.B(n_496),
.C(n_493),
.D(n_495),
.Y(n_4518)
);

AOI21xp5_ASAP7_75t_L g4519 ( 
.A1(n_4408),
.A2(n_496),
.B(n_497),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_4415),
.Y(n_4520)
);

NOR2xp33_ASAP7_75t_L g4521 ( 
.A(n_4359),
.B(n_500),
.Y(n_4521)
);

AOI221xp5_ASAP7_75t_L g4522 ( 
.A1(n_4395),
.A2(n_503),
.B1(n_500),
.B2(n_501),
.C(n_504),
.Y(n_4522)
);

NAND4xp25_ASAP7_75t_L g4523 ( 
.A(n_4398),
.B(n_1019),
.C(n_508),
.D(n_501),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4368),
.Y(n_4524)
);

AND2x2_ASAP7_75t_L g4525 ( 
.A(n_4402),
.B(n_507),
.Y(n_4525)
);

AOI21xp33_ASAP7_75t_L g4526 ( 
.A1(n_4369),
.A2(n_507),
.B(n_509),
.Y(n_4526)
);

NAND4xp75_ASAP7_75t_L g4527 ( 
.A(n_4372),
.B(n_512),
.C(n_510),
.D(n_511),
.Y(n_4527)
);

AOI22xp33_ASAP7_75t_L g4528 ( 
.A1(n_4393),
.A2(n_515),
.B1(n_512),
.B2(n_514),
.Y(n_4528)
);

AOI322xp5_ASAP7_75t_L g4529 ( 
.A1(n_4353),
.A2(n_1002),
.A3(n_523),
.B1(n_518),
.B2(n_521),
.C1(n_516),
.C2(n_517),
.Y(n_4529)
);

NAND3xp33_ASAP7_75t_L g4530 ( 
.A(n_4381),
.B(n_517),
.C(n_520),
.Y(n_4530)
);

NOR3xp33_ASAP7_75t_L g4531 ( 
.A(n_4326),
.B(n_521),
.C(n_524),
.Y(n_4531)
);

OAI22xp5_ASAP7_75t_L g4532 ( 
.A1(n_4320),
.A2(n_526),
.B1(n_524),
.B2(n_525),
.Y(n_4532)
);

AOI221xp5_ASAP7_75t_L g4533 ( 
.A1(n_4406),
.A2(n_528),
.B1(n_525),
.B2(n_526),
.C(n_530),
.Y(n_4533)
);

OAI211xp5_ASAP7_75t_SL g4534 ( 
.A1(n_4322),
.A2(n_531),
.B(n_528),
.C(n_530),
.Y(n_4534)
);

OAI21xp33_ASAP7_75t_L g4535 ( 
.A1(n_4344),
.A2(n_532),
.B(n_535),
.Y(n_4535)
);

AOI22xp5_ASAP7_75t_L g4536 ( 
.A1(n_4412),
.A2(n_538),
.B1(n_532),
.B2(n_536),
.Y(n_4536)
);

OAI211xp5_ASAP7_75t_SL g4537 ( 
.A1(n_4325),
.A2(n_541),
.B(n_538),
.C(n_539),
.Y(n_4537)
);

OAI21xp33_ASAP7_75t_L g4538 ( 
.A1(n_4355),
.A2(n_539),
.B(n_542),
.Y(n_4538)
);

AOI22xp5_ASAP7_75t_L g4539 ( 
.A1(n_4363),
.A2(n_544),
.B1(n_542),
.B2(n_543),
.Y(n_4539)
);

AOI22xp5_ASAP7_75t_L g4540 ( 
.A1(n_4363),
.A2(n_547),
.B1(n_544),
.B2(n_545),
.Y(n_4540)
);

AOI21xp33_ASAP7_75t_L g4541 ( 
.A1(n_4328),
.A2(n_545),
.B(n_547),
.Y(n_4541)
);

NAND3xp33_ASAP7_75t_L g4542 ( 
.A(n_4325),
.B(n_548),
.C(n_550),
.Y(n_4542)
);

OAI211xp5_ASAP7_75t_SL g4543 ( 
.A1(n_4325),
.A2(n_553),
.B(n_551),
.C(n_552),
.Y(n_4543)
);

OAI21xp33_ASAP7_75t_L g4544 ( 
.A1(n_4355),
.A2(n_554),
.B(n_555),
.Y(n_4544)
);

OAI321xp33_ASAP7_75t_L g4545 ( 
.A1(n_4313),
.A2(n_556),
.A3(n_561),
.B1(n_554),
.B2(n_555),
.C(n_558),
.Y(n_4545)
);

AOI21xp5_ASAP7_75t_L g4546 ( 
.A1(n_4340),
.A2(n_561),
.B(n_562),
.Y(n_4546)
);

A2O1A1Ixp33_ASAP7_75t_L g4547 ( 
.A1(n_4340),
.A2(n_568),
.B(n_566),
.C(n_567),
.Y(n_4547)
);

NOR2xp33_ASAP7_75t_L g4548 ( 
.A(n_4409),
.B(n_567),
.Y(n_4548)
);

AOI222xp33_ASAP7_75t_L g4549 ( 
.A1(n_4355),
.A2(n_574),
.B1(n_576),
.B2(n_568),
.C1(n_569),
.C2(n_575),
.Y(n_4549)
);

NAND2xp5_ASAP7_75t_L g4550 ( 
.A(n_4363),
.B(n_574),
.Y(n_4550)
);

AOI21xp33_ASAP7_75t_L g4551 ( 
.A1(n_4328),
.A2(n_575),
.B(n_577),
.Y(n_4551)
);

OAI22xp5_ASAP7_75t_L g4552 ( 
.A1(n_4312),
.A2(n_581),
.B1(n_578),
.B2(n_580),
.Y(n_4552)
);

AOI221xp5_ASAP7_75t_L g4553 ( 
.A1(n_4371),
.A2(n_583),
.B1(n_580),
.B2(n_582),
.C(n_584),
.Y(n_4553)
);

OAI211xp5_ASAP7_75t_L g4554 ( 
.A1(n_4333),
.A2(n_586),
.B(n_584),
.C(n_585),
.Y(n_4554)
);

INVx3_ASAP7_75t_SL g4555 ( 
.A(n_4420),
.Y(n_4555)
);

AND2x2_ASAP7_75t_L g4556 ( 
.A(n_4363),
.B(n_585),
.Y(n_4556)
);

NOR2xp33_ASAP7_75t_L g4557 ( 
.A(n_4409),
.B(n_586),
.Y(n_4557)
);

AOI22xp5_ASAP7_75t_L g4558 ( 
.A1(n_4363),
.A2(n_590),
.B1(n_587),
.B2(n_589),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_4363),
.B(n_589),
.Y(n_4559)
);

OAI221xp5_ASAP7_75t_SL g4560 ( 
.A1(n_4333),
.A2(n_592),
.B1(n_590),
.B2(n_591),
.C(n_593),
.Y(n_4560)
);

OAI221xp5_ASAP7_75t_L g4561 ( 
.A1(n_4325),
.A2(n_593),
.B1(n_591),
.B2(n_592),
.C(n_596),
.Y(n_4561)
);

NAND2xp5_ASAP7_75t_SL g4562 ( 
.A(n_4377),
.B(n_597),
.Y(n_4562)
);

O2A1O1Ixp33_ASAP7_75t_L g4563 ( 
.A1(n_4340),
.A2(n_599),
.B(n_597),
.C(n_598),
.Y(n_4563)
);

NAND2xp5_ASAP7_75t_L g4564 ( 
.A(n_4363),
.B(n_600),
.Y(n_4564)
);

NOR3xp33_ASAP7_75t_L g4565 ( 
.A(n_4333),
.B(n_600),
.C(n_601),
.Y(n_4565)
);

AOI322xp5_ASAP7_75t_L g4566 ( 
.A1(n_4371),
.A2(n_990),
.A3(n_607),
.B1(n_603),
.B2(n_606),
.C1(n_601),
.C2(n_602),
.Y(n_4566)
);

AOI22xp5_ASAP7_75t_L g4567 ( 
.A1(n_4363),
.A2(n_606),
.B1(n_602),
.B2(n_605),
.Y(n_4567)
);

OAI311xp33_ASAP7_75t_L g4568 ( 
.A1(n_4418),
.A2(n_609),
.A3(n_607),
.B1(n_608),
.C1(n_610),
.Y(n_4568)
);

AOI21xp5_ASAP7_75t_L g4569 ( 
.A1(n_4340),
.A2(n_608),
.B(n_609),
.Y(n_4569)
);

AOI221x1_ASAP7_75t_L g4570 ( 
.A1(n_4340),
.A2(n_613),
.B1(n_611),
.B2(n_612),
.C(n_615),
.Y(n_4570)
);

AOI22xp5_ASAP7_75t_L g4571 ( 
.A1(n_4363),
.A2(n_616),
.B1(n_611),
.B2(n_613),
.Y(n_4571)
);

AOI322xp5_ASAP7_75t_L g4572 ( 
.A1(n_4371),
.A2(n_623),
.A3(n_622),
.B1(n_620),
.B2(n_618),
.C1(n_619),
.C2(n_621),
.Y(n_4572)
);

OAI32xp33_ASAP7_75t_L g4573 ( 
.A1(n_4363),
.A2(n_622),
.A3(n_619),
.B1(n_621),
.B2(n_623),
.Y(n_4573)
);

AOI322xp5_ASAP7_75t_L g4574 ( 
.A1(n_4371),
.A2(n_631),
.A3(n_629),
.B1(n_626),
.B2(n_624),
.C1(n_625),
.C2(n_627),
.Y(n_4574)
);

NAND3xp33_ASAP7_75t_L g4575 ( 
.A(n_4325),
.B(n_625),
.C(n_627),
.Y(n_4575)
);

AOI21xp5_ASAP7_75t_L g4576 ( 
.A1(n_4340),
.A2(n_632),
.B(n_633),
.Y(n_4576)
);

OAI211xp5_ASAP7_75t_L g4577 ( 
.A1(n_4431),
.A2(n_634),
.B(n_632),
.C(n_633),
.Y(n_4577)
);

OAI221xp5_ASAP7_75t_L g4578 ( 
.A1(n_4565),
.A2(n_638),
.B1(n_635),
.B2(n_637),
.C(n_639),
.Y(n_4578)
);

NOR3xp33_ASAP7_75t_L g4579 ( 
.A(n_4436),
.B(n_635),
.C(n_638),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_4556),
.Y(n_4580)
);

AOI221xp5_ASAP7_75t_L g4581 ( 
.A1(n_4560),
.A2(n_641),
.B1(n_639),
.B2(n_640),
.C(n_642),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_L g4582 ( 
.A(n_4555),
.B(n_644),
.Y(n_4582)
);

OAI211xp5_ASAP7_75t_L g4583 ( 
.A1(n_4554),
.A2(n_646),
.B(n_644),
.C(n_645),
.Y(n_4583)
);

A2O1A1Ixp33_ASAP7_75t_L g4584 ( 
.A1(n_4563),
.A2(n_988),
.B(n_647),
.C(n_645),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4511),
.Y(n_4585)
);

AOI21xp33_ASAP7_75t_L g4586 ( 
.A1(n_4506),
.A2(n_976),
.B(n_646),
.Y(n_4586)
);

AOI21xp33_ASAP7_75t_L g4587 ( 
.A1(n_4429),
.A2(n_647),
.B(n_648),
.Y(n_4587)
);

AND2x2_ASAP7_75t_L g4588 ( 
.A(n_4459),
.B(n_4446),
.Y(n_4588)
);

NAND4xp25_ASAP7_75t_SL g4589 ( 
.A(n_4458),
.B(n_650),
.C(n_648),
.D(n_649),
.Y(n_4589)
);

OAI22xp5_ASAP7_75t_L g4590 ( 
.A1(n_4539),
.A2(n_653),
.B1(n_651),
.B2(n_652),
.Y(n_4590)
);

AOI221xp5_ASAP7_75t_SL g4591 ( 
.A1(n_4430),
.A2(n_654),
.B1(n_652),
.B2(n_653),
.C(n_657),
.Y(n_4591)
);

OAI22xp5_ASAP7_75t_L g4592 ( 
.A1(n_4540),
.A2(n_659),
.B1(n_654),
.B2(n_658),
.Y(n_4592)
);

INVx1_ASAP7_75t_L g4593 ( 
.A(n_4550),
.Y(n_4593)
);

AOI21xp5_ASAP7_75t_L g4594 ( 
.A1(n_4503),
.A2(n_659),
.B(n_660),
.Y(n_4594)
);

NAND3xp33_ASAP7_75t_L g4595 ( 
.A(n_4542),
.B(n_976),
.C(n_660),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_4559),
.Y(n_4596)
);

NOR2x1_ASAP7_75t_L g4597 ( 
.A(n_4575),
.B(n_662),
.Y(n_4597)
);

AOI21xp5_ASAP7_75t_L g4598 ( 
.A1(n_4500),
.A2(n_665),
.B(n_666),
.Y(n_4598)
);

NOR4xp25_ASAP7_75t_L g4599 ( 
.A(n_4428),
.B(n_670),
.C(n_668),
.D(n_669),
.Y(n_4599)
);

AOI21xp33_ASAP7_75t_L g4600 ( 
.A1(n_4478),
.A2(n_975),
.B(n_668),
.Y(n_4600)
);

INVx1_ASAP7_75t_SL g4601 ( 
.A(n_4456),
.Y(n_4601)
);

OAI21xp33_ASAP7_75t_SL g4602 ( 
.A1(n_4452),
.A2(n_669),
.B(n_671),
.Y(n_4602)
);

INVxp67_ASAP7_75t_L g4603 ( 
.A(n_4548),
.Y(n_4603)
);

INVx1_ASAP7_75t_L g4604 ( 
.A(n_4564),
.Y(n_4604)
);

INVxp33_ASAP7_75t_L g4605 ( 
.A(n_4437),
.Y(n_4605)
);

AOI22xp5_ASAP7_75t_L g4606 ( 
.A1(n_4434),
.A2(n_673),
.B1(n_671),
.B2(n_672),
.Y(n_4606)
);

AOI221xp5_ASAP7_75t_L g4607 ( 
.A1(n_4504),
.A2(n_975),
.B1(n_678),
.B2(n_673),
.C(n_676),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4451),
.Y(n_4608)
);

NAND2xp5_ASAP7_75t_L g4609 ( 
.A(n_4485),
.B(n_676),
.Y(n_4609)
);

O2A1O1Ixp5_ASAP7_75t_L g4610 ( 
.A1(n_4568),
.A2(n_680),
.B(n_678),
.C(n_679),
.Y(n_4610)
);

INVx2_ASAP7_75t_SL g4611 ( 
.A(n_4460),
.Y(n_4611)
);

OAI31xp33_ASAP7_75t_SL g4612 ( 
.A1(n_4537),
.A2(n_681),
.A3(n_679),
.B(n_680),
.Y(n_4612)
);

OAI221xp5_ASAP7_75t_L g4613 ( 
.A1(n_4448),
.A2(n_684),
.B1(n_682),
.B2(n_683),
.C(n_685),
.Y(n_4613)
);

AOI221xp5_ASAP7_75t_L g4614 ( 
.A1(n_4543),
.A2(n_974),
.B1(n_685),
.B2(n_682),
.C(n_684),
.Y(n_4614)
);

OAI21xp5_ASAP7_75t_L g4615 ( 
.A1(n_4470),
.A2(n_4569),
.B(n_4546),
.Y(n_4615)
);

AOI21xp5_ASAP7_75t_L g4616 ( 
.A1(n_4444),
.A2(n_687),
.B(n_688),
.Y(n_4616)
);

NOR3xp33_ASAP7_75t_L g4617 ( 
.A(n_4433),
.B(n_973),
.C(n_687),
.Y(n_4617)
);

INVxp67_ASAP7_75t_L g4618 ( 
.A(n_4557),
.Y(n_4618)
);

OAI21xp5_ASAP7_75t_L g4619 ( 
.A1(n_4576),
.A2(n_688),
.B(n_690),
.Y(n_4619)
);

NAND2xp5_ASAP7_75t_L g4620 ( 
.A(n_4486),
.B(n_690),
.Y(n_4620)
);

INVx1_ASAP7_75t_L g4621 ( 
.A(n_4507),
.Y(n_4621)
);

NOR2x1_ASAP7_75t_L g4622 ( 
.A(n_4518),
.B(n_4462),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_4441),
.Y(n_4623)
);

OA211x2_ASAP7_75t_L g4624 ( 
.A1(n_4538),
.A2(n_693),
.B(n_691),
.C(n_692),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4482),
.Y(n_4625)
);

NOR2xp33_ASAP7_75t_L g4626 ( 
.A(n_4561),
.B(n_691),
.Y(n_4626)
);

NAND2x1_ASAP7_75t_L g4627 ( 
.A(n_4497),
.B(n_694),
.Y(n_4627)
);

OR2x2_ASAP7_75t_L g4628 ( 
.A(n_4499),
.B(n_694),
.Y(n_4628)
);

NAND2xp5_ASAP7_75t_L g4629 ( 
.A(n_4549),
.B(n_4566),
.Y(n_4629)
);

AND2x2_ASAP7_75t_L g4630 ( 
.A(n_4491),
.B(n_695),
.Y(n_4630)
);

AOI22xp5_ASAP7_75t_SL g4631 ( 
.A1(n_4471),
.A2(n_698),
.B1(n_696),
.B2(n_697),
.Y(n_4631)
);

INVxp67_ASAP7_75t_SL g4632 ( 
.A(n_4450),
.Y(n_4632)
);

AOI21xp5_ASAP7_75t_L g4633 ( 
.A1(n_4494),
.A2(n_696),
.B(n_697),
.Y(n_4633)
);

AOI21xp5_ASAP7_75t_L g4634 ( 
.A1(n_4442),
.A2(n_698),
.B(n_700),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4481),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4432),
.Y(n_4636)
);

AND2x2_ASAP7_75t_L g4637 ( 
.A(n_4501),
.B(n_701),
.Y(n_4637)
);

NAND2x1_ASAP7_75t_L g4638 ( 
.A(n_4493),
.B(n_703),
.Y(n_4638)
);

OAI21xp33_ASAP7_75t_L g4639 ( 
.A1(n_4435),
.A2(n_704),
.B(n_705),
.Y(n_4639)
);

NOR2x1_ASAP7_75t_L g4640 ( 
.A(n_4477),
.B(n_705),
.Y(n_4640)
);

OAI21xp33_ASAP7_75t_L g4641 ( 
.A1(n_4476),
.A2(n_706),
.B(n_707),
.Y(n_4641)
);

A2O1A1Ixp33_ASAP7_75t_L g4642 ( 
.A1(n_4440),
.A2(n_709),
.B(n_706),
.C(n_707),
.Y(n_4642)
);

AND2x2_ASAP7_75t_L g4643 ( 
.A(n_4558),
.B(n_710),
.Y(n_4643)
);

AOI22xp33_ASAP7_75t_SL g4644 ( 
.A1(n_4479),
.A2(n_712),
.B1(n_710),
.B2(n_711),
.Y(n_4644)
);

INVx1_ASAP7_75t_L g4645 ( 
.A(n_4525),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_4572),
.B(n_711),
.Y(n_4646)
);

INVxp67_ASAP7_75t_L g4647 ( 
.A(n_4457),
.Y(n_4647)
);

OAI21xp5_ASAP7_75t_L g4648 ( 
.A1(n_4547),
.A2(n_713),
.B(n_714),
.Y(n_4648)
);

OAI22xp33_ASAP7_75t_L g4649 ( 
.A1(n_4567),
.A2(n_717),
.B1(n_714),
.B2(n_715),
.Y(n_4649)
);

INVx1_ASAP7_75t_L g4650 ( 
.A(n_4571),
.Y(n_4650)
);

AOI211xp5_ASAP7_75t_L g4651 ( 
.A1(n_4487),
.A2(n_721),
.B(n_717),
.C(n_718),
.Y(n_4651)
);

AOI222xp33_ASAP7_75t_L g4652 ( 
.A1(n_4562),
.A2(n_722),
.B1(n_724),
.B2(n_718),
.C1(n_721),
.C2(n_723),
.Y(n_4652)
);

A2O1A1Ixp33_ASAP7_75t_L g4653 ( 
.A1(n_4515),
.A2(n_972),
.B(n_725),
.C(n_723),
.Y(n_4653)
);

HB1xp67_ASAP7_75t_L g4654 ( 
.A(n_4505),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4573),
.Y(n_4655)
);

NAND2xp5_ASAP7_75t_L g4656 ( 
.A(n_4574),
.B(n_724),
.Y(n_4656)
);

OAI211xp5_ASAP7_75t_L g4657 ( 
.A1(n_4570),
.A2(n_4468),
.B(n_4439),
.C(n_4553),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4454),
.Y(n_4658)
);

NAND2x1_ASAP7_75t_SL g4659 ( 
.A(n_4536),
.B(n_725),
.Y(n_4659)
);

INVx1_ASAP7_75t_L g4660 ( 
.A(n_4438),
.Y(n_4660)
);

AOI22xp5_ASAP7_75t_L g4661 ( 
.A1(n_4447),
.A2(n_728),
.B1(n_726),
.B2(n_727),
.Y(n_4661)
);

OAI211xp5_ASAP7_75t_L g4662 ( 
.A1(n_4464),
.A2(n_729),
.B(n_726),
.C(n_728),
.Y(n_4662)
);

OAI22xp33_ASAP7_75t_L g4663 ( 
.A1(n_4523),
.A2(n_732),
.B1(n_729),
.B2(n_731),
.Y(n_4663)
);

AOI311xp33_ASAP7_75t_L g4664 ( 
.A1(n_4495),
.A2(n_733),
.A3(n_731),
.B(n_732),
.C(n_734),
.Y(n_4664)
);

AOI22xp5_ASAP7_75t_L g4665 ( 
.A1(n_4589),
.A2(n_4531),
.B1(n_4517),
.B2(n_4445),
.Y(n_4665)
);

AOI22xp5_ASAP7_75t_L g4666 ( 
.A1(n_4655),
.A2(n_4535),
.B1(n_4552),
.B2(n_4524),
.Y(n_4666)
);

NAND2xp5_ASAP7_75t_L g4667 ( 
.A(n_4654),
.B(n_4632),
.Y(n_4667)
);

AOI221xp5_ASAP7_75t_L g4668 ( 
.A1(n_4599),
.A2(n_4443),
.B1(n_4502),
.B2(n_4526),
.C(n_4473),
.Y(n_4668)
);

NOR2x1_ASAP7_75t_SL g4669 ( 
.A(n_4621),
.B(n_4623),
.Y(n_4669)
);

AO22x2_ASAP7_75t_L g4670 ( 
.A1(n_4638),
.A2(n_4519),
.B1(n_4514),
.B2(n_4510),
.Y(n_4670)
);

XOR2x2_ASAP7_75t_L g4671 ( 
.A(n_4622),
.B(n_4527),
.Y(n_4671)
);

INVxp67_ASAP7_75t_L g4672 ( 
.A(n_4627),
.Y(n_4672)
);

AOI21xp33_ASAP7_75t_L g4673 ( 
.A1(n_4605),
.A2(n_4513),
.B(n_4520),
.Y(n_4673)
);

AOI21xp33_ASAP7_75t_L g4674 ( 
.A1(n_4628),
.A2(n_4480),
.B(n_4483),
.Y(n_4674)
);

AOI221xp5_ASAP7_75t_SL g4675 ( 
.A1(n_4602),
.A2(n_4472),
.B1(n_4498),
.B2(n_4461),
.C(n_4544),
.Y(n_4675)
);

INVxp67_ASAP7_75t_L g4676 ( 
.A(n_4588),
.Y(n_4676)
);

INVx2_ASAP7_75t_L g4677 ( 
.A(n_4637),
.Y(n_4677)
);

AOI22xp33_ASAP7_75t_L g4678 ( 
.A1(n_4579),
.A2(n_4534),
.B1(n_4530),
.B2(n_4509),
.Y(n_4678)
);

OAI21xp33_ASAP7_75t_L g4679 ( 
.A1(n_4629),
.A2(n_4455),
.B(n_4528),
.Y(n_4679)
);

AOI21xp5_ASAP7_75t_L g4680 ( 
.A1(n_4615),
.A2(n_4508),
.B(n_4449),
.Y(n_4680)
);

AOI221xp5_ASAP7_75t_L g4681 ( 
.A1(n_4610),
.A2(n_4545),
.B1(n_4551),
.B2(n_4541),
.C(n_4488),
.Y(n_4681)
);

AOI22xp5_ASAP7_75t_L g4682 ( 
.A1(n_4660),
.A2(n_4522),
.B1(n_4516),
.B2(n_4521),
.Y(n_4682)
);

INVx2_ASAP7_75t_L g4683 ( 
.A(n_4630),
.Y(n_4683)
);

INVx1_ASAP7_75t_SL g4684 ( 
.A(n_4659),
.Y(n_4684)
);

AOI22xp5_ASAP7_75t_L g4685 ( 
.A1(n_4580),
.A2(n_4490),
.B1(n_4489),
.B2(n_4512),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_4582),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_L g4687 ( 
.A(n_4631),
.B(n_4453),
.Y(n_4687)
);

INVx2_ASAP7_75t_L g4688 ( 
.A(n_4645),
.Y(n_4688)
);

AOI221xp5_ASAP7_75t_L g4689 ( 
.A1(n_4662),
.A2(n_4532),
.B1(n_4533),
.B2(n_4469),
.C(n_4475),
.Y(n_4689)
);

AOI22xp5_ASAP7_75t_L g4690 ( 
.A1(n_4650),
.A2(n_4465),
.B1(n_4474),
.B2(n_4467),
.Y(n_4690)
);

INVx1_ASAP7_75t_L g4691 ( 
.A(n_4609),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4585),
.Y(n_4692)
);

NOR4xp25_ASAP7_75t_L g4693 ( 
.A(n_4657),
.B(n_4466),
.C(n_4484),
.D(n_4492),
.Y(n_4693)
);

NOR2xp33_ASAP7_75t_L g4694 ( 
.A(n_4639),
.B(n_4496),
.Y(n_4694)
);

AOI21xp33_ASAP7_75t_SL g4695 ( 
.A1(n_4612),
.A2(n_4463),
.B(n_4529),
.Y(n_4695)
);

OAI21xp33_ASAP7_75t_L g4696 ( 
.A1(n_4640),
.A2(n_733),
.B(n_735),
.Y(n_4696)
);

AOI22xp5_ASAP7_75t_L g4697 ( 
.A1(n_4641),
.A2(n_739),
.B1(n_737),
.B2(n_738),
.Y(n_4697)
);

O2A1O1Ixp33_ASAP7_75t_L g4698 ( 
.A1(n_4653),
.A2(n_4642),
.B(n_4584),
.C(n_4646),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4597),
.Y(n_4699)
);

AOI22xp5_ASAP7_75t_L g4700 ( 
.A1(n_4617),
.A2(n_739),
.B1(n_737),
.B2(n_738),
.Y(n_4700)
);

NAND2xp5_ASAP7_75t_L g4701 ( 
.A(n_4644),
.B(n_740),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4608),
.Y(n_4702)
);

INVxp67_ASAP7_75t_L g4703 ( 
.A(n_4626),
.Y(n_4703)
);

INVxp67_ASAP7_75t_L g4704 ( 
.A(n_4656),
.Y(n_4704)
);

AOI221xp5_ASAP7_75t_L g4705 ( 
.A1(n_4600),
.A2(n_743),
.B1(n_740),
.B2(n_742),
.C(n_745),
.Y(n_4705)
);

AOI221xp5_ASAP7_75t_L g4706 ( 
.A1(n_4577),
.A2(n_745),
.B1(n_742),
.B2(n_743),
.C(n_746),
.Y(n_4706)
);

OAI21xp33_ASAP7_75t_L g4707 ( 
.A1(n_4658),
.A2(n_746),
.B(n_747),
.Y(n_4707)
);

AOI221xp5_ASAP7_75t_L g4708 ( 
.A1(n_4607),
.A2(n_749),
.B1(n_747),
.B2(n_748),
.C(n_750),
.Y(n_4708)
);

NOR2xp33_ASAP7_75t_R g4709 ( 
.A(n_4611),
.B(n_4593),
.Y(n_4709)
);

AOI221xp5_ASAP7_75t_L g4710 ( 
.A1(n_4598),
.A2(n_751),
.B1(n_748),
.B2(n_750),
.C(n_752),
.Y(n_4710)
);

AOI221xp5_ASAP7_75t_L g4711 ( 
.A1(n_4587),
.A2(n_755),
.B1(n_753),
.B2(n_754),
.C(n_756),
.Y(n_4711)
);

OAI221xp5_ASAP7_75t_L g4712 ( 
.A1(n_4651),
.A2(n_4591),
.B1(n_4648),
.B2(n_4619),
.C(n_4606),
.Y(n_4712)
);

NAND2xp5_ASAP7_75t_L g4713 ( 
.A(n_4643),
.B(n_753),
.Y(n_4713)
);

AOI211xp5_ASAP7_75t_L g4714 ( 
.A1(n_4583),
.A2(n_760),
.B(n_754),
.C(n_759),
.Y(n_4714)
);

INVxp67_ASAP7_75t_L g4715 ( 
.A(n_4620),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_4624),
.Y(n_4716)
);

AND2x2_ASAP7_75t_L g4717 ( 
.A(n_4601),
.B(n_759),
.Y(n_4717)
);

XNOR2x1_ASAP7_75t_L g4718 ( 
.A(n_4590),
.B(n_760),
.Y(n_4718)
);

O2A1O1Ixp33_ASAP7_75t_L g4719 ( 
.A1(n_4578),
.A2(n_763),
.B(n_761),
.C(n_762),
.Y(n_4719)
);

AOI211xp5_ASAP7_75t_L g4720 ( 
.A1(n_4613),
.A2(n_764),
.B(n_761),
.C(n_763),
.Y(n_4720)
);

INVxp67_ASAP7_75t_L g4721 ( 
.A(n_4595),
.Y(n_4721)
);

AOI211xp5_ASAP7_75t_L g4722 ( 
.A1(n_4663),
.A2(n_768),
.B(n_766),
.C(n_767),
.Y(n_4722)
);

OAI21xp5_ASAP7_75t_L g4723 ( 
.A1(n_4672),
.A2(n_4634),
.B(n_4594),
.Y(n_4723)
);

OAI221xp5_ASAP7_75t_L g4724 ( 
.A1(n_4667),
.A2(n_4581),
.B1(n_4603),
.B2(n_4618),
.C(n_4661),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_L g4725 ( 
.A(n_4684),
.B(n_4614),
.Y(n_4725)
);

NAND2xp5_ASAP7_75t_L g4726 ( 
.A(n_4693),
.B(n_4652),
.Y(n_4726)
);

AOI211xp5_ASAP7_75t_L g4727 ( 
.A1(n_4695),
.A2(n_4649),
.B(n_4636),
.C(n_4604),
.Y(n_4727)
);

AOI32xp33_ASAP7_75t_L g4728 ( 
.A1(n_4716),
.A2(n_4596),
.A3(n_4664),
.B1(n_4635),
.B2(n_4625),
.Y(n_4728)
);

OR2x2_ASAP7_75t_L g4729 ( 
.A(n_4687),
.B(n_4647),
.Y(n_4729)
);

OAI211xp5_ASAP7_75t_SL g4730 ( 
.A1(n_4679),
.A2(n_4633),
.B(n_4616),
.C(n_4586),
.Y(n_4730)
);

NOR3xp33_ASAP7_75t_L g4731 ( 
.A(n_4673),
.B(n_4674),
.C(n_4696),
.Y(n_4731)
);

OAI321xp33_ASAP7_75t_L g4732 ( 
.A1(n_4665),
.A2(n_4592),
.A3(n_768),
.B1(n_769),
.B2(n_770),
.C(n_771),
.Y(n_4732)
);

NOR2xp33_ASAP7_75t_L g4733 ( 
.A(n_4676),
.B(n_767),
.Y(n_4733)
);

AOI21xp33_ASAP7_75t_SL g4734 ( 
.A1(n_4670),
.A2(n_770),
.B(n_771),
.Y(n_4734)
);

AOI22xp5_ASAP7_75t_L g4735 ( 
.A1(n_4694),
.A2(n_774),
.B1(n_772),
.B2(n_773),
.Y(n_4735)
);

INVx2_ASAP7_75t_L g4736 ( 
.A(n_4669),
.Y(n_4736)
);

OA22x2_ASAP7_75t_L g4737 ( 
.A1(n_4666),
.A2(n_776),
.B1(n_773),
.B2(n_775),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4670),
.Y(n_4738)
);

AOI221xp5_ASAP7_75t_SL g4739 ( 
.A1(n_4680),
.A2(n_781),
.B1(n_776),
.B2(n_778),
.C(n_782),
.Y(n_4739)
);

OAI21xp5_ASAP7_75t_L g4740 ( 
.A1(n_4698),
.A2(n_781),
.B(n_783),
.Y(n_4740)
);

AND2x4_ASAP7_75t_L g4741 ( 
.A(n_4699),
.B(n_783),
.Y(n_4741)
);

NOR2xp33_ASAP7_75t_R g4742 ( 
.A(n_4692),
.B(n_784),
.Y(n_4742)
);

AOI221xp5_ASAP7_75t_L g4743 ( 
.A1(n_4681),
.A2(n_786),
.B1(n_784),
.B2(n_785),
.C(n_787),
.Y(n_4743)
);

OAI22xp5_ASAP7_75t_L g4744 ( 
.A1(n_4678),
.A2(n_4682),
.B1(n_4690),
.B2(n_4697),
.Y(n_4744)
);

OAI22xp5_ASAP7_75t_L g4745 ( 
.A1(n_4685),
.A2(n_4700),
.B1(n_4721),
.B2(n_4704),
.Y(n_4745)
);

AND2x2_ASAP7_75t_L g4746 ( 
.A(n_4688),
.B(n_785),
.Y(n_4746)
);

NAND2xp5_ASAP7_75t_L g4747 ( 
.A(n_4675),
.B(n_788),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4717),
.Y(n_4748)
);

NOR2x1_ASAP7_75t_L g4749 ( 
.A(n_4701),
.B(n_789),
.Y(n_4749)
);

OAI22xp33_ASAP7_75t_SL g4750 ( 
.A1(n_4712),
.A2(n_4702),
.B1(n_4715),
.B2(n_4703),
.Y(n_4750)
);

INVxp67_ASAP7_75t_L g4751 ( 
.A(n_4713),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4671),
.Y(n_4752)
);

NOR3xp33_ASAP7_75t_L g4753 ( 
.A(n_4686),
.B(n_789),
.C(n_790),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4677),
.Y(n_4754)
);

OAI22xp5_ASAP7_75t_L g4755 ( 
.A1(n_4714),
.A2(n_4722),
.B1(n_4720),
.B2(n_4683),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4718),
.Y(n_4756)
);

CKINVDCx5p33_ASAP7_75t_R g4757 ( 
.A(n_4709),
.Y(n_4757)
);

NOR2x1_ASAP7_75t_L g4758 ( 
.A(n_4736),
.B(n_4691),
.Y(n_4758)
);

INVxp67_ASAP7_75t_L g4759 ( 
.A(n_4733),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_L g4760 ( 
.A(n_4741),
.B(n_4706),
.Y(n_4760)
);

BUFx6f_ASAP7_75t_L g4761 ( 
.A(n_4741),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4737),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_4746),
.Y(n_4763)
);

AOI22xp5_ASAP7_75t_L g4764 ( 
.A1(n_4757),
.A2(n_4668),
.B1(n_4689),
.B2(n_4708),
.Y(n_4764)
);

NOR2x1_ASAP7_75t_L g4765 ( 
.A(n_4749),
.B(n_4707),
.Y(n_4765)
);

INVx1_ASAP7_75t_SL g4766 ( 
.A(n_4742),
.Y(n_4766)
);

INVx2_ASAP7_75t_L g4767 ( 
.A(n_4729),
.Y(n_4767)
);

INVx1_ASAP7_75t_L g4768 ( 
.A(n_4747),
.Y(n_4768)
);

OR2x2_ASAP7_75t_L g4769 ( 
.A(n_4726),
.B(n_4725),
.Y(n_4769)
);

OAI22xp33_ASAP7_75t_L g4770 ( 
.A1(n_4752),
.A2(n_4705),
.B1(n_4711),
.B2(n_4710),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4738),
.Y(n_4771)
);

INVx2_ASAP7_75t_L g4772 ( 
.A(n_4748),
.Y(n_4772)
);

NOR2x1p5_ASAP7_75t_L g4773 ( 
.A(n_4754),
.B(n_4719),
.Y(n_4773)
);

HB1xp67_ASAP7_75t_L g4774 ( 
.A(n_4740),
.Y(n_4774)
);

AND2x2_ASAP7_75t_L g4775 ( 
.A(n_4723),
.B(n_790),
.Y(n_4775)
);

AND2x4_ASAP7_75t_L g4776 ( 
.A(n_4772),
.B(n_4751),
.Y(n_4776)
);

OR2x2_ASAP7_75t_L g4777 ( 
.A(n_4761),
.B(n_4755),
.Y(n_4777)
);

AOI22xp5_ASAP7_75t_L g4778 ( 
.A1(n_4762),
.A2(n_4731),
.B1(n_4744),
.B2(n_4730),
.Y(n_4778)
);

INVx1_ASAP7_75t_L g4779 ( 
.A(n_4761),
.Y(n_4779)
);

INVx2_ASAP7_75t_L g4780 ( 
.A(n_4773),
.Y(n_4780)
);

XNOR2xp5_ASAP7_75t_L g4781 ( 
.A(n_4764),
.B(n_4727),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4760),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4775),
.Y(n_4783)
);

NOR3xp33_ASAP7_75t_L g4784 ( 
.A(n_4767),
.B(n_4724),
.C(n_4750),
.Y(n_4784)
);

XNOR2x1_ASAP7_75t_L g4785 ( 
.A(n_4769),
.B(n_4745),
.Y(n_4785)
);

AND2x2_ASAP7_75t_L g4786 ( 
.A(n_4766),
.B(n_4756),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_L g4787 ( 
.A(n_4771),
.B(n_4734),
.Y(n_4787)
);

AND2x4_ASAP7_75t_L g4788 ( 
.A(n_4779),
.B(n_4758),
.Y(n_4788)
);

XNOR2x1_ASAP7_75t_L g4789 ( 
.A(n_4785),
.B(n_4765),
.Y(n_4789)
);

O2A1O1Ixp33_ASAP7_75t_L g4790 ( 
.A1(n_4784),
.A2(n_4787),
.B(n_4774),
.C(n_4770),
.Y(n_4790)
);

NOR4xp25_ASAP7_75t_L g4791 ( 
.A(n_4782),
.B(n_4728),
.C(n_4768),
.D(n_4763),
.Y(n_4791)
);

NAND2xp5_ASAP7_75t_L g4792 ( 
.A(n_4776),
.B(n_4739),
.Y(n_4792)
);

AOI22x1_ASAP7_75t_L g4793 ( 
.A1(n_4781),
.A2(n_4759),
.B1(n_4732),
.B2(n_4743),
.Y(n_4793)
);

AOI222xp33_ASAP7_75t_L g4794 ( 
.A1(n_4786),
.A2(n_4753),
.B1(n_4735),
.B2(n_795),
.C1(n_796),
.C2(n_799),
.Y(n_4794)
);

NAND3xp33_ASAP7_75t_SL g4795 ( 
.A(n_4778),
.B(n_4777),
.C(n_4780),
.Y(n_4795)
);

OAI22xp5_ASAP7_75t_L g4796 ( 
.A1(n_4783),
.A2(n_796),
.B1(n_792),
.B2(n_794),
.Y(n_4796)
);

XNOR2x1_ASAP7_75t_L g4797 ( 
.A(n_4789),
.B(n_792),
.Y(n_4797)
);

OR2x2_ASAP7_75t_L g4798 ( 
.A(n_4791),
.B(n_799),
.Y(n_4798)
);

HB1xp67_ASAP7_75t_L g4799 ( 
.A(n_4788),
.Y(n_4799)
);

AND2x2_ASAP7_75t_L g4800 ( 
.A(n_4794),
.B(n_800),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4798),
.Y(n_4801)
);

HB1xp67_ASAP7_75t_L g4802 ( 
.A(n_4797),
.Y(n_4802)
);

AND2x2_ASAP7_75t_SL g4803 ( 
.A(n_4799),
.B(n_4792),
.Y(n_4803)
);

AOI222xp33_ASAP7_75t_L g4804 ( 
.A1(n_4803),
.A2(n_4795),
.B1(n_4800),
.B2(n_4796),
.C1(n_4793),
.C2(n_4790),
.Y(n_4804)
);

XOR2x2_ASAP7_75t_L g4805 ( 
.A(n_4804),
.B(n_4802),
.Y(n_4805)
);

XOR2xp5_ASAP7_75t_L g4806 ( 
.A(n_4805),
.B(n_4801),
.Y(n_4806)
);

AOI22xp5_ASAP7_75t_L g4807 ( 
.A1(n_4806),
.A2(n_802),
.B1(n_800),
.B2(n_801),
.Y(n_4807)
);

NOR2xp33_ASAP7_75t_L g4808 ( 
.A(n_4807),
.B(n_801),
.Y(n_4808)
);

OA21x2_ASAP7_75t_L g4809 ( 
.A1(n_4808),
.A2(n_803),
.B(n_804),
.Y(n_4809)
);

AOI22xp5_ASAP7_75t_L g4810 ( 
.A1(n_4809),
.A2(n_806),
.B1(n_803),
.B2(n_804),
.Y(n_4810)
);

AOI22xp5_ASAP7_75t_L g4811 ( 
.A1(n_4809),
.A2(n_811),
.B1(n_806),
.B2(n_807),
.Y(n_4811)
);

AOI22x1_ASAP7_75t_L g4812 ( 
.A1(n_4810),
.A2(n_813),
.B1(n_807),
.B2(n_812),
.Y(n_4812)
);

OR2x6_ASAP7_75t_L g4813 ( 
.A(n_4811),
.B(n_812),
.Y(n_4813)
);

AOI22xp5_ASAP7_75t_L g4814 ( 
.A1(n_4813),
.A2(n_4812),
.B1(n_815),
.B2(n_813),
.Y(n_4814)
);

AOI211xp5_ASAP7_75t_L g4815 ( 
.A1(n_4814),
.A2(n_970),
.B(n_817),
.C(n_814),
.Y(n_4815)
);


endmodule