module fake_jpeg_457_n_210 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_210);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_210;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_16),
.B(n_2),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_13),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_24),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_20),
.Y(n_67)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_13),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_10),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_73),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_81),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_81),
.A2(n_61),
.B1(n_63),
.B2(n_67),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_95),
.B1(n_80),
.B2(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_91),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_51),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_88),
.B(n_55),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_65),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_80),
.B(n_51),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_72),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_61),
.B1(n_63),
.B2(n_67),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_108),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_100),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_58),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_85),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_102),
.B(n_103),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_69),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_106),
.B(n_113),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_59),
.B1(n_58),
.B2(n_70),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_110),
.B1(n_68),
.B2(n_62),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_82),
.A2(n_64),
.B1(n_57),
.B2(n_66),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_112),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_59),
.B1(n_70),
.B2(n_66),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_74),
.Y(n_111)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_71),
.B(n_64),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_0),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_124),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_101),
.A2(n_85),
.B1(n_94),
.B2(n_93),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_119),
.A2(n_122),
.B1(n_111),
.B2(n_107),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_100),
.A2(n_94),
.B1(n_83),
.B2(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_86),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_89),
.B1(n_111),
.B2(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_23),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_97),
.B(n_0),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_131),
.B(n_112),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_1),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_43),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_134),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_140),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_138),
.B(n_148),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_89),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_146),
.C(n_133),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_115),
.A2(n_68),
.B1(n_62),
.B2(n_53),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_53),
.B1(n_50),
.B2(n_49),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_142),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_48),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_45),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_40),
.Y(n_169)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_145),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_44),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_3),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_120),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_152),
.B(n_154),
.Y(n_162)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_4),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_123),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_SL g172 ( 
.A1(n_156),
.A2(n_38),
.A3(n_36),
.B1(n_34),
.B2(n_31),
.C1(n_30),
.C2(n_29),
.Y(n_172)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_166),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_118),
.Y(n_166)
);

OAI32xp33_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_119),
.A3(n_129),
.B1(n_120),
.B2(n_122),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_172),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_164),
.C(n_174),
.Y(n_184)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_173),
.B(n_174),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_130),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_175),
.B(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_142),
.B(n_8),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_139),
.C(n_146),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_184),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_144),
.B(n_140),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_182),
.A2(n_186),
.B(n_169),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_161),
.B(n_141),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_183),
.B(n_185),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_134),
.C(n_145),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_28),
.B(n_27),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_187),
.A2(n_159),
.B1(n_167),
.B2(n_162),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_193),
.B(n_195),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_189),
.A2(n_194),
.B1(n_178),
.B2(n_11),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_160),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_190),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_177),
.A2(n_167),
.B(n_157),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_180),
.Y(n_194)
);

AO221x1_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_163),
.B1(n_175),
.B2(n_168),
.C(n_157),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_179),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_200),
.C(n_14),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_199),
.A2(n_9),
.B1(n_12),
.B2(n_14),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_26),
.C(n_12),
.Y(n_200)
);

AOI21x1_ASAP7_75t_L g201 ( 
.A1(n_197),
.A2(n_192),
.B(n_189),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_201),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_196),
.B(n_200),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_206),
.A2(n_198),
.B1(n_203),
.B2(n_204),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g208 ( 
.A1(n_207),
.A2(n_15),
.A3(n_16),
.B1(n_17),
.B2(n_18),
.C1(n_19),
.C2(n_20),
.Y(n_208)
);

A2O1A1O1Ixp25_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_15),
.B(n_18),
.C(n_19),
.D(n_21),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_21),
.Y(n_210)
);


endmodule