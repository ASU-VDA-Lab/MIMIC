module fake_jpeg_27751_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_0),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_44),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_7),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_34),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_49),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_17),
.B(n_7),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_48),
.B(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_16),
.B(n_9),
.Y(n_49)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_20),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_72),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_58),
.B(n_67),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

INVx5_ASAP7_75t_SL g104 ( 
.A(n_60),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_29),
.C(n_34),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_64),
.Y(n_103)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_62),
.Y(n_89)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_32),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

OR2x2_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_46),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

AO22x1_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_18),
.B1(n_45),
.B2(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_37),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_61),
.A2(n_41),
.B1(n_36),
.B2(n_18),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_78),
.A2(n_99),
.B1(n_110),
.B2(n_26),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_80),
.B(n_91),
.Y(n_140)
);

AND2x4_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_47),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_86),
.Y(n_116)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

BUFx16f_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_49),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_18),
.B1(n_25),
.B2(n_36),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_93),
.A2(n_102),
.B1(n_108),
.B2(n_30),
.Y(n_137)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_72),
.A2(n_18),
.B1(n_25),
.B2(n_26),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_55),
.A2(n_33),
.B1(n_23),
.B2(n_27),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_58),
.Y(n_105)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_44),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_107),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_69),
.A2(n_22),
.B1(n_27),
.B2(n_31),
.Y(n_108)
);

OR2x2_ASAP7_75t_SL g109 ( 
.A(n_73),
.B(n_22),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_60),
.A2(n_54),
.B1(n_63),
.B2(n_26),
.Y(n_110)
);

CKINVDCx12_ASAP7_75t_R g112 ( 
.A(n_69),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_50),
.B(n_28),
.Y(n_113)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_74),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_21),
.B1(n_74),
.B2(n_43),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_119),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_47),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_131),
.Y(n_150)
);

AO22x2_ASAP7_75t_L g130 ( 
.A1(n_81),
.A2(n_47),
.B1(n_59),
.B2(n_38),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_139),
.B1(n_104),
.B2(n_106),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_50),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_1),
.B(n_2),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_144),
.B(n_94),
.Y(n_168)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_141),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_33),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_96),
.A2(n_20),
.B1(n_21),
.B2(n_31),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_31),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_142),
.B(n_78),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_81),
.A2(n_59),
.B1(n_53),
.B2(n_52),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_95),
.B1(n_76),
.B2(n_104),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_86),
.A2(n_21),
.B(n_35),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_147),
.B(n_148),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_135),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_140),
.B(n_87),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_149),
.B(n_153),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_154),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_133),
.B(n_126),
.Y(n_153)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_77),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_155),
.A2(n_37),
.B1(n_118),
.B2(n_38),
.Y(n_204)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_156),
.A2(n_165),
.B1(n_172),
.B2(n_176),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_109),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_162),
.B1(n_89),
.B2(n_127),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_97),
.B1(n_82),
.B2(n_75),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_163),
.A2(n_167),
.B1(n_120),
.B2(n_117),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_84),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_166),
.B(n_168),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_97),
.B1(n_101),
.B2(n_98),
.Y(n_167)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_14),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_174),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_79),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_170),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_128),
.B(n_94),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_171),
.Y(n_184)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_125),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_90),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_115),
.B(n_43),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_116),
.C(n_144),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_111),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_SL g230 ( 
.A(n_179),
.B(n_38),
.C(n_83),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_180),
.A2(n_161),
.B1(n_176),
.B2(n_154),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_160),
.A2(n_119),
.B1(n_120),
.B2(n_129),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_201),
.B1(n_204),
.B2(n_205),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_192),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_146),
.B(n_116),
.C(n_122),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_116),
.C(n_90),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_195),
.Y(n_222)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_196),
.B(n_199),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_158),
.A2(n_118),
.B(n_2),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_197),
.A2(n_209),
.B(n_3),
.Y(n_234)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_89),
.B1(n_123),
.B2(n_121),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_121),
.C(n_85),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_203),
.B(n_210),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_155),
.A2(n_33),
.B1(n_29),
.B2(n_34),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_92),
.Y(n_207)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_168),
.Y(n_208)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_152),
.A2(n_1),
.B(n_2),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_157),
.B(n_85),
.C(n_92),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_111),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_187),
.B(n_169),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_212),
.B(n_233),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_214),
.A2(n_225),
.B1(n_234),
.B2(n_202),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_191),
.Y(n_215)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

INVxp33_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_216),
.A2(n_217),
.B1(n_224),
.B2(n_229),
.Y(n_261)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

INVx13_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_196),
.A2(n_206),
.B1(n_200),
.B2(n_195),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_189),
.A2(n_178),
.B1(n_165),
.B2(n_164),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_236),
.B1(n_238),
.B2(n_184),
.Y(n_246)
);

OAI22x1_ASAP7_75t_SL g229 ( 
.A1(n_208),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_230),
.A2(n_186),
.B1(n_199),
.B2(n_197),
.Y(n_245)
);

OA22x2_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_83),
.B1(n_19),
.B2(n_35),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_231),
.Y(n_259)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_181),
.B(n_28),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_200),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_235),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_189),
.A2(n_28),
.B1(n_51),
.B2(n_5),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_188),
.A2(n_51),
.B1(n_4),
.B2(n_5),
.Y(n_238)
);

INVx13_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_183),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_203),
.C(n_192),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_221),
.C(n_227),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_245),
.A2(n_246),
.B1(n_231),
.B2(n_224),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_182),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_250),
.Y(n_268)
);

XNOR2x1_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_182),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_190),
.C(n_223),
.Y(n_267)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_210),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_251),
.A2(n_234),
.B1(n_239),
.B2(n_231),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_207),
.Y(n_252)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_SL g254 ( 
.A(n_229),
.B(n_194),
.Y(n_254)
);

HAxp5_ASAP7_75t_SL g266 ( 
.A(n_254),
.B(n_238),
.CON(n_266),
.SN(n_266)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_256),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_209),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_213),
.B(n_187),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_262),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_219),
.A2(n_194),
.B1(n_179),
.B2(n_193),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_258),
.A2(n_222),
.B1(n_214),
.B2(n_223),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_226),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_265),
.A2(n_255),
.B1(n_243),
.B2(n_259),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_266),
.A2(n_259),
.B1(n_242),
.B2(n_246),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_274),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_241),
.Y(n_269)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_250),
.C(n_245),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_253),
.B(n_212),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_272),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_243),
.A2(n_235),
.B1(n_230),
.B2(n_217),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_273),
.A2(n_279),
.B1(n_256),
.B2(n_262),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_236),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_221),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_278),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_183),
.Y(n_276)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_276),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_239),
.Y(n_277)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_227),
.Y(n_278)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

XOR2x2_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_265),
.Y(n_282)
);

AO21x1_ASAP7_75t_L g305 ( 
.A1(n_282),
.A2(n_287),
.B(n_296),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_290),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_267),
.C(n_268),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_287),
.B(n_291),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_264),
.A2(n_248),
.B1(n_261),
.B2(n_252),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_280),
.A2(n_271),
.B1(n_266),
.B2(n_279),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_297),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_294),
.A2(n_270),
.B1(n_274),
.B2(n_278),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_263),
.A2(n_249),
.B(n_231),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_268),
.Y(n_302)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

BUFx12_ASAP7_75t_L g298 ( 
.A(n_282),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_298),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_305),
.C(n_306),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_302),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_224),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_304),
.A2(n_307),
.B(n_284),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_217),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_57),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_310),
.C(n_292),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_311),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_316),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_293),
.C(n_290),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_318),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_293),
.C(n_285),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_40),
.C(n_42),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_57),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_303),
.C(n_307),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_325),
.C(n_326),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_324),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_303),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_42),
.C(n_40),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_323),
.A2(n_313),
.B1(n_10),
.B2(n_11),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_326),
.Y(n_332)
);

AOI31xp67_ASAP7_75t_L g329 ( 
.A1(n_320),
.A2(n_10),
.A3(n_13),
.B(n_12),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_329),
.A2(n_10),
.B(n_11),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_331),
.Y(n_333)
);

AOI322xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_332),
.A3(n_330),
.B1(n_328),
.B2(n_321),
.C1(n_9),
.C2(n_11),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_328),
.C(n_6),
.Y(n_335)
);

AOI322xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_42),
.C2(n_329),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_6),
.C(n_4),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_3),
.B(n_5),
.Y(n_339)
);


endmodule