module fake_jpeg_23834_n_333 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_47),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_31),
.B1(n_24),
.B2(n_25),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_53),
.A2(n_77),
.B1(n_9),
.B2(n_15),
.Y(n_123)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_61),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_68),
.Y(n_99)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_28),
.Y(n_62)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_71),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_25),
.B1(n_44),
.B2(n_20),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_64),
.A2(n_66),
.B1(n_78),
.B2(n_84),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_24),
.B1(n_31),
.B2(n_35),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_65),
.A2(n_69),
.B1(n_82),
.B2(n_22),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_17),
.B1(n_20),
.B2(n_23),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_39),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_35),
.B1(n_36),
.B2(n_26),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_76),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_35),
.B1(n_21),
.B2(n_22),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_30),
.B1(n_23),
.B2(n_28),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_14),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_18),
.Y(n_89)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_85),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_36),
.B1(n_32),
.B2(n_26),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_45),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_48),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_48),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_86),
.Y(n_110)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_0),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_89),
.B(n_10),
.Y(n_151)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_60),
.A2(n_29),
.B1(n_21),
.B2(n_33),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_94),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_96),
.B(n_97),
.Y(n_159)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_100),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_38),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_38),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_54),
.A2(n_18),
.B1(n_33),
.B2(n_11),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_52),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_111),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_60),
.A2(n_18),
.B1(n_33),
.B2(n_10),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_52),
.Y(n_111)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_58),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_114),
.B(n_116),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_56),
.B(n_52),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_119),
.B(n_120),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_56),
.B(n_48),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_121),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_75),
.B1(n_80),
.B2(n_59),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_61),
.B(n_8),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_124),
.Y(n_132)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_126),
.B(n_137),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_119),
.A2(n_53),
.B1(n_87),
.B2(n_73),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_130),
.B1(n_142),
.B2(n_144),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_L g133 ( 
.A1(n_90),
.A2(n_79),
.B1(n_71),
.B2(n_73),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_133),
.A2(n_121),
.B1(n_97),
.B2(n_118),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_110),
.Y(n_137)
);

AO22x1_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_73),
.B1(n_80),
.B2(n_74),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_120),
.B1(n_116),
.B2(n_111),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_76),
.B1(n_72),
.B2(n_85),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_102),
.A2(n_85),
.B1(n_83),
.B2(n_75),
.Y(n_144)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_154),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_103),
.A2(n_83),
.B1(n_70),
.B2(n_3),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_158),
.B1(n_10),
.B2(n_16),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_13),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_70),
.C(n_2),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_118),
.C(n_12),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_110),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_115),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_157),
.Y(n_189)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_105),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_134),
.A2(n_98),
.B1(n_113),
.B2(n_92),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_161),
.A2(n_178),
.B1(n_180),
.B2(n_186),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_141),
.B1(n_130),
.B2(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_165),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_147),
.B(n_99),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_99),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_168),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_167),
.B(n_185),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_137),
.B(n_96),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_101),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_170),
.Y(n_203)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_104),
.B(n_106),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_171),
.A2(n_183),
.B(n_187),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_154),
.B(n_112),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_140),
.A2(n_89),
.B1(n_91),
.B2(n_117),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_152),
.B(n_91),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

AO21x2_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_125),
.B(n_158),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_184),
.Y(n_213)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_145),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_156),
.B(n_109),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_193),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_109),
.Y(n_191)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_7),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_192),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_135),
.B(n_94),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_135),
.B(n_1),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g224 ( 
.A(n_194),
.B(n_1),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_196),
.B(n_221),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_188),
.A2(n_141),
.B1(n_146),
.B2(n_129),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_197),
.A2(n_208),
.B1(n_222),
.B2(n_173),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_129),
.B1(n_127),
.B2(n_136),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_200),
.A2(n_180),
.B1(n_164),
.B2(n_170),
.Y(n_227)
);

OAI32xp33_ASAP7_75t_L g204 ( 
.A1(n_163),
.A2(n_180),
.A3(n_187),
.B1(n_179),
.B2(n_166),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_224),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_132),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_211),
.C(n_220),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_162),
.A2(n_131),
.B1(n_127),
.B2(n_136),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_132),
.C(n_139),
.Y(n_211)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_175),
.Y(n_226)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_150),
.C(n_148),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_131),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_162),
.A2(n_143),
.B1(n_2),
.B2(n_3),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_14),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_225),
.C(n_183),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_15),
.Y(n_225)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_227),
.A2(n_217),
.B1(n_224),
.B2(n_212),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_198),
.B(n_184),
.Y(n_228)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_203),
.B(n_182),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_232),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_231),
.A2(n_243),
.B1(n_246),
.B2(n_248),
.Y(n_256)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_216),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_235),
.Y(n_259)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_199),
.Y(n_236)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_224),
.C(n_197),
.Y(n_265)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_206),
.A2(n_195),
.B(n_171),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_241),
.B(n_242),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_211),
.B(n_194),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_240),
.A2(n_244),
.B(n_245),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_207),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_208),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_225),
.B(n_194),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_221),
.B(n_176),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_189),
.B(n_167),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_218),
.A2(n_186),
.B(n_143),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_214),
.B1(n_202),
.B2(n_215),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_251),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_239),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_254),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_232),
.A2(n_218),
.B1(n_204),
.B2(n_196),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_255),
.A2(n_258),
.B1(n_227),
.B2(n_256),
.Y(n_278)
);

XNOR2x1_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_202),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_262),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_205),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_269),
.C(n_237),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_267),
.A2(n_231),
.B1(n_249),
.B2(n_248),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_201),
.C(n_223),
.Y(n_269)
);

AOI21xp33_ASAP7_75t_L g270 ( 
.A1(n_268),
.A2(n_234),
.B(n_233),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_270),
.A2(n_278),
.B1(n_286),
.B2(n_254),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_259),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_276),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_282),
.C(n_287),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_247),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_264),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_267),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_253),
.A2(n_233),
.B(n_243),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_277),
.A2(n_242),
.B(n_260),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_257),
.B(n_241),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_281),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_250),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_245),
.C(n_236),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_244),
.C(n_266),
.Y(n_300)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_263),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_275),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_201),
.Y(n_302)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_291),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_277),
.B(n_273),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_269),
.C(n_272),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_294),
.C(n_300),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_265),
.C(n_264),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_298),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_278),
.B(n_255),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_290),
.A2(n_287),
.B1(n_286),
.B2(n_284),
.Y(n_301)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_302),
.B(n_300),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_296),
.A2(n_280),
.B(n_235),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_304),
.Y(n_313)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_273),
.C(n_281),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_304),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_212),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_296),
.Y(n_314)
);

OA21x2_ASAP7_75t_L g310 ( 
.A1(n_292),
.A2(n_280),
.B(n_268),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_266),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_314),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_297),
.B1(n_288),
.B2(n_298),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_315),
.A2(n_318),
.B1(n_301),
.B2(n_230),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_316),
.A2(n_317),
.B(n_310),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_306),
.A2(n_252),
.B1(n_238),
.B2(n_228),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_308),
.C(n_305),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_319),
.B(n_322),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_310),
.Y(n_321)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_321),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_323),
.A2(n_311),
.B1(n_317),
.B2(n_240),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_325),
.A2(n_321),
.B(n_318),
.Y(n_327)
);

OAI321xp33_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_328),
.A3(n_324),
.B1(n_325),
.B2(n_305),
.C(n_219),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_326),
.A2(n_320),
.B(n_308),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_16),
.B1(n_4),
.B2(n_5),
.Y(n_330)
);

OAI31xp33_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_1),
.A3(n_4),
.B(n_5),
.Y(n_331)
);

NAND2xp33_ASAP7_75t_R g332 ( 
.A(n_331),
.B(n_4),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_16),
.Y(n_333)
);


endmodule