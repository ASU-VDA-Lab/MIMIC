module fake_ibex_663_n_1241 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_201, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_195, n_163, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_202, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1241);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_195;
input n_163;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1241;

wire n_1084;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_280;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_875;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_242;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_235;
wire n_538;
wire n_1155;
wire n_459;
wire n_518;
wire n_852;
wire n_1133;
wire n_904;
wire n_355;
wire n_646;
wire n_448;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_230;
wire n_917;
wire n_968;
wire n_352;
wire n_558;
wire n_666;
wire n_219;
wire n_1071;
wire n_793;
wire n_937;
wire n_234;
wire n_973;
wire n_1038;
wire n_618;
wire n_662;
wire n_979;
wire n_209;
wire n_1215;
wire n_629;
wire n_573;
wire n_359;
wire n_433;
wire n_262;
wire n_439;
wire n_1007;
wire n_643;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_369;
wire n_257;
wire n_869;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_562;
wire n_564;
wire n_795;
wire n_592;
wire n_762;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_397;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_499;
wire n_702;
wire n_971;
wire n_451;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1190;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1108;
wire n_382;
wire n_1239;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_695;
wire n_639;
wire n_482;
wire n_282;
wire n_870;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1154;
wire n_345;
wire n_455;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_252;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_241;
wire n_231;
wire n_657;
wire n_1156;
wire n_749;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1031;
wire n_372;
wire n_256;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1015;
wire n_663;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_258;
wire n_1129;
wire n_449;
wire n_421;
wire n_738;
wire n_1217;
wire n_236;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_840;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_574;
wire n_515;
wire n_1229;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_944;
wire n_623;
wire n_585;
wire n_483;
wire n_1137;
wire n_222;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_207;
wire n_1028;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_267;
wire n_1009;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_413;
wire n_1069;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_998;
wire n_1115;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_227;
wire n_1087;
wire n_757;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_517;
wire n_211;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_291;
wire n_318;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_997;
wire n_891;
wire n_303;
wire n_717;
wire n_668;
wire n_871;
wire n_266;
wire n_485;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_460;
wire n_461;
wire n_903;
wire n_1095;
wire n_1048;
wire n_774;
wire n_588;
wire n_528;
wire n_260;
wire n_836;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_213;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_920;
wire n_664;
wire n_1067;
wire n_255;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_578;
wire n_432;
wire n_403;
wire n_423;
wire n_357;
wire n_226;
wire n_216;
wire n_996;
wire n_915;
wire n_1174;
wire n_542;
wire n_900;
wire n_377;
wire n_647;
wire n_317;
wire n_326;
wire n_270;
wire n_259;
wire n_276;
wire n_339;
wire n_348;
wire n_220;
wire n_674;
wire n_287;
wire n_552;
wire n_251;
wire n_1112;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_224;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_838;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_1191;
wire n_221;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_246;
wire n_922;
wire n_851;
wire n_993;
wire n_253;
wire n_208;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_245;
wire n_571;
wire n_229;
wire n_648;
wire n_830;
wire n_473;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_768;
wire n_839;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_976;
wire n_1063;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_804;
wire n_484;
wire n_480;
wire n_1057;
wire n_354;
wire n_516;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_248;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_218;
wire n_277;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_247;
wire n_237;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_782;
wire n_616;
wire n_833;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1221;
wire n_284;
wire n_1047;
wire n_792;
wire n_575;
wire n_313;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_302;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_587;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_232;
wire n_1050;
wire n_599;
wire n_1060;
wire n_756;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_249;
wire n_478;
wire n_239;
wire n_336;
wire n_861;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_753;
wire n_747;
wire n_645;
wire n_1147;
wire n_1098;
wire n_584;
wire n_1187;
wire n_698;
wire n_1061;
wire n_682;
wire n_327;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_265;
wire n_1029;
wire n_470;
wire n_770;
wire n_210;
wire n_941;
wire n_243;
wire n_228;
wire n_632;
wire n_373;
wire n_854;
wire n_244;
wire n_343;
wire n_714;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_333;
wire n_967;
wire n_736;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_215;
wire n_987;
wire n_750;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1023;
wire n_568;
wire n_813;
wire n_1211;
wire n_1116;
wire n_791;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1074;
wire n_759;
wire n_953;
wire n_1180;
wire n_536;
wire n_1220;
wire n_467;
wire n_427;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_263;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_735;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1089;
wire n_392;
wire n_206;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1033;
wire n_627;
wire n_990;
wire n_322;
wire n_888;
wire n_582;
wire n_653;
wire n_1205;
wire n_238;
wire n_214;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_225;
wire n_511;
wire n_223;
wire n_381;
wire n_1002;
wire n_1111;
wire n_405;
wire n_612;
wire n_955;
wire n_440;
wire n_342;
wire n_233;
wire n_414;
wire n_378;
wire n_952;
wire n_264;
wire n_1145;
wire n_217;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1016;
wire n_240;
wire n_680;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_493;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_212;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_254;
wire n_908;
wire n_565;
wire n_1123;
wire n_271;
wire n_984;
wire n_394;
wire n_364;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_SL g206 ( 
.A(n_185),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_97),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_25),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_201),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_177),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_109),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_175),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_61),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_135),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_116),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_96),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_39),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_134),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_7),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_58),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_98),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_111),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_176),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_103),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_158),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_131),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_143),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_17),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_159),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_18),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_192),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_91),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_104),
.Y(n_234)
);

BUFx8_ASAP7_75t_SL g235 ( 
.A(n_174),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_165),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_53),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_29),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_62),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_133),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_164),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_166),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_75),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_27),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_128),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_92),
.Y(n_247)
);

NOR2xp67_ASAP7_75t_L g248 ( 
.A(n_24),
.B(n_203),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_112),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_120),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_83),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_22),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_30),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_18),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_141),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_118),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_160),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_108),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_L g259 ( 
.A(n_51),
.B(n_198),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_95),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_2),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_52),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_188),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_145),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_55),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_171),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_101),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_9),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_44),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_138),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_78),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_190),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_127),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_113),
.Y(n_274)
);

BUFx5_ASAP7_75t_L g275 ( 
.A(n_146),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_181),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_48),
.B(n_2),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_73),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_173),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_21),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_69),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_178),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_1),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_85),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_155),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_4),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_152),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_117),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_204),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_193),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_87),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_26),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_191),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_140),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_12),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_12),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_19),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_182),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_139),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_184),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_100),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_24),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_202),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_105),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_66),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_50),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_163),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_90),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_106),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_102),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_55),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_162),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_68),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_114),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_63),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_183),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_46),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_147),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_115),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_46),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_20),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_34),
.B(n_170),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_161),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_144),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_79),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_59),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_80),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_172),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_1),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_136),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_126),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_41),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_0),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_8),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_110),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_130),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_5),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_44),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_93),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_39),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_132),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_107),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_194),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_63),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_167),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_179),
.Y(n_346)
);

INVxp33_ASAP7_75t_SL g347 ( 
.A(n_99),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_32),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_38),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_35),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_72),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_57),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_169),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_9),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_129),
.Y(n_355)
);

BUFx10_ASAP7_75t_L g356 ( 
.A(n_84),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_137),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_195),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_255),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_228),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_317),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_255),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_213),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_228),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_213),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_222),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_222),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_317),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_218),
.B(n_0),
.Y(n_369)
);

OA21x2_ASAP7_75t_L g370 ( 
.A1(n_282),
.A2(n_76),
.B(n_74),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_247),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_228),
.Y(n_372)
);

OA21x2_ASAP7_75t_L g373 ( 
.A1(n_282),
.A2(n_81),
.B(n_77),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_238),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_222),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_269),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_222),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_255),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_356),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_269),
.B(n_3),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_255),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_222),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_289),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_247),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_207),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_222),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_215),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_308),
.B(n_4),
.Y(n_388)
);

BUFx8_ASAP7_75t_L g389 ( 
.A(n_236),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_216),
.Y(n_390)
);

OAI21x1_ASAP7_75t_L g391 ( 
.A1(n_284),
.A2(n_86),
.B(n_82),
.Y(n_391)
);

BUFx8_ASAP7_75t_SL g392 ( 
.A(n_239),
.Y(n_392)
);

OA21x2_ASAP7_75t_L g393 ( 
.A1(n_284),
.A2(n_328),
.B(n_298),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_219),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_222),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_289),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_231),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_275),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_289),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_223),
.Y(n_400)
);

BUFx8_ASAP7_75t_SL g401 ( 
.A(n_239),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_224),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_208),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_226),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_275),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_261),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_230),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_356),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_289),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_356),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_272),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_229),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_221),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_310),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_310),
.Y(n_415)
);

BUFx8_ASAP7_75t_SL g416 ( 
.A(n_261),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_275),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_235),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_310),
.Y(n_419)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_272),
.Y(n_420)
);

AND2x6_ASAP7_75t_L g421 ( 
.A(n_273),
.B(n_316),
.Y(n_421)
);

BUFx12f_ASAP7_75t_L g422 ( 
.A(n_227),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_275),
.Y(n_423)
);

BUFx8_ASAP7_75t_SL g424 ( 
.A(n_305),
.Y(n_424)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_298),
.A2(n_89),
.B(n_88),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_310),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_273),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_275),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_234),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_240),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_316),
.Y(n_431)
);

INVx5_ASAP7_75t_L g432 ( 
.A(n_312),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_330),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_235),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_237),
.B(n_13),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_330),
.B(n_14),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_252),
.B(n_15),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_358),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_220),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_358),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_275),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_253),
.B(n_15),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_242),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_246),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_229),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_254),
.B(n_16),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_360),
.B(n_249),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_433),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_436),
.B(n_275),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_433),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_433),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_418),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_369),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_369),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_360),
.B(n_291),
.Y(n_455)
);

CKINVDCx6p67_ASAP7_75t_R g456 ( 
.A(n_418),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_369),
.Y(n_457)
);

AND3x2_ASAP7_75t_L g458 ( 
.A(n_397),
.B(n_277),
.C(n_265),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_360),
.B(n_291),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_380),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_360),
.B(n_251),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_396),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_438),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_364),
.B(n_244),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_364),
.B(n_268),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_380),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_380),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_410),
.B(n_278),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_380),
.Y(n_469)
);

CKINVDCx6p67_ASAP7_75t_R g470 ( 
.A(n_422),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_436),
.Y(n_471)
);

NAND3xp33_ASAP7_75t_L g472 ( 
.A(n_388),
.B(n_295),
.C(n_286),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_438),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_410),
.B(n_296),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_438),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_422),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_364),
.B(n_297),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_436),
.B(n_256),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_361),
.B(n_302),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_366),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_361),
.B(n_311),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_368),
.B(n_315),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_403),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_368),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_385),
.B(n_257),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_440),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_440),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_396),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_434),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_435),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_437),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_440),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_440),
.Y(n_493)
);

INVxp33_ASAP7_75t_SL g494 ( 
.A(n_439),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_392),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_385),
.B(n_258),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_427),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_437),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_430),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_427),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_379),
.B(n_320),
.Y(n_501)
);

AO21x2_ASAP7_75t_L g502 ( 
.A1(n_391),
.A2(n_322),
.B(n_263),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_430),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_427),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_363),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_427),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_379),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_427),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_363),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_387),
.B(n_260),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_421),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_365),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_431),
.Y(n_513)
);

NOR2x1p5_ASAP7_75t_L g514 ( 
.A(n_408),
.B(n_292),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_SL g515 ( 
.A(n_413),
.B(n_210),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_408),
.B(n_267),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_408),
.B(n_329),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_387),
.B(n_271),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_431),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_401),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_372),
.B(n_274),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_431),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_421),
.B(n_209),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_366),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_393),
.Y(n_525)
);

INVx8_ASAP7_75t_L g526 ( 
.A(n_421),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_393),
.Y(n_527)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_390),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_367),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_393),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_416),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_374),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_393),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_374),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_376),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_390),
.B(n_288),
.Y(n_536)
);

OR2x6_ASAP7_75t_L g537 ( 
.A(n_442),
.B(n_306),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_375),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_394),
.B(n_400),
.Y(n_539)
);

NAND3xp33_ASAP7_75t_L g540 ( 
.A(n_389),
.B(n_334),
.C(n_332),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_394),
.B(n_337),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_400),
.B(n_340),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_402),
.B(n_293),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_404),
.B(n_349),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_377),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_432),
.B(n_294),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_377),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_404),
.B(n_351),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_382),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_446),
.Y(n_550)
);

OR2x6_ASAP7_75t_L g551 ( 
.A(n_425),
.B(n_313),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_386),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_407),
.B(n_303),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_395),
.Y(n_554)
);

INVxp33_ASAP7_75t_L g555 ( 
.A(n_424),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_407),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_432),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_395),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_398),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_429),
.B(n_354),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_398),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_429),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_405),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_443),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_405),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_417),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_417),
.Y(n_567)
);

AO22x2_ASAP7_75t_L g568 ( 
.A1(n_444),
.A2(n_333),
.B1(n_338),
.B2(n_321),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_423),
.Y(n_569)
);

AO22x2_ASAP7_75t_L g570 ( 
.A1(n_420),
.A2(n_348),
.B1(n_350),
.B2(n_344),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_428),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_432),
.B(n_307),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_389),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_L g574 ( 
.A(n_441),
.B(n_211),
.Y(n_574)
);

INVx5_ASAP7_75t_L g575 ( 
.A(n_420),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_371),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_432),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_420),
.B(n_347),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_550),
.B(n_389),
.Y(n_579)
);

NAND2xp33_ASAP7_75t_SL g580 ( 
.A(n_573),
.B(n_210),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_528),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_515),
.A2(n_389),
.B1(n_212),
.B2(n_250),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_528),
.B(n_539),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_464),
.B(n_371),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_465),
.B(n_371),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_501),
.B(n_384),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_483),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_495),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_455),
.B(n_384),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_515),
.A2(n_212),
.B1(n_250),
.B2(n_217),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_477),
.B(n_384),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_505),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_495),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_459),
.B(n_411),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_452),
.B(n_406),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_479),
.B(n_262),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_541),
.B(n_411),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_542),
.B(n_411),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_544),
.B(n_214),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_548),
.B(n_225),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_509),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_560),
.B(n_232),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_556),
.B(n_233),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_512),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_SL g605 ( 
.A(n_511),
.B(n_217),
.Y(n_605)
);

NOR3xp33_ASAP7_75t_L g606 ( 
.A(n_472),
.B(n_406),
.C(n_283),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_568),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_517),
.B(n_309),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_471),
.A2(n_373),
.B1(n_370),
.B2(n_229),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_481),
.B(n_281),
.Y(n_610)
);

BUFx8_ASAP7_75t_L g611 ( 
.A(n_468),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_514),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_562),
.B(n_241),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_532),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_482),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_456),
.B(n_476),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_521),
.B(n_314),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_521),
.B(n_323),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_568),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_537),
.A2(n_279),
.B1(n_318),
.B2(n_266),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_564),
.B(n_245),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_525),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_499),
.B(n_324),
.Y(n_623)
);

AO221x1_ASAP7_75t_L g624 ( 
.A1(n_570),
.A2(n_318),
.B1(n_342),
.B2(n_266),
.C(n_279),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_568),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_503),
.B(n_331),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_534),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_573),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_447),
.B(n_264),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_537),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_535),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_494),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_447),
.B(n_270),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_461),
.B(n_276),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_576),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_474),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_516),
.B(n_285),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_537),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_525),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_490),
.B(n_287),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_527),
.Y(n_641)
);

AND2x6_ASAP7_75t_L g642 ( 
.A(n_527),
.B(n_335),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_491),
.B(n_336),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_516),
.B(n_290),
.Y(n_644)
);

INVxp67_ASAP7_75t_SL g645 ( 
.A(n_530),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_578),
.B(n_507),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_453),
.Y(n_647)
);

BUFx8_ASAP7_75t_L g648 ( 
.A(n_484),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_498),
.B(n_341),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_478),
.B(n_300),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_454),
.A2(n_373),
.B1(n_370),
.B2(n_280),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_570),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_457),
.A2(n_373),
.B1(n_370),
.B2(n_280),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_540),
.B(n_301),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_478),
.B(n_304),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g656 ( 
.A(n_494),
.B(n_342),
.Y(n_656)
);

NAND2xp33_ASAP7_75t_SL g657 ( 
.A(n_489),
.B(n_305),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_460),
.B(n_319),
.Y(n_658)
);

AND2x6_ASAP7_75t_L g659 ( 
.A(n_533),
.B(n_343),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_466),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_570),
.A2(n_467),
.B1(n_469),
.B2(n_449),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_470),
.B(n_326),
.Y(n_662)
);

NOR2xp67_ASAP7_75t_L g663 ( 
.A(n_520),
.B(n_489),
.Y(n_663)
);

NOR2xp67_ASAP7_75t_L g664 ( 
.A(n_485),
.B(n_496),
.Y(n_664)
);

BUFx6f_ASAP7_75t_SL g665 ( 
.A(n_555),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_449),
.B(n_325),
.Y(n_666)
);

INVx8_ASAP7_75t_L g667 ( 
.A(n_526),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_551),
.Y(n_668)
);

BUFx8_ASAP7_75t_L g669 ( 
.A(n_555),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_551),
.A2(n_373),
.B1(n_370),
.B2(n_280),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_485),
.B(n_339),
.Y(n_671)
);

NOR3xp33_ASAP7_75t_L g672 ( 
.A(n_496),
.B(n_346),
.C(n_243),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_510),
.B(n_345),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_458),
.B(n_326),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_510),
.B(n_206),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_518),
.Y(n_676)
);

NOR2x1p5_ASAP7_75t_L g677 ( 
.A(n_531),
.B(n_352),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_518),
.B(n_353),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_536),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_536),
.B(n_357),
.Y(n_680)
);

AOI221xp5_ASAP7_75t_L g681 ( 
.A1(n_543),
.A2(n_352),
.B1(n_280),
.B2(n_299),
.C(n_327),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_575),
.B(n_355),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_575),
.B(n_248),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_543),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_553),
.B(n_259),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_574),
.B(n_412),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_480),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_546),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_524),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_546),
.B(n_445),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_572),
.B(n_445),
.Y(n_691)
);

OAI22xp33_ASAP7_75t_SL g692 ( 
.A1(n_551),
.A2(n_16),
.B1(n_17),
.B2(n_20),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_529),
.B(n_21),
.Y(n_693)
);

NAND2xp33_ASAP7_75t_L g694 ( 
.A(n_557),
.B(n_359),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_538),
.B(n_359),
.Y(n_695)
);

NOR2xp67_ASAP7_75t_L g696 ( 
.A(n_497),
.B(n_22),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_L g697 ( 
.A(n_577),
.B(n_359),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_545),
.B(n_362),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_502),
.B(n_23),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_587),
.B(n_523),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_632),
.B(n_547),
.Y(n_701)
);

O2A1O1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_607),
.A2(n_571),
.B(n_569),
.C(n_567),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_619),
.A2(n_571),
.B(n_569),
.C(n_567),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_583),
.B(n_549),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_587),
.B(n_25),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_581),
.Y(n_706)
);

OR2x6_ASAP7_75t_L g707 ( 
.A(n_620),
.B(n_549),
.Y(n_707)
);

BUFx4f_ASAP7_75t_L g708 ( 
.A(n_616),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_588),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_579),
.B(n_552),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_639),
.A2(n_554),
.B(n_552),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_652),
.A2(n_566),
.B1(n_565),
.B2(n_563),
.Y(n_712)
);

OAI21xp33_ASAP7_75t_L g713 ( 
.A1(n_605),
.A2(n_558),
.B(n_554),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_579),
.B(n_558),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_641),
.A2(n_561),
.B(n_559),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_630),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_652),
.A2(n_565),
.B1(n_563),
.B2(n_561),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_617),
.B(n_26),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_617),
.B(n_27),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_661),
.A2(n_500),
.B1(n_522),
.B2(n_504),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_618),
.B(n_28),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_668),
.Y(n_722)
);

A2O1A1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_608),
.A2(n_506),
.B(n_522),
.C(n_508),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_656),
.B(n_28),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_667),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_615),
.B(n_638),
.Y(n_726)
);

AND2x4_ASAP7_75t_SL g727 ( 
.A(n_662),
.B(n_513),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_589),
.A2(n_594),
.B(n_646),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_608),
.B(n_29),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_595),
.B(n_30),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_596),
.B(n_31),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_636),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_610),
.B(n_31),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_L g734 ( 
.A(n_663),
.B(n_32),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_597),
.A2(n_519),
.B(n_448),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_668),
.B(n_463),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_598),
.A2(n_670),
.B(n_586),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_668),
.B(n_463),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_667),
.Y(n_739)
);

O2A1O1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_606),
.A2(n_473),
.B(n_493),
.C(n_492),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_648),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_647),
.A2(n_660),
.B(n_585),
.C(n_591),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_SL g743 ( 
.A(n_667),
.B(n_450),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_592),
.Y(n_744)
);

NOR2x1p5_ASAP7_75t_SL g745 ( 
.A(n_699),
.B(n_451),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_643),
.B(n_33),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_582),
.A2(n_493),
.B1(n_487),
.B2(n_475),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_601),
.Y(n_748)
);

NOR3xp33_ASAP7_75t_L g749 ( 
.A(n_657),
.B(n_486),
.C(n_475),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_643),
.B(n_649),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_670),
.A2(n_651),
.B(n_609),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_649),
.B(n_35),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_612),
.B(n_36),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_604),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_623),
.B(n_36),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_584),
.A2(n_399),
.B(n_419),
.C(n_426),
.Y(n_756)
);

AND2x6_ASAP7_75t_SL g757 ( 
.A(n_674),
.B(n_669),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_653),
.A2(n_585),
.B(n_584),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_590),
.A2(n_362),
.B1(n_378),
.B2(n_381),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_653),
.A2(n_488),
.B(n_462),
.Y(n_760)
);

A2O1A1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_591),
.A2(n_399),
.B(n_419),
.C(n_426),
.Y(n_761)
);

OAI21xp33_ASAP7_75t_L g762 ( 
.A1(n_681),
.A2(n_381),
.B(n_378),
.Y(n_762)
);

AOI22x1_ASAP7_75t_L g763 ( 
.A1(n_688),
.A2(n_635),
.B1(n_614),
.B2(n_627),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_669),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_676),
.A2(n_378),
.B1(n_381),
.B2(n_383),
.Y(n_765)
);

OAI321xp33_ASAP7_75t_L g766 ( 
.A1(n_685),
.A2(n_414),
.A3(n_381),
.B1(n_383),
.B2(n_409),
.C(n_378),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_593),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_648),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_628),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_631),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_623),
.B(n_37),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_672),
.A2(n_681),
.B1(n_675),
.B2(n_664),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_626),
.B(n_40),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_640),
.B(n_41),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_687),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_693),
.Y(n_776)
);

A2O1A1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_626),
.A2(n_426),
.B(n_419),
.C(n_399),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_599),
.B(n_600),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_672),
.B(n_42),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_675),
.B(n_42),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_602),
.B(n_43),
.Y(n_781)
);

A2O1A1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_679),
.A2(n_419),
.B(n_399),
.C(n_414),
.Y(n_782)
);

OAI21xp33_ASAP7_75t_L g783 ( 
.A1(n_629),
.A2(n_634),
.B(n_633),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_689),
.Y(n_784)
);

O2A1O1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_692),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_684),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_611),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_580),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_603),
.B(n_383),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_624),
.B(n_677),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_637),
.A2(n_415),
.B1(n_383),
.B2(n_50),
.Y(n_791)
);

OAI21xp33_ASAP7_75t_L g792 ( 
.A1(n_644),
.A2(n_383),
.B(n_49),
.Y(n_792)
);

INVx1_ASAP7_75t_SL g793 ( 
.A(n_642),
.Y(n_793)
);

NOR2x1p5_ASAP7_75t_L g794 ( 
.A(n_665),
.B(n_49),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_650),
.A2(n_655),
.B1(n_666),
.B2(n_621),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_658),
.B(n_54),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_613),
.B(n_56),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_642),
.B(n_57),
.Y(n_798)
);

NOR2x1p5_ASAP7_75t_L g799 ( 
.A(n_665),
.B(n_58),
.Y(n_799)
);

OR2x6_ASAP7_75t_L g800 ( 
.A(n_654),
.B(n_60),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_642),
.B(n_60),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_642),
.Y(n_802)
);

NAND3xp33_ASAP7_75t_L g803 ( 
.A(n_686),
.B(n_61),
.C(n_62),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_671),
.Y(n_804)
);

AO21x1_ASAP7_75t_L g805 ( 
.A1(n_690),
.A2(n_64),
.B(n_65),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_642),
.A2(n_659),
.B1(n_673),
.B2(n_680),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_659),
.B(n_64),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_678),
.B(n_65),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_659),
.B(n_67),
.Y(n_809)
);

BUFx4f_ASAP7_75t_L g810 ( 
.A(n_659),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_683),
.B(n_70),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_682),
.B(n_71),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_695),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_686),
.A2(n_142),
.B(n_94),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_696),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_751),
.A2(n_690),
.B(n_691),
.Y(n_816)
);

NAND3xp33_ASAP7_75t_L g817 ( 
.A(n_758),
.B(n_803),
.C(n_742),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_725),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_725),
.Y(n_819)
);

AO31x2_ASAP7_75t_L g820 ( 
.A1(n_805),
.A2(n_698),
.A3(n_697),
.B(n_694),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_708),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_737),
.A2(n_698),
.B(n_124),
.Y(n_822)
);

OAI21x1_ASAP7_75t_SL g823 ( 
.A1(n_802),
.A2(n_123),
.B(n_125),
.Y(n_823)
);

INVx6_ASAP7_75t_L g824 ( 
.A(n_764),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_744),
.Y(n_825)
);

OAI22x1_ASAP7_75t_L g826 ( 
.A1(n_794),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_708),
.B(n_151),
.Y(n_827)
);

AO31x2_ASAP7_75t_L g828 ( 
.A1(n_720),
.A2(n_153),
.A3(n_154),
.B(n_156),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_772),
.B(n_168),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_757),
.Y(n_830)
);

INVx1_ASAP7_75t_SL g831 ( 
.A(n_706),
.Y(n_831)
);

INVx4_ASAP7_75t_L g832 ( 
.A(n_739),
.Y(n_832)
);

OR2x6_ASAP7_75t_L g833 ( 
.A(n_787),
.B(n_180),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_804),
.B(n_730),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_748),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_776),
.A2(n_187),
.B1(n_189),
.B2(n_196),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_718),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_790),
.B(n_726),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_783),
.A2(n_781),
.B(n_808),
.C(n_762),
.Y(n_839)
);

AND2x2_ASAP7_75t_SL g840 ( 
.A(n_810),
.B(n_802),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_711),
.A2(n_715),
.B(n_795),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_735),
.A2(n_714),
.B(n_710),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_700),
.A2(n_719),
.B(n_721),
.C(n_780),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_731),
.B(n_733),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_754),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_706),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_810),
.A2(n_746),
.B1(n_752),
.B2(n_793),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_704),
.B(n_705),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_707),
.B(n_724),
.Y(n_849)
);

OAI22x1_ASAP7_75t_L g850 ( 
.A1(n_799),
.A2(n_741),
.B1(n_768),
.B2(n_774),
.Y(n_850)
);

OAI22x1_ASAP7_75t_L g851 ( 
.A1(n_774),
.A2(n_769),
.B1(n_767),
.B2(n_709),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_707),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_745),
.A2(n_773),
.B(n_771),
.C(n_755),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_775),
.Y(n_854)
);

AO31x2_ASAP7_75t_L g855 ( 
.A1(n_756),
.A2(n_761),
.A3(n_723),
.B(n_777),
.Y(n_855)
);

CKINVDCx14_ASAP7_75t_R g856 ( 
.A(n_800),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_707),
.B(n_716),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_702),
.A2(n_789),
.B(n_738),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_797),
.B(n_786),
.Y(n_859)
);

AO31x2_ASAP7_75t_L g860 ( 
.A1(n_782),
.A2(n_815),
.A3(n_703),
.B(n_791),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_727),
.B(n_753),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_736),
.A2(n_712),
.B(n_717),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_813),
.Y(n_863)
);

OR2x6_ASAP7_75t_L g864 ( 
.A(n_800),
.B(n_734),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_796),
.A2(n_779),
.B(n_806),
.C(n_785),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_811),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_722),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_749),
.B(n_759),
.Y(n_868)
);

BUFx10_ASAP7_75t_L g869 ( 
.A(n_813),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_798),
.A2(n_801),
.B(n_807),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_809),
.A2(n_792),
.B(n_812),
.Y(n_871)
);

INVx5_ASAP7_75t_L g872 ( 
.A(n_784),
.Y(n_872)
);

AOI21x1_ASAP7_75t_L g873 ( 
.A1(n_765),
.A2(n_766),
.B(n_793),
.Y(n_873)
);

INVx5_ASAP7_75t_L g874 ( 
.A(n_743),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_750),
.B(n_579),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_725),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_744),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_750),
.B(n_579),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_750),
.B(n_579),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_744),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_750),
.B(n_579),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_750),
.B(n_579),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_750),
.B(n_579),
.Y(n_883)
);

OA22x2_ASAP7_75t_L g884 ( 
.A1(n_790),
.A2(n_590),
.B1(n_582),
.B2(n_620),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_732),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_778),
.A2(n_783),
.B(n_728),
.C(n_750),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_708),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_750),
.B(n_579),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_744),
.Y(n_889)
);

NOR2xp67_ASAP7_75t_L g890 ( 
.A(n_802),
.B(n_652),
.Y(n_890)
);

AOI21xp33_ASAP7_75t_L g891 ( 
.A1(n_740),
.A2(n_762),
.B(n_747),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_708),
.Y(n_892)
);

AOI21xp33_ASAP7_75t_L g893 ( 
.A1(n_740),
.A2(n_762),
.B(n_747),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_751),
.A2(n_645),
.B(n_622),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_750),
.B(n_579),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_770),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_778),
.A2(n_783),
.B(n_728),
.C(n_750),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_744),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_744),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_750),
.B(n_579),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_751),
.A2(n_645),
.B(n_622),
.Y(n_901)
);

OAI21xp33_ASAP7_75t_SL g902 ( 
.A1(n_751),
.A2(n_814),
.B(n_619),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_708),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_701),
.B(n_632),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_SL g905 ( 
.A1(n_788),
.A2(n_239),
.B1(n_305),
.B2(n_261),
.Y(n_905)
);

NOR2x1_ASAP7_75t_SL g906 ( 
.A(n_725),
.B(n_739),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_750),
.B(n_778),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_769),
.B(n_632),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_764),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_750),
.A2(n_607),
.B1(n_625),
.B2(n_619),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_744),
.Y(n_911)
);

OAI21xp33_ASAP7_75t_L g912 ( 
.A1(n_750),
.A2(n_778),
.B(n_762),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_R g913 ( 
.A(n_709),
.B(n_573),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_750),
.A2(n_607),
.B1(n_625),
.B2(n_619),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_764),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_764),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_725),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_750),
.B(n_579),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_701),
.B(n_632),
.Y(n_919)
);

AOI21xp33_ASAP7_75t_L g920 ( 
.A1(n_740),
.A2(n_762),
.B(n_747),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_725),
.B(n_739),
.Y(n_921)
);

OAI21x1_ASAP7_75t_SL g922 ( 
.A1(n_802),
.A2(n_814),
.B(n_763),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_701),
.B(n_632),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_770),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_725),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_708),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_750),
.B(n_579),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_778),
.A2(n_783),
.B(n_728),
.C(n_750),
.Y(n_928)
);

O2A1O1Ixp5_ASAP7_75t_L g929 ( 
.A1(n_758),
.A2(n_751),
.B(n_737),
.C(n_729),
.Y(n_929)
);

AOI221x1_ASAP7_75t_L g930 ( 
.A1(n_751),
.A2(n_792),
.B1(n_760),
.B2(n_758),
.C(n_713),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_725),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_725),
.B(n_739),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_750),
.B(n_579),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_744),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_913),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_825),
.Y(n_936)
);

INVxp67_ASAP7_75t_SL g937 ( 
.A(n_831),
.Y(n_937)
);

OAI21xp33_ASAP7_75t_SL g938 ( 
.A1(n_833),
.A2(n_864),
.B(n_907),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_830),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_835),
.Y(n_940)
);

NAND2x1p5_ASAP7_75t_L g941 ( 
.A(n_832),
.B(n_831),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_846),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_921),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_902),
.A2(n_929),
.B(n_897),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_846),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_845),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_877),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_932),
.Y(n_948)
);

AOI21x1_ASAP7_75t_L g949 ( 
.A1(n_930),
.A2(n_922),
.B(n_873),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_896),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_824),
.Y(n_951)
);

OR2x6_ASAP7_75t_L g952 ( 
.A(n_833),
.B(n_864),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_932),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_886),
.A2(n_928),
.B(n_843),
.Y(n_954)
);

INVx4_ASAP7_75t_L g955 ( 
.A(n_818),
.Y(n_955)
);

INVx4_ASAP7_75t_L g956 ( 
.A(n_819),
.Y(n_956)
);

BUFx2_ASAP7_75t_R g957 ( 
.A(n_915),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_841),
.A2(n_839),
.B(n_853),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_904),
.B(n_919),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_884),
.A2(n_882),
.B1(n_933),
.B2(n_895),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_890),
.B(n_833),
.Y(n_961)
);

NAND2x1p5_ASAP7_75t_L g962 ( 
.A(n_819),
.B(n_876),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_902),
.A2(n_901),
.B(n_894),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_867),
.Y(n_964)
);

NOR2x1_ASAP7_75t_SL g965 ( 
.A(n_874),
.B(n_864),
.Y(n_965)
);

BUFx12f_ASAP7_75t_L g966 ( 
.A(n_916),
.Y(n_966)
);

INVx1_ASAP7_75t_SL g967 ( 
.A(n_923),
.Y(n_967)
);

AO21x1_ASAP7_75t_L g968 ( 
.A1(n_836),
.A2(n_837),
.B(n_910),
.Y(n_968)
);

OA21x2_ASAP7_75t_L g969 ( 
.A1(n_817),
.A2(n_893),
.B(n_891),
.Y(n_969)
);

AO21x2_ASAP7_75t_L g970 ( 
.A1(n_920),
.A2(n_817),
.B(n_871),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_875),
.B(n_878),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_842),
.A2(n_822),
.B(n_912),
.Y(n_972)
);

OR2x6_ASAP7_75t_L g973 ( 
.A(n_892),
.B(n_903),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_880),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_889),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_879),
.B(n_881),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_890),
.B(n_906),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_898),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_824),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_821),
.B(n_887),
.Y(n_980)
);

NOR2xp67_ASAP7_75t_SL g981 ( 
.A(n_874),
.B(n_909),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_899),
.Y(n_982)
);

CKINVDCx16_ASAP7_75t_R g983 ( 
.A(n_856),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_926),
.B(n_911),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_924),
.Y(n_985)
);

AO21x2_ASAP7_75t_L g986 ( 
.A1(n_870),
.A2(n_862),
.B(n_816),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_SL g987 ( 
.A(n_840),
.B(n_827),
.Y(n_987)
);

AO31x2_ASAP7_75t_L g988 ( 
.A1(n_910),
.A2(n_914),
.A3(n_847),
.B(n_865),
.Y(n_988)
);

AO21x2_ASAP7_75t_L g989 ( 
.A1(n_829),
.A2(n_868),
.B(n_858),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_908),
.B(n_834),
.Y(n_990)
);

NAND2x1p5_ASAP7_75t_L g991 ( 
.A(n_917),
.B(n_925),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_869),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_883),
.A2(n_927),
.B(n_918),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_SL g994 ( 
.A(n_836),
.B(n_852),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_934),
.Y(n_995)
);

OR2x6_ASAP7_75t_L g996 ( 
.A(n_850),
.B(n_905),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_854),
.Y(n_997)
);

OAI21x1_ASAP7_75t_SL g998 ( 
.A1(n_823),
.A2(n_914),
.B(n_837),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_888),
.A2(n_900),
.B(n_844),
.C(n_848),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_869),
.Y(n_1000)
);

BUFx12f_ASAP7_75t_L g1001 ( 
.A(n_917),
.Y(n_1001)
);

OA21x2_ASAP7_75t_L g1002 ( 
.A1(n_849),
.A2(n_859),
.B(n_828),
.Y(n_1002)
);

AOI221xp5_ASAP7_75t_L g1003 ( 
.A1(n_905),
.A2(n_851),
.B1(n_838),
.B2(n_885),
.C(n_826),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_857),
.B(n_866),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_855),
.Y(n_1005)
);

BUFx8_ASAP7_75t_L g1006 ( 
.A(n_931),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_L g1007 ( 
.A1(n_855),
.A2(n_860),
.B(n_863),
.Y(n_1007)
);

INVxp67_ASAP7_75t_L g1008 ( 
.A(n_861),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_860),
.A2(n_820),
.B(n_872),
.Y(n_1009)
);

BUFx2_ASAP7_75t_SL g1010 ( 
.A(n_872),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_820),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_913),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_825),
.Y(n_1013)
);

CKINVDCx16_ASAP7_75t_R g1014 ( 
.A(n_913),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_904),
.B(n_919),
.Y(n_1015)
);

INVx3_ASAP7_75t_SL g1016 ( 
.A(n_915),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_884),
.A2(n_624),
.B1(n_878),
.B2(n_875),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_904),
.B(n_919),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_825),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_967),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_967),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_936),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_940),
.Y(n_1023)
);

BUFx4f_ASAP7_75t_L g1024 ( 
.A(n_952),
.Y(n_1024)
);

OR2x6_ASAP7_75t_L g1025 ( 
.A(n_952),
.B(n_961),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_946),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_950),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_SL g1028 ( 
.A1(n_965),
.A2(n_998),
.B(n_968),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_950),
.Y(n_1029)
);

AOI221xp5_ASAP7_75t_L g1030 ( 
.A1(n_976),
.A2(n_999),
.B1(n_960),
.B2(n_971),
.C(n_1017),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_937),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_1006),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_976),
.A2(n_990),
.B1(n_1003),
.B2(n_996),
.Y(n_1033)
);

CKINVDCx16_ASAP7_75t_R g1034 ( 
.A(n_1014),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_1003),
.A2(n_996),
.B1(n_952),
.B2(n_1017),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_1006),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_947),
.Y(n_1037)
);

INVx4_ASAP7_75t_L g1038 ( 
.A(n_1001),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_974),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_975),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_978),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_977),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_982),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_985),
.B(n_997),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_1015),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_959),
.B(n_942),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_960),
.A2(n_996),
.B1(n_993),
.B2(n_999),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_985),
.Y(n_1048)
);

INVx4_ASAP7_75t_L g1049 ( 
.A(n_977),
.Y(n_1049)
);

OR2x2_ASAP7_75t_L g1050 ( 
.A(n_942),
.B(n_945),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_997),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_SL g1052 ( 
.A1(n_938),
.A2(n_994),
.B1(n_987),
.B2(n_961),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1011),
.Y(n_1053)
);

BUFx2_ASAP7_75t_R g1054 ( 
.A(n_939),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_995),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_941),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1013),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_1018),
.Y(n_1058)
);

AOI21x1_ASAP7_75t_L g1059 ( 
.A1(n_949),
.A2(n_972),
.B(n_958),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_971),
.B(n_1019),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1009),
.Y(n_1061)
);

AOI21x1_ASAP7_75t_L g1062 ( 
.A1(n_972),
.A2(n_958),
.B(n_954),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_964),
.Y(n_1063)
);

OA21x2_ASAP7_75t_L g1064 ( 
.A1(n_944),
.A2(n_954),
.B(n_963),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_945),
.B(n_1002),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_984),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_984),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_964),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_1016),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_1016),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_935),
.A2(n_1004),
.B1(n_1012),
.B2(n_973),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1002),
.B(n_988),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_994),
.A2(n_987),
.B1(n_1008),
.B2(n_935),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1007),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1053),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1060),
.B(n_992),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1044),
.B(n_1005),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1030),
.A2(n_983),
.B1(n_1008),
.B2(n_1010),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_1033),
.A2(n_1047),
.B1(n_1035),
.B2(n_1024),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1024),
.A2(n_1000),
.B1(n_992),
.B2(n_989),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1060),
.B(n_1000),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1027),
.B(n_988),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1029),
.B(n_988),
.Y(n_1083)
);

BUFx10_ASAP7_75t_L g1084 ( 
.A(n_1032),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1048),
.B(n_988),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_1042),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1074),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1051),
.B(n_970),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1072),
.B(n_970),
.Y(n_1089)
);

INVx4_ASAP7_75t_L g1090 ( 
.A(n_1042),
.Y(n_1090)
);

NAND2xp33_ASAP7_75t_R g1091 ( 
.A(n_1056),
.B(n_939),
.Y(n_1091)
);

OR2x2_ASAP7_75t_L g1092 ( 
.A(n_1046),
.B(n_986),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_1031),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1072),
.B(n_1064),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1055),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_1025),
.B(n_1061),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_1042),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_1020),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_1021),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_1045),
.A2(n_953),
.B1(n_948),
.B2(n_943),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_1046),
.B(n_986),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1022),
.B(n_969),
.Y(n_1102)
);

NAND2x1p5_ASAP7_75t_L g1103 ( 
.A(n_1086),
.B(n_1049),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1094),
.B(n_1089),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1087),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1075),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1094),
.B(n_1064),
.Y(n_1107)
);

OR2x6_ASAP7_75t_L g1108 ( 
.A(n_1086),
.B(n_1090),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1089),
.B(n_1065),
.Y(n_1109)
);

CKINVDCx6p67_ASAP7_75t_R g1110 ( 
.A(n_1086),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1082),
.B(n_1083),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_1097),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_SL g1113 ( 
.A1(n_1086),
.A2(n_1028),
.B1(n_1025),
.B2(n_1063),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1082),
.B(n_1065),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_1096),
.B(n_1061),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1083),
.B(n_1062),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_1093),
.Y(n_1117)
);

BUFx12f_ASAP7_75t_L g1118 ( 
.A(n_1084),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_1097),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1085),
.B(n_1077),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_1079),
.A2(n_1052),
.B1(n_1058),
.B2(n_1073),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1077),
.B(n_1059),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1102),
.B(n_1068),
.Y(n_1123)
);

INVxp67_ASAP7_75t_L g1124 ( 
.A(n_1093),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_1092),
.B(n_1050),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1104),
.B(n_1088),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1107),
.B(n_1102),
.Y(n_1127)
);

NAND4xp25_ASAP7_75t_SL g1128 ( 
.A(n_1113),
.B(n_1078),
.C(n_1079),
.D(n_1069),
.Y(n_1128)
);

BUFx2_ASAP7_75t_SL g1129 ( 
.A(n_1112),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1107),
.B(n_1095),
.Y(n_1130)
);

INVxp67_ASAP7_75t_SL g1131 ( 
.A(n_1117),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1105),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_1115),
.B(n_1096),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1108),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_1115),
.B(n_1107),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1104),
.B(n_1088),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_1108),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1116),
.B(n_1123),
.Y(n_1138)
);

INVxp67_ASAP7_75t_SL g1139 ( 
.A(n_1117),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_1104),
.B(n_1101),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1106),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1108),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1111),
.B(n_1109),
.Y(n_1143)
);

INVx6_ASAP7_75t_L g1144 ( 
.A(n_1108),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1116),
.B(n_1095),
.Y(n_1145)
);

NAND3xp33_ASAP7_75t_L g1146 ( 
.A(n_1134),
.B(n_1078),
.C(n_1098),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1143),
.B(n_1109),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_1144),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_1131),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1143),
.B(n_1111),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1126),
.B(n_1116),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1141),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1141),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1145),
.B(n_1120),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1138),
.B(n_1125),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1132),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1145),
.B(n_1120),
.Y(n_1157)
);

OR2x2_ASAP7_75t_L g1158 ( 
.A(n_1138),
.B(n_1125),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1126),
.B(n_1114),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1136),
.B(n_1114),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1136),
.B(n_1114),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1130),
.B(n_1070),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1130),
.B(n_1034),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1135),
.B(n_1122),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1132),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1151),
.B(n_1164),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_1155),
.B(n_1140),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1156),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1150),
.B(n_1127),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1162),
.B(n_1054),
.Y(n_1170)
);

OAI32xp33_ASAP7_75t_L g1171 ( 
.A1(n_1149),
.A2(n_1142),
.A3(n_1103),
.B1(n_1137),
.B2(n_1090),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1151),
.B(n_1135),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1163),
.A2(n_1128),
.B1(n_1146),
.B2(n_1144),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_1164),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_1155),
.B(n_1140),
.Y(n_1175)
);

INVxp67_ASAP7_75t_SL g1176 ( 
.A(n_1165),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1150),
.B(n_1127),
.Y(n_1177)
);

NOR2xp67_ASAP7_75t_L g1178 ( 
.A(n_1146),
.B(n_1142),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1158),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1158),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1167),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1167),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1174),
.B(n_1166),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1175),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1179),
.B(n_1154),
.Y(n_1185)
);

XOR2x2_ASAP7_75t_L g1186 ( 
.A(n_1170),
.B(n_1036),
.Y(n_1186)
);

XOR2x2_ASAP7_75t_L g1187 ( 
.A(n_1173),
.B(n_1036),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1174),
.B(n_1134),
.Y(n_1188)
);

OAI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1178),
.A2(n_1144),
.B1(n_1142),
.B2(n_1137),
.Y(n_1189)
);

AOI322xp5_ASAP7_75t_L g1190 ( 
.A1(n_1181),
.A2(n_1180),
.A3(n_1177),
.B1(n_1169),
.B2(n_1147),
.C1(n_1166),
.C2(n_1159),
.Y(n_1190)
);

AOI221xp5_ASAP7_75t_L g1191 ( 
.A1(n_1189),
.A2(n_1171),
.B1(n_1128),
.B2(n_1176),
.C(n_1121),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1187),
.A2(n_1108),
.B(n_1142),
.Y(n_1192)
);

NOR4xp25_ASAP7_75t_L g1193 ( 
.A(n_1189),
.B(n_1071),
.C(n_1175),
.D(n_1023),
.Y(n_1193)
);

OA22x2_ASAP7_75t_L g1194 ( 
.A1(n_1188),
.A2(n_1148),
.B1(n_1172),
.B2(n_1108),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1182),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1183),
.A2(n_1144),
.B1(n_1172),
.B2(n_1110),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1184),
.A2(n_1148),
.B1(n_1144),
.B2(n_1135),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1185),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1188),
.A2(n_1135),
.B1(n_1133),
.B2(n_1139),
.Y(n_1199)
);

NOR3xp33_ASAP7_75t_L g1200 ( 
.A(n_1191),
.B(n_979),
.C(n_951),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1198),
.B(n_1185),
.Y(n_1201)
);

NAND3xp33_ASAP7_75t_SL g1202 ( 
.A(n_1193),
.B(n_1103),
.C(n_1113),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1194),
.B(n_1196),
.Y(n_1203)
);

AOI222xp33_ASAP7_75t_L g1204 ( 
.A1(n_1195),
.A2(n_1186),
.B1(n_1147),
.B2(n_1124),
.C1(n_1099),
.C2(n_1160),
.Y(n_1204)
);

OAI211xp5_ASAP7_75t_SL g1205 ( 
.A1(n_1190),
.A2(n_1032),
.B(n_1080),
.C(n_1100),
.Y(n_1205)
);

AOI311xp33_ASAP7_75t_L g1206 ( 
.A1(n_1192),
.A2(n_1067),
.A3(n_1066),
.B(n_1153),
.C(n_1152),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1199),
.A2(n_1103),
.B(n_1090),
.Y(n_1207)
);

AOI211x1_ASAP7_75t_L g1208 ( 
.A1(n_1202),
.A2(n_1160),
.B(n_1161),
.C(n_1159),
.Y(n_1208)
);

NAND4xp75_ASAP7_75t_L g1209 ( 
.A(n_1203),
.B(n_1197),
.C(n_957),
.D(n_1080),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1201),
.Y(n_1210)
);

INVx2_ASAP7_75t_SL g1211 ( 
.A(n_1200),
.Y(n_1211)
);

NOR4xp75_ASAP7_75t_L g1212 ( 
.A(n_1204),
.B(n_957),
.C(n_1157),
.D(n_1028),
.Y(n_1212)
);

NOR3xp33_ASAP7_75t_L g1213 ( 
.A(n_1205),
.B(n_1038),
.C(n_980),
.Y(n_1213)
);

NOR2x1p5_ASAP7_75t_L g1214 ( 
.A(n_1206),
.B(n_966),
.Y(n_1214)
);

NAND4xp75_ASAP7_75t_L g1215 ( 
.A(n_1208),
.B(n_1207),
.C(n_1038),
.D(n_1091),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1210),
.B(n_1168),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1211),
.A2(n_1038),
.B(n_1025),
.Y(n_1217)
);

NOR3xp33_ASAP7_75t_L g1218 ( 
.A(n_1213),
.B(n_980),
.C(n_956),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1213),
.A2(n_1025),
.B1(n_1110),
.B2(n_1129),
.Y(n_1219)
);

AND3x4_ASAP7_75t_L g1220 ( 
.A(n_1212),
.B(n_1119),
.C(n_1112),
.Y(n_1220)
);

NOR3xp33_ASAP7_75t_L g1221 ( 
.A(n_1209),
.B(n_956),
.C(n_955),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1214),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1222),
.B(n_1084),
.Y(n_1223)
);

NOR4xp75_ASAP7_75t_L g1224 ( 
.A(n_1215),
.B(n_1076),
.C(n_1081),
.D(n_1084),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_1216),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1225),
.Y(n_1226)
);

OAI322xp33_ASAP7_75t_L g1227 ( 
.A1(n_1223),
.A2(n_1217),
.A3(n_1219),
.B1(n_1218),
.B2(n_1220),
.C1(n_1057),
.C2(n_1026),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1224),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1226),
.Y(n_1229)
);

OA22x2_ASAP7_75t_L g1230 ( 
.A1(n_1228),
.A2(n_1221),
.B1(n_973),
.B2(n_1129),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1229),
.A2(n_1227),
.B(n_973),
.Y(n_1231)
);

INVxp67_ASAP7_75t_SL g1232 ( 
.A(n_1230),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1229),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1232),
.A2(n_1084),
.B1(n_981),
.B2(n_1118),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1233),
.B(n_1037),
.Y(n_1235)
);

AOI31xp33_ASAP7_75t_L g1236 ( 
.A1(n_1231),
.A2(n_1103),
.A3(n_991),
.B(n_962),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1234),
.Y(n_1237)
);

AOI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1237),
.A2(n_1235),
.B1(n_1236),
.B2(n_1118),
.Y(n_1238)
);

OA21x2_ASAP7_75t_L g1239 ( 
.A1(n_1238),
.A2(n_1040),
.B(n_1039),
.Y(n_1239)
);

OR2x6_ASAP7_75t_L g1240 ( 
.A(n_1239),
.B(n_1118),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1240),
.A2(n_1043),
.B(n_1041),
.Y(n_1241)
);


endmodule