module fake_jpeg_26248_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_22),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_45),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_23),
.B1(n_30),
.B2(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_52),
.B1(n_59),
.B2(n_32),
.Y(n_75)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_26),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_17),
.B1(n_16),
.B2(n_19),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_21),
.B1(n_17),
.B2(n_19),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_25),
.B1(n_20),
.B2(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_28),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_33),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_25),
.B1(n_20),
.B2(n_16),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g88 ( 
.A(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_28),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_71),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_32),
.B1(n_27),
.B2(n_28),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_67),
.A2(n_77),
.B1(n_53),
.B2(n_1),
.Y(n_108)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_28),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_81),
.Y(n_100)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_1),
.Y(n_114)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_32),
.B1(n_27),
.B2(n_18),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_54),
.B(n_47),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_44),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_18),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_89),
.A2(n_3),
.B(n_4),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_61),
.B(n_49),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_88),
.B(n_83),
.Y(n_127)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_97),
.Y(n_134)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_55),
.C(n_33),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_88),
.C(n_66),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_72),
.B(n_18),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_53),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_107),
.B1(n_100),
.B2(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_70),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_0),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_0),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_111),
.B(n_2),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_113),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_114),
.A2(n_77),
.B1(n_71),
.B2(n_82),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_85),
.B(n_75),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_115),
.A2(n_119),
.B(n_96),
.Y(n_153)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_125),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_108),
.B1(n_94),
.B2(n_105),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_117),
.A2(n_123),
.B1(n_124),
.B2(n_138),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_118),
.A2(n_121),
.B(n_126),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_87),
.B(n_82),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_136),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_89),
.B(n_63),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_108),
.A2(n_63),
.B1(n_68),
.B2(n_74),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_89),
.B(n_76),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_129),
.B(n_133),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_100),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_128),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_131),
.Y(n_142)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_103),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_141),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_109),
.B(n_83),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_88),
.C(n_83),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_137),
.B(n_110),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_90),
.B1(n_94),
.B2(n_111),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_144),
.B(n_160),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_131),
.A2(n_104),
.B1(n_114),
.B2(n_95),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_146),
.A2(n_152),
.B1(n_98),
.B2(n_112),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_135),
.Y(n_181)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_154),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_118),
.A2(n_114),
.B1(n_95),
.B2(n_97),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_165),
.B(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_102),
.Y(n_184)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_166),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_112),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_163),
.B(n_169),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_98),
.B1(n_91),
.B2(n_92),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_167),
.B1(n_126),
.B2(n_121),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_91),
.B(n_112),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_125),
.B1(n_116),
.B2(n_122),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_170),
.A2(n_182),
.B1(n_152),
.B2(n_168),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_126),
.C(n_136),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_191),
.C(n_146),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_172),
.A2(n_176),
.B(n_180),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_158),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_174),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_157),
.A2(n_126),
.B(n_121),
.Y(n_176)
);

NOR2xp67_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_121),
.Y(n_178)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_117),
.B(n_137),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_143),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_154),
.A2(n_129),
.B1(n_98),
.B2(n_92),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_186),
.Y(n_201)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_142),
.B(n_145),
.Y(n_187)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_189),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_150),
.A2(n_102),
.B(n_92),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_148),
.B(n_168),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_78),
.Y(n_191)
);

BUFx24_ASAP7_75t_SL g193 ( 
.A(n_149),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_193),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_198),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_153),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_162),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_177),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_150),
.B1(n_159),
.B2(n_166),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_208),
.B1(n_183),
.B2(n_172),
.Y(n_216)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_206),
.C(n_212),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_148),
.C(n_147),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_209),
.Y(n_227)
);

INVxp67_ASAP7_75t_SL g211 ( 
.A(n_185),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_179),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_155),
.C(n_78),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_189),
.A2(n_102),
.B1(n_4),
.B2(n_5),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_213),
.A2(n_186),
.B1(n_175),
.B2(n_188),
.Y(n_223)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_174),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_220),
.Y(n_234)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_181),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_229),
.C(n_206),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_182),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_224),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_225),
.B1(n_209),
.B2(n_207),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_197),
.A2(n_190),
.B1(n_175),
.B2(n_176),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_229),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_177),
.C(n_5),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_200),
.C(n_214),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_227),
.Y(n_248)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_198),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_235),
.A2(n_213),
.B(n_7),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_237),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_195),
.C(n_207),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_241),
.C(n_226),
.Y(n_244)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_223),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_226),
.C(n_215),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_246),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_233),
.B(n_214),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_249),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_237),
.B(n_196),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_8),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_3),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_252),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_7),
.C(n_8),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_253),
.B(n_257),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_245),
.A2(n_242),
.B1(n_238),
.B2(n_234),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_248),
.A2(n_235),
.B1(n_241),
.B2(n_252),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_257),
.Y(n_262)
);

AO21x1_ASAP7_75t_L g260 ( 
.A1(n_255),
.A2(n_247),
.B(n_244),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_260),
.B(n_262),
.Y(n_265)
);

OAI21xp33_ASAP7_75t_SL g263 ( 
.A1(n_254),
.A2(n_258),
.B(n_259),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_263),
.A2(n_9),
.B(n_11),
.Y(n_266)
);

AOI322xp5_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_9),
.A3(n_11),
.B1(n_12),
.B2(n_14),
.C1(n_15),
.C2(n_249),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_9),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_266),
.A2(n_267),
.B(n_261),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_268),
.A2(n_269),
.B(n_12),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_265),
.Y(n_269)
);

BUFx24_ASAP7_75t_SL g271 ( 
.A(n_270),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_271),
.B(n_15),
.Y(n_272)
);


endmodule