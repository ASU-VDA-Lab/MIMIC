module fake_aes_6479_n_709 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_709);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_709;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_4), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_48), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_38), .Y(n_81) );
CKINVDCx14_ASAP7_75t_R g82 ( .A(n_17), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_9), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_64), .Y(n_84) );
INVx4_ASAP7_75t_R g85 ( .A(n_58), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_32), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_6), .Y(n_87) );
CKINVDCx16_ASAP7_75t_R g88 ( .A(n_4), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_34), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_59), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_42), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_37), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_40), .Y(n_93) );
INVx2_ASAP7_75t_SL g94 ( .A(n_27), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_46), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_13), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_70), .Y(n_97) );
INVx1_ASAP7_75t_SL g98 ( .A(n_61), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_45), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_51), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_17), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_26), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_10), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_31), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_72), .Y(n_105) );
BUFx2_ASAP7_75t_L g106 ( .A(n_1), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_2), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_35), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_8), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_14), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_75), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_33), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_11), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_49), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_73), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_30), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_60), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_39), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_47), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_24), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_50), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_6), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_43), .Y(n_124) );
INVxp67_ASAP7_75t_L g125 ( .A(n_18), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_57), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_82), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_126), .Y(n_128) );
INVx5_ASAP7_75t_L g129 ( .A(n_94), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_86), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_126), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_94), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_84), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_86), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_90), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_106), .B(n_0), .Y(n_136) );
BUFx3_ASAP7_75t_L g137 ( .A(n_112), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_90), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_106), .B(n_1), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_92), .Y(n_140) );
AND2x2_ASAP7_75t_SL g141 ( .A(n_112), .B(n_29), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_92), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_97), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_97), .Y(n_144) );
OA21x2_ASAP7_75t_L g145 ( .A1(n_120), .A2(n_28), .B(n_77), .Y(n_145) );
NOR2xp33_ASAP7_75t_SL g146 ( .A(n_81), .B(n_25), .Y(n_146) );
AND2x6_ASAP7_75t_L g147 ( .A(n_120), .B(n_36), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_121), .Y(n_148) );
INVxp67_ASAP7_75t_L g149 ( .A(n_79), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_121), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_115), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_124), .Y(n_152) );
AND2x2_ASAP7_75t_SL g153 ( .A(n_104), .B(n_78), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_81), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_124), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_109), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_80), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_83), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_88), .B(n_2), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_109), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_99), .Y(n_161) );
CKINVDCx11_ASAP7_75t_R g162 ( .A(n_87), .Y(n_162) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_83), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_125), .B(n_3), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_100), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_105), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_108), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_111), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_116), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_153), .A2(n_101), .B1(n_122), .B2(n_107), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_137), .B(n_123), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_132), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_137), .B(n_101), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_131), .Y(n_174) );
BUFx10_ASAP7_75t_L g175 ( .A(n_154), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_131), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_137), .B(n_102), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_138), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_158), .B(n_91), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_138), .Y(n_181) );
AND2x2_ASAP7_75t_SL g182 ( .A(n_141), .B(n_119), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_131), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_132), .Y(n_184) );
XNOR2x2_ASAP7_75t_SL g185 ( .A(n_136), .B(n_123), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_147), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_158), .B(n_102), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_138), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_138), .Y(n_189) );
NAND2x1p5_ASAP7_75t_L g190 ( .A(n_141), .B(n_118), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_138), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_131), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_161), .B(n_114), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_138), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_163), .Y(n_195) );
AOI22xp5_ASAP7_75t_SL g196 ( .A1(n_133), .A2(n_95), .B1(n_114), .B2(n_89), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_141), .B(n_89), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_132), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_161), .B(n_95), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_166), .B(n_113), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_153), .B(n_149), .Y(n_201) );
AND2x6_ASAP7_75t_L g202 ( .A(n_136), .B(n_96), .Y(n_202) );
INVx5_ASAP7_75t_L g203 ( .A(n_147), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_131), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_139), .A2(n_96), .B1(n_103), .B2(n_87), .Y(n_205) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_139), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_140), .Y(n_207) );
OR2x2_ASAP7_75t_L g208 ( .A(n_159), .B(n_103), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_166), .B(n_110), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_167), .B(n_93), .Y(n_210) );
INVx4_ASAP7_75t_L g211 ( .A(n_147), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_132), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_167), .B(n_117), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_130), .B(n_98), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_130), .B(n_3), .Y(n_215) );
AND2x6_ASAP7_75t_L g216 ( .A(n_134), .B(n_85), .Y(n_216) );
CKINVDCx14_ASAP7_75t_R g217 ( .A(n_127), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_140), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_132), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_134), .B(n_5), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_143), .B(n_5), .Y(n_221) );
BUFx10_ASAP7_75t_L g222 ( .A(n_153), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_143), .B(n_7), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_132), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_140), .Y(n_225) );
INVx4_ASAP7_75t_L g226 ( .A(n_147), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_144), .B(n_41), .Y(n_227) );
INVx6_ASAP7_75t_L g228 ( .A(n_129), .Y(n_228) );
BUFx3_ASAP7_75t_L g229 ( .A(n_147), .Y(n_229) );
INVxp33_ASAP7_75t_L g230 ( .A(n_162), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_144), .B(n_7), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_152), .B(n_8), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_186), .B(n_129), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_199), .B(n_152), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_223), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_223), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_223), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_193), .B(n_155), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_182), .A2(n_164), .B1(n_155), .B2(n_147), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_171), .B(n_157), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_186), .B(n_129), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_177), .B(n_157), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_229), .Y(n_243) );
INVx2_ASAP7_75t_SL g244 ( .A(n_206), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_221), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_214), .B(n_142), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_173), .B(n_142), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_171), .B(n_135), .Y(n_248) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_203), .A2(n_147), .B(n_145), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_171), .B(n_156), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_202), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_221), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_212), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_231), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_213), .B(n_135), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_182), .A2(n_147), .B1(n_168), .B2(n_150), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_187), .B(n_168), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_186), .B(n_129), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_212), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_202), .B(n_156), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_180), .B(n_168), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_202), .B(n_150), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_231), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_211), .B(n_129), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_208), .B(n_129), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_232), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_202), .B(n_150), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_202), .B(n_160), .Y(n_268) );
NAND2x2_ASAP7_75t_L g269 ( .A(n_208), .B(n_151), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_202), .B(n_160), .Y(n_270) );
INVx5_ASAP7_75t_L g271 ( .A(n_202), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_217), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_219), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_229), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_211), .B(n_148), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_195), .B(n_128), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_210), .B(n_128), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_182), .A2(n_146), .B1(n_128), .B2(n_169), .Y(n_278) );
O2A1O1Ixp33_ASAP7_75t_L g279 ( .A1(n_201), .A2(n_145), .B(n_148), .C(n_140), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_195), .B(n_148), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_211), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_232), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_215), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_172), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_190), .B(n_169), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_190), .B(n_169), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_219), .Y(n_287) );
INVx2_ASAP7_75t_SL g288 ( .A(n_175), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_224), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_226), .B(n_148), .Y(n_290) );
NOR2x2_ASAP7_75t_L g291 ( .A(n_185), .B(n_9), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_226), .B(n_148), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_220), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_200), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_172), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_190), .A2(n_169), .B1(n_165), .B2(n_148), .Y(n_296) );
BUFx12f_ASAP7_75t_L g297 ( .A(n_175), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_197), .B(n_169), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_170), .A2(n_140), .B1(n_165), .B2(n_169), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_244), .B(n_170), .Y(n_300) );
AOI222xp33_ASAP7_75t_L g301 ( .A1(n_294), .A2(n_276), .B1(n_245), .B2(n_252), .C1(n_254), .C2(n_263), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_281), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_288), .B(n_196), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_250), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_250), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_235), .A2(n_222), .B1(n_205), .B2(n_175), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_266), .A2(n_282), .B1(n_222), .B2(n_236), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_271), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_246), .B(n_222), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_284), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_237), .A2(n_226), .B1(n_209), .B2(n_203), .Y(n_311) );
INVx5_ASAP7_75t_L g312 ( .A(n_271), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_297), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_271), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_281), .Y(n_315) );
BUFx8_ASAP7_75t_L g316 ( .A(n_297), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_260), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_250), .Y(n_318) );
INVx5_ASAP7_75t_L g319 ( .A(n_271), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_260), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_281), .B(n_203), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_256), .A2(n_203), .B1(n_230), .B2(n_140), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_284), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_260), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_240), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_279), .A2(n_203), .B(n_145), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_240), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_240), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_248), .Y(n_329) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_251), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_280), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_281), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_268), .Y(n_333) );
BUFx6f_ASAP7_75t_SL g334 ( .A(n_283), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_249), .A2(n_145), .B(n_227), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_265), .B(n_216), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_251), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_293), .B(n_216), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_265), .B(n_216), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_272), .Y(n_340) );
AO22x1_ASAP7_75t_L g341 ( .A1(n_291), .A2(n_262), .B1(n_267), .B2(n_216), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_261), .B(n_165), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_275), .A2(n_224), .B(n_225), .Y(n_343) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_274), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g345 ( .A1(n_285), .A2(n_286), .B(n_239), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_238), .B(n_216), .Y(n_346) );
OR2x6_ASAP7_75t_L g347 ( .A(n_270), .B(n_165), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_278), .A2(n_165), .B1(n_228), .B2(n_184), .Y(n_348) );
NAND3xp33_ASAP7_75t_L g349 ( .A(n_296), .B(n_184), .C(n_198), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_234), .A2(n_257), .B1(n_255), .B2(n_247), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_295), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_302), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_350), .B(n_242), .Y(n_353) );
NAND2x1p5_ASAP7_75t_L g354 ( .A(n_312), .B(n_243), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_329), .Y(n_355) );
OA21x2_ASAP7_75t_L g356 ( .A1(n_326), .A2(n_298), .B(n_181), .Y(n_356) );
OAI21x1_ASAP7_75t_L g357 ( .A1(n_326), .A2(n_299), .B(n_298), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g358 ( .A1(n_345), .A2(n_292), .B(n_290), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_333), .Y(n_359) );
NAND2xp33_ASAP7_75t_L g360 ( .A(n_302), .B(n_243), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_300), .B(n_303), .Y(n_361) );
AOI21xp5_ASAP7_75t_SL g362 ( .A1(n_348), .A2(n_274), .B(n_243), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_334), .A2(n_269), .B1(n_242), .B2(n_216), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_316), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g365 ( .A1(n_335), .A2(n_346), .B(n_336), .Y(n_365) );
BUFx4f_ASAP7_75t_SL g366 ( .A(n_316), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_324), .B(n_275), .Y(n_367) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_302), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_303), .B(n_277), .Y(n_369) );
AO21x2_ASAP7_75t_L g370 ( .A1(n_335), .A2(n_290), .B(n_292), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_342), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_339), .A2(n_233), .B(n_241), .Y(n_372) );
INVx2_ASAP7_75t_SL g373 ( .A(n_312), .Y(n_373) );
OAI21xp5_ASAP7_75t_L g374 ( .A1(n_343), .A2(n_258), .B(n_233), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_302), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_307), .A2(n_269), .B1(n_165), .B2(n_291), .Y(n_376) );
CKINVDCx8_ASAP7_75t_R g377 ( .A(n_313), .Y(n_377) );
OAI21x1_ASAP7_75t_L g378 ( .A1(n_343), .A2(n_258), .B(n_241), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_334), .B(n_216), .Y(n_379) );
AOI21xp33_ASAP7_75t_L g380 ( .A1(n_301), .A2(n_198), .B(n_178), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_315), .Y(n_381) );
OAI21xp5_ASAP7_75t_L g382 ( .A1(n_338), .A2(n_264), .B(n_289), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_324), .B(n_243), .Y(n_383) );
INVx3_ASAP7_75t_L g384 ( .A(n_312), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_361), .A2(n_307), .B1(n_309), .B2(n_331), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_376), .A2(n_355), .B1(n_353), .B2(n_363), .C(n_369), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_376), .A2(n_322), .B1(n_304), .B2(n_318), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_369), .A2(n_305), .B1(n_306), .B2(n_320), .Y(n_388) );
AO21x2_ASAP7_75t_L g389 ( .A1(n_365), .A2(n_311), .B(n_218), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_355), .A2(n_325), .B1(n_327), .B2(n_328), .C(n_341), .Y(n_390) );
OAI211xp5_ASAP7_75t_L g391 ( .A1(n_377), .A2(n_340), .B(n_317), .C(n_337), .Y(n_391) );
A2O1A1Ixp33_ASAP7_75t_L g392 ( .A1(n_353), .A2(n_330), .B(n_337), .C(n_310), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_371), .A2(n_347), .B1(n_330), .B2(n_308), .Y(n_393) );
BUFx3_ASAP7_75t_L g394 ( .A(n_354), .Y(n_394) );
OAI22xp33_ASAP7_75t_L g395 ( .A1(n_366), .A2(n_319), .B1(n_312), .B2(n_308), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_359), .Y(n_396) );
INVx2_ASAP7_75t_SL g397 ( .A(n_384), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_359), .A2(n_178), .B1(n_225), .B2(n_218), .C(n_194), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_371), .A2(n_347), .B1(n_344), .B2(n_315), .Y(n_399) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_365), .A2(n_264), .B(n_321), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g401 ( .A1(n_358), .A2(n_347), .B1(n_351), .B2(n_323), .C(n_314), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_364), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_367), .Y(n_403) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_377), .A2(n_319), .B1(n_332), .B2(n_315), .Y(n_404) );
OAI211xp5_ASAP7_75t_L g405 ( .A1(n_379), .A2(n_314), .B(n_194), .C(n_191), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_367), .B(n_315), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_356), .A2(n_332), .B(n_349), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_367), .A2(n_344), .B1(n_332), .B2(n_319), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_367), .B(n_332), .Y(n_409) );
OA21x2_ASAP7_75t_L g410 ( .A1(n_357), .A2(n_192), .B(n_183), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_383), .B(n_319), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_368), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_396), .B(n_357), .Y(n_413) );
BUFx2_ASAP7_75t_L g414 ( .A(n_394), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_396), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_403), .B(n_352), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_403), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_406), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_394), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_410), .Y(n_420) );
INVxp67_ASAP7_75t_L g421 ( .A(n_402), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_410), .Y(n_422) );
INVx5_ASAP7_75t_L g423 ( .A(n_394), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_406), .Y(n_424) );
INVxp67_ASAP7_75t_L g425 ( .A(n_411), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_409), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_409), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_397), .B(n_356), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_397), .B(n_356), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_411), .B(n_352), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_386), .B(n_352), .Y(n_431) );
BUFx3_ASAP7_75t_L g432 ( .A(n_412), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_386), .B(n_375), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_387), .B(n_357), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_399), .B(n_356), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_399), .B(n_373), .Y(n_436) );
OAI21xp5_ASAP7_75t_L g437 ( .A1(n_400), .A2(n_358), .B(n_380), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_410), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_410), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_391), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_412), .Y(n_441) );
BUFx2_ASAP7_75t_L g442 ( .A(n_404), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_388), .B(n_373), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_385), .B(n_375), .Y(n_444) );
INVx3_ASAP7_75t_L g445 ( .A(n_389), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_392), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_390), .A2(n_380), .B1(n_383), .B2(n_370), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_407), .Y(n_448) );
OAI211xp5_ASAP7_75t_SL g449 ( .A1(n_421), .A2(n_390), .B(n_393), .C(n_408), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_420), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_415), .B(n_395), .Y(n_451) );
INVx4_ASAP7_75t_L g452 ( .A(n_423), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_415), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_420), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_440), .B(n_10), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g456 ( .A1(n_418), .A2(n_401), .B1(n_398), .B2(n_407), .C(n_374), .Y(n_456) );
INVx2_ASAP7_75t_SL g457 ( .A(n_423), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_418), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_426), .B(n_389), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_420), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_426), .B(n_401), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_427), .B(n_389), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_427), .B(n_389), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_422), .Y(n_464) );
NAND2xp33_ASAP7_75t_L g465 ( .A(n_423), .B(n_368), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_443), .A2(n_383), .B1(n_384), .B2(n_370), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_424), .B(n_375), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_425), .B(n_11), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_417), .B(n_381), .Y(n_469) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_448), .B(n_405), .C(n_398), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_417), .B(n_381), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_430), .B(n_381), .Y(n_472) );
AO21x2_ASAP7_75t_L g473 ( .A1(n_437), .A2(n_362), .B(n_374), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_416), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_436), .A2(n_384), .B(n_383), .C(n_382), .Y(n_475) );
NOR2xp33_ASAP7_75t_SL g476 ( .A(n_423), .B(n_384), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_416), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_430), .Y(n_478) );
AOI222xp33_ASAP7_75t_L g479 ( .A1(n_431), .A2(n_382), .B1(n_13), .B2(n_14), .C1(n_15), .C2(n_16), .Y(n_479) );
AOI22xp33_ASAP7_75t_SL g480 ( .A1(n_442), .A2(n_368), .B1(n_354), .B2(n_370), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_423), .B(n_368), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_423), .Y(n_482) );
INVxp67_ASAP7_75t_SL g483 ( .A(n_428), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_443), .B(n_370), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_431), .B(n_12), .Y(n_485) );
OAI33xp33_ASAP7_75t_L g486 ( .A1(n_448), .A2(n_191), .A3(n_189), .B1(n_188), .B2(n_181), .B3(n_12), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_433), .B(n_368), .Y(n_487) );
OAI33xp33_ASAP7_75t_L g488 ( .A1(n_413), .A2(n_189), .A3(n_188), .B1(n_18), .B2(n_19), .B3(n_15), .Y(n_488) );
BUFx2_ASAP7_75t_L g489 ( .A(n_414), .Y(n_489) );
OAI221xp5_ASAP7_75t_L g490 ( .A1(n_447), .A2(n_362), .B1(n_354), .B2(n_360), .C(n_204), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_433), .B(n_368), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_441), .B(n_16), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_422), .Y(n_493) );
AND2x4_ASAP7_75t_L g494 ( .A(n_423), .B(n_378), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_441), .B(n_19), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_419), .Y(n_496) );
INVx3_ASAP7_75t_SL g497 ( .A(n_436), .Y(n_497) );
NAND4xp25_ASAP7_75t_SL g498 ( .A(n_435), .B(n_20), .C(n_21), .D(n_22), .Y(n_498) );
NAND4xp25_ASAP7_75t_L g499 ( .A(n_434), .B(n_204), .C(n_176), .D(n_179), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_484), .B(n_413), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_450), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_459), .B(n_445), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_483), .B(n_434), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_450), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_459), .B(n_445), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_489), .Y(n_506) );
INVx1_ASAP7_75t_SL g507 ( .A(n_482), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_478), .B(n_414), .Y(n_508) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_470), .A2(n_437), .B(n_439), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_453), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_458), .B(n_444), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_454), .Y(n_512) );
INVx1_ASAP7_75t_SL g513 ( .A(n_482), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_497), .B(n_435), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_463), .B(n_445), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_463), .B(n_445), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_455), .B(n_444), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_497), .B(n_428), .Y(n_518) );
INVx3_ASAP7_75t_L g519 ( .A(n_452), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_487), .B(n_429), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_454), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_460), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_460), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_487), .B(n_429), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_464), .Y(n_525) );
OAI33xp33_ASAP7_75t_L g526 ( .A1(n_485), .A2(n_446), .A3(n_439), .B1(n_438), .B2(n_422), .B3(n_179), .Y(n_526) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_452), .B(n_442), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_464), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_493), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_493), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_491), .B(n_438), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_491), .B(n_438), .Y(n_532) );
NOR3xp33_ASAP7_75t_L g533 ( .A(n_488), .B(n_449), .C(n_468), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_462), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_462), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_474), .B(n_432), .Y(n_536) );
AOI33xp33_ASAP7_75t_L g537 ( .A1(n_466), .A2(n_446), .A3(n_176), .B1(n_192), .B2(n_183), .B3(n_289), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_477), .B(n_432), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_469), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_469), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_465), .A2(n_432), .B(n_378), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_494), .B(n_174), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_492), .B(n_372), .Y(n_543) );
NOR2x1p5_ASAP7_75t_L g544 ( .A(n_482), .B(n_344), .Y(n_544) );
OAI211xp5_ASAP7_75t_L g545 ( .A1(n_479), .A2(n_174), .B(n_207), .C(n_344), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_494), .B(n_174), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_452), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_494), .B(n_174), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_471), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_473), .B(n_174), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_473), .B(n_461), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_473), .B(n_372), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_461), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_496), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_475), .B(n_23), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_451), .A2(n_207), .B1(n_295), .B2(n_273), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_492), .B(n_44), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_495), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_553), .B(n_467), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_502), .B(n_475), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_502), .B(n_480), .Y(n_561) );
NAND2x1p5_ASAP7_75t_L g562 ( .A(n_544), .B(n_457), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_554), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_554), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_505), .B(n_515), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_501), .Y(n_566) );
A2O1A1Ixp33_ASAP7_75t_L g567 ( .A1(n_545), .A2(n_457), .B(n_495), .C(n_476), .Y(n_567) );
NAND2xp33_ASAP7_75t_SL g568 ( .A(n_547), .B(n_481), .Y(n_568) );
AND2x4_ASAP7_75t_L g569 ( .A(n_519), .B(n_481), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_501), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_519), .B(n_481), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_553), .B(n_472), .Y(n_572) );
NOR2x1_ASAP7_75t_L g573 ( .A(n_519), .B(n_498), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_505), .B(n_456), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_510), .Y(n_575) );
AOI211xp5_ASAP7_75t_L g576 ( .A1(n_533), .A2(n_465), .B(n_490), .C(n_499), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_515), .B(n_52), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_510), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_539), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_516), .B(n_53), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_516), .B(n_54), .Y(n_581) );
INVxp33_ASAP7_75t_SL g582 ( .A(n_547), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_539), .Y(n_583) );
OR2x6_ASAP7_75t_L g584 ( .A(n_527), .B(n_486), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_540), .B(n_55), .Y(n_585) );
AOI22xp33_ASAP7_75t_SL g586 ( .A1(n_506), .A2(n_207), .B1(n_62), .B2(n_63), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_540), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_551), .B(n_56), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_551), .B(n_65), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_520), .B(n_66), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_520), .B(n_67), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_549), .Y(n_592) );
INVx3_ASAP7_75t_L g593 ( .A(n_546), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_524), .B(n_68), .Y(n_594) );
NAND2xp33_ASAP7_75t_SL g595 ( .A(n_514), .B(n_69), .Y(n_595) );
INVx2_ASAP7_75t_SL g596 ( .A(n_506), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_503), .B(n_71), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_549), .B(n_74), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_558), .B(n_76), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_518), .B(n_253), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_517), .B(n_253), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_507), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_524), .B(n_259), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_535), .B(n_259), .Y(n_604) );
INVxp67_ASAP7_75t_L g605 ( .A(n_518), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_531), .B(n_273), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_504), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_535), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_531), .B(n_287), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_511), .B(n_287), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_534), .B(n_228), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_608), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_575), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_605), .B(n_503), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_582), .A2(n_514), .B1(n_527), .B2(n_508), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_596), .B(n_500), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_567), .A2(n_555), .B(n_537), .Y(n_617) );
INVxp67_ASAP7_75t_L g618 ( .A(n_596), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_578), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_582), .A2(n_538), .B1(n_513), .B2(n_555), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_566), .Y(n_621) );
NAND2xp67_ASAP7_75t_L g622 ( .A(n_574), .B(n_536), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_566), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_602), .B(n_500), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_570), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_595), .A2(n_526), .B(n_541), .Y(n_626) );
NAND3xp33_ASAP7_75t_L g627 ( .A(n_576), .B(n_552), .C(n_550), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_574), .A2(n_534), .B1(n_536), .B2(n_552), .C(n_557), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_592), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_579), .Y(n_630) );
OAI21xp5_ASAP7_75t_L g631 ( .A1(n_567), .A2(n_556), .B(n_550), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_565), .B(n_543), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_565), .B(n_532), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_572), .B(n_532), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_583), .Y(n_635) );
AOI321xp33_ASAP7_75t_L g636 ( .A1(n_561), .A2(n_525), .A3(n_530), .B1(n_529), .B2(n_528), .C(n_521), .Y(n_636) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_563), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_587), .Y(n_638) );
OAI21xp33_ASAP7_75t_L g639 ( .A1(n_561), .A2(n_573), .B(n_560), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_569), .B(n_571), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_564), .Y(n_641) );
OAI22xp33_ASAP7_75t_SL g642 ( .A1(n_562), .A2(n_525), .B1(n_530), .B2(n_529), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_572), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_560), .A2(n_509), .B1(n_548), .B2(n_542), .Y(n_644) );
OR2x6_ASAP7_75t_L g645 ( .A(n_562), .B(n_544), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_559), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_570), .B(n_509), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_603), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_628), .B(n_603), .Y(n_649) );
AOI211xp5_ASAP7_75t_SL g650 ( .A1(n_639), .A2(n_594), .B(n_591), .C(n_590), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_617), .A2(n_584), .B(n_599), .C(n_597), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_637), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_620), .A2(n_584), .B1(n_593), .B2(n_571), .Y(n_653) );
NOR2xp67_ASAP7_75t_L g654 ( .A(n_615), .B(n_593), .Y(n_654) );
OAI21xp33_ASAP7_75t_L g655 ( .A1(n_622), .A2(n_584), .B(n_589), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_643), .B(n_593), .Y(n_656) );
AOI21xp33_ASAP7_75t_L g657 ( .A1(n_627), .A2(n_584), .B(n_601), .Y(n_657) );
A2O1A1Ixp33_ASAP7_75t_L g658 ( .A1(n_636), .A2(n_568), .B(n_617), .C(n_595), .Y(n_658) );
O2A1O1Ixp33_ASAP7_75t_L g659 ( .A1(n_642), .A2(n_597), .B(n_588), .C(n_589), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_614), .Y(n_660) );
AOI211xp5_ASAP7_75t_SL g661 ( .A1(n_620), .A2(n_590), .B(n_591), .C(n_594), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_629), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_632), .B(n_509), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_616), .Y(n_664) );
XOR2xp5_ASAP7_75t_L g665 ( .A(n_648), .B(n_600), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_615), .A2(n_568), .B1(n_588), .B2(n_577), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_646), .B(n_571), .Y(n_667) );
NAND3x2_ASAP7_75t_L g668 ( .A(n_640), .B(n_569), .C(n_581), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_624), .B(n_609), .Y(n_669) );
INVx1_ASAP7_75t_SL g670 ( .A(n_634), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_612), .Y(n_671) );
INVx1_ASAP7_75t_SL g672 ( .A(n_670), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_652), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_656), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_662), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_653), .A2(n_644), .B1(n_618), .B2(n_630), .C(n_638), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_668), .A2(n_631), .B1(n_635), .B2(n_619), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_658), .A2(n_645), .B(n_626), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_649), .B(n_641), .Y(n_679) );
OAI321xp33_ASAP7_75t_L g680 ( .A1(n_658), .A2(n_631), .A3(n_645), .B1(n_647), .B2(n_581), .C(n_580), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_654), .A2(n_613), .B1(n_645), .B2(n_577), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_666), .A2(n_633), .B1(n_569), .B2(n_580), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_671), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_660), .Y(n_684) );
OAI221xp5_ASAP7_75t_L g685 ( .A1(n_655), .A2(n_647), .B1(n_586), .B2(n_621), .C(n_625), .Y(n_685) );
AOI321xp33_ASAP7_75t_L g686 ( .A1(n_680), .A2(n_651), .A3(n_659), .B1(n_657), .B2(n_661), .C(n_650), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_678), .A2(n_663), .B1(n_664), .B2(n_665), .C(n_669), .Y(n_687) );
AOI211x1_ASAP7_75t_L g688 ( .A1(n_685), .A2(n_667), .B(n_656), .C(n_598), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_676), .A2(n_667), .B1(n_623), .B2(n_585), .C(n_610), .Y(n_689) );
O2A1O1Ixp33_ASAP7_75t_L g690 ( .A1(n_672), .A2(n_604), .B(n_611), .C(n_542), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_672), .A2(n_609), .B1(n_606), .B2(n_548), .Y(n_691) );
NOR4xp25_ASAP7_75t_L g692 ( .A(n_679), .B(n_606), .C(n_607), .D(n_523), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_677), .A2(n_607), .B1(n_528), .B2(n_523), .C(n_521), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_693), .B(n_673), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_691), .B(n_681), .Y(n_695) );
NAND4xp25_ASAP7_75t_L g696 ( .A(n_686), .B(n_682), .C(n_684), .D(n_683), .Y(n_696) );
NOR3xp33_ASAP7_75t_L g697 ( .A(n_687), .B(n_675), .C(n_546), .Y(n_697) );
OR2x2_ASAP7_75t_L g698 ( .A(n_692), .B(n_674), .Y(n_698) );
NAND4xp25_ASAP7_75t_L g699 ( .A(n_696), .B(n_688), .C(n_689), .D(n_690), .Y(n_699) );
NAND3xp33_ASAP7_75t_SL g700 ( .A(n_697), .B(n_504), .C(n_512), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_698), .A2(n_512), .B1(n_522), .B2(n_546), .C(n_228), .Y(n_701) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_701), .Y(n_702) );
INVx1_ASAP7_75t_SL g703 ( .A(n_699), .Y(n_703) );
INVx4_ASAP7_75t_L g704 ( .A(n_702), .Y(n_704) );
OA22x2_ASAP7_75t_L g705 ( .A1(n_703), .A2(n_695), .B1(n_700), .B2(n_694), .Y(n_705) );
INVx4_ASAP7_75t_L g706 ( .A(n_704), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_706), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_707), .B(n_705), .C(n_546), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_708), .A2(n_522), .B(n_228), .Y(n_709) );
endmodule