module fake_jpeg_23465_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_9),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_42),
.A2(n_45),
.B(n_34),
.C(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_0),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_32),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_51),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_50),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_53),
.B(n_58),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_56),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_57),
.B(n_71),
.Y(n_85)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_27),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_68),
.Y(n_108)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_38),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_73),
.Y(n_121)
);

OR2x4_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_25),
.Y(n_89)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_40),
.B(n_34),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_43),
.A2(n_19),
.B1(n_37),
.B2(n_25),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_78),
.A2(n_79),
.B1(n_20),
.B2(n_17),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_30),
.B1(n_26),
.B2(n_37),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_36),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_43),
.A2(n_30),
.B1(n_26),
.B2(n_27),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_19),
.B1(n_35),
.B2(n_28),
.Y(n_93)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_20),
.B1(n_44),
.B2(n_47),
.Y(n_104)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_79),
.B1(n_70),
.B2(n_64),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_87),
.A2(n_114),
.B1(n_5),
.B2(n_6),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_35),
.B(n_26),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_88),
.A2(n_120),
.B(n_10),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_89),
.B(n_91),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_30),
.B1(n_19),
.B2(n_37),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_90),
.A2(n_100),
.B1(n_105),
.B2(n_62),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_25),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_93),
.A2(n_62),
.B1(n_70),
.B2(n_60),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_94),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_97),
.B(n_114),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_31),
.B1(n_29),
.B2(n_24),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_20),
.B1(n_31),
.B2(n_29),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_111),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_55),
.A2(n_47),
.B(n_44),
.C(n_31),
.Y(n_113)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_80),
.A2(n_29),
.B1(n_24),
.B2(n_21),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_117),
.Y(n_148)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_2),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_58),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_66),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_127),
.Y(n_164)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_132),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_126),
.B(n_129),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_47),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_24),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_21),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_134),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_119),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_131),
.Y(n_182)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_84),
.C(n_75),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_133),
.B(n_138),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_21),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_154),
.B1(n_157),
.B2(n_98),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_63),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_147),
.B1(n_90),
.B2(n_100),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_0),
.Y(n_140)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_146),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_1),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_107),
.CI(n_118),
.CON(n_178),
.SN(n_178)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_87),
.A2(n_2),
.B(n_4),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_151),
.B(n_115),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_4),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_102),
.B(n_4),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_152),
.B(n_7),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_86),
.B(n_5),
.Y(n_155)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_121),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_158),
.A2(n_174),
.B1(n_135),
.B2(n_137),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_126),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_168),
.A2(n_12),
.B(n_13),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_169),
.A2(n_177),
.B1(n_183),
.B2(n_184),
.Y(n_204)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_171),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_148),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_172),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_173),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_107),
.B1(n_98),
.B2(n_111),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_132),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_176),
.Y(n_202)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_136),
.A2(n_141),
.B1(n_157),
.B2(n_124),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_123),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_136),
.A2(n_121),
.B1(n_99),
.B2(n_116),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_124),
.A2(n_92),
.B1(n_95),
.B2(n_94),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_125),
.B(n_95),
.Y(n_185)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_189),
.A2(n_191),
.B(n_140),
.Y(n_207)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_134),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_127),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_194),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_129),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_195),
.A2(n_201),
.B1(n_212),
.B2(n_215),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_130),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_199),
.A2(n_203),
.B(n_216),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_169),
.A2(n_154),
.B1(n_122),
.B2(n_138),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_200),
.A2(n_214),
.B1(n_218),
.B2(n_181),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_188),
.A2(n_122),
.B1(n_154),
.B2(n_131),
.Y(n_201)
);

NOR2xp67_ASAP7_75t_SL g203 ( 
.A(n_172),
.B(n_151),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_167),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_206),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_189),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_163),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_175),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_142),
.B1(n_143),
.B2(n_146),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_177),
.A2(n_153),
.B1(n_144),
.B2(n_155),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_164),
.A2(n_144),
.B1(n_152),
.B2(n_151),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_166),
.A2(n_191),
.B1(n_165),
.B2(n_168),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_184),
.A2(n_110),
.B1(n_103),
.B2(n_10),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_161),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_219),
.A2(n_162),
.B1(n_159),
.B2(n_190),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_183),
.A2(n_9),
.B(n_12),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_160),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_160),
.B(n_13),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_162),
.C(n_159),
.Y(n_234)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_224),
.A2(n_245),
.B(n_16),
.Y(n_265)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_227),
.Y(n_249)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_229),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_230),
.A2(n_218),
.B1(n_192),
.B2(n_216),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_178),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_238),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_182),
.Y(n_233)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_240),
.C(n_222),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_196),
.B(n_170),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_235),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_243),
.B1(n_220),
.B2(n_219),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_178),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_173),
.C(n_190),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_212),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_210),
.B(n_13),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_244),
.Y(n_257)
);

OAI21xp33_ASAP7_75t_L g245 ( 
.A1(n_203),
.A2(n_14),
.B(n_15),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_204),
.A2(n_192),
.B1(n_200),
.B2(n_214),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_247),
.A2(n_201),
.B1(n_195),
.B2(n_215),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_250),
.C(n_260),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_237),
.C(n_224),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_255),
.A2(n_259),
.B1(n_261),
.B2(n_263),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_258),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_232),
.A2(n_199),
.B1(n_208),
.B2(n_213),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_231),
.B(n_199),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_208),
.B1(n_213),
.B2(n_217),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_262),
.B(n_246),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_236),
.A2(n_217),
.B1(n_221),
.B2(n_205),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_16),
.C(n_237),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_250),
.C(n_234),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_230),
.B(n_227),
.Y(n_283)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_261),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_273),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_233),
.Y(n_270)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_265),
.B(n_240),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_271),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_252),
.B(n_233),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_276),
.Y(n_298)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_281),
.B1(n_284),
.B2(n_252),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_248),
.C(n_254),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_225),
.B(n_247),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_280),
.A2(n_282),
.B(n_256),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_251),
.A2(n_225),
.B(n_242),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_283),
.A2(n_285),
.B(n_260),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_251),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_253),
.B(n_238),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_274),
.A2(n_258),
.B1(n_264),
.B2(n_249),
.Y(n_287)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_288),
.A2(n_290),
.B(n_299),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_289),
.B(n_271),
.CI(n_285),
.CON(n_304),
.SN(n_304)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_294),
.C(n_295),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_254),
.C(n_256),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_257),
.C(n_279),
.Y(n_295)
);

XOR2x1_ASAP7_75t_SL g296 ( 
.A(n_283),
.B(n_280),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_296),
.B(n_290),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_270),
.A2(n_269),
.B(n_276),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_277),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_308),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_278),
.C(n_282),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_295),
.C(n_292),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_304),
.B(n_306),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_297),
.B(n_275),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_281),
.Y(n_307)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_307),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_298),
.A2(n_292),
.B(n_299),
.Y(n_309)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_309),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_300),
.C(n_291),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_293),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_300),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_289),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_287),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_308),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_317),
.B(n_302),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_315),
.A2(n_301),
.B(n_298),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_318),
.B(n_316),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_320),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_322),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_310),
.C(n_314),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_327),
.C(n_312),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_312),
.Y(n_327)
);

OA21x2_ASAP7_75t_SL g329 ( 
.A1(n_328),
.A2(n_324),
.B(n_311),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_319),
.C(n_291),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_330),
.B(n_304),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_304),
.Y(n_332)
);


endmodule