module real_aes_6306_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g482 ( .A1(n_0), .A2(n_186), .B(n_483), .C(n_486), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_1), .B(n_477), .Y(n_488) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
INVx1_ASAP7_75t_L g235 ( .A(n_3), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_4), .B(n_174), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_5), .A2(n_461), .B(n_531), .Y(n_530) );
OAI22xp5_ASAP7_75t_SL g756 ( .A1(n_6), .A2(n_9), .B1(n_444), .B2(n_757), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_6), .Y(n_757) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_7), .A2(n_191), .B(n_540), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_8), .A2(n_38), .B1(n_147), .B2(n_159), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_9), .A2(n_131), .B1(n_132), .B2(n_444), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_9), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_10), .B(n_191), .Y(n_224) );
AND2x6_ASAP7_75t_L g162 ( .A(n_11), .B(n_163), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_12), .A2(n_162), .B(n_464), .C(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g106 ( .A(n_13), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_13), .B(n_39), .Y(n_125) );
INVx1_ASAP7_75t_L g143 ( .A(n_14), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_15), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g229 ( .A(n_16), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_17), .B(n_174), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_18), .B(n_189), .Y(n_207) );
AO32x2_ASAP7_75t_L g183 ( .A1(n_19), .A2(n_184), .A3(n_188), .B1(n_190), .B2(n_191), .Y(n_183) );
AOI222xp33_ASAP7_75t_SL g127 ( .A1(n_20), .A2(n_92), .B1(n_128), .B2(n_742), .C1(n_743), .C2(n_745), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_20), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_21), .B(n_147), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_22), .B(n_189), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_23), .A2(n_54), .B1(n_147), .B2(n_159), .Y(n_187) );
AOI22xp33_ASAP7_75t_SL g200 ( .A1(n_24), .A2(n_79), .B1(n_147), .B2(n_151), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_25), .B(n_147), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g463 ( .A1(n_26), .A2(n_190), .B(n_464), .C(n_466), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_27), .A2(n_190), .B(n_464), .C(n_543), .Y(n_542) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_28), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_29), .B(n_139), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_30), .A2(n_461), .B(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_31), .B(n_139), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_32), .A2(n_101), .B1(n_114), .B2(n_760), .Y(n_100) );
INVx2_ASAP7_75t_L g149 ( .A(n_33), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_34), .A2(n_495), .B(n_496), .C(n_500), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_35), .B(n_147), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_36), .B(n_139), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_37), .B(n_154), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_39), .B(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_40), .B(n_460), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_41), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_42), .B(n_174), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_43), .B(n_461), .Y(n_541) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_44), .A2(n_495), .B(n_500), .C(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_45), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_46), .B(n_147), .Y(n_217) );
INVx1_ASAP7_75t_L g484 ( .A(n_47), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_48), .A2(n_88), .B1(n_159), .B2(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g523 ( .A(n_49), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_50), .B(n_147), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_51), .B(n_147), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_52), .B(n_461), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_53), .B(n_222), .Y(n_221) );
AOI22xp33_ASAP7_75t_SL g211 ( .A1(n_55), .A2(n_59), .B1(n_147), .B2(n_151), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_56), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_57), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_58), .B(n_147), .Y(n_248) );
INVx1_ASAP7_75t_L g163 ( .A(n_60), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_61), .B(n_461), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_62), .B(n_477), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_63), .A2(n_222), .B(n_232), .C(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_64), .B(n_147), .Y(n_236) );
INVx1_ASAP7_75t_L g142 ( .A(n_65), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_66), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_67), .B(n_174), .Y(n_498) );
AO32x2_ASAP7_75t_L g196 ( .A1(n_68), .A2(n_190), .A3(n_191), .B1(n_197), .B2(n_201), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_69), .B(n_175), .Y(n_554) );
INVx1_ASAP7_75t_L g247 ( .A(n_70), .Y(n_247) );
INVx1_ASAP7_75t_L g172 ( .A(n_71), .Y(n_172) );
CKINVDCx16_ASAP7_75t_R g480 ( .A(n_72), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_73), .B(n_468), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_74), .A2(n_464), .B(n_500), .C(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_75), .B(n_151), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g532 ( .A(n_76), .Y(n_532) );
INVx1_ASAP7_75t_L g113 ( .A(n_77), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_78), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_80), .B(n_159), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_81), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_82), .B(n_151), .Y(n_178) );
INVx2_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_84), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_85), .B(n_161), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_86), .B(n_151), .Y(n_218) );
INVx2_ASAP7_75t_L g110 ( .A(n_87), .Y(n_110) );
OR2x2_ASAP7_75t_L g122 ( .A(n_87), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g447 ( .A(n_87), .B(n_124), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_89), .A2(n_99), .B1(n_151), .B2(n_152), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_90), .B(n_461), .Y(n_493) );
INVx1_ASAP7_75t_L g497 ( .A(n_91), .Y(n_497) );
INVxp67_ASAP7_75t_L g535 ( .A(n_93), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_94), .B(n_151), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_95), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g510 ( .A(n_96), .Y(n_510) );
INVx1_ASAP7_75t_L g550 ( .A(n_97), .Y(n_550) );
AND2x2_ASAP7_75t_L g525 ( .A(n_98), .B(n_139), .Y(n_525) );
INVx1_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g762 ( .A(n_103), .Y(n_762) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx14_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_110), .C(n_111), .Y(n_108) );
AND2x2_ASAP7_75t_L g124 ( .A(n_109), .B(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g741 ( .A(n_110), .B(n_124), .Y(n_741) );
NOR2x2_ASAP7_75t_L g747 ( .A(n_110), .B(n_123), .Y(n_747) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
AOI22x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_127), .B1(n_748), .B2(n_749), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_120), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g748 ( .A(n_118), .Y(n_748) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g749 ( .A1(n_120), .A2(n_750), .B(n_758), .Y(n_749) );
NOR2xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_126), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g759 ( .A(n_122), .Y(n_759) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22x1_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_445), .B1(n_448), .B2(n_739), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_130), .A2(n_449), .B1(n_739), .B2(n_744), .Y(n_743) );
OAI22xp5_ASAP7_75t_SL g754 ( .A1(n_131), .A2(n_132), .B1(n_755), .B2(n_756), .Y(n_754) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OR2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_366), .Y(n_132) );
NAND5xp2_ASAP7_75t_L g133 ( .A(n_134), .B(n_285), .C(n_300), .D(n_326), .E(n_348), .Y(n_133) );
NOR2xp33_ASAP7_75t_SL g134 ( .A(n_135), .B(n_265), .Y(n_134) );
OAI221xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_202), .B1(n_238), .B2(n_254), .C(n_255), .Y(n_135) );
NOR2xp33_ASAP7_75t_SL g136 ( .A(n_137), .B(n_192), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_137), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_SL g442 ( .A(n_137), .Y(n_442) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_165), .Y(n_137) );
INVx1_ASAP7_75t_L g282 ( .A(n_138), .Y(n_282) );
AND2x2_ASAP7_75t_L g284 ( .A(n_138), .B(n_183), .Y(n_284) );
AND2x2_ASAP7_75t_L g294 ( .A(n_138), .B(n_182), .Y(n_294) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_138), .Y(n_312) );
INVx1_ASAP7_75t_L g322 ( .A(n_138), .Y(n_322) );
OR2x2_ASAP7_75t_L g360 ( .A(n_138), .B(n_259), .Y(n_360) );
INVx2_ASAP7_75t_L g410 ( .A(n_138), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_138), .B(n_258), .Y(n_427) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_144), .B(n_164), .Y(n_138) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_139), .A2(n_169), .B(n_181), .Y(n_168) );
INVx2_ASAP7_75t_L g201 ( .A(n_139), .Y(n_201) );
INVx1_ASAP7_75t_L g474 ( .A(n_139), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_139), .A2(n_493), .B(n_494), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_139), .A2(n_520), .B(n_521), .Y(n_519) );
AND2x2_ASAP7_75t_SL g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_L g189 ( .A(n_140), .B(n_141), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
OAI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_156), .B(n_162), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_150), .B(n_153), .Y(n_145) );
INVx3_ASAP7_75t_L g171 ( .A(n_147), .Y(n_171) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_147), .Y(n_512) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g159 ( .A(n_148), .Y(n_159) );
BUFx3_ASAP7_75t_L g199 ( .A(n_148), .Y(n_199) );
AND2x6_ASAP7_75t_L g464 ( .A(n_148), .B(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g152 ( .A(n_149), .Y(n_152) );
INVx1_ASAP7_75t_L g223 ( .A(n_149), .Y(n_223) );
INVx2_ASAP7_75t_L g230 ( .A(n_151), .Y(n_230) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_155), .Y(n_161) );
INVx3_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
AND2x2_ASAP7_75t_L g462 ( .A(n_155), .B(n_223), .Y(n_462) );
INVx1_ASAP7_75t_L g465 ( .A(n_155), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_160), .Y(n_156) );
O2A1O1Ixp5_ASAP7_75t_L g246 ( .A1(n_160), .A2(n_234), .B(n_247), .C(n_248), .Y(n_246) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_161), .A2(n_185), .B1(n_186), .B2(n_187), .Y(n_184) );
OAI22xp5_ASAP7_75t_SL g197 ( .A1(n_161), .A2(n_175), .B1(n_198), .B2(n_200), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g209 ( .A1(n_161), .A2(n_186), .B1(n_210), .B2(n_211), .Y(n_209) );
INVx4_ASAP7_75t_L g485 ( .A(n_161), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g169 ( .A1(n_162), .A2(n_170), .B(n_176), .Y(n_169) );
BUFx3_ASAP7_75t_L g190 ( .A(n_162), .Y(n_190) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_162), .A2(n_216), .B(n_219), .Y(n_215) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_162), .A2(n_228), .B(n_233), .Y(n_227) );
AND2x4_ASAP7_75t_L g461 ( .A(n_162), .B(n_462), .Y(n_461) );
INVx4_ASAP7_75t_SL g487 ( .A(n_162), .Y(n_487) );
NAND2x1p5_ASAP7_75t_L g551 ( .A(n_162), .B(n_462), .Y(n_551) );
NOR2xp67_ASAP7_75t_L g165 ( .A(n_166), .B(n_182), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_167), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_167), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_SL g342 ( .A(n_167), .B(n_282), .Y(n_342) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_168), .Y(n_194) );
INVx2_ASAP7_75t_L g259 ( .A(n_168), .Y(n_259) );
OR2x2_ASAP7_75t_L g321 ( .A(n_168), .B(n_322), .Y(n_321) );
O2A1O1Ixp5_ASAP7_75t_SL g170 ( .A1(n_171), .A2(n_172), .B(n_173), .C(n_174), .Y(n_170) );
INVx2_ASAP7_75t_L g186 ( .A(n_174), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_174), .A2(n_217), .B(n_218), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_174), .A2(n_244), .B(n_245), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_174), .B(n_535), .Y(n_534) );
INVx5_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_179), .Y(n_176) );
INVx1_ASAP7_75t_L g232 ( .A(n_179), .Y(n_232) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g468 ( .A(n_180), .Y(n_468) );
AND2x2_ASAP7_75t_L g260 ( .A(n_182), .B(n_196), .Y(n_260) );
AND2x2_ASAP7_75t_L g277 ( .A(n_182), .B(n_257), .Y(n_277) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g195 ( .A(n_183), .B(n_196), .Y(n_195) );
BUFx2_ASAP7_75t_L g280 ( .A(n_183), .Y(n_280) );
AND2x2_ASAP7_75t_L g409 ( .A(n_183), .B(n_410), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_186), .A2(n_220), .B(n_221), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_186), .A2(n_234), .B(n_235), .C(n_236), .Y(n_233) );
INVx2_ASAP7_75t_L g226 ( .A(n_188), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_188), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_189), .Y(n_191) );
NAND3xp33_ASAP7_75t_L g208 ( .A(n_190), .B(n_209), .C(n_212), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g242 ( .A1(n_190), .A2(n_243), .B(n_246), .Y(n_242) );
INVx4_ASAP7_75t_L g212 ( .A(n_191), .Y(n_212) );
OA21x2_ASAP7_75t_L g214 ( .A1(n_191), .A2(n_215), .B(n_224), .Y(n_214) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_191), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_191), .A2(n_541), .B(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g254 ( .A(n_192), .Y(n_254) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_195), .Y(n_192) );
AND2x2_ASAP7_75t_L g372 ( .A(n_193), .B(n_260), .Y(n_372) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g373 ( .A(n_194), .B(n_284), .Y(n_373) );
O2A1O1Ixp33_ASAP7_75t_L g340 ( .A1(n_195), .A2(n_341), .B(n_343), .C(n_345), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_195), .B(n_341), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_195), .A2(n_271), .B1(n_414), .B2(n_415), .C(n_417), .Y(n_413) );
INVx1_ASAP7_75t_L g257 ( .A(n_196), .Y(n_257) );
INVx1_ASAP7_75t_L g293 ( .A(n_196), .Y(n_293) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_196), .Y(n_302) );
INVx2_ASAP7_75t_L g486 ( .A(n_199), .Y(n_486) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_199), .Y(n_499) );
INVx1_ASAP7_75t_L g471 ( .A(n_201), .Y(n_471) );
INVx1_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_213), .Y(n_203) );
AND2x2_ASAP7_75t_L g319 ( .A(n_204), .B(n_264), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_204), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_205), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g411 ( .A(n_205), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g443 ( .A(n_205), .Y(n_443) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx3_ASAP7_75t_L g273 ( .A(n_206), .Y(n_273) );
AND2x2_ASAP7_75t_L g299 ( .A(n_206), .B(n_253), .Y(n_299) );
NOR2x1_ASAP7_75t_L g308 ( .A(n_206), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g315 ( .A(n_206), .B(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
INVx1_ASAP7_75t_L g251 ( .A(n_207), .Y(n_251) );
AO21x1_ASAP7_75t_L g250 ( .A1(n_209), .A2(n_212), .B(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g477 ( .A(n_212), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_212), .B(n_502), .Y(n_501) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_212), .A2(n_507), .B(n_514), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_212), .B(n_515), .Y(n_514) );
AO21x2_ASAP7_75t_L g548 ( .A1(n_212), .A2(n_549), .B(n_556), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_213), .B(n_355), .Y(n_390) );
INVx1_ASAP7_75t_SL g394 ( .A(n_213), .Y(n_394) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_225), .Y(n_213) );
INVx3_ASAP7_75t_L g253 ( .A(n_214), .Y(n_253) );
AND2x2_ASAP7_75t_L g264 ( .A(n_214), .B(n_241), .Y(n_264) );
AND2x2_ASAP7_75t_L g286 ( .A(n_214), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g331 ( .A(n_214), .B(n_325), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_214), .B(n_263), .Y(n_412) );
INVx2_ASAP7_75t_L g234 ( .A(n_222), .Y(n_234) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g252 ( .A(n_225), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g263 ( .A(n_225), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_225), .B(n_241), .Y(n_288) );
AND2x2_ASAP7_75t_L g324 ( .A(n_225), .B(n_325), .Y(n_324) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_237), .Y(n_225) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_226), .A2(n_242), .B(n_249), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_231), .C(n_232), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_230), .A2(n_544), .B(n_545), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_230), .A2(n_554), .B(n_555), .Y(n_553) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_232), .A2(n_510), .B(n_511), .C(n_512), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_234), .A2(n_467), .B(n_469), .Y(n_466) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_252), .Y(n_239) );
INVx1_ASAP7_75t_L g304 ( .A(n_240), .Y(n_304) );
AND2x2_ASAP7_75t_L g346 ( .A(n_240), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_240), .B(n_267), .Y(n_352) );
AOI21xp5_ASAP7_75t_SL g426 ( .A1(n_240), .A2(n_258), .B(n_281), .Y(n_426) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_250), .Y(n_240) );
OR2x2_ASAP7_75t_L g269 ( .A(n_241), .B(n_250), .Y(n_269) );
AND2x2_ASAP7_75t_L g316 ( .A(n_241), .B(n_253), .Y(n_316) );
INVx2_ASAP7_75t_L g325 ( .A(n_241), .Y(n_325) );
INVx1_ASAP7_75t_L g431 ( .A(n_241), .Y(n_431) );
AND2x2_ASAP7_75t_L g355 ( .A(n_250), .B(n_325), .Y(n_355) );
INVx1_ASAP7_75t_L g380 ( .A(n_250), .Y(n_380) );
AND2x2_ASAP7_75t_L g289 ( .A(n_252), .B(n_273), .Y(n_289) );
AND2x2_ASAP7_75t_L g301 ( .A(n_252), .B(n_302), .Y(n_301) );
INVx2_ASAP7_75t_SL g419 ( .A(n_252), .Y(n_419) );
INVx2_ASAP7_75t_L g309 ( .A(n_253), .Y(n_309) );
AND2x2_ASAP7_75t_L g347 ( .A(n_253), .B(n_263), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_253), .B(n_431), .Y(n_430) );
OAI21xp33_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_260), .B(n_261), .Y(n_255) );
AND2x2_ASAP7_75t_L g362 ( .A(n_256), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g416 ( .A(n_256), .Y(n_416) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g336 ( .A(n_257), .Y(n_336) );
BUFx2_ASAP7_75t_L g435 ( .A(n_257), .Y(n_435) );
BUFx2_ASAP7_75t_L g306 ( .A(n_258), .Y(n_306) );
AND2x2_ASAP7_75t_L g408 ( .A(n_258), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g391 ( .A(n_259), .Y(n_391) );
AND2x4_ASAP7_75t_L g318 ( .A(n_260), .B(n_281), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_260), .B(n_342), .Y(n_354) );
AOI32xp33_ASAP7_75t_L g278 ( .A1(n_261), .A2(n_279), .A3(n_281), .B1(n_283), .B2(n_284), .Y(n_278) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
INVx3_ASAP7_75t_L g267 ( .A(n_262), .Y(n_267) );
OR2x2_ASAP7_75t_L g403 ( .A(n_262), .B(n_359), .Y(n_403) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g272 ( .A(n_263), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g379 ( .A(n_263), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g271 ( .A(n_264), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g283 ( .A(n_264), .B(n_273), .Y(n_283) );
INVx1_ASAP7_75t_L g404 ( .A(n_264), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_264), .B(n_379), .Y(n_437) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_270), .B(n_274), .C(n_278), .Y(n_265) );
OAI322xp33_ASAP7_75t_L g374 ( .A1(n_266), .A2(n_311), .A3(n_375), .B1(n_377), .B2(n_381), .C1(n_382), .C2(n_386), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVxp67_ASAP7_75t_L g339 ( .A(n_267), .Y(n_339) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g393 ( .A(n_269), .B(n_394), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_269), .B(n_309), .Y(n_440) );
INVxp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g332 ( .A(n_272), .Y(n_332) );
OR2x2_ASAP7_75t_L g418 ( .A(n_273), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_276), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g327 ( .A(n_277), .B(n_306), .Y(n_327) );
AND2x2_ASAP7_75t_L g398 ( .A(n_277), .B(n_311), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_277), .B(n_385), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g285 ( .A1(n_279), .A2(n_286), .B1(n_289), .B2(n_290), .C(n_295), .Y(n_285) );
OR2x2_ASAP7_75t_L g296 ( .A(n_279), .B(n_292), .Y(n_296) );
AND2x2_ASAP7_75t_L g384 ( .A(n_279), .B(n_385), .Y(n_384) );
AOI32xp33_ASAP7_75t_L g423 ( .A1(n_279), .A2(n_309), .A3(n_424), .B1(n_425), .B2(n_428), .Y(n_423) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND3xp33_ASAP7_75t_L g357 ( .A(n_280), .B(n_316), .C(n_339), .Y(n_357) );
AND2x2_ASAP7_75t_L g383 ( .A(n_280), .B(n_376), .Y(n_383) );
INVxp67_ASAP7_75t_L g363 ( .A(n_281), .Y(n_363) );
BUFx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_284), .B(n_336), .Y(n_392) );
INVx2_ASAP7_75t_L g402 ( .A(n_284), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_284), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g371 ( .A(n_287), .Y(n_371) );
OR2x2_ASAP7_75t_L g297 ( .A(n_288), .B(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_290), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_294), .Y(n_290) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_293), .Y(n_376) );
AND2x2_ASAP7_75t_L g335 ( .A(n_294), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g381 ( .A(n_294), .Y(n_381) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_294), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AOI21xp33_ASAP7_75t_SL g320 ( .A1(n_296), .A2(n_321), .B(n_323), .Y(n_320) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g414 ( .A(n_299), .B(n_324), .Y(n_414) );
AOI211xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_303), .B(n_313), .C(n_320), .Y(n_300) );
AND2x2_ASAP7_75t_L g344 ( .A(n_302), .B(n_312), .Y(n_344) );
INVx2_ASAP7_75t_L g359 ( .A(n_302), .Y(n_359) );
OR2x2_ASAP7_75t_L g397 ( .A(n_302), .B(n_360), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_302), .B(n_440), .Y(n_439) );
AOI211xp5_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_305), .B(n_307), .C(n_310), .Y(n_303) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_306), .B(n_344), .Y(n_343) );
OAI211xp5_ASAP7_75t_L g425 ( .A1(n_307), .A2(n_402), .B(n_426), .C(n_427), .Y(n_425) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2x1p5_ASAP7_75t_L g323 ( .A(n_308), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g365 ( .A(n_309), .B(n_355), .Y(n_365) );
INVx1_ASAP7_75t_L g370 ( .A(n_309), .Y(n_370) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_314), .B(n_317), .Y(n_313) );
INVxp33_ASAP7_75t_L g421 ( .A(n_315), .Y(n_421) );
AND2x2_ASAP7_75t_L g400 ( .A(n_316), .B(n_379), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_321), .A2(n_383), .B(n_384), .Y(n_382) );
OAI322xp33_ASAP7_75t_L g401 ( .A1(n_323), .A2(n_402), .A3(n_403), .B1(n_404), .B2(n_405), .C1(n_407), .C2(n_411), .Y(n_401) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_328), .B1(n_333), .B2(n_337), .C(n_340), .Y(n_326) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g378 ( .A(n_331), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g422 ( .A(n_335), .Y(n_422) );
INVxp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_338), .B(n_358), .Y(n_424) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g387 ( .A(n_347), .B(n_355), .Y(n_387) );
AOI221xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_351), .B1(n_353), .B2(n_355), .C(n_356), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_351), .A2(n_368), .B1(n_372), .B2(n_373), .C(n_374), .Y(n_367) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVxp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_355), .B(n_370), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_358), .B1(n_361), .B2(n_364), .Y(n_356) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx2_ASAP7_75t_SL g385 ( .A(n_360), .Y(n_385) );
INVxp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND5xp2_ASAP7_75t_L g366 ( .A(n_367), .B(n_388), .C(n_413), .D(n_423), .E(n_433), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_369), .B(n_371), .Y(n_368) );
NOR4xp25_ASAP7_75t_L g441 ( .A(n_370), .B(n_376), .C(n_442), .D(n_443), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_373), .A2(n_434), .B1(n_436), .B2(n_438), .C(n_441), .Y(n_433) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g432 ( .A(n_379), .Y(n_432) );
OAI322xp33_ASAP7_75t_L g389 ( .A1(n_383), .A2(n_390), .A3(n_391), .B1(n_392), .B2(n_393), .C1(n_395), .C2(n_399), .Y(n_389) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_401), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g434 ( .A(n_409), .B(n_435), .Y(n_434) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_420), .B1(n_421), .B2(n_422), .Y(n_417) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g744 ( .A(n_446), .Y(n_744) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_450), .B(n_694), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_629), .Y(n_450) );
NAND4xp25_ASAP7_75t_SL g451 ( .A(n_452), .B(n_574), .C(n_598), .D(n_621), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_516), .B1(n_546), .B2(n_558), .C(n_561), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_489), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_455), .A2(n_475), .B1(n_517), .B2(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_455), .B(n_490), .Y(n_632) );
AND2x2_ASAP7_75t_L g651 ( .A(n_455), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_455), .B(n_635), .Y(n_721) );
AND2x4_ASAP7_75t_L g455 ( .A(n_456), .B(n_475), .Y(n_455) );
AND2x2_ASAP7_75t_L g589 ( .A(n_456), .B(n_490), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_456), .B(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g612 ( .A(n_456), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g617 ( .A(n_456), .B(n_476), .Y(n_617) );
INVx2_ASAP7_75t_L g649 ( .A(n_456), .Y(n_649) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_456), .Y(n_693) );
AND2x2_ASAP7_75t_L g710 ( .A(n_456), .B(n_587), .Y(n_710) );
INVx5_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g628 ( .A(n_457), .B(n_587), .Y(n_628) );
AND2x4_ASAP7_75t_L g642 ( .A(n_457), .B(n_475), .Y(n_642) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_457), .Y(n_646) );
AND2x2_ASAP7_75t_L g666 ( .A(n_457), .B(n_581), .Y(n_666) );
AND2x2_ASAP7_75t_L g716 ( .A(n_457), .B(n_491), .Y(n_716) );
AND2x2_ASAP7_75t_L g726 ( .A(n_457), .B(n_476), .Y(n_726) );
OR2x6_ASAP7_75t_L g457 ( .A(n_458), .B(n_472), .Y(n_457) );
AOI21xp5_ASAP7_75t_SL g458 ( .A1(n_459), .A2(n_463), .B(n_471), .Y(n_458) );
BUFx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx5_ASAP7_75t_L g481 ( .A(n_464), .Y(n_481) );
INVx2_ASAP7_75t_L g470 ( .A(n_468), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_470), .A2(n_497), .B(n_498), .C(n_499), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_470), .A2(n_499), .B(n_523), .C(n_524), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
AND2x2_ASAP7_75t_L g582 ( .A(n_475), .B(n_490), .Y(n_582) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_475), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_475), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g672 ( .A(n_475), .Y(n_672) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g560 ( .A(n_476), .B(n_505), .Y(n_560) );
AND2x2_ASAP7_75t_L g587 ( .A(n_476), .B(n_506), .Y(n_587) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B(n_488), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_SL g479 ( .A1(n_480), .A2(n_481), .B(n_482), .C(n_487), .Y(n_479) );
INVx2_ASAP7_75t_L g495 ( .A(n_481), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_481), .A2(n_487), .B(n_532), .C(n_533), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVx1_ASAP7_75t_L g500 ( .A(n_487), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_489), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_503), .Y(n_489) );
OR2x2_ASAP7_75t_L g613 ( .A(n_490), .B(n_504), .Y(n_613) );
AND2x2_ASAP7_75t_L g650 ( .A(n_490), .B(n_560), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_490), .B(n_581), .Y(n_661) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_490), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_490), .B(n_617), .Y(n_734) );
INVx5_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g559 ( .A(n_491), .Y(n_559) );
AND2x2_ASAP7_75t_L g568 ( .A(n_491), .B(n_504), .Y(n_568) );
AND2x2_ASAP7_75t_L g684 ( .A(n_491), .B(n_579), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_491), .B(n_617), .Y(n_706) );
OR2x6_ASAP7_75t_L g491 ( .A(n_492), .B(n_501), .Y(n_491) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_504), .Y(n_652) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_505), .Y(n_604) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_L g581 ( .A(n_506), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_513), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_517), .B(n_526), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_517), .B(n_594), .Y(n_713) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_518), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g565 ( .A(n_518), .B(n_566), .Y(n_565) );
INVx5_ASAP7_75t_SL g573 ( .A(n_518), .Y(n_573) );
OR2x2_ASAP7_75t_L g596 ( .A(n_518), .B(n_566), .Y(n_596) );
OR2x2_ASAP7_75t_L g606 ( .A(n_518), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g669 ( .A(n_518), .B(n_528), .Y(n_669) );
AND2x2_ASAP7_75t_SL g707 ( .A(n_518), .B(n_527), .Y(n_707) );
NOR4xp25_ASAP7_75t_L g728 ( .A(n_518), .B(n_649), .C(n_729), .D(n_730), .Y(n_728) );
AND2x2_ASAP7_75t_L g738 ( .A(n_518), .B(n_570), .Y(n_738) );
OR2x6_ASAP7_75t_L g518 ( .A(n_519), .B(n_525), .Y(n_518) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g563 ( .A(n_527), .B(n_559), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_527), .B(n_565), .Y(n_732) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_537), .Y(n_527) );
OR2x2_ASAP7_75t_L g572 ( .A(n_528), .B(n_573), .Y(n_572) );
INVx3_ASAP7_75t_L g579 ( .A(n_528), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_528), .B(n_548), .Y(n_591) );
INVxp67_ASAP7_75t_L g594 ( .A(n_528), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_528), .B(n_566), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_528), .B(n_538), .Y(n_660) );
AND2x2_ASAP7_75t_L g675 ( .A(n_528), .B(n_570), .Y(n_675) );
OR2x2_ASAP7_75t_L g704 ( .A(n_528), .B(n_538), .Y(n_704) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B(n_536), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_537), .B(n_609), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_537), .B(n_573), .Y(n_712) );
OR2x2_ASAP7_75t_L g733 ( .A(n_537), .B(n_610), .Y(n_733) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g547 ( .A(n_538), .B(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g570 ( .A(n_538), .B(n_566), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_538), .B(n_548), .Y(n_585) );
AND2x2_ASAP7_75t_L g655 ( .A(n_538), .B(n_579), .Y(n_655) );
AND2x2_ASAP7_75t_L g689 ( .A(n_538), .B(n_573), .Y(n_689) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_539), .B(n_573), .Y(n_592) );
AND2x2_ASAP7_75t_L g620 ( .A(n_539), .B(n_548), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_546), .B(n_628), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_547), .A2(n_635), .B1(n_671), .B2(n_688), .C(n_690), .Y(n_687) );
INVx5_ASAP7_75t_SL g566 ( .A(n_548), .Y(n_566) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_551), .B(n_552), .Y(n_549) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
OAI33xp33_ASAP7_75t_L g586 ( .A1(n_559), .A2(n_587), .A3(n_588), .B1(n_590), .B2(n_593), .B3(n_597), .Y(n_586) );
OR2x2_ASAP7_75t_L g602 ( .A(n_559), .B(n_603), .Y(n_602) );
AOI322xp5_ASAP7_75t_L g711 ( .A1(n_559), .A2(n_628), .A3(n_635), .B1(n_712), .B2(n_713), .C1(n_714), .C2(n_717), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_559), .B(n_587), .Y(n_729) );
A2O1A1Ixp33_ASAP7_75t_SL g735 ( .A1(n_559), .A2(n_587), .B(n_736), .C(n_738), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g574 ( .A1(n_560), .A2(n_575), .B1(n_580), .B2(n_583), .C(n_586), .Y(n_574) );
INVx1_ASAP7_75t_L g667 ( .A(n_560), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_560), .B(n_716), .Y(n_715) );
OAI22xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_564), .B1(n_567), .B2(n_569), .Y(n_561) );
INVx1_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g644 ( .A(n_565), .B(n_579), .Y(n_644) );
AND2x2_ASAP7_75t_L g702 ( .A(n_565), .B(n_703), .Y(n_702) );
OR2x2_ASAP7_75t_L g610 ( .A(n_566), .B(n_573), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_566), .B(n_579), .Y(n_638) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_568), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_568), .B(n_646), .Y(n_700) );
OAI321xp33_ASAP7_75t_L g719 ( .A1(n_568), .A2(n_641), .A3(n_720), .B1(n_721), .B2(n_722), .C(n_723), .Y(n_719) );
INVx1_ASAP7_75t_L g686 ( .A(n_569), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_570), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g625 ( .A(n_570), .B(n_573), .Y(n_625) );
AOI321xp33_ASAP7_75t_L g683 ( .A1(n_570), .A2(n_587), .A3(n_684), .B1(n_685), .B2(n_686), .C(n_687), .Y(n_683) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g600 ( .A(n_572), .B(n_585), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_573), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_573), .B(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_573), .B(n_659), .Y(n_696) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x4_ASAP7_75t_L g619 ( .A(n_577), .B(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g584 ( .A(n_578), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g692 ( .A(n_579), .Y(n_692) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_582), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g615 ( .A(n_587), .Y(n_615) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_589), .B(n_624), .Y(n_673) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
OR2x2_ASAP7_75t_L g637 ( .A(n_592), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_SL g682 ( .A(n_592), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_593), .A2(n_640), .B1(n_643), .B2(n_645), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g737 ( .A(n_596), .B(n_660), .Y(n_737) );
AOI221xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_601), .B1(n_605), .B2(n_611), .C(n_614), .Y(n_598) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx2_ASAP7_75t_L g635 ( .A(n_604), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVx1_ASAP7_75t_SL g681 ( .A(n_607), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_609), .B(n_659), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_609), .A2(n_677), .B(n_679), .Y(n_676) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g722 ( .A(n_610), .B(n_704), .Y(n_722) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_SL g624 ( .A(n_613), .Y(n_624) );
AOI21xp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_616), .B(n_618), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g668 ( .A(n_620), .B(n_669), .Y(n_668) );
INVxp67_ASAP7_75t_L g730 ( .A(n_620), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_625), .B(n_626), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_624), .B(n_642), .Y(n_678) );
INVxp67_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g699 ( .A(n_628), .Y(n_699) );
NAND5xp2_ASAP7_75t_L g629 ( .A(n_630), .B(n_647), .C(n_656), .D(n_676), .E(n_683), .Y(n_629) );
O2A1O1Ixp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_633), .B(n_636), .C(n_639), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g671 ( .A(n_635), .Y(n_671) );
CKINVDCx16_ASAP7_75t_R g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_643), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g685 ( .A(n_645), .Y(n_685) );
OAI21xp5_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_651), .B(n_653), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_648), .A2(n_702), .B1(n_705), .B2(n_707), .C(n_708), .Y(n_701) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
AOI321xp33_ASAP7_75t_L g656 ( .A1(n_649), .A2(n_657), .A3(n_661), .B1(n_662), .B2(n_668), .C(n_670), .Y(n_656) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g727 ( .A(n_661), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_663), .B(n_667), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g679 ( .A(n_664), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
NOR2xp67_ASAP7_75t_SL g691 ( .A(n_665), .B(n_672), .Y(n_691) );
AOI321xp33_ASAP7_75t_SL g723 ( .A1(n_668), .A2(n_724), .A3(n_725), .B1(n_726), .B2(n_727), .C(n_728), .Y(n_723) );
O2A1O1Ixp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .B(n_673), .C(n_674), .Y(n_670) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_681), .B(n_689), .Y(n_718) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND3xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .C(n_693), .Y(n_690) );
NOR3xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_719), .C(n_731), .Y(n_694) );
OAI211xp5_ASAP7_75t_SL g695 ( .A1(n_696), .A2(n_697), .B(n_701), .C(n_711), .Y(n_695) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_699), .B(n_700), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g731 ( .A1(n_700), .A2(n_732), .B1(n_733), .B2(n_734), .C(n_735), .Y(n_731) );
INVx1_ASAP7_75t_L g720 ( .A(n_702), .Y(n_720) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g724 ( .A(n_722), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
CKINVDCx14_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
endmodule