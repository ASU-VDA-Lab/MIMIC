module fake_netlist_5_1626_n_29 (n_8, n_4, n_5, n_7, n_0, n_9, n_2, n_3, n_6, n_1, n_29);

input n_8;
input n_4;
input n_5;
input n_7;
input n_0;
input n_9;
input n_2;
input n_3;
input n_6;
input n_1;

output n_29;

wire n_16;
wire n_12;
wire n_25;
wire n_18;
wire n_27;
wire n_22;
wire n_10;
wire n_24;
wire n_28;
wire n_21;
wire n_11;
wire n_17;
wire n_19;
wire n_15;
wire n_26;
wire n_20;
wire n_14;
wire n_23;
wire n_13;

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_0),
.Y(n_10)
);

NAND3x1_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_8),
.C(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_9),
.A2(n_4),
.B1(n_6),
.B2(n_3),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_2),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_0),
.Y(n_17)
);

OAI21x1_ASAP7_75t_L g18 ( 
.A1(n_12),
.A2(n_2),
.B(n_3),
.Y(n_18)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx11_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

OAI221xp5_ASAP7_75t_L g21 ( 
.A1(n_17),
.A2(n_10),
.B1(n_15),
.B2(n_16),
.C(n_13),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_16),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g23 ( 
.A1(n_21),
.A2(n_17),
.B(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

AOI211xp5_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_18),
.B(n_11),
.C(n_20),
.Y(n_25)
);

AOI211xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_18),
.B(n_16),
.C(n_5),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_18),
.B1(n_27),
.B2(n_24),
.Y(n_29)
);


endmodule