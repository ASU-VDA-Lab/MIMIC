module fake_netlist_5_2025_n_250 (n_54, n_29, n_16, n_43, n_0, n_12, n_9, n_47, n_58, n_67, n_69, n_36, n_25, n_53, n_18, n_27, n_42, n_64, n_22, n_1, n_8, n_45, n_10, n_24, n_28, n_46, n_21, n_44, n_40, n_34, n_62, n_70, n_38, n_71, n_61, n_68, n_72, n_4, n_32, n_35, n_41, n_65, n_56, n_51, n_63, n_73, n_11, n_17, n_19, n_57, n_7, n_37, n_59, n_15, n_26, n_30, n_20, n_5, n_33, n_55, n_14, n_48, n_2, n_31, n_23, n_13, n_50, n_66, n_3, n_49, n_52, n_60, n_6, n_39, n_250);

input n_54;
input n_29;
input n_16;
input n_43;
input n_0;
input n_12;
input n_9;
input n_47;
input n_58;
input n_67;
input n_69;
input n_36;
input n_25;
input n_53;
input n_18;
input n_27;
input n_42;
input n_64;
input n_22;
input n_1;
input n_8;
input n_45;
input n_10;
input n_24;
input n_28;
input n_46;
input n_21;
input n_44;
input n_40;
input n_34;
input n_62;
input n_70;
input n_38;
input n_71;
input n_61;
input n_68;
input n_72;
input n_4;
input n_32;
input n_35;
input n_41;
input n_65;
input n_56;
input n_51;
input n_63;
input n_73;
input n_11;
input n_17;
input n_19;
input n_57;
input n_7;
input n_37;
input n_59;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_55;
input n_14;
input n_48;
input n_2;
input n_31;
input n_23;
input n_13;
input n_50;
input n_66;
input n_3;
input n_49;
input n_52;
input n_60;
input n_6;
input n_39;

output n_250;

wire n_137;
wire n_210;
wire n_168;
wire n_164;
wire n_91;
wire n_208;
wire n_122;
wire n_82;
wire n_194;
wire n_142;
wire n_176;
wire n_214;
wire n_140;
wire n_248;
wire n_124;
wire n_136;
wire n_146;
wire n_86;
wire n_182;
wire n_143;
wire n_83;
wire n_132;
wire n_237;
wire n_90;
wire n_241;
wire n_127;
wire n_75;
wire n_101;
wire n_180;
wire n_184;
wire n_226;
wire n_235;
wire n_78;
wire n_74;
wire n_144;
wire n_207;
wire n_240;
wire n_114;
wire n_96;
wire n_189;
wire n_220;
wire n_165;
wire n_111;
wire n_229;
wire n_108;
wire n_231;
wire n_213;
wire n_129;
wire n_98;
wire n_177;
wire n_155;
wire n_152;
wire n_197;
wire n_107;
wire n_236;
wire n_116;
wire n_195;
wire n_227;
wire n_117;
wire n_249;
wire n_233;
wire n_94;
wire n_203;
wire n_245;
wire n_205;
wire n_123;
wire n_113;
wire n_139;
wire n_105;
wire n_246;
wire n_80;
wire n_179;
wire n_125;
wire n_167;
wire n_128;
wire n_234;
wire n_92;
wire n_149;
wire n_120;
wire n_232;
wire n_135;
wire n_156;
wire n_126;
wire n_225;
wire n_84;
wire n_202;
wire n_130;
wire n_219;
wire n_157;
wire n_79;
wire n_193;
wire n_151;
wire n_131;
wire n_192;
wire n_173;
wire n_244;
wire n_160;
wire n_198;
wire n_223;
wire n_247;
wire n_188;
wire n_190;
wire n_201;
wire n_158;
wire n_224;
wire n_154;
wire n_100;
wire n_138;
wire n_148;
wire n_228;
wire n_109;
wire n_112;
wire n_212;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_185;
wire n_183;
wire n_243;
wire n_239;
wire n_175;
wire n_169;
wire n_133;
wire n_238;
wire n_215;
wire n_196;
wire n_99;
wire n_211;
wire n_218;
wire n_181;
wire n_147;
wire n_178;
wire n_221;
wire n_121;
wire n_242;
wire n_76;
wire n_200;
wire n_87;
wire n_150;
wire n_162;
wire n_170;
wire n_77;
wire n_106;
wire n_161;
wire n_102;
wire n_209;
wire n_222;
wire n_230;
wire n_81;
wire n_118;
wire n_89;
wire n_115;
wire n_93;
wire n_174;
wire n_186;
wire n_199;
wire n_134;
wire n_187;
wire n_104;
wire n_191;
wire n_172;
wire n_103;
wire n_97;
wire n_141;
wire n_166;
wire n_217;
wire n_206;
wire n_171;
wire n_153;
wire n_145;
wire n_204;
wire n_88;
wire n_110;
wire n_216;

INVx2_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVxp67_ASAP7_75t_SL g83 ( 
.A(n_24),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_7),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_11),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_10),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_12),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_15),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_21),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_33),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

CKINVDCx11_ASAP7_75t_R g105 ( 
.A(n_72),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_13),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_36),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_25),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_14),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_42),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_20),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_9),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_105),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_0),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

BUFx8_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_80),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_4),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

AND2x4_ASAP7_75t_L g130 ( 
.A(n_79),
.B(n_74),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_5),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_6),
.Y(n_136)
);

AND3x2_ASAP7_75t_L g137 ( 
.A(n_83),
.B(n_6),
.C(n_8),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_8),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_107),
.Y(n_148)
);

BUFx10_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

OR2x6_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_82),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_134),
.B(n_88),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_R g154 ( 
.A(n_117),
.B(n_113),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

BUFx4f_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_128),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_SL g161 ( 
.A(n_153),
.B(n_119),
.C(n_136),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_123),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_153),
.B1(n_140),
.B2(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_131),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

NOR3xp33_ASAP7_75t_SL g168 ( 
.A(n_145),
.B(n_101),
.C(n_108),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_99),
.B(n_84),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_135),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

AND2x4_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

NAND2xp33_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_114),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_100),
.B1(n_86),
.B2(n_87),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_135),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_149),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

AND2x4_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_85),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_111),
.B1(n_92),
.B2(n_93),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_112),
.B1(n_95),
.B2(n_96),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_156),
.B(n_139),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_149),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_170),
.A2(n_139),
.B(n_159),
.Y(n_193)
);

OR2x6_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_91),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_157),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_127),
.B(n_132),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_181),
.B1(n_178),
.B2(n_102),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

AO31x2_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_116),
.A3(n_115),
.B(n_110),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_190),
.Y(n_204)
);

OAI21x1_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_109),
.B(n_179),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

OAI21x1_ASAP7_75t_L g208 ( 
.A1(n_193),
.A2(n_176),
.B(n_175),
.Y(n_208)
);

OA21x2_ASAP7_75t_L g209 ( 
.A1(n_195),
.A2(n_168),
.B(n_175),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_198),
.B(n_183),
.Y(n_214)
);

OAI22x1_ASAP7_75t_L g215 ( 
.A1(n_204),
.A2(n_196),
.B1(n_192),
.B2(n_189),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_207),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_71),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_209),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_218),
.Y(n_223)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

AND2x4_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

OAI33xp33_ASAP7_75t_L g229 ( 
.A1(n_227),
.A2(n_200),
.A3(n_219),
.B1(n_206),
.B2(n_203),
.B3(n_212),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_225),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_224),
.Y(n_231)
);

OAI33xp33_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_219),
.A3(n_203),
.B1(n_220),
.B2(n_207),
.B3(n_222),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_228),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_226),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_35),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_238),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_239),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_240),
.A2(n_232),
.B1(n_229),
.B2(n_236),
.Y(n_241)
);

NOR4xp25_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_232),
.C(n_229),
.D(n_237),
.Y(n_242)
);

AND3x1_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_231),
.C(n_41),
.Y(n_243)
);

OR4x2_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_45),
.C(n_47),
.D(n_48),
.Y(n_244)
);

OAI21x1_ASAP7_75t_L g245 ( 
.A1(n_244),
.A2(n_50),
.B(n_53),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_245),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_246),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_247),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_248),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_249),
.A2(n_63),
.B1(n_66),
.B2(n_70),
.Y(n_250)
);


endmodule