module fake_jpeg_15137_n_145 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_145);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx8_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_15),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_20),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_43),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_22),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_33),
.B(n_11),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_52),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_27),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_28),
.B1(n_17),
.B2(n_18),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_36),
.B1(n_11),
.B2(n_21),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_18),
.B1(n_17),
.B2(n_15),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_61),
.B1(n_45),
.B2(n_19),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_36),
.B1(n_32),
.B2(n_15),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_58),
.B1(n_53),
.B2(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_12),
.B1(n_21),
.B2(n_19),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_64),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_71),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_65),
.A2(n_48),
.B1(n_42),
.B2(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_65),
.B(n_44),
.C(n_58),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_75),
.B(n_48),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_55),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_74),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_62),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_57),
.B(n_63),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_79),
.B(n_74),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_63),
.B(n_29),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_76),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_83),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_51),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_72),
.B1(n_32),
.B2(n_38),
.Y(n_100)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_87),
.B(n_71),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_88),
.B(n_14),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_90),
.B1(n_95),
.B2(n_40),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_85),
.B1(n_82),
.B2(n_86),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_93),
.Y(n_106)
);

AOI221xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_12),
.B1(n_20),
.B2(n_19),
.C(n_16),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_14),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_82),
.A2(n_80),
.B1(n_79),
.B2(n_88),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_78),
.B(n_16),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_98),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_47),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_25),
.C(n_37),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_50),
.B1(n_40),
.B2(n_16),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_SL g101 ( 
.A1(n_92),
.A2(n_47),
.B(n_50),
.C(n_37),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_107),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_104),
.Y(n_117)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_91),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_97),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_98),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_14),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_111),
.C(n_94),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_110),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_30),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_114),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_113),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_102),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_116),
.B(n_119),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_10),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_0),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_101),
.B1(n_1),
.B2(n_2),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_101),
.B(n_1),
.Y(n_121)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_0),
.B(n_3),
.Y(n_123)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_3),
.B(n_4),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_126),
.B(n_117),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_125),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_5),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_115),
.B1(n_5),
.B2(n_6),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_131),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_135),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_131),
.B(n_127),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_138),
.C(n_133),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_7),
.B(n_8),
.Y(n_138)
);

XNOR2x2_ASAP7_75t_SL g142 ( 
.A(n_139),
.B(n_141),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_132),
.C(n_9),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_25),
.C(n_8),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_143),
.B(n_9),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_142),
.Y(n_145)
);


endmodule