module fake_ariane_321_n_109 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_10, n_109);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_109;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_40;
wire n_106;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_108;
wire n_102;
wire n_22;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVxp67_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVxp33_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVxp67_ASAP7_75t_SL g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

NAND2x1_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_32),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_23),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_29),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_21),
.B(n_30),
.C(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_31),
.Y(n_52)
);

OAI221xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_42),
.C(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_27),
.B1(n_30),
.B2(n_17),
.Y(n_56)
);

AO22x2_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_18),
.B1(n_27),
.B2(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_38),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_56),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_37),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_57),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_49),
.Y(n_66)
);

NAND2x1p5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_55),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_59),
.B1(n_63),
.B2(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

OA21x2_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_58),
.B(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_64),
.B(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_65),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_70),
.B(n_72),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_74),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_71),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

OAI21x1_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_78),
.B(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_88),
.B(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_71),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_83),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_86),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_86),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_95),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_85),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_87),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_100),
.A3(n_63),
.B1(n_96),
.B2(n_66),
.C1(n_68),
.C2(n_85),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_103),
.B1(n_102),
.B2(n_85),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_102),
.B1(n_74),
.B2(n_68),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_74),
.B(n_66),
.Y(n_108)
);

AOI31xp33_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_61),
.A3(n_67),
.B(n_107),
.Y(n_109)
);


endmodule