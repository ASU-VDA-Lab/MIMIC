module real_jpeg_5373_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_1),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_1),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_1),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_1),
.B(n_109),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_2),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_3),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_3),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_3),
.B(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_3),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_3),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_4),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_4),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_4),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_4),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_4),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_4),
.B(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_5),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_5),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_5),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_5),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_5),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_5),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_5),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_5),
.B(n_295),
.Y(n_294)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_7),
.Y(n_105)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_7),
.Y(n_141)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_7),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_7),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_7),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_8),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_8),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_8),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_8),
.B(n_42),
.Y(n_271)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_8),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_8),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_8),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_8),
.B(n_371),
.Y(n_370)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_9),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_9),
.Y(n_157)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_9),
.Y(n_197)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_11),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_11),
.B(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_11),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_11),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_11),
.B(n_367),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_12),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_12),
.Y(n_111)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_12),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_12),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_13),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_13),
.B(n_196),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_13),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_13),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_13),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_13),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_14),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_14),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_14),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_14),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_14),
.B(n_235),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_15),
.Y(n_96)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_15),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g329 ( 
.A(n_15),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_212),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_211),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_173),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_19),
.B(n_173),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_19),
.B(n_215),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_19),
.B(n_215),
.Y(n_417)
);

FAx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_64),
.CI(n_127),
.CON(n_19),
.SN(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_52),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_35),
.B1(n_50),
.B2(n_51),
.Y(n_21)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_22),
.B(n_51),
.C(n_52),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_27),
.C(n_32),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_23),
.A2(n_57),
.B1(n_58),
.B2(n_62),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_23),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_23),
.A2(n_32),
.B1(n_62),
.B2(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_23),
.B(n_54),
.C(n_58),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_23),
.A2(n_62),
.B1(n_278),
.B2(n_279),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

OR2x2_ASAP7_75t_SL g87 ( 
.A(n_24),
.B(n_88),
.Y(n_87)
);

OR2x2_ASAP7_75t_SL g106 ( 
.A(n_24),
.B(n_107),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_24),
.B(n_83),
.Y(n_185)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_27),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_66)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_29),
.Y(n_192)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_30),
.Y(n_369)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_31),
.Y(n_281)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_32),
.B(n_185),
.C(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_32),
.A2(n_69),
.B1(n_184),
.B2(n_185),
.Y(n_352)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g257 ( 
.A(n_34),
.Y(n_257)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_40),
.B2(n_49),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_36),
.A2(n_37),
.B1(n_146),
.B2(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_37),
.B(n_143),
.C(n_146),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_37),
.B(n_41),
.C(n_44),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_39),
.Y(n_274)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_43),
.Y(n_150)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_48),
.Y(n_145)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_48),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_63),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_57),
.A2(n_58),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_57),
.A2(n_58),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_58),
.B(n_270),
.C(n_275),
.Y(n_354)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_62),
.B(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_98),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_65),
.B(n_99),
.C(n_115),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_71),
.C(n_85),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_66),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_71),
.B(n_85),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.C(n_81),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_72),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_76),
.Y(n_289)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_77),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_81),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_78),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_78),
.Y(n_194)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_84),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_90),
.B2(n_97),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_125),
.C(n_126),
.Y(n_124)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_95),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_115),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_110),
.C(n_112),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_101),
.B(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.C(n_108),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_102),
.A2(n_108),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_102),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_102),
.A2(n_243),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_106),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_106),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_108),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_110),
.B(n_112),
.Y(n_172)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_124),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_116)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_120),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_120),
.B(n_122),
.C(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_120),
.A2(n_123),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_124),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_151),
.C(n_171),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_128),
.B(n_218),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.C(n_142),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_129),
.B(n_142),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_131),
.B(n_406),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.C(n_138),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_132),
.B(n_138),
.Y(n_224)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_135),
.B(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_137),
.Y(n_372)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_141),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_143),
.A2(n_385),
.B1(n_386),
.B2(n_388),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_143),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_144),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_145),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_145),
.Y(n_262)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_146),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_151),
.B(n_171),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_162),
.C(n_169),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_152),
.B(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_152),
.A2(n_153),
.B(n_158),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.Y(n_152)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_170),
.Y(n_169)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_161),
.B(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_162),
.B(n_169),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_166),
.Y(n_305)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_167),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_170),
.B(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_170),
.B(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_170),
.B(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_199),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_186),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_183),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_195),
.B2(n_198),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_191),
.Y(n_193)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_210),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_246),
.B(n_417),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.C(n_221),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_219),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_221),
.B(n_411),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_238),
.C(n_244),
.Y(n_221)
);

FAx1_ASAP7_75t_L g402 ( 
.A(n_222),
.B(n_238),
.CI(n_244),
.CON(n_402),
.SN(n_402)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.C(n_231),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_223),
.B(n_394),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_225),
.A2(n_231),
.B1(n_232),
.B2(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_225),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_226),
.B(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_355)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_243),
.B(n_287),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_398),
.B(n_413),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_376),
.B(n_397),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_346),
.B(n_375),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_300),
.B(n_345),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_290),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_252),
.B(n_290),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_276),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_267),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_254),
.B(n_267),
.C(n_276),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.C(n_263),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_255),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_292)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_257),
.Y(n_331)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_263),
.B(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_275),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_272),
.Y(n_275)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_282),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_277),
.B(n_359),
.C(n_360),
.Y(n_358)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_283),
.Y(n_359)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_286),
.Y(n_360)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.C(n_299),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_291),
.B(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_293),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_293),
.A2(n_299),
.B1(n_337),
.B2(n_343),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_297),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_294),
.Y(n_335)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_297),
.Y(n_336)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_299),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_339),
.B(n_344),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_325),
.B(n_338),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_310),
.B(n_324),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_321),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_321),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_316),
.B(n_320),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_316),
.Y(n_320)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_320),
.A2(n_327),
.B1(n_332),
.B2(n_333),
.Y(n_326)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_320),
.Y(n_332)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_334),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_334),
.Y(n_338)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_327),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_328),
.A2(n_330),
.B(n_332),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_335),
.A2(n_336),
.B(n_337),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_340),
.B(n_341),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_347),
.B(n_348),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_356),
.B2(n_357),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_349),
.B(n_358),
.C(n_361),
.Y(n_377)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_353),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_351),
.B(n_354),
.C(n_355),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_364),
.B2(n_374),
.Y(n_361)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_362),
.Y(n_374)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_366),
.B1(n_370),
.B2(n_373),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_373),
.C(n_374),
.Y(n_381)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx5_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_370),
.Y(n_373)
);

INVx5_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_377),
.B(n_378),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_380),
.B1(n_391),
.B2(n_396),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_379),
.B(n_392),
.C(n_393),
.Y(n_407)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_381),
.B(n_384),
.C(n_389),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_383),
.A2(n_384),
.B1(n_389),
.B2(n_390),
.Y(n_382)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_383),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_384),
.Y(n_390)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_386),
.Y(n_388)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_391),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_408),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_401),
.B(n_407),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_401),
.B(n_407),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_402),
.B(n_404),
.C(n_405),
.Y(n_409)
);

BUFx24_ASAP7_75t_SL g419 ( 
.A(n_402),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_408),
.A2(n_415),
.B(n_416),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_409),
.B(n_410),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);


endmodule