module fake_jpeg_20227_n_338 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_15),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_38),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_9),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_44),
.Y(n_60)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_9),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_61),
.Y(n_81)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_28),
.B1(n_32),
.B2(n_38),
.Y(n_75)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_70),
.Y(n_90)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_44),
.B1(n_65),
.B2(n_33),
.Y(n_88)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_26),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_68),
.A2(n_23),
.B1(n_29),
.B2(n_31),
.Y(n_97)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_47),
.Y(n_72)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_72),
.Y(n_117)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_69),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_69),
.Y(n_111)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_75),
.A2(n_51),
.B1(n_67),
.B2(n_63),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_55),
.B1(n_60),
.B2(n_43),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_77),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_78),
.B(n_87),
.Y(n_102)
);

HAxp5_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_61),
.CON(n_80),
.SN(n_80)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_88),
.B1(n_44),
.B2(n_65),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_45),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_95),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_48),
.Y(n_87)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_45),
.Y(n_92)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_31),
.C(n_29),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_23),
.Y(n_107)
);

OAI22x1_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_37),
.B1(n_46),
.B2(n_39),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_126),
.B1(n_53),
.B2(n_52),
.Y(n_134)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_111),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_25),
.Y(n_112)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_83),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_119),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_77),
.A2(n_44),
.B(n_51),
.C(n_67),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_114),
.A2(n_120),
.B(n_73),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_52),
.B1(n_82),
.B2(n_91),
.Y(n_139)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_70),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_66),
.B(n_1),
.Y(n_120)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_125),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_81),
.B(n_49),
.CI(n_51),
.CON(n_125),
.SN(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_79),
.A2(n_71),
.B1(n_63),
.B2(n_53),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_108),
.A2(n_75),
.B1(n_90),
.B2(n_81),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_127),
.A2(n_134),
.B1(n_147),
.B2(n_151),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_97),
.B(n_87),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_142),
.B(n_149),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_84),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_96),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_144),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_139),
.A2(n_145),
.B1(n_104),
.B2(n_116),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_82),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_99),
.A2(n_119),
.B1(n_118),
.B2(n_102),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_114),
.A2(n_52),
.B1(n_85),
.B2(n_79),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_85),
.B(n_69),
.C(n_58),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_100),
.A2(n_103),
.B1(n_117),
.B2(n_107),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_101),
.B(n_46),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_26),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_156),
.A2(n_163),
.B1(n_171),
.B2(n_182),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_123),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_158),
.B(n_138),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_159),
.B(n_165),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_124),
.B(n_110),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_162),
.B(n_164),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_121),
.B(n_98),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_145),
.A2(n_122),
.B1(n_84),
.B2(n_59),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_106),
.B(n_83),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_106),
.B(n_83),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_170),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_46),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_174),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_144),
.B(n_130),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_84),
.B1(n_25),
.B2(n_30),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_151),
.B(n_46),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_0),
.B(n_1),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_176),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_139),
.B(n_143),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_154),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_179),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_132),
.B(n_39),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_26),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_136),
.A2(n_59),
.B1(n_37),
.B2(n_30),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_17),
.B(n_22),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_183),
.A2(n_135),
.B1(n_153),
.B2(n_129),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_SL g234 ( 
.A(n_185),
.B(n_186),
.C(n_193),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_146),
.Y(n_186)
);

BUFx24_ASAP7_75t_SL g187 ( 
.A(n_158),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_201),
.Y(n_217)
);

OAI21xp33_ASAP7_75t_SL g193 ( 
.A1(n_157),
.A2(n_17),
.B(n_22),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_165),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_170),
.C(n_174),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_198),
.C(n_199),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_129),
.C(n_128),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_150),
.C(n_131),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_180),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_138),
.Y(n_202)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_203),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_156),
.A2(n_59),
.B1(n_37),
.B2(n_13),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_204),
.A2(n_175),
.B1(n_169),
.B2(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_209),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_26),
.C(n_34),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_210),
.C(n_168),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_160),
.B(n_27),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_34),
.C(n_21),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_160),
.Y(n_213)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_188),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_220),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_216),
.A2(n_222),
.B1(n_206),
.B2(n_191),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_171),
.Y(n_219)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_219),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_206),
.A2(n_164),
.B1(n_166),
.B2(n_163),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_159),
.Y(n_223)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_179),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_227),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_226),
.B(n_198),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_168),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_183),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_237),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_233),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_167),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_231),
.B(n_236),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_189),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_235),
.B(n_213),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_207),
.B(n_167),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_190),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_239),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_242),
.A2(n_251),
.B1(n_256),
.B2(n_218),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_199),
.C(n_208),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_230),
.C(n_226),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_222),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_214),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_229),
.A2(n_192),
.B1(n_204),
.B2(n_210),
.Y(n_246)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_216),
.A2(n_191),
.B1(n_192),
.B2(n_155),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_191),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_254),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_20),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_232),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_255),
.A2(n_217),
.B1(n_34),
.B2(n_21),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_220),
.A2(n_11),
.B1(n_16),
.B2(n_15),
.Y(n_256)
);

NAND3xp33_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_12),
.C(n_16),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_258),
.B(n_10),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_233),
.A2(n_10),
.B(n_15),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_260),
.A2(n_212),
.B(n_225),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_264),
.C(n_271),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_252),
.B(n_234),
.Y(n_264)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_259),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_269),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_234),
.B(n_224),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_268),
.A2(n_278),
.B(n_256),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_212),
.C(n_218),
.Y(n_271)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

INVx13_ASAP7_75t_L g287 ( 
.A(n_275),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_248),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_238),
.B(n_20),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_244),
.C(n_242),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_L g278 ( 
.A1(n_250),
.A2(n_7),
.B(n_14),
.Y(n_278)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_273),
.B1(n_266),
.B2(n_278),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_274),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_251),
.B(n_253),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

XNOR2x2_ASAP7_75t_SL g289 ( 
.A(n_264),
.B(n_239),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_277),
.Y(n_295)
);

OAI322xp33_ASAP7_75t_L g291 ( 
.A1(n_262),
.A2(n_241),
.A3(n_244),
.B1(n_254),
.B2(n_247),
.C1(n_13),
.C2(n_6),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_7),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_34),
.C(n_21),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_293),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_0),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_263),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_294),
.B(n_295),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_274),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_297),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_286),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_305),
.Y(n_310)
);

AOI211xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_284),
.B(n_279),
.C(n_283),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_303),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_261),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_261),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_14),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_293),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_14),
.B1(n_9),
.B2(n_6),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_287),
.B1(n_2),
.B2(n_3),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_304),
.A2(n_290),
.B1(n_283),
.B2(n_280),
.Y(n_308)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_308),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_314),
.B(n_303),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_282),
.C(n_281),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_27),
.C(n_3),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_299),
.A2(n_282),
.B(n_289),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_0),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_317),
.A2(n_298),
.B1(n_304),
.B2(n_295),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_318),
.A2(n_323),
.B1(n_320),
.B2(n_325),
.Y(n_329)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_319),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_321),
.A2(n_308),
.B1(n_309),
.B2(n_5),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_325),
.C(n_311),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_2),
.C(n_4),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_326),
.A2(n_328),
.B(n_330),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_322),
.B(n_310),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_329),
.A2(n_324),
.B(n_323),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_327),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_331),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_330),
.B(n_311),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_2),
.C(n_4),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_2),
.B(n_5),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_5),
.C(n_293),
.Y(n_338)
);


endmodule