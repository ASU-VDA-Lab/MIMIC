module fake_jpeg_18178_n_284 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_284);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_27),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_38),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_36),
.B1(n_19),
.B2(n_37),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_50),
.A2(n_53),
.B1(n_66),
.B2(n_67),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_36),
.B1(n_19),
.B2(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_54),
.B(n_27),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_27),
.C(n_28),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_56),
.B(n_4),
.C(n_5),
.Y(n_117)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_36),
.B1(n_19),
.B2(n_38),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_29),
.B1(n_23),
.B2(n_24),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_43),
.B1(n_47),
.B2(n_44),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_69),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_35),
.B1(n_33),
.B2(n_31),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_30),
.B1(n_23),
.B2(n_22),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_72),
.B1(n_2),
.B2(n_3),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_29),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_79),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_22),
.B1(n_24),
.B2(n_30),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_35),
.B1(n_25),
.B2(n_33),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_80),
.B1(n_55),
.B2(n_52),
.Y(n_96)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_31),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_45),
.A2(n_25),
.B1(n_34),
.B2(n_18),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_28),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_48),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_39),
.B(n_43),
.C(n_48),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_82),
.A2(n_90),
.B1(n_108),
.B2(n_55),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_83),
.B(n_117),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_92),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_88),
.B(n_105),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_48),
.B1(n_28),
.B2(n_32),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_3),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_3),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_101),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_72),
.Y(n_101)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_65),
.A2(n_34),
.B1(n_18),
.B2(n_28),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_104),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_34),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_21),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_106),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_56),
.A2(n_32),
.B1(n_21),
.B2(n_6),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_111),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_32),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_115),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_69),
.A2(n_21),
.B1(n_5),
.B2(n_6),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_4),
.B1(n_7),
.B2(n_9),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_73),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

AND2x6_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_73),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_130),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_124),
.A2(n_136),
.B1(n_143),
.B2(n_123),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_59),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_131),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_78),
.B1(n_77),
.B2(n_55),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_132),
.B1(n_140),
.B2(n_82),
.Y(n_151)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_74),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_64),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_63),
.B1(n_60),
.B2(n_51),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_97),
.A2(n_51),
.B(n_57),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_137),
.A2(n_91),
.B(n_87),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_94),
.A2(n_4),
.B1(n_7),
.B2(n_9),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_138),
.A2(n_146),
.B1(n_114),
.B2(n_107),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_76),
.B1(n_57),
.B2(n_11),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_83),
.B(n_76),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_95),
.Y(n_147)
);

OAI22x1_ASAP7_75t_SL g143 ( 
.A1(n_106),
.A2(n_76),
.B1(n_10),
.B2(n_11),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_156),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_110),
.B(n_112),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_149),
.A2(n_150),
.B(n_155),
.Y(n_193)
);

XOR2x2_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_106),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_151),
.A2(n_153),
.B1(n_161),
.B2(n_163),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_103),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_154),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_84),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_125),
.B(n_117),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_160),
.B(n_165),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_90),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_164),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_124),
.A2(n_108),
.B1(n_89),
.B2(n_107),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_102),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_118),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_89),
.B1(n_87),
.B2(n_100),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_168),
.A2(n_172),
.B1(n_174),
.B2(n_143),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_119),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_169),
.A2(n_170),
.B(n_176),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_119),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_86),
.Y(n_171)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_134),
.A2(n_100),
.B1(n_86),
.B2(n_93),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_126),
.A2(n_93),
.B1(n_13),
.B2(n_14),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_119),
.Y(n_175)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_126),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_159),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_177),
.B(n_180),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_163),
.B1(n_161),
.B2(n_165),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_166),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_167),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_181),
.A2(n_182),
.B(n_186),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_137),
.B(n_141),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_137),
.Y(n_183)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_129),
.Y(n_186)
);

AO22x1_ASAP7_75t_SL g188 ( 
.A1(n_150),
.A2(n_144),
.B1(n_121),
.B2(n_141),
.Y(n_188)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_148),
.A2(n_122),
.B(n_145),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_194),
.B(n_175),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_158),
.A2(n_122),
.B(n_145),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_149),
.A2(n_144),
.B(n_121),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_196),
.A2(n_174),
.B(n_152),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_183),
.A2(n_156),
.B1(n_162),
.B2(n_147),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_205),
.B1(n_207),
.B2(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_206),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_183),
.A2(n_171),
.B1(n_151),
.B2(n_172),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_208),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_214),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_152),
.C(n_169),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_182),
.C(n_178),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_121),
.B1(n_144),
.B2(n_135),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_178),
.B(n_180),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_191),
.B(n_170),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_216),
.B(n_221),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_135),
.B1(n_157),
.B2(n_175),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_220),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_186),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_99),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_196),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_199),
.A2(n_109),
.B1(n_127),
.B2(n_116),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_224),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_219),
.B(n_203),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_228),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_193),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_200),
.C(n_192),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_235),
.C(n_213),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_207),
.B(n_192),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_233),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_209),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_197),
.C(n_195),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_243),
.C(n_244),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_226),
.A2(n_205),
.B1(n_208),
.B2(n_215),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

OAI31xp33_ASAP7_75t_L g241 ( 
.A1(n_238),
.A2(n_210),
.A3(n_188),
.B(n_202),
.Y(n_241)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_179),
.B1(n_186),
.B2(n_210),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_250),
.B1(n_251),
.B2(n_232),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_230),
.C(n_224),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_202),
.C(n_222),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_245),
.A2(n_225),
.B(n_236),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_206),
.C(n_195),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_190),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_237),
.B(n_185),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_177),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_256),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_227),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_261),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_249),
.A2(n_233),
.B(n_231),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_173),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_244),
.A2(n_220),
.B1(n_181),
.B2(n_188),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_259),
.A2(n_260),
.B1(n_247),
.B2(n_248),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_246),
.A2(n_248),
.B1(n_239),
.B2(n_243),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_263),
.B(n_264),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_201),
.C(n_187),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_SL g266 ( 
.A(n_259),
.B(n_187),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_266),
.A2(n_268),
.B(n_256),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_201),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_254),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_255),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_261),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_273),
.Y(n_277)
);

AOI21x1_ASAP7_75t_L g275 ( 
.A1(n_269),
.A2(n_262),
.B(n_258),
.Y(n_275)
);

AOI322xp5_ASAP7_75t_L g279 ( 
.A1(n_275),
.A2(n_276),
.A3(n_173),
.B1(n_116),
.B2(n_99),
.C1(n_16),
.C2(n_12),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_270),
.A2(n_253),
.B1(n_264),
.B2(n_257),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_275),
.Y(n_278)
);

AO221x1_ASAP7_75t_L g281 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_173),
.C(n_15),
.Y(n_281)
);

AOI322xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_173),
.A3(n_99),
.B1(n_116),
.B2(n_17),
.C1(n_15),
.C2(n_16),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_13),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_17),
.B1(n_99),
.B2(n_274),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_17),
.Y(n_284)
);


endmodule