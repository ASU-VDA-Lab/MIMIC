module fake_jpeg_16591_n_55 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_55);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_55;

wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_36),
.B1(n_6),
.B2(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

CKINVDCx10_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_34),
.Y(n_39)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_26),
.B1(n_0),
.B2(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_5),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_37),
.Y(n_42)
);

OA21x2_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_15),
.B(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_17),
.Y(n_47)
);

OAI32xp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_45),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_47),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_50),
.B(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_19),
.Y(n_53)
);

MAJx2_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_20),
.C(n_22),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_42),
.Y(n_55)
);


endmodule