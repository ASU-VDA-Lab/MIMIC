module real_jpeg_15930_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_0),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_1),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_1),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_1),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_1),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_1),
.B(n_175),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_2),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_2),
.Y(n_164)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_3),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_3),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_3),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_4),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_4),
.B(n_72),
.Y(n_142)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_5),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_6),
.Y(n_128)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_6),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_7),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_7),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_7),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_7),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_7),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_7),
.B(n_127),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_7),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_8),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_8),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_8),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_8),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_8),
.B(n_197),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_8),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_9),
.Y(n_110)
);

AOI22x1_ASAP7_75t_SL g113 ( 
.A1(n_9),
.A2(n_11),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_10),
.Y(n_94)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_10),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_11),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_11),
.B(n_58),
.Y(n_57)
);

AOI31xp33_ASAP7_75t_L g105 ( 
.A1(n_11),
.A2(n_106),
.A3(n_109),
.B(n_113),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_11),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_11),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_11),
.B(n_85),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_12),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_12),
.B(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

BUFx4f_ASAP7_75t_L g83 ( 
.A(n_13),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_13),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_14),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_153),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_151),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_101),
.Y(n_17)
);

NOR2xp67_ASAP7_75t_L g152 ( 
.A(n_18),
.B(n_101),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_66),
.C(n_87),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_19),
.A2(n_20),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_21),
.B(n_149),
.C(n_150),
.Y(n_148)
);

XOR2x2_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_22),
.B(n_29),
.C(n_34),
.Y(n_147)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_29),
.A2(n_37),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_29),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_51),
.Y(n_38)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_39),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_40),
.B(n_45),
.Y(n_146)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_51),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.C(n_61),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_52),
.A2(n_61),
.B1(n_62),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_52),
.Y(n_184)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

XOR2x2_ASAP7_75t_L g182 ( 
.A(n_57),
.B(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_66),
.A2(n_88),
.B1(n_89),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_66),
.Y(n_233)
);

MAJx2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_73),
.C(n_78),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_67),
.B(n_73),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_71),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_71),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_71),
.A2(n_202),
.B1(n_203),
.B2(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_72),
.Y(n_173)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_78),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_84),
.Y(n_78)
);

AO22x1_ASAP7_75t_SL g177 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_84),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_86),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_95),
.C(n_99),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_91)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_130),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_118),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx2_ASAP7_75t_SL g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_125),
.B1(n_126),
.B2(n_129),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_125),
.B(n_160),
.C(n_165),
.Y(n_181)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2x2_ASAP7_75t_SL g158 ( 
.A(n_126),
.B(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_148),
.Y(n_130)
);

XNOR2x1_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_145),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_138),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_142),
.Y(n_143)
);

XNOR2x1_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AOI21x1_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_229),
.B(n_235),
.Y(n_154)
);

OAI21x1_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_187),
.B(n_228),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_179),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_157),
.B(n_179),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_169),
.C(n_177),
.Y(n_157)
);

XOR2x1_ASAP7_75t_L g222 ( 
.A(n_158),
.B(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_165),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_169),
.A2(n_170),
.B1(n_177),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_171),
.B(n_174),
.Y(n_192)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_185),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_181),
.B(n_182),
.C(n_185),
.Y(n_234)
);

AOI21x1_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_221),
.B(n_227),
.Y(n_187)
);

OAI21x1_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_204),
.B(n_220),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_201),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_201),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_195),
.C(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_203),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_212),
.B(n_219),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_210),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_209),
.B(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

NOR2xp67_ASAP7_75t_SL g227 ( 
.A(n_222),
.B(n_225),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_234),
.Y(n_229)
);

NOR2xp67_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_234),
.Y(n_235)
);

INVxp33_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);


endmodule