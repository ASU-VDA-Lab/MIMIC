module real_aes_14803_n_7 (n_4, n_0, n_3, n_5, n_2, n_6, n_1, n_7);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_6;
input n_1;
output n_7;
wire n_17;
wire n_13;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_9;
wire n_20;
wire n_18;
wire n_21;
wire n_8;
wire n_10;
BUFx10_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
BUFx6f_ASAP7_75t_SL g15 ( .A(n_1), .Y(n_15) );
OAI22xp33_ASAP7_75t_SL g13 ( .A1(n_2), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_13) );
INVx1_ASAP7_75t_L g16 ( .A(n_2), .Y(n_16) );
INVx1_ASAP7_75t_L g21 ( .A(n_3), .Y(n_21) );
INVx1_ASAP7_75t_L g10 ( .A(n_4), .Y(n_10) );
AOI221xp5_ASAP7_75t_L g7 ( .A1(n_5), .A2(n_8), .B1(n_12), .B2(n_13), .C(n_17), .Y(n_7) );
AND2x4_ASAP7_75t_L g20 ( .A(n_6), .B(n_21), .Y(n_20) );
INVx2_ASAP7_75t_L g12 ( .A(n_8), .Y(n_12) );
AND2x2_ASAP7_75t_L g8 ( .A(n_9), .B(n_11), .Y(n_8) );
BUFx2_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
CKINVDCx16_ASAP7_75t_R g14 ( .A(n_15), .Y(n_14) );
INVx1_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
endmodule