module fake_netlist_5_183_n_107 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_107);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_107;

wire n_91;
wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_78;
wire n_65;
wire n_74;
wire n_57;
wire n_96;
wire n_37;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_94;
wire n_38;
wire n_105;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_85;
wire n_95;
wire n_59;
wire n_26;
wire n_55;
wire n_99;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx11_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVxp67_ASAP7_75t_SL g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_48),
.Y(n_53)
);

AO22x2_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_32),
.B1(n_34),
.B2(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_24),
.Y(n_55)
);

OAI221xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_24),
.B1(n_33),
.B2(n_23),
.C(n_21),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_41),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_43),
.B1(n_42),
.B2(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_36),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

NOR2xp67_ASAP7_75t_SL g65 ( 
.A(n_60),
.B(n_31),
.Y(n_65)
);

OAI21x1_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_52),
.B(n_51),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_49),
.B(n_38),
.C(n_54),
.Y(n_67)
);

O2A1O1Ixp5_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_38),
.B(n_54),
.C(n_31),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_58),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_37),
.B1(n_39),
.B2(n_31),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_69),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_71),
.A2(n_37),
.B1(n_69),
.B2(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

AO31x2_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_66),
.A3(n_67),
.B(n_68),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_70),
.Y(n_78)
);

NAND4xp25_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_72),
.C(n_68),
.D(n_74),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_73),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_77),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_11),
.Y(n_85)
);

OR2x6_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_61),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_0),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_19),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_85),
.C(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

AOI321xp33_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_83),
.A3(n_5),
.B1(n_6),
.B2(n_4),
.C(n_13),
.Y(n_97)
);

AOI31xp33_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_83),
.A3(n_6),
.B(n_86),
.Y(n_98)
);

AOI221xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_65),
.B1(n_83),
.B2(n_50),
.C(n_86),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

BUFx4f_ASAP7_75t_SL g102 ( 
.A(n_101),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_102),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_100),
.B1(n_97),
.B2(n_94),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_96),
.B1(n_86),
.B2(n_65),
.Y(n_107)
);


endmodule