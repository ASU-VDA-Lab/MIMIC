module fake_jpeg_17670_n_242 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_27),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_8),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_27),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_47),
.Y(n_79)
);

CKINVDCx12_ASAP7_75t_R g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_52),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_34),
.Y(n_47)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_34),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_64),
.Y(n_80)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_19),
.B1(n_28),
.B2(n_29),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_54),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_29),
.B1(n_22),
.B2(n_31),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_58),
.B1(n_20),
.B2(n_30),
.Y(n_84)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_29),
.B1(n_22),
.B2(n_31),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_63),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_21),
.B1(n_23),
.B2(n_30),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_32),
.B1(n_20),
.B2(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_32),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_47),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_89),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_37),
.C(n_41),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_76),
.Y(n_117)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_74),
.Y(n_108)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_64),
.B(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_73),
.B(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_77),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_41),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_63),
.B(n_36),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_35),
.B1(n_43),
.B2(n_42),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_92),
.B1(n_52),
.B2(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_20),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_24),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_84),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_128)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_23),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_94),
.Y(n_118)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_1),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_44),
.C(n_37),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_90),
.B(n_100),
.Y(n_124)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_60),
.B(n_21),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_93),
.B(n_95),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_44),
.B(n_30),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_46),
.B(n_17),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_98),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_26),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_58),
.A2(n_26),
.B(n_24),
.C(n_18),
.Y(n_101)
);

A2O1A1O1Ixp25_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_18),
.B(n_17),
.C(n_3),
.D(n_4),
.Y(n_113)
);

NAND2xp33_ASAP7_75t_SL g102 ( 
.A(n_49),
.B(n_42),
.Y(n_102)
);

NOR2xp67_ASAP7_75t_SL g110 ( 
.A(n_102),
.B(n_103),
.Y(n_110)
);

NAND2x1p5_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_25),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_106),
.B1(n_84),
.B2(n_94),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_67),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_107),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_52),
.B1(n_26),
.B2(n_24),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_109),
.B(n_122),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_18),
.B1(n_17),
.B2(n_3),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_131),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_125),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_68),
.B(n_1),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_2),
.Y(n_127)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_89),
.B1(n_80),
.B2(n_101),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_5),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_79),
.B(n_5),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_90),
.C(n_69),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_143),
.C(n_111),
.Y(n_174)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_103),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_134),
.A2(n_126),
.B(n_11),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_83),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_147),
.B(n_126),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_142),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_124),
.A2(n_80),
.B(n_85),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_139),
.A2(n_150),
.B(n_155),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_141),
.B(n_145),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_115),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_76),
.C(n_79),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_80),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_115),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_151),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_89),
.B(n_102),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_118),
.A2(n_91),
.B(n_72),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_91),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_152),
.A2(n_157),
.B1(n_131),
.B2(n_127),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_154),
.Y(n_177)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

AND2x6_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_82),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_106),
.A2(n_118),
.B1(n_129),
.B2(n_109),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_98),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_105),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_166),
.Y(n_184)
);

AOI221xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_145),
.B1(n_141),
.B2(n_144),
.C(n_156),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_114),
.Y(n_161)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_122),
.C(n_108),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_174),
.C(n_161),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_155),
.A2(n_92),
.B1(n_130),
.B2(n_125),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_114),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_116),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_168),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_116),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_119),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_170),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_119),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_72),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_178),
.B(n_180),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_148),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_153),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_182),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_183),
.A2(n_175),
.B(n_167),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_174),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_187),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_134),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_192),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_144),
.C(n_156),
.Y(n_192)
);

AO221x1_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_153),
.B1(n_138),
.B2(n_142),
.C(n_146),
.Y(n_193)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_171),
.A2(n_149),
.B(n_135),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_194),
.A2(n_164),
.B(n_177),
.Y(n_213)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_150),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_133),
.C(n_140),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_179),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_195),
.A2(n_172),
.B1(n_171),
.B2(n_165),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_203),
.A2(n_209),
.B1(n_210),
.B2(n_214),
.Y(n_224)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_186),
.A2(n_172),
.B1(n_182),
.B2(n_178),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_168),
.B1(n_164),
.B2(n_176),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_SL g211 ( 
.A1(n_200),
.A2(n_160),
.A3(n_175),
.B1(n_170),
.B2(n_167),
.C1(n_159),
.C2(n_163),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_211),
.B(n_212),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_188),
.B(n_191),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_194),
.A2(n_186),
.B1(n_189),
.B2(n_191),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_218),
.Y(n_226)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_220),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_190),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_185),
.C(n_204),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_221),
.B(n_201),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_206),
.A2(n_200),
.B1(n_173),
.B2(n_179),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_202),
.A2(n_184),
.B1(n_192),
.B2(n_179),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_228),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_203),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_223),
.A2(n_213),
.B(n_205),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_SL g230 ( 
.A1(n_229),
.A2(n_224),
.B(n_217),
.C(n_219),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_230),
.A2(n_233),
.B(n_226),
.Y(n_234)
);

AOI322xp5_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_215),
.A3(n_224),
.B1(n_218),
.B2(n_222),
.C1(n_221),
.C2(n_11),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_226),
.A2(n_227),
.B(n_12),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_234),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_13),
.B(n_14),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_236),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_230),
.A2(n_14),
.B(n_15),
.Y(n_236)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_232),
.C(n_231),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_240),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_237),
.A2(n_15),
.B(n_16),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_16),
.Y(n_242)
);


endmodule