module fake_ibex_429_n_188 (n_49, n_7, n_20, n_40, n_17, n_25, n_36, n_41, n_48, n_43, n_18, n_3, n_22, n_28, n_32, n_39, n_53, n_4, n_33, n_54, n_5, n_11, n_30, n_6, n_50, n_29, n_13, n_2, n_8, n_26, n_35, n_14, n_0, n_9, n_34, n_12, n_38, n_42, n_15, n_37, n_24, n_52, n_47, n_31, n_44, n_10, n_23, n_21, n_51, n_27, n_46, n_45, n_19, n_16, n_1, n_188);

input n_49;
input n_7;
input n_20;
input n_40;
input n_17;
input n_25;
input n_36;
input n_41;
input n_48;
input n_43;
input n_18;
input n_3;
input n_22;
input n_28;
input n_32;
input n_39;
input n_53;
input n_4;
input n_33;
input n_54;
input n_5;
input n_11;
input n_30;
input n_6;
input n_50;
input n_29;
input n_13;
input n_2;
input n_8;
input n_26;
input n_35;
input n_14;
input n_0;
input n_9;
input n_34;
input n_12;
input n_38;
input n_42;
input n_15;
input n_37;
input n_24;
input n_52;
input n_47;
input n_31;
input n_44;
input n_10;
input n_23;
input n_21;
input n_51;
input n_27;
input n_46;
input n_45;
input n_19;
input n_16;
input n_1;

output n_188;

wire n_151;
wire n_147;
wire n_85;
wire n_167;
wire n_128;
wire n_84;
wire n_64;
wire n_73;
wire n_152;
wire n_171;
wire n_145;
wire n_65;
wire n_103;
wire n_95;
wire n_139;
wire n_55;
wire n_130;
wire n_63;
wire n_98;
wire n_129;
wire n_161;
wire n_143;
wire n_106;
wire n_177;
wire n_148;
wire n_76;
wire n_118;
wire n_183;
wire n_67;
wire n_164;
wire n_124;
wire n_110;
wire n_169;
wire n_108;
wire n_82;
wire n_165;
wire n_78;
wire n_60;
wire n_86;
wire n_70;
wire n_87;
wire n_109;
wire n_69;
wire n_75;
wire n_121;
wire n_127;
wire n_175;
wire n_137;
wire n_57;
wire n_59;
wire n_125;
wire n_178;
wire n_62;
wire n_71;
wire n_153;
wire n_173;
wire n_120;
wire n_93;
wire n_168;
wire n_155;
wire n_162;
wire n_180;
wire n_122;
wire n_116;
wire n_61;
wire n_94;
wire n_134;
wire n_77;
wire n_112;
wire n_150;
wire n_88;
wire n_133;
wire n_142;
wire n_80;
wire n_172;
wire n_66;
wire n_90;
wire n_74;
wire n_176;
wire n_58;
wire n_140;
wire n_136;
wire n_119;
wire n_100;
wire n_179;
wire n_72;
wire n_166;
wire n_163;
wire n_114;
wire n_97;
wire n_102;
wire n_181;
wire n_131;
wire n_123;
wire n_99;
wire n_135;
wire n_105;
wire n_156;
wire n_126;
wire n_187;
wire n_154;
wire n_182;
wire n_111;
wire n_104;
wire n_141;
wire n_89;
wire n_83;
wire n_107;
wire n_115;
wire n_149;
wire n_186;
wire n_92;
wire n_144;
wire n_170;
wire n_101;
wire n_113;
wire n_138;
wire n_96;
wire n_185;
wire n_68;
wire n_117;
wire n_79;
wire n_81;
wire n_159;
wire n_158;
wire n_132;
wire n_174;
wire n_157;
wire n_160;
wire n_184;
wire n_56;
wire n_146;
wire n_91;

BUFx10_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_32),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_4),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

BUFx2_ASAP7_75t_SL g63 ( 
.A(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_11),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_0),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

OA21x2_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_57),
.B(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_59),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_60),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_80),
.B(n_68),
.Y(n_87)
);

OR2x6_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_63),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_67),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_92),
.Y(n_97)
);

AND2x4_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_87),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_65),
.B(n_64),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_1),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

BUFx4f_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

OR2x6_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_2),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

BUFx4f_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_5),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

NAND2x1p5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_10),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

AO32x2_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_17),
.A3(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_125)
);

OAI21x1_ASAP7_75t_L g126 ( 
.A1(n_119),
.A2(n_121),
.B(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_21),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

BUFx8_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_116),
.B1(n_117),
.B2(n_113),
.Y(n_132)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_130),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

AND2x4_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_132),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_138),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_135),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_143),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_136),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_145),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_146),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_149),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_150),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

AND2x4_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_147),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_151),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_154),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_155),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_156),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_23),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_159),
.Y(n_162)
);

NOR2x1_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_25),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_26),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_27),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_164),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_28),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_29),
.B(n_30),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_33),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

NAND3x1_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_34),
.C(n_35),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_178),
.A2(n_175),
.B1(n_43),
.B2(n_41),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_179),
.A2(n_42),
.B(n_43),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_44),
.Y(n_182)
);

AO21x1_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_44),
.B(n_45),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_181),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_184),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_183),
.Y(n_186)
);

OAI221xp5_ASAP7_75t_R g187 ( 
.A1(n_185),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.C(n_49),
.Y(n_187)
);

AOI211xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_186),
.B(n_50),
.C(n_48),
.Y(n_188)
);


endmodule