module fake_netlist_6_4093_n_1936 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1936);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1936;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_84),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_194),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_31),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_128),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_154),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_180),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_171),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_132),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_42),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_34),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_130),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_105),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_7),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_56),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_55),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_15),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_64),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_13),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_145),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_131),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_50),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_129),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_159),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_70),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_18),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_134),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_55),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_53),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_48),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_186),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_46),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_12),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_124),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_16),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_177),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_35),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_133),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_69),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_118),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_23),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_15),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_100),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_101),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_57),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_74),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_64),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_81),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_96),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_71),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_80),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_99),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_49),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_172),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_85),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_188),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_183),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_91),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_167),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_76),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_53),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_83),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_150),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_52),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_113),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_144),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_135),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_2),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_39),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_191),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_26),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_59),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_95),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_87),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_37),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_89),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_157),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_161),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_143),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_68),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_123),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_176),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_90),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_11),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_13),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_148),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_119),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_187),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_149),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_9),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_178),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_137),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_33),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_16),
.Y(n_291)
);

BUFx8_ASAP7_75t_SL g292 ( 
.A(n_86),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_52),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_28),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_136),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_9),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_170),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_26),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_110),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_184),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_93),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_37),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_50),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_46),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_139),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_97),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_82),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_61),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_8),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_17),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_147),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_35),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_1),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_56),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_182),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_107),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_98),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_5),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_104),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_65),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_33),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_75),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_0),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_79),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_3),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_51),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_121),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_48),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_195),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_28),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_108),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_31),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_22),
.Y(n_333)
);

BUFx10_ASAP7_75t_L g334 ( 
.A(n_32),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_36),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_18),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_179),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_103),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_102),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_122),
.Y(n_340)
);

BUFx5_ASAP7_75t_L g341 ( 
.A(n_40),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_5),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_22),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_12),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_189),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_54),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_45),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_10),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_169),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_163),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_44),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_2),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_120),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_138),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_1),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_67),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_117),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_49),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_146),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_4),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_3),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_11),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_126),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_141),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_192),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_162),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_114),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_60),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_57),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_25),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_142),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_175),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_156),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_62),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_116),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_8),
.Y(n_376)
);

BUFx10_ASAP7_75t_L g377 ( 
.A(n_109),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_62),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_6),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_21),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_168),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_173),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_165),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_65),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_61),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_92),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_127),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_44),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_51),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_10),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_166),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_63),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_25),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_153),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_341),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_210),
.B(n_0),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_202),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_206),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_228),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_216),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_341),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_228),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_341),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_266),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_341),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_235),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_341),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_263),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_258),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_281),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_246),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_292),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_372),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_271),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_341),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_287),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_290),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_341),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_271),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_336),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_336),
.Y(n_422)
);

INVxp33_ASAP7_75t_SL g423 ( 
.A(n_205),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_307),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_211),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_211),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_291),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_248),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_249),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_294),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_302),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_282),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_198),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g434 ( 
.A(n_282),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_293),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_293),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_342),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_251),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_299),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_208),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_342),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_208),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_255),
.B(n_4),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_303),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_351),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_304),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_336),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_312),
.Y(n_448)
);

BUFx2_ASAP7_75t_SL g449 ( 
.A(n_255),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_256),
.B(n_6),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_351),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_320),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_252),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_358),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_321),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_299),
.Y(n_456)
);

NOR2xp67_ASAP7_75t_L g457 ( 
.A(n_241),
.B(n_7),
.Y(n_457)
);

INVxp33_ASAP7_75t_SL g458 ( 
.A(n_205),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_323),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_259),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_262),
.Y(n_461)
);

BUFx10_ASAP7_75t_L g462 ( 
.A(n_336),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_358),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_336),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_204),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_325),
.Y(n_466)
);

NOR2xp67_ASAP7_75t_L g467 ( 
.A(n_241),
.B(n_14),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_209),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_213),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_215),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_328),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_256),
.B(n_14),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_223),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_264),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_330),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_270),
.Y(n_476)
);

INVxp33_ASAP7_75t_L g477 ( 
.A(n_229),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_234),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_242),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_274),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_214),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_261),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_275),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_241),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_214),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_218),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_244),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_269),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_218),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_272),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_298),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_261),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_225),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_225),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_391),
.B(n_17),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_408),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_408),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_421),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_421),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_447),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_413),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_422),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_422),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_428),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_447),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_401),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_464),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_397),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_484),
.B(n_391),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_R g510 ( 
.A(n_424),
.B(n_429),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_402),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_438),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_399),
.B(n_265),
.Y(n_513)
);

CKINVDCx8_ASAP7_75t_R g514 ( 
.A(n_412),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_453),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_398),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_433),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_434),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_395),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_395),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_419),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_460),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_419),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_461),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_403),
.B(n_420),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_404),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_439),
.B(n_220),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_456),
.B(n_220),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_457),
.B(n_203),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_406),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_416),
.Y(n_531)
);

NOR2xp67_ASAP7_75t_L g532 ( 
.A(n_434),
.B(n_207),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_410),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_410),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_474),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_482),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_495),
.B(n_196),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_405),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_476),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_480),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_415),
.B(n_425),
.Y(n_541)
);

BUFx8_ASAP7_75t_L g542 ( 
.A(n_415),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_400),
.Y(n_543)
);

NAND2x1p5_ASAP7_75t_L g544 ( 
.A(n_467),
.B(n_237),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_411),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_482),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_492),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_462),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_483),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_492),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_411),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_407),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_405),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_462),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_449),
.B(n_267),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_462),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_417),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_417),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_465),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_409),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_468),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_469),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_414),
.Y(n_563)
);

OA21x2_ASAP7_75t_L g564 ( 
.A1(n_443),
.A2(n_219),
.B(n_212),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_470),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_473),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_478),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_418),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_479),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_449),
.B(n_224),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_418),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_427),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_487),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_488),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_490),
.Y(n_575)
);

BUFx4f_ASAP7_75t_L g576 ( 
.A(n_564),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_513),
.B(n_525),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_519),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_565),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_520),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_571),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_544),
.B(n_364),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_517),
.B(n_481),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_496),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_520),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_518),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_537),
.B(n_481),
.Y(n_587)
);

INVx4_ASAP7_75t_SL g588 ( 
.A(n_521),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_537),
.B(n_423),
.Y(n_589)
);

INVx4_ASAP7_75t_SL g590 ( 
.A(n_521),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_496),
.Y(n_591)
);

INVx6_ASAP7_75t_L g592 ( 
.A(n_542),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_554),
.B(n_450),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_523),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_496),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_497),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_513),
.B(n_491),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_525),
.B(n_509),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_497),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_497),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_509),
.B(n_426),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_554),
.B(n_472),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_556),
.B(n_458),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_533),
.A2(n_396),
.B1(n_430),
.B2(n_427),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_564),
.A2(n_296),
.B1(n_318),
.B2(n_265),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_541),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_544),
.B(n_364),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_556),
.B(n_430),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_541),
.B(n_432),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_554),
.B(n_431),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_565),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_509),
.B(n_431),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_523),
.Y(n_613)
);

INVx6_ASAP7_75t_L g614 ( 
.A(n_542),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_500),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_509),
.B(n_435),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_564),
.A2(n_529),
.B1(n_528),
.B2(n_527),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_565),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_555),
.B(n_444),
.Y(n_619)
);

INVxp67_ASAP7_75t_SL g620 ( 
.A(n_530),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_536),
.B(n_436),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_534),
.B(n_444),
.Y(n_622)
);

AO22x2_ASAP7_75t_L g623 ( 
.A1(n_529),
.A2(n_318),
.B1(n_390),
.B2(n_296),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_564),
.A2(n_390),
.B1(n_355),
.B2(n_308),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_557),
.B(n_446),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_530),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_529),
.B(n_437),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_559),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_565),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_529),
.B(n_446),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_544),
.B(n_364),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_500),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_559),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_567),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_548),
.B(n_448),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_570),
.A2(n_494),
.B1(n_493),
.B2(n_489),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_565),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_567),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_500),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_574),
.Y(n_640)
);

INVx5_ASAP7_75t_L g641 ( 
.A(n_574),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_558),
.B(n_485),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_505),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_536),
.B(n_441),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_548),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_569),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_548),
.B(n_448),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_505),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_505),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_569),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_542),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_551),
.B(n_452),
.Y(n_652)
);

BUFx6f_ASAP7_75t_SL g653 ( 
.A(n_573),
.Y(n_653)
);

BUFx4f_ASAP7_75t_L g654 ( 
.A(n_574),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_573),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_506),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_542),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_506),
.B(n_452),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_506),
.Y(n_659)
);

INVx6_ASAP7_75t_L g660 ( 
.A(n_574),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_546),
.B(n_445),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_511),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_532),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_575),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_568),
.B(n_455),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_572),
.B(n_455),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_511),
.B(n_459),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_575),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_511),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_526),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_526),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_546),
.B(n_547),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_526),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_574),
.B(n_364),
.Y(n_674)
);

AND2x2_ASAP7_75t_SL g675 ( 
.A(n_558),
.B(n_364),
.Y(n_675)
);

INVx5_ASAP7_75t_L g676 ( 
.A(n_574),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_531),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_538),
.B(n_485),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_531),
.B(n_459),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_531),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_498),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_498),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_561),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_499),
.B(n_466),
.Y(n_684)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_561),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_507),
.Y(n_686)
);

AND2x2_ASAP7_75t_SL g687 ( 
.A(n_545),
.B(n_236),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_507),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_561),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_532),
.B(n_466),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_499),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_562),
.B(n_471),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_502),
.B(n_471),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_502),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_503),
.B(n_562),
.Y(n_695)
);

AND3x2_ASAP7_75t_L g696 ( 
.A(n_538),
.B(n_442),
.C(n_440),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_510),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_566),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_503),
.B(n_475),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_562),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_566),
.B(n_475),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_566),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_547),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_553),
.B(n_243),
.Y(n_704)
);

INVx4_ASAP7_75t_L g705 ( 
.A(n_550),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_553),
.B(n_247),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_550),
.B(n_295),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_514),
.B(n_253),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_504),
.B(n_383),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_514),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_512),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_515),
.B(n_277),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_522),
.B(n_486),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_524),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_535),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_539),
.B(n_254),
.Y(n_716)
);

INVx4_ASAP7_75t_L g717 ( 
.A(n_540),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_549),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_501),
.B(n_486),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_508),
.Y(n_720)
);

XOR2xp5_ASAP7_75t_L g721 ( 
.A(n_516),
.B(n_489),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_563),
.B(n_278),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_543),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_552),
.B(n_493),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_560),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_517),
.B(n_494),
.Y(n_726)
);

BUFx4_ASAP7_75t_L g727 ( 
.A(n_711),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_598),
.B(n_257),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_672),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_672),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_598),
.B(n_260),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_606),
.B(n_451),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_589),
.A2(n_687),
.B1(n_675),
.B2(n_577),
.Y(n_733)
);

NOR2x1_ASAP7_75t_L g734 ( 
.A(n_587),
.B(n_722),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_675),
.B(n_276),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_577),
.B(n_280),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_681),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_620),
.B(n_593),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_681),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_609),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_586),
.B(n_477),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_628),
.Y(n_742)
);

BUFx4f_ASAP7_75t_L g743 ( 
.A(n_614),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_602),
.B(n_283),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_705),
.B(n_288),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_687),
.B(n_289),
.Y(n_746)
);

INVx8_ASAP7_75t_L g747 ( 
.A(n_653),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_705),
.B(n_300),
.Y(n_748)
);

A2O1A1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_576),
.A2(n_326),
.B(n_376),
.C(n_309),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_603),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_605),
.A2(n_346),
.B1(n_313),
.B2(n_380),
.Y(n_751)
);

O2A1O1Ixp5_ASAP7_75t_L g752 ( 
.A1(n_576),
.A2(n_306),
.B(n_311),
.C(n_394),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_587),
.B(n_463),
.C(n_454),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_682),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_578),
.B(n_316),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_682),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_SL g757 ( 
.A(n_697),
.B(n_268),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_624),
.A2(n_361),
.B1(n_392),
.B2(n_374),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_580),
.B(n_585),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_594),
.B(n_319),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_633),
.Y(n_761)
);

INVxp67_ASAP7_75t_SL g762 ( 
.A(n_662),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_576),
.B(n_322),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_617),
.B(n_327),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_634),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_612),
.B(n_331),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_609),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_606),
.B(n_619),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_638),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_613),
.B(n_340),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_658),
.B(n_385),
.Y(n_771)
);

AND2x2_ASAP7_75t_SL g772 ( 
.A(n_616),
.B(n_349),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_626),
.B(n_350),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_646),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_694),
.B(n_353),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_584),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_583),
.B(n_393),
.Y(n_777)
);

A2O1A1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_601),
.A2(n_314),
.B(n_388),
.C(n_363),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_694),
.B(n_365),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_683),
.B(n_366),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_683),
.B(n_367),
.Y(n_781)
);

AO221x1_ASAP7_75t_L g782 ( 
.A1(n_623),
.A2(n_387),
.B1(n_386),
.B2(n_371),
.C(n_377),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_683),
.B(n_279),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_685),
.B(n_286),
.Y(n_784)
);

NOR3xp33_ASAP7_75t_L g785 ( 
.A(n_636),
.B(n_393),
.C(n_389),
.Y(n_785)
);

O2A1O1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_582),
.A2(n_332),
.B(n_384),
.C(n_310),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_650),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_685),
.B(n_297),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_685),
.B(n_301),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_623),
.A2(n_389),
.B1(n_379),
.B2(n_378),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_689),
.B(n_315),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_689),
.B(n_317),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_689),
.B(n_324),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_655),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_609),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_664),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_584),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_668),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_591),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_621),
.Y(n_800)
);

O2A1O1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_582),
.A2(n_329),
.B(n_382),
.C(n_199),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_698),
.B(n_196),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_621),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_698),
.B(n_197),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_591),
.Y(n_805)
);

NOR2xp67_ASAP7_75t_L g806 ( 
.A(n_697),
.B(n_197),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_623),
.A2(n_379),
.B1(n_378),
.B2(n_226),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_662),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_616),
.B(n_601),
.Y(n_809)
);

INVxp67_ASAP7_75t_SL g810 ( 
.A(n_662),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_583),
.B(n_226),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_667),
.A2(n_382),
.B1(n_381),
.B2(n_200),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_703),
.B(n_199),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_679),
.B(n_200),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_630),
.A2(n_381),
.B1(n_217),
.B2(n_375),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_691),
.B(n_627),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_597),
.B(n_208),
.Y(n_817)
);

OAI221xp5_ASAP7_75t_L g818 ( 
.A1(n_707),
.A2(n_335),
.B1(n_227),
.B2(n_230),
.C(n_370),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_595),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_701),
.B(n_201),
.Y(n_820)
);

NOR2x1_ASAP7_75t_L g821 ( 
.A(n_645),
.B(n_712),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_627),
.B(n_201),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_627),
.B(n_217),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_595),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_644),
.Y(n_825)
);

OAI22xp33_ASAP7_75t_L g826 ( 
.A1(n_610),
.A2(n_227),
.B1(n_230),
.B2(n_232),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_597),
.A2(n_338),
.B1(n_375),
.B2(n_231),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_644),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_599),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_SL g830 ( 
.A1(n_721),
.A2(n_232),
.B1(n_238),
.B2(n_370),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_698),
.B(n_221),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_597),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_579),
.Y(n_833)
);

BUFx10_ASAP7_75t_L g834 ( 
.A(n_652),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_607),
.B(n_221),
.Y(n_835)
);

BUFx8_ASAP7_75t_L g836 ( 
.A(n_653),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_686),
.B(n_231),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_688),
.B(n_233),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_684),
.B(n_233),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_693),
.B(n_240),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_615),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_608),
.B(n_250),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_720),
.Y(n_843)
);

OAI22xp33_ASAP7_75t_L g844 ( 
.A1(n_699),
.A2(n_347),
.B1(n_238),
.B2(n_369),
.Y(n_844)
);

NOR2xp67_ASAP7_75t_SL g845 ( 
.A(n_592),
.B(n_240),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_635),
.B(n_250),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_607),
.B(n_631),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_647),
.B(n_245),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_700),
.B(n_245),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_661),
.Y(n_850)
);

OAI22xp33_ASAP7_75t_L g851 ( 
.A1(n_726),
.A2(n_642),
.B1(n_604),
.B2(n_709),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_623),
.A2(n_344),
.B1(n_239),
.B2(n_369),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_654),
.A2(n_285),
.B(n_337),
.Y(n_853)
);

NOR2xp67_ASAP7_75t_L g854 ( 
.A(n_710),
.B(n_284),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_599),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_702),
.B(n_284),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_692),
.B(n_285),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_631),
.B(n_337),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_692),
.B(n_338),
.Y(n_859)
);

NAND2x1_ASAP7_75t_L g860 ( 
.A(n_660),
.B(n_72),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_622),
.B(n_339),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_665),
.B(n_666),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_695),
.B(n_663),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_596),
.B(n_339),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_L g865 ( 
.A(n_710),
.B(n_719),
.Y(n_865)
);

NOR2xp67_ASAP7_75t_L g866 ( 
.A(n_710),
.B(n_345),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_625),
.B(n_345),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_596),
.B(n_354),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_596),
.B(n_354),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_661),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_704),
.B(n_357),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_600),
.B(n_357),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_704),
.B(n_359),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_656),
.B(n_359),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_600),
.B(n_222),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_SL g876 ( 
.A(n_717),
.B(n_222),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_632),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_639),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_716),
.A2(n_377),
.B1(n_373),
.B2(n_273),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_600),
.B(n_222),
.Y(n_880)
);

O2A1O1Ixp5_ASAP7_75t_L g881 ( 
.A1(n_674),
.A2(n_377),
.B(n_373),
.C(n_273),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_639),
.Y(n_882)
);

NOR3xp33_ASAP7_75t_L g883 ( 
.A(n_716),
.B(n_344),
.C(n_368),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_706),
.B(n_239),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_643),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_645),
.B(n_273),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_642),
.B(n_250),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_656),
.B(n_373),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_678),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_669),
.B(n_305),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_659),
.B(n_305),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_678),
.B(n_334),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_706),
.A2(n_305),
.B(n_362),
.C(n_360),
.Y(n_893)
);

BUFx8_ASAP7_75t_L g894 ( 
.A(n_653),
.Y(n_894)
);

BUFx2_ASAP7_75t_L g895 ( 
.A(n_714),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_L g896 ( 
.A(n_851),
.B(n_713),
.C(n_724),
.Y(n_896)
);

INVx11_ASAP7_75t_L g897 ( 
.A(n_836),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_738),
.B(n_690),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_763),
.A2(n_673),
.B(n_670),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_768),
.B(n_690),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_847),
.A2(n_654),
.B(n_640),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_847),
.A2(n_654),
.B(n_640),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_750),
.B(n_726),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_733),
.B(n_719),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_771),
.B(n_659),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_771),
.B(n_670),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_763),
.A2(n_764),
.B(n_809),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_861),
.B(n_671),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_764),
.A2(n_611),
.B(n_640),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_746),
.A2(n_708),
.B(n_674),
.C(n_671),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_SL g911 ( 
.A(n_879),
.B(n_581),
.C(n_725),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_884),
.A2(n_708),
.B(n_651),
.C(n_657),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_737),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_861),
.B(n_677),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_741),
.B(n_862),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_889),
.B(n_723),
.Y(n_916)
);

INVx1_ASAP7_75t_SL g917 ( 
.A(n_895),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_841),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_772),
.A2(n_867),
.B1(n_729),
.B2(n_730),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_884),
.A2(n_651),
.B(n_657),
.C(n_343),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_786),
.A2(n_873),
.B(n_871),
.C(n_857),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_762),
.A2(n_618),
.B(n_579),
.Y(n_922)
);

NAND2x1p5_ASAP7_75t_L g923 ( 
.A(n_743),
.B(n_717),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_735),
.A2(n_680),
.B(n_677),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_867),
.B(n_680),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_814),
.B(n_615),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_832),
.B(n_715),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_808),
.A2(n_637),
.B(n_579),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_814),
.B(n_615),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_820),
.B(n_588),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_772),
.B(n_715),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_734),
.B(n_718),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_810),
.A2(n_618),
.B(n_629),
.Y(n_933)
);

INVx1_ASAP7_75t_SL g934 ( 
.A(n_843),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_863),
.B(n_777),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_836),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_841),
.A2(n_648),
.B(n_643),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_811),
.B(n_717),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_865),
.B(n_718),
.Y(n_939)
);

AND2x6_ASAP7_75t_SL g940 ( 
.A(n_857),
.B(n_696),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_816),
.A2(n_592),
.B1(n_614),
.B2(n_660),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_887),
.B(n_614),
.Y(n_942)
);

AO22x1_ASAP7_75t_L g943 ( 
.A1(n_883),
.A2(n_333),
.B1(n_368),
.B2(n_335),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_783),
.A2(n_618),
.B(n_637),
.Y(n_944)
);

AO21x1_ASAP7_75t_L g945 ( 
.A1(n_746),
.A2(n_648),
.B(n_649),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_892),
.B(n_592),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_788),
.A2(n_618),
.B(n_637),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_817),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_739),
.B(n_588),
.Y(n_949)
);

BUFx2_ASAP7_75t_SL g950 ( 
.A(n_806),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_789),
.A2(n_629),
.B(n_637),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_820),
.A2(n_592),
.B1(n_660),
.B2(n_629),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_739),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_744),
.B(n_588),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_791),
.A2(n_793),
.B(n_792),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_728),
.A2(n_629),
.B(n_676),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_731),
.A2(n_676),
.B(n_641),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_754),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_848),
.B(n_588),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_736),
.B(n_590),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_751),
.A2(n_334),
.B1(n_333),
.B2(n_352),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_871),
.A2(n_352),
.B(n_343),
.C(n_347),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_842),
.B(n_334),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_735),
.A2(n_752),
.B(n_748),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_759),
.A2(n_676),
.B(n_641),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_756),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_742),
.B(n_590),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_761),
.B(n_765),
.Y(n_968)
);

CKINVDCx6p67_ASAP7_75t_R g969 ( 
.A(n_747),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_833),
.A2(n_780),
.B(n_784),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_833),
.A2(n_676),
.B(n_641),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_833),
.A2(n_676),
.B(n_641),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_778),
.A2(n_649),
.B(n_590),
.C(n_360),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_756),
.B(n_800),
.Y(n_974)
);

AO21x1_ASAP7_75t_L g975 ( 
.A1(n_859),
.A2(n_590),
.B(n_660),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_769),
.B(n_641),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_774),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_745),
.A2(n_362),
.B(n_356),
.Y(n_978)
);

AOI21x1_ASAP7_75t_L g979 ( 
.A1(n_781),
.A2(n_151),
.B(n_77),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_859),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_833),
.A2(n_356),
.B(n_348),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_740),
.A2(n_348),
.B1(n_190),
.B2(n_185),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_787),
.B(n_794),
.Y(n_983)
);

NAND2x1p5_ASAP7_75t_L g984 ( 
.A(n_743),
.B(n_181),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_776),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_796),
.B(n_19),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_846),
.B(n_19),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_751),
.A2(n_164),
.B1(n_160),
.B2(n_158),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_821),
.A2(n_155),
.B(n_152),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_798),
.B(n_20),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_803),
.B(n_20),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_839),
.B(n_21),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_776),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_825),
.B(n_828),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_850),
.B(n_23),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_797),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_864),
.A2(n_140),
.B(n_125),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_868),
.A2(n_872),
.B(n_869),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_870),
.B(n_24),
.Y(n_999)
);

AO22x1_ASAP7_75t_L g1000 ( 
.A1(n_873),
.A2(n_24),
.B1(n_27),
.B2(n_29),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_840),
.A2(n_115),
.B1(n_112),
.B2(n_106),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_781),
.A2(n_94),
.B(n_88),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_766),
.A2(n_78),
.B(n_73),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_732),
.B(n_834),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_732),
.B(n_27),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_775),
.B(n_29),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_779),
.A2(n_30),
.B(n_32),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_766),
.A2(n_30),
.B(n_34),
.Y(n_1008)
);

BUFx4f_ASAP7_75t_L g1009 ( 
.A(n_747),
.Y(n_1009)
);

CKINVDCx10_ASAP7_75t_R g1010 ( 
.A(n_727),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_834),
.B(n_36),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_797),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_758),
.B(n_38),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_767),
.B(n_38),
.Y(n_1014)
);

BUFx4f_ASAP7_75t_L g1015 ( 
.A(n_747),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_795),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_749),
.A2(n_41),
.B(n_42),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_758),
.B(n_43),
.Y(n_1018)
);

AOI21x1_ASAP7_75t_L g1019 ( 
.A1(n_877),
.A2(n_43),
.B(n_45),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_826),
.B(n_47),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_773),
.B(n_47),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_854),
.B(n_866),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_755),
.B(n_54),
.Y(n_1023)
);

CKINVDCx11_ASAP7_75t_R g1024 ( 
.A(n_894),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_853),
.A2(n_58),
.B(n_59),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_760),
.B(n_58),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_822),
.A2(n_60),
.B(n_63),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_770),
.B(n_66),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_799),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_799),
.B(n_66),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_805),
.B(n_67),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_823),
.A2(n_878),
.B(n_882),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_805),
.B(n_829),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_819),
.Y(n_1034)
);

CKINVDCx10_ASAP7_75t_R g1035 ( 
.A(n_894),
.Y(n_1035)
);

OAI321xp33_ASAP7_75t_L g1036 ( 
.A1(n_818),
.A2(n_844),
.A3(n_830),
.B1(n_807),
.B2(n_852),
.C(n_790),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_824),
.B(n_829),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_858),
.A2(n_886),
.B1(n_807),
.B2(n_852),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_855),
.B(n_885),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_813),
.B(n_837),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_838),
.B(n_856),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_860),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_875),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_753),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_802),
.A2(n_831),
.B(n_804),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_802),
.A2(n_831),
.B(n_804),
.Y(n_1046)
);

NOR3xp33_ASAP7_75t_L g1047 ( 
.A(n_785),
.B(n_893),
.C(n_891),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_880),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_757),
.B(n_876),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_849),
.A2(n_835),
.B(n_874),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_835),
.A2(n_874),
.B(n_890),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_827),
.B(n_815),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_749),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_790),
.B(n_812),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_801),
.A2(n_778),
.B(n_888),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_888),
.A2(n_891),
.B(n_881),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_782),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_845),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_763),
.A2(n_576),
.B(n_764),
.Y(n_1059)
);

NOR3xp33_ASAP7_75t_L g1060 ( 
.A(n_851),
.B(n_713),
.C(n_724),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_847),
.A2(n_576),
.B(n_654),
.Y(n_1061)
);

NOR3xp33_ASAP7_75t_L g1062 ( 
.A(n_851),
.B(n_713),
.C(n_724),
.Y(n_1062)
);

INVxp67_ASAP7_75t_L g1063 ( 
.A(n_741),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_737),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_889),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_889),
.B(n_642),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_738),
.B(n_768),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_833),
.Y(n_1068)
);

INVxp67_ASAP7_75t_SL g1069 ( 
.A(n_833),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_847),
.A2(n_576),
.B(n_654),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_738),
.B(n_768),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_746),
.A2(n_735),
.B(n_764),
.C(n_738),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_738),
.B(n_768),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_741),
.B(n_768),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_733),
.A2(n_884),
.B(n_786),
.C(n_589),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_738),
.B(n_768),
.Y(n_1076)
);

CKINVDCx10_ASAP7_75t_R g1077 ( 
.A(n_727),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_733),
.A2(n_738),
.B1(n_750),
.B2(n_764),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_847),
.A2(n_576),
.B(n_654),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_741),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_917),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_1068),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_1059),
.A2(n_921),
.B(n_1061),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_977),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1067),
.B(n_1071),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_915),
.B(n_1074),
.Y(n_1086)
);

AOI21xp33_ASAP7_75t_L g1087 ( 
.A1(n_921),
.A2(n_1038),
.B(n_1054),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_955),
.A2(n_970),
.B(n_1070),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1079),
.A2(n_907),
.B(n_998),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_909),
.A2(n_902),
.B(n_901),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_944),
.A2(n_951),
.B(n_947),
.Y(n_1091)
);

AOI221xp5_ASAP7_75t_L g1092 ( 
.A1(n_1036),
.A2(n_961),
.B1(n_1020),
.B2(n_896),
.C(n_1062),
.Y(n_1092)
);

AO21x1_ASAP7_75t_L g1093 ( 
.A1(n_1025),
.A2(n_1078),
.B(n_1046),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_1060),
.A2(n_992),
.B1(n_904),
.B2(n_1052),
.Y(n_1094)
);

AO21x2_ASAP7_75t_L g1095 ( 
.A1(n_964),
.A2(n_1045),
.B(n_1056),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_1075),
.A2(n_992),
.B(n_1072),
.C(n_980),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1073),
.B(n_1076),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_948),
.B(n_927),
.Y(n_1098)
);

BUFx8_ASAP7_75t_SL g1099 ( 
.A(n_936),
.Y(n_1099)
);

AOI21xp33_ASAP7_75t_L g1100 ( 
.A1(n_1075),
.A2(n_904),
.B(n_898),
.Y(n_1100)
);

AO31x2_ASAP7_75t_L g1101 ( 
.A1(n_945),
.A2(n_975),
.A3(n_1053),
.B(n_912),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1040),
.B(n_1041),
.Y(n_1102)
);

AOI21xp33_ASAP7_75t_L g1103 ( 
.A1(n_935),
.A2(n_900),
.B(n_1049),
.Y(n_1103)
);

AOI21x1_ASAP7_75t_L g1104 ( 
.A1(n_926),
.A2(n_929),
.B(n_930),
.Y(n_1104)
);

NOR2x1_ASAP7_75t_SL g1105 ( 
.A(n_1068),
.B(n_1058),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_935),
.B(n_927),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_927),
.B(n_942),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1043),
.B(n_1048),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_1068),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1043),
.B(n_1048),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_908),
.A2(n_925),
.B(n_914),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_905),
.B(n_906),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_919),
.A2(n_1050),
.B(n_924),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1032),
.A2(n_956),
.B(n_899),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_922),
.A2(n_928),
.B(n_933),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_903),
.B(n_987),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_1068),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_903),
.B(n_968),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_1049),
.A2(n_1051),
.B(n_910),
.C(n_1055),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_1009),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_1065),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_960),
.A2(n_959),
.B(n_954),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_1080),
.B(n_1066),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_957),
.A2(n_1033),
.B(n_1039),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1009),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_938),
.A2(n_1047),
.B(n_912),
.C(n_1044),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1037),
.A2(n_972),
.B(n_971),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_983),
.B(n_994),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1042),
.A2(n_1069),
.B(n_1022),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_963),
.B(n_1063),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_913),
.A2(n_958),
.B(n_1064),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_1065),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_938),
.B(n_1004),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1015),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_913),
.A2(n_1064),
.B(n_958),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_978),
.A2(n_1020),
.B(n_931),
.C(n_1017),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_946),
.B(n_1005),
.Y(n_1137)
);

AO21x1_ASAP7_75t_L g1138 ( 
.A1(n_1003),
.A2(n_931),
.B(n_1001),
.Y(n_1138)
);

O2A1O1Ixp5_ASAP7_75t_L g1139 ( 
.A1(n_1006),
.A2(n_932),
.B(n_1028),
.C(n_1026),
.Y(n_1139)
);

AND2x6_ASAP7_75t_L g1140 ( 
.A(n_1058),
.B(n_1042),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_962),
.A2(n_991),
.B(n_995),
.C(n_999),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_974),
.B(n_986),
.Y(n_1142)
);

INVx5_ASAP7_75t_L g1143 ( 
.A(n_1058),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_993),
.A2(n_1029),
.B(n_1034),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_974),
.A2(n_962),
.B(n_1029),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_934),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_990),
.B(n_939),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_939),
.B(n_966),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_SL g1149 ( 
.A1(n_961),
.A2(n_936),
.B1(n_1016),
.B2(n_916),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_993),
.A2(n_1034),
.B(n_1030),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1013),
.A2(n_1018),
.B(n_973),
.C(n_920),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_965),
.A2(n_985),
.B(n_953),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_1011),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_950),
.B(n_943),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1031),
.A2(n_996),
.B(n_1012),
.Y(n_1155)
);

AO31x2_ASAP7_75t_L g1156 ( 
.A1(n_1057),
.A2(n_920),
.A3(n_1021),
.B(n_1023),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_952),
.A2(n_941),
.B(n_967),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_918),
.B(n_932),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1014),
.A2(n_988),
.B1(n_982),
.B2(n_918),
.Y(n_1159)
);

INVx1_ASAP7_75t_SL g1160 ( 
.A(n_1014),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_976),
.A2(n_949),
.B(n_985),
.Y(n_1161)
);

INVxp67_ASAP7_75t_L g1162 ( 
.A(n_981),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_923),
.B(n_1027),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_911),
.B(n_940),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_979),
.A2(n_997),
.B(n_989),
.Y(n_1165)
);

INVx1_ASAP7_75t_SL g1166 ( 
.A(n_923),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_SL g1167 ( 
.A1(n_1008),
.A2(n_1019),
.B(n_1002),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_984),
.Y(n_1168)
);

NAND3xp33_ASAP7_75t_L g1169 ( 
.A(n_1000),
.B(n_1007),
.C(n_1058),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_984),
.A2(n_1015),
.B(n_969),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_897),
.A2(n_1024),
.B(n_1035),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1024),
.A2(n_1010),
.B(n_1077),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1059),
.A2(n_921),
.B(n_1061),
.Y(n_1173)
);

BUFx10_ASAP7_75t_L g1174 ( 
.A(n_1049),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1067),
.B(n_1071),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1059),
.A2(n_921),
.B(n_1061),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_945),
.A2(n_975),
.A3(n_749),
.B(n_921),
.Y(n_1177)
);

AO31x2_ASAP7_75t_L g1178 ( 
.A1(n_945),
.A2(n_975),
.A3(n_749),
.B(n_921),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1068),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1067),
.B(n_1071),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_985),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_915),
.B(n_1074),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1067),
.B(n_1071),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1059),
.A2(n_921),
.B(n_1061),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_985),
.Y(n_1185)
);

NAND2x1_ASAP7_75t_L g1186 ( 
.A(n_1068),
.B(n_985),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1059),
.A2(n_921),
.B(n_1061),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1067),
.B(n_1071),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_977),
.Y(n_1189)
);

INVx4_ASAP7_75t_L g1190 ( 
.A(n_1068),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1068),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_937),
.A2(n_947),
.B(n_944),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_1068),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_937),
.A2(n_947),
.B(n_944),
.Y(n_1194)
);

AO21x1_ASAP7_75t_L g1195 ( 
.A1(n_1025),
.A2(n_1078),
.B(n_1046),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1068),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1068),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_917),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1059),
.A2(n_921),
.B(n_1061),
.Y(n_1199)
);

OAI22x1_ASAP7_75t_L g1200 ( 
.A1(n_1049),
.A2(n_879),
.B1(n_733),
.B2(n_980),
.Y(n_1200)
);

AOI21xp33_ASAP7_75t_L g1201 ( 
.A1(n_921),
.A2(n_1038),
.B(n_1054),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_937),
.A2(n_947),
.B(n_944),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_937),
.A2(n_947),
.B(n_944),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_921),
.A2(n_1075),
.B(n_733),
.C(n_992),
.Y(n_1204)
);

INVx4_ASAP7_75t_L g1205 ( 
.A(n_1068),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1059),
.A2(n_921),
.B(n_1061),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1067),
.B(n_1071),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1067),
.B(n_1071),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_980),
.B(n_750),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1059),
.A2(n_921),
.B(n_1061),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_937),
.A2(n_947),
.B(n_944),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1067),
.B(n_1071),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1059),
.A2(n_921),
.B(n_1061),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1067),
.B(n_1071),
.Y(n_1214)
);

HAxp5_ASAP7_75t_L g1215 ( 
.A(n_1010),
.B(n_830),
.CON(n_1215),
.SN(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_955),
.A2(n_576),
.B(n_1059),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_921),
.A2(n_1075),
.B(n_733),
.C(n_992),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_937),
.A2(n_947),
.B(n_944),
.Y(n_1218)
);

AOI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1061),
.A2(n_764),
.B(n_1070),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_921),
.A2(n_733),
.B1(n_1075),
.B2(n_1054),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_985),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_937),
.A2(n_947),
.B(n_944),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_937),
.A2(n_947),
.B(n_944),
.Y(n_1223)
);

AOI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1061),
.A2(n_764),
.B(n_1070),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_937),
.A2(n_947),
.B(n_944),
.Y(n_1225)
);

AOI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1061),
.A2(n_764),
.B(n_1070),
.Y(n_1226)
);

NAND2x1_ASAP7_75t_L g1227 ( 
.A(n_1068),
.B(n_985),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1068),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_937),
.A2(n_947),
.B(n_944),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1054),
.A2(n_1038),
.B1(n_1060),
.B2(n_896),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_937),
.A2(n_947),
.B(n_944),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_915),
.B(n_1074),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1081),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1102),
.B(n_1118),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1097),
.B(n_1175),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_1123),
.B(n_1116),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1085),
.B(n_1207),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1086),
.B(n_1182),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1097),
.B(n_1175),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1120),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1232),
.B(n_1153),
.Y(n_1241)
);

INVx8_ASAP7_75t_L g1242 ( 
.A(n_1082),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1180),
.B(n_1183),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1081),
.B(n_1198),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1121),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1153),
.B(n_1130),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1190),
.Y(n_1247)
);

NAND2x1p5_ASAP7_75t_L g1248 ( 
.A(n_1198),
.B(n_1120),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1107),
.B(n_1098),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1180),
.B(n_1183),
.Y(n_1250)
);

AOI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1230),
.A2(n_1106),
.B1(n_1164),
.B2(n_1188),
.Y(n_1251)
);

BUFx12f_ASAP7_75t_L g1252 ( 
.A(n_1120),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1188),
.B(n_1208),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1103),
.B(n_1209),
.Y(n_1254)
);

INVx4_ASAP7_75t_L g1255 ( 
.A(n_1125),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1212),
.B(n_1214),
.Y(n_1256)
);

INVx4_ASAP7_75t_L g1257 ( 
.A(n_1125),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1133),
.B(n_1128),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1204),
.A2(n_1217),
.B1(n_1096),
.B2(n_1220),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1132),
.B(n_1146),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1107),
.B(n_1160),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1132),
.B(n_1108),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_1108),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1112),
.B(n_1110),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1200),
.A2(n_1149),
.B1(n_1100),
.B2(n_1220),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1112),
.B(n_1110),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1189),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1160),
.B(n_1111),
.Y(n_1268)
);

OR2x2_ASAP7_75t_SL g1269 ( 
.A(n_1125),
.B(n_1134),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1100),
.A2(n_1087),
.B1(n_1201),
.B2(n_1138),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1126),
.B(n_1137),
.Y(n_1271)
);

INVx3_ASAP7_75t_SL g1272 ( 
.A(n_1134),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1098),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1174),
.B(n_1147),
.Y(n_1274)
);

OAI21xp33_ASAP7_75t_L g1275 ( 
.A1(n_1087),
.A2(n_1201),
.B(n_1141),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1154),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1134),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1093),
.A2(n_1195),
.B1(n_1159),
.B2(n_1169),
.Y(n_1278)
);

AOI21x1_ASAP7_75t_SL g1279 ( 
.A1(n_1163),
.A2(n_1142),
.B(n_1158),
.Y(n_1279)
);

OR2x6_ASAP7_75t_L g1280 ( 
.A(n_1170),
.B(n_1168),
.Y(n_1280)
);

AOI221xp5_ASAP7_75t_L g1281 ( 
.A1(n_1159),
.A2(n_1151),
.B1(n_1083),
.B2(n_1187),
.C(n_1199),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1181),
.Y(n_1282)
);

INVx4_ASAP7_75t_L g1283 ( 
.A(n_1082),
.Y(n_1283)
);

OR2x6_ASAP7_75t_L g1284 ( 
.A(n_1082),
.B(n_1191),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1191),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1174),
.B(n_1215),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1162),
.A2(n_1083),
.B1(n_1187),
.B2(n_1210),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1191),
.Y(n_1288)
);

AOI221xp5_ASAP7_75t_L g1289 ( 
.A1(n_1173),
.A2(n_1199),
.B1(n_1176),
.B2(n_1184),
.C(n_1213),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_1099),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1171),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1119),
.A2(n_1143),
.B1(n_1206),
.B2(n_1176),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1216),
.A2(n_1089),
.B(n_1088),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1193),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1185),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1148),
.Y(n_1296)
);

NOR2xp67_ASAP7_75t_L g1297 ( 
.A(n_1143),
.B(n_1190),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1166),
.B(n_1145),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1156),
.B(n_1221),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1193),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1143),
.B(n_1166),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1171),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1113),
.A2(n_1129),
.B(n_1184),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1156),
.B(n_1145),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1109),
.B(n_1197),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1193),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1156),
.B(n_1109),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_1172),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1117),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1117),
.B(n_1179),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_SL g1311 ( 
.A(n_1205),
.B(n_1140),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1139),
.A2(n_1206),
.B(n_1173),
.C(n_1213),
.Y(n_1312)
);

OR2x6_ASAP7_75t_L g1313 ( 
.A(n_1196),
.B(n_1228),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1179),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1140),
.B(n_1155),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1197),
.B(n_1105),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1228),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1095),
.B(n_1155),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1228),
.B(n_1140),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1210),
.A2(n_1113),
.B1(n_1150),
.B2(n_1157),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1101),
.B(n_1178),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1090),
.A2(n_1122),
.B(n_1091),
.Y(n_1322)
);

NAND3xp33_ASAP7_75t_SL g1323 ( 
.A(n_1150),
.B(n_1161),
.C(n_1186),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1140),
.B(n_1101),
.Y(n_1324)
);

INVx5_ASAP7_75t_L g1325 ( 
.A(n_1227),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1219),
.B(n_1226),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1152),
.Y(n_1327)
);

NOR2xp67_ASAP7_75t_L g1328 ( 
.A(n_1224),
.B(n_1104),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1127),
.B(n_1115),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1124),
.Y(n_1330)
);

INVxp67_ASAP7_75t_L g1331 ( 
.A(n_1167),
.Y(n_1331)
);

AOI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1192),
.A2(n_1231),
.B(n_1203),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1177),
.B(n_1178),
.Y(n_1333)
);

OR2x6_ASAP7_75t_L g1334 ( 
.A(n_1114),
.B(n_1165),
.Y(n_1334)
);

BUFx12f_ASAP7_75t_L g1335 ( 
.A(n_1178),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1194),
.B(n_1222),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1202),
.Y(n_1337)
);

OR2x2_ASAP7_75t_L g1338 ( 
.A(n_1211),
.B(n_1218),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1223),
.A2(n_921),
.B(n_1092),
.C(n_1136),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1225),
.B(n_1229),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1190),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1121),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1086),
.B(n_915),
.Y(n_1343)
);

CKINVDCx8_ASAP7_75t_R g1344 ( 
.A(n_1120),
.Y(n_1344)
);

NAND2x1_ASAP7_75t_L g1345 ( 
.A(n_1140),
.B(n_1068),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1107),
.B(n_1098),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1102),
.B(n_1123),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1084),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1086),
.B(n_915),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1107),
.B(n_1098),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1086),
.B(n_915),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1102),
.B(n_1097),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1107),
.B(n_1098),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1121),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1131),
.A2(n_1144),
.B(n_1135),
.Y(n_1355)
);

INVx3_ASAP7_75t_SL g1356 ( 
.A(n_1081),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1120),
.Y(n_1357)
);

CKINVDCx8_ASAP7_75t_R g1358 ( 
.A(n_1120),
.Y(n_1358)
);

INVxp67_ASAP7_75t_L g1359 ( 
.A(n_1121),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1190),
.Y(n_1360)
);

CKINVDCx16_ASAP7_75t_R g1361 ( 
.A(n_1171),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1102),
.B(n_750),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1102),
.B(n_1097),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1107),
.B(n_1098),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1102),
.B(n_1097),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1121),
.Y(n_1366)
);

INVx4_ASAP7_75t_L g1367 ( 
.A(n_1120),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1102),
.A2(n_1094),
.B1(n_1136),
.B2(n_733),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1086),
.B(n_915),
.Y(n_1369)
);

INVx2_ASAP7_75t_SL g1370 ( 
.A(n_1121),
.Y(n_1370)
);

NAND2x1p5_ASAP7_75t_L g1371 ( 
.A(n_1081),
.B(n_1198),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1086),
.B(n_915),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1102),
.B(n_1097),
.Y(n_1373)
);

OA21x2_ASAP7_75t_L g1374 ( 
.A1(n_1339),
.A2(n_1322),
.B(n_1293),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1238),
.B(n_1343),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1269),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1344),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_SL g1378 ( 
.A1(n_1361),
.A2(n_1259),
.B1(n_1368),
.B2(n_1254),
.Y(n_1378)
);

AOI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1302),
.A2(n_1362),
.B1(n_1251),
.B2(n_1258),
.Y(n_1379)
);

AOI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1274),
.A2(n_1368),
.B1(n_1349),
.B2(n_1351),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1237),
.B(n_1256),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1267),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1369),
.B(n_1372),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1263),
.Y(n_1384)
);

NAND2x1p5_ASAP7_75t_L g1385 ( 
.A(n_1263),
.B(n_1301),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1348),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1356),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1308),
.A2(n_1265),
.B1(n_1291),
.B2(n_1276),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_SL g1389 ( 
.A1(n_1259),
.A2(n_1292),
.B1(n_1253),
.B2(n_1234),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1233),
.Y(n_1390)
);

AO21x1_ASAP7_75t_L g1391 ( 
.A1(n_1271),
.A2(n_1292),
.B(n_1268),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1244),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1288),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1352),
.B(n_1363),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1253),
.A2(n_1235),
.B1(n_1250),
.B2(n_1239),
.Y(n_1395)
);

NAND2x1p5_ASAP7_75t_L g1396 ( 
.A(n_1301),
.B(n_1345),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1281),
.A2(n_1275),
.B1(n_1289),
.B2(n_1270),
.Y(n_1397)
);

BUFx4f_ASAP7_75t_SL g1398 ( 
.A(n_1252),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1358),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1261),
.B(n_1249),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1249),
.B(n_1346),
.Y(n_1401)
);

OR2x6_ASAP7_75t_L g1402 ( 
.A(n_1280),
.B(n_1315),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1352),
.B(n_1363),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1262),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1365),
.B(n_1373),
.Y(n_1405)
);

INVx4_ASAP7_75t_L g1406 ( 
.A(n_1240),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1282),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1241),
.B(n_1246),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1245),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1299),
.Y(n_1410)
);

CKINVDCx8_ASAP7_75t_R g1411 ( 
.A(n_1240),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1286),
.A2(n_1350),
.B1(n_1364),
.B2(n_1346),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1295),
.Y(n_1413)
);

OAI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1365),
.A2(n_1373),
.B1(n_1235),
.B2(n_1239),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1355),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1317),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1296),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1264),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1347),
.B(n_1236),
.Y(n_1419)
);

AO21x1_ASAP7_75t_L g1420 ( 
.A1(n_1315),
.A2(n_1320),
.B(n_1298),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1266),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1243),
.B(n_1250),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1309),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1275),
.A2(n_1243),
.B1(n_1287),
.B2(n_1278),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1314),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1317),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1350),
.B(n_1353),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1310),
.Y(n_1428)
);

NOR2xp67_ASAP7_75t_L g1429 ( 
.A(n_1260),
.B(n_1359),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1353),
.A2(n_1364),
.B1(n_1273),
.B2(n_1354),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1366),
.A2(n_1370),
.B1(n_1342),
.B2(n_1272),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1306),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1326),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1305),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1371),
.B(n_1248),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1307),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1285),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1240),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1290),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1333),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1320),
.A2(n_1303),
.B1(n_1318),
.B2(n_1335),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1277),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1304),
.A2(n_1333),
.B1(n_1321),
.B2(n_1331),
.Y(n_1443)
);

INVx4_ASAP7_75t_SL g1444 ( 
.A(n_1284),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1294),
.B(n_1300),
.Y(n_1445)
);

INVx6_ASAP7_75t_L g1446 ( 
.A(n_1255),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_SL g1447 ( 
.A1(n_1311),
.A2(n_1357),
.B1(n_1367),
.B2(n_1255),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1257),
.B(n_1367),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1338),
.A2(n_1279),
.B(n_1336),
.Y(n_1449)
);

BUFx12f_ASAP7_75t_L g1450 ( 
.A(n_1357),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1312),
.B(n_1257),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1357),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1327),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1316),
.B(n_1360),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1247),
.B(n_1360),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1334),
.Y(n_1456)
);

AOI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1328),
.A2(n_1329),
.B(n_1334),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1334),
.Y(n_1458)
);

NAND2x1p5_ASAP7_75t_L g1459 ( 
.A(n_1297),
.B(n_1341),
.Y(n_1459)
);

CKINVDCx20_ASAP7_75t_R g1460 ( 
.A(n_1242),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1313),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1330),
.Y(n_1462)
);

BUFx2_ASAP7_75t_SL g1463 ( 
.A(n_1297),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1247),
.B(n_1341),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1317),
.Y(n_1465)
);

AOI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1329),
.A2(n_1324),
.B(n_1280),
.Y(n_1466)
);

OAI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1311),
.A2(n_1325),
.B1(n_1323),
.B2(n_1283),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_SL g1468 ( 
.A1(n_1325),
.A2(n_1242),
.B1(n_1330),
.B2(n_1340),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1337),
.Y(n_1469)
);

CKINVDCx11_ASAP7_75t_R g1470 ( 
.A(n_1242),
.Y(n_1470)
);

INVx6_ASAP7_75t_L g1471 ( 
.A(n_1325),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1337),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_1269),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1263),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1237),
.B(n_1256),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1368),
.A2(n_1092),
.B1(n_1094),
.B2(n_896),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1234),
.A2(n_1094),
.B1(n_1363),
.B2(n_1352),
.Y(n_1477)
);

CKINVDCx6p67_ASAP7_75t_R g1478 ( 
.A(n_1356),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1263),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1368),
.A2(n_1092),
.B1(n_1094),
.B2(n_896),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1263),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1234),
.A2(n_1094),
.B1(n_1363),
.B2(n_1352),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1355),
.A2(n_1332),
.B(n_1194),
.Y(n_1483)
);

OAI22xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1234),
.A2(n_876),
.B1(n_980),
.B2(n_1049),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1269),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1368),
.A2(n_1092),
.B1(n_1094),
.B2(n_896),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1355),
.A2(n_1332),
.B(n_1194),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1234),
.A2(n_1094),
.B1(n_1363),
.B2(n_1352),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1319),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1237),
.B(n_1256),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1269),
.Y(n_1491)
);

INVx6_ASAP7_75t_L g1492 ( 
.A(n_1252),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1402),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1436),
.B(n_1443),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1384),
.Y(n_1495)
);

BUFx2_ASAP7_75t_SL g1496 ( 
.A(n_1429),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1457),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1478),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1384),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1410),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1385),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1410),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1443),
.B(n_1441),
.Y(n_1503)
);

AO22x1_ASAP7_75t_L g1504 ( 
.A1(n_1394),
.A2(n_1418),
.B1(n_1421),
.B2(n_1376),
.Y(n_1504)
);

AO21x1_ASAP7_75t_SL g1505 ( 
.A1(n_1476),
.A2(n_1486),
.B(n_1480),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1462),
.Y(n_1506)
);

OA21x2_ASAP7_75t_L g1507 ( 
.A1(n_1441),
.A2(n_1487),
.B(n_1483),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1474),
.Y(n_1508)
);

AO21x2_ASAP7_75t_L g1509 ( 
.A1(n_1467),
.A2(n_1415),
.B(n_1391),
.Y(n_1509)
);

INVx2_ASAP7_75t_SL g1510 ( 
.A(n_1474),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1394),
.B(n_1419),
.Y(n_1511)
);

AO31x2_ASAP7_75t_L g1512 ( 
.A1(n_1420),
.A2(n_1415),
.A3(n_1453),
.B(n_1440),
.Y(n_1512)
);

OAI21xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1397),
.A2(n_1480),
.B(n_1476),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1385),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1456),
.B(n_1458),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1449),
.A2(n_1466),
.B(n_1458),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1439),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1456),
.B(n_1479),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1481),
.B(n_1453),
.Y(n_1519)
);

BUFx12f_ASAP7_75t_L g1520 ( 
.A(n_1470),
.Y(n_1520)
);

AOI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1451),
.A2(n_1477),
.B(n_1488),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1481),
.Y(n_1522)
);

AO21x2_ASAP7_75t_L g1523 ( 
.A1(n_1467),
.A2(n_1414),
.B(n_1469),
.Y(n_1523)
);

AO21x2_ASAP7_75t_L g1524 ( 
.A1(n_1414),
.A2(n_1469),
.B(n_1472),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1486),
.A2(n_1378),
.B1(n_1379),
.B2(n_1397),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1374),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1433),
.B(n_1408),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1383),
.B(n_1375),
.Y(n_1528)
);

AO21x2_ASAP7_75t_L g1529 ( 
.A1(n_1472),
.A2(n_1482),
.B(n_1380),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1381),
.B(n_1475),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1404),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1395),
.B(n_1490),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1382),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1403),
.B(n_1405),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1386),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1439),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1392),
.B(n_1388),
.Y(n_1537)
);

INVxp33_ASAP7_75t_L g1538 ( 
.A(n_1409),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1418),
.B(n_1421),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1444),
.B(n_1400),
.Y(n_1540)
);

INVx3_ASAP7_75t_L g1541 ( 
.A(n_1396),
.Y(n_1541)
);

CKINVDCx14_ASAP7_75t_R g1542 ( 
.A(n_1387),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1470),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1396),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1428),
.B(n_1389),
.Y(n_1545)
);

INVx3_ASAP7_75t_L g1546 ( 
.A(n_1471),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1424),
.B(n_1417),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1471),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1424),
.A2(n_1423),
.B(n_1425),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1422),
.B(n_1390),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1435),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1471),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1434),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1461),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1376),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1468),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1407),
.B(n_1413),
.Y(n_1557)
);

INVxp67_ASAP7_75t_SL g1558 ( 
.A(n_1432),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1437),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1444),
.Y(n_1560)
);

BUFx12f_ASAP7_75t_L g1561 ( 
.A(n_1452),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1454),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1455),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1444),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1464),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1459),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1400),
.B(n_1484),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1459),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1473),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1463),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1400),
.A2(n_1485),
.B1(n_1473),
.B2(n_1491),
.Y(n_1571)
);

INVx5_ASAP7_75t_SL g1572 ( 
.A(n_1401),
.Y(n_1572)
);

AOI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1465),
.A2(n_1448),
.B(n_1401),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_1446),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1489),
.Y(n_1575)
);

OA21x2_ASAP7_75t_L g1576 ( 
.A1(n_1412),
.A2(n_1430),
.B(n_1445),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1431),
.A2(n_1452),
.B(n_1427),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1512),
.B(n_1491),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1547),
.B(n_1485),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1512),
.B(n_1426),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1500),
.B(n_1426),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1547),
.B(n_1447),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1522),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1512),
.B(n_1526),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1512),
.B(n_1416),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1512),
.B(n_1416),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1493),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1499),
.B(n_1416),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1500),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1502),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1502),
.Y(n_1591)
);

BUFx4f_ASAP7_75t_SL g1592 ( 
.A(n_1520),
.Y(n_1592)
);

AOI221xp5_ASAP7_75t_L g1593 ( 
.A1(n_1513),
.A2(n_1377),
.B1(n_1399),
.B2(n_1442),
.C(n_1427),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1494),
.B(n_1426),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1530),
.B(n_1377),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1533),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1509),
.B(n_1393),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1577),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1508),
.B(n_1393),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1509),
.B(n_1393),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1509),
.B(n_1438),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1524),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1507),
.B(n_1438),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1505),
.A2(n_1399),
.B1(n_1492),
.B2(n_1398),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1507),
.B(n_1516),
.Y(n_1605)
);

INVxp67_ASAP7_75t_SL g1606 ( 
.A(n_1519),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1507),
.B(n_1406),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1518),
.B(n_1411),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1507),
.B(n_1492),
.Y(n_1609)
);

BUFx8_ASAP7_75t_L g1610 ( 
.A(n_1520),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1516),
.B(n_1492),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1503),
.B(n_1446),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1495),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1503),
.B(n_1446),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1495),
.B(n_1450),
.Y(n_1615)
);

AOI211xp5_ASAP7_75t_SL g1616 ( 
.A1(n_1556),
.A2(n_1460),
.B(n_1398),
.C(n_1450),
.Y(n_1616)
);

NOR2x1p5_ASAP7_75t_L g1617 ( 
.A(n_1521),
.B(n_1460),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1510),
.B(n_1519),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1515),
.B(n_1524),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1578),
.B(n_1577),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1578),
.B(n_1577),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1618),
.B(n_1510),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1618),
.B(n_1531),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1579),
.B(n_1532),
.Y(n_1624)
);

NAND3xp33_ASAP7_75t_L g1625 ( 
.A(n_1593),
.B(n_1525),
.C(n_1513),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1593),
.A2(n_1504),
.B(n_1534),
.Y(n_1626)
);

NAND4xp25_ASAP7_75t_L g1627 ( 
.A(n_1595),
.B(n_1567),
.C(n_1550),
.D(n_1537),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1617),
.A2(n_1505),
.B1(n_1545),
.B2(n_1537),
.Y(n_1628)
);

NAND3xp33_ASAP7_75t_L g1629 ( 
.A(n_1601),
.B(n_1556),
.C(n_1545),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_SL g1630 ( 
.A(n_1592),
.B(n_1498),
.Y(n_1630)
);

OAI21xp33_ASAP7_75t_L g1631 ( 
.A1(n_1579),
.A2(n_1521),
.B(n_1562),
.Y(n_1631)
);

OAI221xp5_ASAP7_75t_SL g1632 ( 
.A1(n_1604),
.A2(n_1571),
.B1(n_1511),
.B2(n_1553),
.C(n_1542),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1617),
.A2(n_1529),
.B1(n_1576),
.B2(n_1496),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1606),
.B(n_1562),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1606),
.B(n_1518),
.Y(n_1635)
);

NAND3xp33_ASAP7_75t_L g1636 ( 
.A(n_1601),
.B(n_1576),
.C(n_1504),
.Y(n_1636)
);

AOI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1582),
.A2(n_1553),
.B1(n_1528),
.B2(n_1558),
.C(n_1565),
.Y(n_1637)
);

NAND3xp33_ASAP7_75t_L g1638 ( 
.A(n_1601),
.B(n_1576),
.C(n_1570),
.Y(n_1638)
);

NAND3xp33_ASAP7_75t_L g1639 ( 
.A(n_1616),
.B(n_1600),
.C(n_1597),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1594),
.B(n_1563),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_L g1641 ( 
.A(n_1616),
.B(n_1576),
.C(n_1570),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1582),
.B(n_1496),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1619),
.B(n_1523),
.Y(n_1643)
);

OAI21xp33_ASAP7_75t_L g1644 ( 
.A1(n_1598),
.A2(n_1515),
.B(n_1527),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1611),
.B(n_1497),
.Y(n_1645)
);

NAND3xp33_ASAP7_75t_L g1646 ( 
.A(n_1597),
.B(n_1568),
.C(n_1554),
.Y(n_1646)
);

OAI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1615),
.A2(n_1555),
.B1(n_1569),
.B2(n_1551),
.C(n_1559),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1594),
.B(n_1554),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1612),
.B(n_1573),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1613),
.B(n_1529),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1613),
.B(n_1583),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1610),
.A2(n_1529),
.B1(n_1523),
.B2(n_1538),
.Y(n_1652)
);

OAI21xp33_ASAP7_75t_L g1653 ( 
.A1(n_1598),
.A2(n_1501),
.B(n_1514),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1592),
.A2(n_1555),
.B1(n_1569),
.B2(n_1561),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1619),
.B(n_1523),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1583),
.B(n_1535),
.Y(n_1656)
);

OAI221xp5_ASAP7_75t_L g1657 ( 
.A1(n_1615),
.A2(n_1555),
.B1(n_1569),
.B2(n_1544),
.C(n_1541),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_SL g1658 ( 
.A1(n_1610),
.A2(n_1540),
.B1(n_1572),
.B2(n_1541),
.Y(n_1658)
);

NAND3xp33_ASAP7_75t_L g1659 ( 
.A(n_1597),
.B(n_1568),
.C(n_1566),
.Y(n_1659)
);

OAI221xp5_ASAP7_75t_SL g1660 ( 
.A1(n_1608),
.A2(n_1557),
.B1(n_1539),
.B2(n_1564),
.C(n_1560),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1612),
.B(n_1573),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1588),
.B(n_1599),
.Y(n_1662)
);

OAI221xp5_ASAP7_75t_L g1663 ( 
.A1(n_1608),
.A2(n_1541),
.B1(n_1544),
.B2(n_1552),
.C(n_1546),
.Y(n_1663)
);

NAND3xp33_ASAP7_75t_L g1664 ( 
.A(n_1600),
.B(n_1566),
.C(n_1575),
.Y(n_1664)
);

NAND3xp33_ASAP7_75t_L g1665 ( 
.A(n_1600),
.B(n_1566),
.C(n_1575),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1614),
.B(n_1608),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1599),
.B(n_1587),
.Y(n_1667)
);

OA21x2_ASAP7_75t_L g1668 ( 
.A1(n_1605),
.A2(n_1549),
.B(n_1506),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1645),
.B(n_1609),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1635),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1643),
.B(n_1655),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1624),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1643),
.B(n_1589),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1620),
.B(n_1621),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1655),
.B(n_1650),
.Y(n_1675)
);

NOR2x1_ASAP7_75t_L g1676 ( 
.A(n_1636),
.B(n_1659),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1656),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1634),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1651),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1668),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1622),
.Y(n_1681)
);

INVx2_ASAP7_75t_SL g1682 ( 
.A(n_1645),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1668),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1668),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1623),
.B(n_1590),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1648),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1664),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1638),
.B(n_1602),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1665),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1649),
.B(n_1584),
.Y(n_1690)
);

AND2x4_ASAP7_75t_L g1691 ( 
.A(n_1639),
.B(n_1611),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1631),
.B(n_1590),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1640),
.B(n_1591),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1649),
.B(n_1605),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1661),
.B(n_1605),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1646),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1662),
.B(n_1591),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1667),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1661),
.B(n_1603),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1629),
.B(n_1596),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1644),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1666),
.B(n_1602),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1666),
.B(n_1603),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1652),
.B(n_1607),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1641),
.B(n_1611),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1674),
.B(n_1633),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1682),
.B(n_1580),
.Y(n_1707)
);

BUFx2_ASAP7_75t_L g1708 ( 
.A(n_1676),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1675),
.B(n_1581),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1672),
.B(n_1630),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1672),
.B(n_1624),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1674),
.B(n_1653),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1677),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1675),
.B(n_1581),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1679),
.B(n_1627),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1678),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1678),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1682),
.B(n_1580),
.Y(n_1718)
);

NOR2xp67_ASAP7_75t_L g1719 ( 
.A(n_1696),
.B(n_1657),
.Y(n_1719)
);

INVxp67_ASAP7_75t_L g1720 ( 
.A(n_1696),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1679),
.B(n_1642),
.Y(n_1721)
);

BUFx2_ASAP7_75t_L g1722 ( 
.A(n_1676),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1673),
.B(n_1581),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1684),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1677),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1682),
.B(n_1585),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1684),
.Y(n_1727)
);

INVxp67_ASAP7_75t_L g1728 ( 
.A(n_1687),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1687),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1684),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1689),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1681),
.B(n_1642),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1684),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1700),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1700),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1697),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1697),
.Y(n_1737)
);

OAI21xp33_ASAP7_75t_L g1738 ( 
.A1(n_1701),
.A2(n_1628),
.B(n_1652),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1685),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1681),
.B(n_1637),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1698),
.B(n_1543),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1674),
.B(n_1585),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1685),
.Y(n_1743)
);

INVx1_ASAP7_75t_SL g1744 ( 
.A(n_1698),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1669),
.B(n_1586),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1693),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1686),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1693),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1706),
.B(n_1694),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1715),
.B(n_1689),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1716),
.Y(n_1751)
);

INVx1_ASAP7_75t_SL g1752 ( 
.A(n_1708),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1713),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1706),
.B(n_1712),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1729),
.B(n_1671),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1725),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1724),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1724),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1716),
.Y(n_1759)
);

NAND2x1p5_ASAP7_75t_L g1760 ( 
.A(n_1708),
.B(n_1705),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1717),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1731),
.B(n_1702),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1720),
.B(n_1702),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1712),
.B(n_1694),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1745),
.B(n_1694),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1727),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1740),
.B(n_1701),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1717),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1747),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1747),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1745),
.B(n_1705),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1734),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1711),
.B(n_1699),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1745),
.B(n_1695),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1735),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1742),
.B(n_1695),
.Y(n_1776)
);

OR2x6_ASAP7_75t_L g1777 ( 
.A(n_1722),
.B(n_1626),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1723),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1727),
.Y(n_1779)
);

NAND2x1p5_ASAP7_75t_L g1780 ( 
.A(n_1722),
.B(n_1705),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1730),
.Y(n_1781)
);

NAND2x2_ASAP7_75t_L g1782 ( 
.A(n_1721),
.B(n_1610),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1742),
.B(n_1695),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1723),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1728),
.B(n_1699),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1709),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1707),
.B(n_1699),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1732),
.B(n_1703),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1707),
.B(n_1690),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1709),
.Y(n_1790)
);

OR2x6_ASAP7_75t_L g1791 ( 
.A(n_1719),
.B(n_1654),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1714),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1736),
.B(n_1702),
.Y(n_1793)
);

BUFx3_ASAP7_75t_L g1794 ( 
.A(n_1710),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1771),
.B(n_1707),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1751),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1755),
.B(n_1737),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1752),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1794),
.B(n_1741),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1751),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1754),
.B(n_1718),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1759),
.Y(n_1802)
);

BUFx2_ASAP7_75t_L g1803 ( 
.A(n_1760),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1759),
.Y(n_1804)
);

BUFx2_ASAP7_75t_L g1805 ( 
.A(n_1760),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1754),
.B(n_1718),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1761),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1762),
.Y(n_1808)
);

NAND2xp33_ASAP7_75t_SL g1809 ( 
.A(n_1750),
.B(n_1628),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1764),
.B(n_1718),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1767),
.B(n_1744),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1777),
.A2(n_1738),
.B1(n_1625),
.B2(n_1691),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1761),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1794),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1791),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1784),
.B(n_1739),
.Y(n_1816)
);

AND2x4_ASAP7_75t_L g1817 ( 
.A(n_1771),
.B(n_1726),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1768),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1760),
.Y(n_1819)
);

INVx1_ASAP7_75t_SL g1820 ( 
.A(n_1791),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1791),
.B(n_1610),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1768),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_1791),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1784),
.B(n_1773),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1778),
.B(n_1743),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1762),
.Y(n_1826)
);

NAND3xp33_ASAP7_75t_L g1827 ( 
.A(n_1777),
.B(n_1688),
.C(n_1632),
.Y(n_1827)
);

INVx1_ASAP7_75t_SL g1828 ( 
.A(n_1763),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_L g1829 ( 
.A(n_1777),
.B(n_1610),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1764),
.B(n_1726),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1753),
.Y(n_1831)
);

OAI32xp33_ASAP7_75t_L g1832 ( 
.A1(n_1827),
.A2(n_1780),
.A3(n_1809),
.B1(n_1815),
.B2(n_1820),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1814),
.B(n_1777),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1796),
.Y(n_1834)
);

INVx1_ASAP7_75t_SL g1835 ( 
.A(n_1823),
.Y(n_1835)
);

INVx2_ASAP7_75t_SL g1836 ( 
.A(n_1801),
.Y(n_1836)
);

OAI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1798),
.A2(n_1780),
.B1(n_1782),
.B2(n_1785),
.Y(n_1837)
);

AOI31xp33_ASAP7_75t_L g1838 ( 
.A1(n_1821),
.A2(n_1780),
.A3(n_1536),
.B(n_1517),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1812),
.A2(n_1775),
.B(n_1772),
.Y(n_1839)
);

AOI221xp5_ASAP7_75t_L g1840 ( 
.A1(n_1828),
.A2(n_1786),
.B1(n_1792),
.B2(n_1790),
.C(n_1775),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1826),
.B(n_1808),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1829),
.A2(n_1782),
.B1(n_1790),
.B2(n_1786),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1799),
.A2(n_1772),
.B(n_1763),
.Y(n_1843)
);

AOI322xp5_ASAP7_75t_L g1844 ( 
.A1(n_1811),
.A2(n_1749),
.A3(n_1704),
.B1(n_1691),
.B2(n_1690),
.C1(n_1789),
.C2(n_1787),
.Y(n_1844)
);

INVxp67_ASAP7_75t_SL g1845 ( 
.A(n_1819),
.Y(n_1845)
);

OR2x6_ASAP7_75t_L g1846 ( 
.A(n_1803),
.B(n_1561),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1831),
.B(n_1749),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1796),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1800),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_R g1850 ( 
.A(n_1803),
.B(n_1574),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1824),
.B(n_1788),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1800),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1802),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1831),
.B(n_1792),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1801),
.B(n_1746),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1802),
.Y(n_1856)
);

BUFx3_ASAP7_75t_L g1857 ( 
.A(n_1805),
.Y(n_1857)
);

AOI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1817),
.A2(n_1771),
.B1(n_1705),
.B2(n_1691),
.Y(n_1858)
);

INVx2_ASAP7_75t_SL g1859 ( 
.A(n_1857),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1843),
.A2(n_1805),
.B1(n_1806),
.B2(n_1819),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1852),
.Y(n_1861)
);

INVx1_ASAP7_75t_SL g1862 ( 
.A(n_1850),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1835),
.B(n_1825),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1852),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1836),
.B(n_1806),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1841),
.B(n_1816),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1838),
.B(n_1832),
.Y(n_1867)
);

AOI221xp5_ASAP7_75t_L g1868 ( 
.A1(n_1840),
.A2(n_1813),
.B1(n_1822),
.B2(n_1818),
.C(n_1804),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1834),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1837),
.A2(n_1817),
.B1(n_1795),
.B2(n_1810),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1851),
.B(n_1810),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1846),
.B(n_1830),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1833),
.B(n_1797),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1839),
.B(n_1830),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1846),
.B(n_1797),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1846),
.B(n_1795),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1847),
.B(n_1755),
.Y(n_1877)
);

BUFx2_ASAP7_75t_L g1878 ( 
.A(n_1845),
.Y(n_1878)
);

BUFx6f_ASAP7_75t_L g1879 ( 
.A(n_1848),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1849),
.Y(n_1880)
);

AOI221xp5_ASAP7_75t_L g1881 ( 
.A1(n_1867),
.A2(n_1837),
.B1(n_1854),
.B2(n_1856),
.C(n_1853),
.Y(n_1881)
);

OAI21x1_ASAP7_75t_L g1882 ( 
.A1(n_1861),
.A2(n_1845),
.B(n_1842),
.Y(n_1882)
);

AND3x1_ASAP7_75t_L g1883 ( 
.A(n_1867),
.B(n_1858),
.C(n_1855),
.Y(n_1883)
);

AOI222xp33_ASAP7_75t_L g1884 ( 
.A1(n_1863),
.A2(n_1813),
.B1(n_1822),
.B2(n_1818),
.C1(n_1804),
.C2(n_1807),
.Y(n_1884)
);

AOI211xp5_ASAP7_75t_L g1885 ( 
.A1(n_1863),
.A2(n_1807),
.B(n_1817),
.C(n_1795),
.Y(n_1885)
);

AOI21xp33_ASAP7_75t_SL g1886 ( 
.A1(n_1859),
.A2(n_1817),
.B(n_1756),
.Y(n_1886)
);

NAND3xp33_ASAP7_75t_L g1887 ( 
.A(n_1860),
.B(n_1844),
.C(n_1758),
.Y(n_1887)
);

AOI211xp5_ASAP7_75t_L g1888 ( 
.A1(n_1875),
.A2(n_1868),
.B(n_1870),
.C(n_1862),
.Y(n_1888)
);

OAI211xp5_ASAP7_75t_L g1889 ( 
.A1(n_1860),
.A2(n_1688),
.B(n_1781),
.C(n_1766),
.Y(n_1889)
);

AOI22x1_ASAP7_75t_L g1890 ( 
.A1(n_1878),
.A2(n_1876),
.B1(n_1872),
.B2(n_1866),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1873),
.B(n_1787),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1865),
.B(n_1765),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1891),
.Y(n_1893)
);

NAND3xp33_ASAP7_75t_L g1894 ( 
.A(n_1888),
.B(n_1879),
.C(n_1864),
.Y(n_1894)
);

NOR2x1_ASAP7_75t_L g1895 ( 
.A(n_1887),
.B(n_1879),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1886),
.B(n_1871),
.Y(n_1896)
);

AOI322xp5_ASAP7_75t_L g1897 ( 
.A1(n_1881),
.A2(n_1874),
.A3(n_1873),
.B1(n_1880),
.B2(n_1869),
.C1(n_1879),
.C2(n_1704),
.Y(n_1897)
);

NAND4xp25_ASAP7_75t_L g1898 ( 
.A(n_1885),
.B(n_1877),
.C(n_1879),
.D(n_1658),
.Y(n_1898)
);

OA22x2_ASAP7_75t_L g1899 ( 
.A1(n_1882),
.A2(n_1781),
.B1(n_1757),
.B2(n_1758),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_1890),
.Y(n_1900)
);

NOR2x1_ASAP7_75t_L g1901 ( 
.A(n_1889),
.B(n_1757),
.Y(n_1901)
);

AOI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1883),
.A2(n_1892),
.B1(n_1884),
.B2(n_1705),
.Y(n_1902)
);

NAND4xp25_ASAP7_75t_L g1903 ( 
.A(n_1896),
.B(n_1897),
.C(n_1895),
.D(n_1894),
.Y(n_1903)
);

AOI21xp5_ASAP7_75t_L g1904 ( 
.A1(n_1900),
.A2(n_1884),
.B(n_1779),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1902),
.B(n_1766),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1893),
.B(n_1793),
.Y(n_1906)
);

AOI322xp5_ASAP7_75t_L g1907 ( 
.A1(n_1901),
.A2(n_1691),
.A3(n_1704),
.B1(n_1690),
.B2(n_1683),
.C1(n_1789),
.C2(n_1776),
.Y(n_1907)
);

NOR3xp33_ASAP7_75t_L g1908 ( 
.A(n_1898),
.B(n_1647),
.C(n_1779),
.Y(n_1908)
);

AOI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1903),
.A2(n_1899),
.B1(n_1765),
.B2(n_1774),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1906),
.Y(n_1910)
);

AOI31xp33_ASAP7_75t_L g1911 ( 
.A1(n_1904),
.A2(n_1774),
.A3(n_1793),
.B(n_1574),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1905),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1908),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1907),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1906),
.Y(n_1915)
);

INVx1_ASAP7_75t_SL g1916 ( 
.A(n_1912),
.Y(n_1916)
);

NOR2x1_ASAP7_75t_L g1917 ( 
.A(n_1910),
.B(n_1769),
.Y(n_1917)
);

AND3x2_ASAP7_75t_L g1918 ( 
.A(n_1915),
.B(n_1691),
.C(n_1776),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1913),
.Y(n_1919)
);

INVxp67_ASAP7_75t_SL g1920 ( 
.A(n_1909),
.Y(n_1920)
);

OAI21xp33_ASAP7_75t_L g1921 ( 
.A1(n_1914),
.A2(n_1770),
.B(n_1769),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1917),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1916),
.B(n_1911),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1919),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1922),
.Y(n_1925)
);

NAND5xp2_ASAP7_75t_L g1926 ( 
.A(n_1925),
.B(n_1920),
.C(n_1924),
.D(n_1921),
.E(n_1923),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1926),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1926),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1928),
.A2(n_1923),
.B(n_1918),
.Y(n_1929)
);

AOI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1927),
.A2(n_1730),
.B1(n_1733),
.B2(n_1770),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1929),
.A2(n_1733),
.B(n_1748),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1930),
.B(n_1783),
.Y(n_1932)
);

OAI21xp5_ASAP7_75t_SL g1933 ( 
.A1(n_1931),
.A2(n_1548),
.B(n_1546),
.Y(n_1933)
);

AOI222xp33_ASAP7_75t_L g1934 ( 
.A1(n_1933),
.A2(n_1932),
.B1(n_1783),
.B2(n_1683),
.C1(n_1670),
.C2(n_1726),
.Y(n_1934)
);

AOI221xp5_ASAP7_75t_L g1935 ( 
.A1(n_1934),
.A2(n_1670),
.B1(n_1692),
.B2(n_1680),
.C(n_1688),
.Y(n_1935)
);

AOI211xp5_ASAP7_75t_L g1936 ( 
.A1(n_1935),
.A2(n_1692),
.B(n_1660),
.C(n_1663),
.Y(n_1936)
);


endmodule