module fake_jpeg_8918_n_312 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_SL g28 ( 
.A(n_8),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_44),
.Y(n_49)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_21),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_47),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_27),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_53),
.Y(n_75)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_61),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_36),
.B1(n_30),
.B2(n_29),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_64),
.B1(n_70),
.B2(n_25),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_30),
.B1(n_31),
.B2(n_29),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_56),
.A2(n_37),
.B1(n_44),
.B2(n_48),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_30),
.B1(n_29),
.B2(n_31),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_73),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_47),
.B1(n_39),
.B2(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_21),
.B(n_20),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_24),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_17),
.B1(n_35),
.B2(n_34),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_24),
.B1(n_20),
.B2(n_35),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_47),
.A2(n_17),
.B1(n_34),
.B2(n_18),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_44),
.A2(n_18),
.B1(n_22),
.B2(n_23),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_74),
.B(n_101),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_76),
.A2(n_84),
.B1(n_88),
.B2(n_109),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_22),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_77),
.B(n_78),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_54),
.B(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_49),
.B(n_23),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_82),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_21),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_86),
.Y(n_116)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_37),
.B1(n_48),
.B2(n_32),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_94),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_74),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_66),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_96),
.Y(n_125)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_72),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_103),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_27),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_105),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_21),
.Y(n_105)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_21),
.Y(n_107)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_64),
.A2(n_43),
.B1(n_27),
.B2(n_26),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_108),
.A2(n_76),
.B1(n_103),
.B2(n_85),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_57),
.A2(n_32),
.B1(n_24),
.B2(n_26),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_43),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_3),
.Y(n_137)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_43),
.C(n_32),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_139),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_24),
.B(n_26),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_120),
.A2(n_123),
.B(n_98),
.Y(n_171)
);

AOI22x1_ASAP7_75t_SL g121 ( 
.A1(n_92),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_121),
.A2(n_99),
.B(n_7),
.Y(n_175)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_1),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_126),
.B(n_130),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_1),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_133),
.C(n_16),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_2),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_138),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_5),
.B(n_6),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_75),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_82),
.B(n_4),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_77),
.B(n_79),
.Y(n_141)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g156 ( 
.A(n_145),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_4),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_5),
.Y(n_147)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_149),
.B(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_153),
.B(n_157),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_131),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_161),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_95),
.Y(n_160)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_86),
.Y(n_162)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_165),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_143),
.A2(n_94),
.B1(n_93),
.B2(n_89),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_167),
.B1(n_127),
.B2(n_89),
.Y(n_191)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

AO22x1_ASAP7_75t_SL g167 ( 
.A1(n_121),
.A2(n_102),
.B1(n_93),
.B2(n_106),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_169),
.Y(n_208)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_134),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_170),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_173),
.B(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_172),
.A2(n_143),
.B1(n_140),
.B2(n_139),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_176),
.Y(n_195)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_177),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_117),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_186),
.C(n_207),
.Y(n_219)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_182),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_191),
.B1(n_193),
.B2(n_148),
.Y(n_215)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_185),
.B(n_189),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_135),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_123),
.Y(n_187)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_156),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_178),
.Y(n_211)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_173),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_176),
.A2(n_130),
.B1(n_126),
.B2(n_133),
.Y(n_193)
);

AND2x2_ASAP7_75t_SL g196 ( 
.A(n_150),
.B(n_123),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_196),
.A2(n_197),
.B(n_203),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_167),
.A2(n_120),
.B1(n_140),
.B2(n_146),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_151),
.A2(n_137),
.B1(n_114),
.B2(n_99),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_167),
.B1(n_151),
.B2(n_148),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_122),
.B(n_8),
.Y(n_203)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_154),
.B(n_128),
.C(n_9),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_209),
.Y(n_247)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_208),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_213),
.Y(n_248)
);

INVx13_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_194),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_216),
.B(n_220),
.Y(n_243)
);

NOR4xp25_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_150),
.C(n_149),
.D(n_158),
.Y(n_217)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_217),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_201),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_179),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_222),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_223),
.A2(n_225),
.B1(n_226),
.B2(n_229),
.Y(n_246)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_195),
.A2(n_192),
.B1(n_189),
.B2(n_200),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_186),
.B(n_159),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_197),
.B(n_207),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_203),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_177),
.C(n_128),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_196),
.C(n_187),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_236),
.C(n_238),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_230),
.B(n_223),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_235),
.B(n_6),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_232),
.C(n_180),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_193),
.C(n_188),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_188),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_245),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_209),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_240),
.Y(n_254)
);

AOI321xp33_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_227),
.A3(n_214),
.B1(n_222),
.B2(n_231),
.C(n_213),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_195),
.C(n_205),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_185),
.C(n_184),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_124),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_225),
.A2(n_198),
.B1(n_199),
.B2(n_179),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_250),
.A2(n_241),
.B1(n_245),
.B2(n_249),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_221),
.B1(n_210),
.B2(n_226),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_255),
.A2(n_256),
.B1(n_259),
.B2(n_244),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_210),
.B1(n_228),
.B2(n_231),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_240),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_260),
.Y(n_278)
);

XNOR2x1_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_235),
.Y(n_273)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_233),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_263),
.Y(n_282)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_241),
.A2(n_227),
.B(n_122),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_270),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_178),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_266),
.C(n_267),
.Y(n_276)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_246),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_117),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_258),
.B1(n_264),
.B2(n_262),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_236),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_10),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_234),
.C(n_238),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_281),
.C(n_270),
.Y(n_284)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_256),
.A2(n_239),
.B1(n_113),
.B2(n_96),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_280),
.B(n_283),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_6),
.C(n_9),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_254),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_285),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_266),
.C(n_261),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_286),
.B(n_290),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_255),
.B(n_11),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_12),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_11),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_281),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_289),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_291),
.B(n_279),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_SL g295 ( 
.A1(n_292),
.A2(n_273),
.B(n_279),
.C(n_272),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_298),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_296),
.B(n_297),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_278),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_285),
.B(n_284),
.Y(n_300)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_300),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_304),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_290),
.B(n_13),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_SL g305 ( 
.A1(n_303),
.A2(n_295),
.B(n_14),
.C(n_15),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_305),
.B(n_12),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_301),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_308),
.B(n_309),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_307),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_14),
.Y(n_312)
);


endmodule