module fake_jpeg_23941_n_264 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_264);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_227;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_48),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_1),
.C(n_2),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_22),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_58),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_29),
.B1(n_28),
.B2(n_36),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_57),
.A2(n_90),
.B1(n_27),
.B2(n_31),
.Y(n_97)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_60),
.B(n_61),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_19),
.B(n_21),
.C(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_62),
.B(n_63),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_29),
.B1(n_28),
.B2(n_32),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_65),
.A2(n_68),
.B1(n_80),
.B2(n_82),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_71),
.Y(n_116)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_37),
.B(n_26),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_75),
.Y(n_117)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_50),
.B(n_25),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_77),
.B(n_88),
.Y(n_102)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_86),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_44),
.B1(n_19),
.B2(n_21),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_26),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_30),
.B1(n_35),
.B2(n_27),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_30),
.B1(n_35),
.B2(n_27),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_84),
.A2(n_20),
.B1(n_18),
.B2(n_4),
.Y(n_114)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_47),
.A2(n_35),
.B1(n_27),
.B2(n_31),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_35),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_104),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_76),
.B(n_89),
.Y(n_127)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_106),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_66),
.B(n_67),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_68),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_34),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_34),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_109),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_34),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_31),
.B1(n_20),
.B2(n_18),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_112),
.A2(n_65),
.B1(n_55),
.B2(n_61),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_108),
.Y(n_139)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_120),
.Y(n_137)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_115),
.A2(n_71),
.B1(n_75),
.B2(n_72),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_127),
.B(n_144),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_118),
.B(n_117),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_123),
.B(n_103),
.Y(n_166)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_125),
.Y(n_153)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_132),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_136),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_91),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_53),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_135),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_91),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_140),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_141),
.Y(n_155)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_142),
.B(n_143),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_83),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_95),
.A2(n_64),
.B1(n_78),
.B2(n_59),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_98),
.Y(n_145)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_108),
.A2(n_59),
.B1(n_55),
.B2(n_62),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_146),
.A2(n_113),
.B1(n_96),
.B2(n_106),
.Y(n_156)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_147),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_83),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_99),
.Y(n_159)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_149),
.B(n_96),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_117),
.B1(n_102),
.B2(n_95),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_107),
.B(n_104),
.C(n_109),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_151),
.A2(n_159),
.B(n_127),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_157),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_156),
.B(n_126),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_134),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_169),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_102),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_171),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_172),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_99),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_132),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_166),
.B(n_120),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

AND2x6_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_99),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_SL g181 ( 
.A(n_170),
.B(n_129),
.C(n_132),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_103),
.C(n_113),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_176),
.Y(n_195)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_149),
.Y(n_184)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_148),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_191),
.C(n_182),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_184),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_181),
.A2(n_188),
.B(n_192),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_131),
.Y(n_182)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_141),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_185),
.B(n_187),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_SL g199 ( 
.A1(n_186),
.A2(n_177),
.B(n_170),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_130),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_146),
.B(n_105),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_165),
.A2(n_172),
.B1(n_152),
.B2(n_155),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_154),
.B1(n_177),
.B2(n_151),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_196),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_126),
.B(n_121),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_194),
.A2(n_192),
.B(n_183),
.Y(n_212)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_197),
.B(n_166),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_195),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_206),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_199),
.A2(n_213),
.B1(n_181),
.B2(n_189),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_208),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_194),
.A2(n_177),
.B(n_152),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_212),
.B(n_214),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_205),
.B(n_178),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_171),
.C(n_160),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_174),
.Y(n_209)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_163),
.C(n_157),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_179),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_186),
.A2(n_156),
.B1(n_169),
.B2(n_163),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_185),
.A2(n_158),
.B(n_174),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_221),
.Y(n_239)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_223),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_228),
.Y(n_231)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_213),
.A2(n_193),
.B1(n_178),
.B2(n_184),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_224),
.A2(n_204),
.B1(n_210),
.B2(n_212),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_227),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_203),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_187),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_200),
.C(n_208),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_233),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_218),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_232),
.A2(n_227),
.B1(n_222),
.B2(n_176),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_216),
.B(n_217),
.Y(n_233)
);

NOR3xp33_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_210),
.C(n_207),
.Y(n_234)
);

OAI31xp33_ASAP7_75t_L g246 ( 
.A1(n_234),
.A2(n_237),
.A3(n_197),
.B(n_235),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_207),
.C(n_196),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_235),
.B(n_236),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_225),
.B(n_173),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_238),
.A2(n_226),
.B1(n_221),
.B2(n_224),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_244),
.B1(n_246),
.B2(n_54),
.Y(n_251)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_245),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_2),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_223),
.Y(n_244)
);

AOI322xp5_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_246),
.A3(n_244),
.B1(n_241),
.B2(n_240),
.C1(n_234),
.C2(n_239),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_249),
.Y(n_254)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_243),
.A2(n_105),
.A3(n_121),
.B1(n_140),
.B2(n_145),
.C1(n_14),
.C2(n_16),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_13),
.B(n_4),
.Y(n_256)
);

AOI322xp5_ASAP7_75t_L g252 ( 
.A1(n_247),
.A2(n_145),
.A3(n_14),
.B1(n_20),
.B2(n_18),
.C1(n_54),
.C2(n_8),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_253),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_257),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_3),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_253),
.Y(n_258)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_258),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_260),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_3),
.C(n_5),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_259),
.B(n_5),
.C(n_7),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_262),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_9),
.Y(n_264)
);


endmodule