module fake_jpeg_24870_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_1),
.B(n_2),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx2_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

AO22x2_ASAP7_75t_L g16 ( 
.A1(n_13),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_16),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_10),
.A2(n_0),
.B1(n_3),
.B2(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_7),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_19),
.Y(n_29)
);

NOR3xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_15),
.C(n_12),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_10),
.A2(n_14),
.B1(n_7),
.B2(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_25),
.C(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_15),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_31),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_6),
.C(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_34),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_36),
.A2(n_16),
.B1(n_28),
.B2(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_26),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_33),
.B(n_16),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_37),
.C(n_16),
.Y(n_41)
);

XNOR2x1_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_16),
.Y(n_40)
);

OAI211xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_41),
.B(n_27),
.C(n_31),
.Y(n_43)
);

AOI322xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_29),
.A3(n_35),
.B1(n_27),
.B2(n_18),
.C1(n_23),
.C2(n_30),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_43),
.C(n_23),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_30),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_30),
.C(n_28),
.Y(n_46)
);


endmodule