module real_jpeg_7384_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g15 ( 
.A1(n_1),
.A2(n_16),
.B1(n_20),
.B2(n_25),
.Y(n_15)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_1),
.A2(n_25),
.B1(n_140),
.B2(n_143),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_2),
.A2(n_87),
.B1(n_149),
.B2(n_153),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_2),
.Y(n_153)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_3),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_4),
.A2(n_33),
.B1(n_35),
.B2(n_39),
.Y(n_32)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_5),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_6),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_7),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_7),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_7),
.A2(n_92),
.B1(n_102),
.B2(n_104),
.Y(n_101)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_8),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_8),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_9),
.B(n_54),
.C(n_59),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_9),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_9),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_9),
.A2(n_27),
.B1(n_101),
.B2(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_9),
.B(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_120),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_97),
.B(n_119),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_45),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_13),
.B(n_45),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_26),
.B1(n_31),
.B2(n_40),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_15),
.A2(n_27),
.B1(n_101),
.B2(n_105),
.Y(n_100)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_27),
.A2(n_32),
.B(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_30),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

BUFx8_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_38),
.Y(n_117)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_44),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_63),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_46),
.B(n_63),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_53),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_52),
.Y(n_131)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_52),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_52),
.Y(n_143)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_70),
.B1(n_89),
.B2(n_91),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_113),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_70),
.A2(n_89),
.B1(n_91),
.B2(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_81),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_74),
.B1(n_77),
.B2(n_79),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_130),
.B1(n_132),
.B2(n_135),
.Y(n_129)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_107),
.B(n_118),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_100),
.Y(n_118)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_155),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_124),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_145),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_138),
.B2(n_144),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_138),
.Y(n_144)
);

INVx4_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_154),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);


endmodule