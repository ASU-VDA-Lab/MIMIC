module fake_jpeg_12752_n_179 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_10),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_45),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_25),
.B(n_0),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_21),
.B(n_1),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_51),
.Y(n_72)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_53),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_3),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_55),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g55 ( 
.A(n_15),
.B(n_1),
.C(n_3),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_27),
.B(n_26),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_61),
.A2(n_68),
.B(n_75),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_16),
.B1(n_24),
.B2(n_30),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_75),
.B1(n_78),
.B2(n_66),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_33),
.A2(n_27),
.B1(n_26),
.B2(n_19),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_22),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_22),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_21),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_73),
.B(n_83),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_19),
.B1(n_24),
.B2(n_30),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_34),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_84),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_16),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_85),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_14),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_48),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_14),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_36),
.B(n_5),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_77),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_79),
.A2(n_37),
.B1(n_40),
.B2(n_7),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_88),
.B(n_96),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_85),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_94),
.Y(n_113)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_92),
.Y(n_124)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_5),
.B1(n_6),
.B2(n_40),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_100),
.B1(n_74),
.B2(n_57),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_8),
.B1(n_11),
.B2(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_11),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_103),
.Y(n_128)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_60),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_74),
.Y(n_116)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_107),
.Y(n_121)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_109),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_64),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_68),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_112),
.B(n_117),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_61),
.A3(n_68),
.B1(n_80),
.B2(n_56),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_127),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_56),
.B(n_57),
.C(n_59),
.Y(n_115)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_116),
.B(n_120),
.Y(n_143)
);

AO22x1_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_64),
.B1(n_100),
.B2(n_94),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_104),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_95),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_120),
.C(n_116),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_64),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_98),
.B1(n_107),
.B2(n_87),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_90),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_135),
.B(n_136),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_89),
.C(n_93),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_124),
.C(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_109),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_109),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_137),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_149),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_151),
.C(n_134),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_141),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_119),
.C(n_122),
.Y(n_151)
);

AOI221xp5_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_143),
.B1(n_134),
.B2(n_138),
.C(n_133),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_153),
.C(n_152),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_160),
.C(n_151),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_145),
.A2(n_138),
.B1(n_130),
.B2(n_131),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_159),
.B1(n_161),
.B2(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_143),
.A3(n_131),
.B1(n_119),
.B2(n_139),
.C1(n_117),
.C2(n_118),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_115),
.B1(n_118),
.B2(n_114),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_165),
.C(n_155),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_164),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_157),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_148),
.C(n_144),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_163),
.B(n_155),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_161),
.C(n_159),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_171),
.B(n_123),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_158),
.B(n_111),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_170),
.B(n_111),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_SL g176 ( 
.A1(n_174),
.A2(n_175),
.B(n_172),
.C(n_92),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_129),
.B(n_106),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_129),
.C(n_105),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_106),
.Y(n_179)
);


endmodule