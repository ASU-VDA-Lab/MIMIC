module fake_ibex_689_n_2106 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_403, n_357, n_88, n_412, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_407, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_199, n_410, n_308, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_385, n_414, n_118, n_378, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_408, n_119, n_361, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_393, n_297, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_2106);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_403;
input n_357;
input n_88;
input n_412;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_407;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_410;
input n_308;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_118;
input n_378;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_393;
input n_297;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;

output n_2106;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_766;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_1930;
wire n_452;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_773;
wire n_2038;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_1391;
wire n_884;
wire n_667;
wire n_850;
wire n_1971;
wire n_879;
wire n_1957;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_557;
wire n_641;
wire n_1937;
wire n_893;
wire n_527;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_2025;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_745;
wire n_447;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1936;
wire n_1717;
wire n_1609;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_1121;
wire n_693;
wire n_737;
wire n_606;
wire n_1571;
wire n_1980;
wire n_462;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2076;
wire n_974;
wire n_1036;
wire n_1831;
wire n_864;
wire n_608;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_1825;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2006;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_585;
wire n_1982;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_607;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_2094;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_2010;
wire n_1756;
wire n_2097;
wire n_1470;
wire n_2098;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_650;
wire n_1575;
wire n_1448;
wire n_2077;
wire n_517;
wire n_817;
wire n_2095;
wire n_555;
wire n_951;
wire n_2053;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1967;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_1925;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2045;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2064;
wire n_1679;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_418;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_1353;
wire n_423;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_1830;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1850;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2087;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_464;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_1725;
wire n_1135;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_826;
wire n_1976;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_804;
wire n_484;
wire n_1455;
wire n_1871;
wire n_1642;
wire n_480;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_2078;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_2067;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_1956;
wire n_681;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_2093;
wire n_786;
wire n_505;
wire n_2043;
wire n_1621;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1433;
wire n_1314;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1893;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1961;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1542;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_753;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_682;
wire n_2061;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_2083;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_2044;
wire n_755;
wire n_2091;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_714;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_2013;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_665;
wire n_1101;
wire n_2079;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_438;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_1868;
wire n_966;
wire n_2104;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2092;
wire n_566;
wire n_581;
wire n_1472;
wire n_1365;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_1916;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_519;
wire n_1843;
wire n_2030;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_2100;
wire n_1902;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;
wire n_425;

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_138),
.B(n_111),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_18),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_362),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_5),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_79),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_330),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_27),
.Y(n_423)
);

BUFx10_ASAP7_75t_L g424 ( 
.A(n_410),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_404),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_338),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_46),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_122),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_116),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_65),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_104),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_110),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_310),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_278),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_394),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_225),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_58),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_7),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_79),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_384),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_316),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_403),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_97),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_329),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_389),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_122),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_252),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_271),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_347),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_196),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_261),
.B(n_300),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_35),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_343),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_148),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_318),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_301),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_167),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_193),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_53),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_94),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_76),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_202),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_89),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_258),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_121),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_257),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_4),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_259),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_307),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_74),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_206),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_123),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_340),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_245),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_167),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_249),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_36),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_352),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_231),
.Y(n_479)
);

NOR2xp67_ASAP7_75t_L g480 ( 
.A(n_285),
.B(n_308),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_276),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_274),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_97),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g484 ( 
.A(n_243),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_293),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_327),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_385),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_96),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_157),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_110),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_302),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_26),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_234),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_407),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_17),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_216),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_236),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_231),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_313),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_261),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_163),
.Y(n_501)
);

BUFx10_ASAP7_75t_L g502 ( 
.A(n_332),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_395),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_64),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_119),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_73),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_408),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_334),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_66),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_179),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_363),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_281),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_89),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_349),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_61),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_396),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_218),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_137),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_40),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_380),
.Y(n_520)
);

BUFx5_ASAP7_75t_L g521 ( 
.A(n_127),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_341),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_402),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_416),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_4),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_182),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_93),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_115),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_82),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_156),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_314),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_61),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_328),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_135),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_350),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_381),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_373),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_10),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_392),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_118),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_270),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_353),
.Y(n_542)
);

BUFx8_ASAP7_75t_SL g543 ( 
.A(n_106),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_85),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_386),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_103),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_279),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_366),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_81),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_96),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_348),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_20),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_74),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_337),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_220),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_367),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_195),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_48),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_346),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_317),
.B(n_356),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_357),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_312),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_166),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_306),
.Y(n_564)
);

BUFx10_ASAP7_75t_L g565 ( 
.A(n_164),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_229),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_213),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_44),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_331),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_414),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_406),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_40),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_280),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_38),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_109),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_372),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_272),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_8),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_103),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_59),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_51),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_239),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_62),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_173),
.Y(n_584)
);

INVxp67_ASAP7_75t_SL g585 ( 
.A(n_275),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_183),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_68),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_185),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_365),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_354),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_125),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_203),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_124),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_265),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_99),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_319),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_169),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_45),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_415),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_283),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_120),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_185),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_178),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_196),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_390),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_351),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_33),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_177),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_80),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_374),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_181),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_320),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_88),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_240),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_200),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_19),
.Y(n_616)
);

CKINVDCx16_ASAP7_75t_R g617 ( 
.A(n_323),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_20),
.Y(n_618)
);

NOR2xp67_ASAP7_75t_L g619 ( 
.A(n_383),
.B(n_45),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_31),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_258),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_136),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_296),
.Y(n_623)
);

BUFx5_ASAP7_75t_L g624 ( 
.A(n_158),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_391),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_88),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_342),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_220),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_147),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_109),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_230),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_315),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_397),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_38),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_66),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_204),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_68),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_188),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_16),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_388),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_39),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_368),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_53),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_137),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_247),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_379),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_190),
.B(n_382),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_393),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_179),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_154),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_129),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_23),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_57),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_176),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_248),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_203),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_377),
.Y(n_657)
);

BUFx10_ASAP7_75t_L g658 ( 
.A(n_413),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_189),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_387),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_364),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_124),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_371),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_193),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_215),
.Y(n_665)
);

BUFx10_ASAP7_75t_L g666 ( 
.A(n_173),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_117),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_170),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_335),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_100),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_398),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_120),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_304),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_199),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_23),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_243),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_305),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_170),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_169),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_221),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_521),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_521),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_468),
.B(n_0),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_529),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_468),
.B(n_0),
.Y(n_685)
);

OA21x2_ASAP7_75t_L g686 ( 
.A1(n_494),
.A2(n_267),
.B(n_266),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_521),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_656),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_521),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_503),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_508),
.B(n_1),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_543),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_SL g693 ( 
.A(n_486),
.B(n_268),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_567),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_521),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_521),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_521),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_624),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_590),
.B(n_2),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_567),
.B(n_3),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_453),
.Y(n_701)
);

OA21x2_ASAP7_75t_L g702 ( 
.A1(n_494),
.A2(n_273),
.B(n_269),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_624),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_631),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_624),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_544),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_542),
.B(n_6),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_629),
.Y(n_708)
);

XNOR2x2_ASAP7_75t_L g709 ( 
.A(n_540),
.B(n_6),
.Y(n_709)
);

NOR2x1_ASAP7_75t_L g710 ( 
.A(n_619),
.B(n_7),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_453),
.Y(n_711)
);

OA21x2_ASAP7_75t_L g712 ( 
.A1(n_512),
.A2(n_282),
.B(n_277),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_453),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_678),
.B(n_8),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_423),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_SL g716 ( 
.A1(n_459),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_453),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_460),
.B(n_9),
.Y(n_718)
);

BUFx8_ASAP7_75t_L g719 ( 
.A(n_542),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_548),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_624),
.Y(n_721)
);

INVx5_ASAP7_75t_L g722 ( 
.A(n_548),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_548),
.Y(n_723)
);

AND2x2_ASAP7_75t_SL g724 ( 
.A(n_560),
.B(n_412),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_624),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_624),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_545),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_727)
);

INVx5_ASAP7_75t_L g728 ( 
.A(n_548),
.Y(n_728)
);

CKINVDCx6p67_ASAP7_75t_R g729 ( 
.A(n_617),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_624),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_SL g731 ( 
.A1(n_459),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_512),
.Y(n_732)
);

INVx5_ASAP7_75t_L g733 ( 
.A(n_642),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_474),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_474),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_492),
.Y(n_736)
);

OAI21x1_ASAP7_75t_L g737 ( 
.A1(n_514),
.A2(n_286),
.B(n_284),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_424),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_514),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_484),
.B(n_16),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_541),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_492),
.Y(n_742)
);

CKINVDCx20_ASAP7_75t_R g743 ( 
.A(n_496),
.Y(n_743)
);

OA21x2_ASAP7_75t_L g744 ( 
.A1(n_516),
.A2(n_288),
.B(n_287),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_578),
.B(n_17),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_418),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_578),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_543),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_642),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_642),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_594),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_516),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_537),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_594),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_597),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_642),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_597),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_618),
.B(n_18),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_541),
.Y(n_759)
);

OA21x2_ASAP7_75t_L g760 ( 
.A1(n_537),
.A2(n_290),
.B(n_289),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_611),
.B(n_19),
.Y(n_761)
);

XNOR2x1_ASAP7_75t_L g762 ( 
.A(n_417),
.B(n_21),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_611),
.Y(n_763)
);

BUFx12f_ASAP7_75t_L g764 ( 
.A(n_424),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_419),
.B(n_21),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_620),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_573),
.B(n_600),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_418),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_620),
.Y(n_769)
);

AOI22x1_ASAP7_75t_SL g770 ( 
.A1(n_472),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_570),
.Y(n_771)
);

OA21x2_ASAP7_75t_L g772 ( 
.A1(n_570),
.A2(n_292),
.B(n_291),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_630),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_625),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_625),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_427),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_427),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_633),
.Y(n_778)
);

INVx8_ASAP7_75t_L g779 ( 
.A(n_764),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_718),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_718),
.Y(n_781)
);

INVx8_ASAP7_75t_L g782 ( 
.A(n_764),
.Y(n_782)
);

OAI21xp33_ASAP7_75t_SL g783 ( 
.A1(n_724),
.A2(n_421),
.B(n_420),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_684),
.A2(n_473),
.B1(n_478),
.B2(n_441),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_767),
.B(n_433),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_L g786 ( 
.A(n_767),
.B(n_433),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_746),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_687),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_738),
.B(n_445),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_687),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_695),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_685),
.B(n_633),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_695),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_724),
.A2(n_429),
.B1(n_431),
.B2(n_430),
.Y(n_794)
);

NAND2xp33_ASAP7_75t_L g795 ( 
.A(n_767),
.B(n_434),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_718),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_R g797 ( 
.A(n_740),
.B(n_692),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_729),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_698),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_767),
.Y(n_800)
);

NAND3xp33_ASAP7_75t_L g801 ( 
.A(n_691),
.B(n_699),
.C(n_707),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_698),
.Y(n_802)
);

INVx1_ASAP7_75t_SL g803 ( 
.A(n_706),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_777),
.Y(n_804)
);

INVx4_ASAP7_75t_L g805 ( 
.A(n_767),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_767),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_685),
.B(n_422),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_703),
.Y(n_808)
);

INVxp33_ASAP7_75t_L g809 ( 
.A(n_708),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_703),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_690),
.B(n_431),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_685),
.B(n_425),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_705),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_745),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_745),
.Y(n_815)
);

NAND2xp33_ASAP7_75t_L g816 ( 
.A(n_767),
.B(n_434),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_706),
.B(n_691),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_721),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_761),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_685),
.B(n_426),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_730),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_724),
.B(n_435),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_730),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_719),
.B(n_449),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_699),
.A2(n_439),
.B1(n_443),
.B2(n_436),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_759),
.Y(n_826)
);

NAND2xp33_ASAP7_75t_L g827 ( 
.A(n_681),
.B(n_440),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_681),
.B(n_442),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_682),
.B(n_444),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_759),
.Y(n_830)
);

NAND2xp33_ASAP7_75t_L g831 ( 
.A(n_682),
.B(n_440),
.Y(n_831)
);

INVxp67_ASAP7_75t_SL g832 ( 
.A(n_694),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_761),
.A2(n_432),
.B1(n_437),
.B2(n_428),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_683),
.Y(n_834)
);

INVxp67_ASAP7_75t_SL g835 ( 
.A(n_694),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_759),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_759),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_700),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_700),
.Y(n_839)
);

INVx1_ASAP7_75t_SL g840 ( 
.A(n_715),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_689),
.B(n_448),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_689),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_700),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_694),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_701),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_696),
.Y(n_846)
);

OAI22xp33_ASAP7_75t_SL g847 ( 
.A1(n_727),
.A2(n_443),
.B1(n_447),
.B2(n_446),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_701),
.Y(n_848)
);

NOR2x1p5_ASAP7_75t_L g849 ( 
.A(n_692),
.B(n_447),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_732),
.A2(n_454),
.B1(n_462),
.B2(n_438),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_697),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_704),
.B(n_637),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_719),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_704),
.B(n_565),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_725),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_748),
.B(n_565),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_743),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_726),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_726),
.Y(n_859)
);

AND3x2_ASAP7_75t_L g860 ( 
.A(n_693),
.B(n_585),
.C(n_465),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_741),
.B(n_455),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_778),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_739),
.Y(n_863)
);

OAI22xp33_ASAP7_75t_SL g864 ( 
.A1(n_688),
.A2(n_452),
.B1(n_457),
.B2(n_450),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_739),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_752),
.A2(n_464),
.B1(n_470),
.B2(n_467),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_747),
.B(n_450),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_686),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_753),
.Y(n_869)
);

INVx4_ASAP7_75t_L g870 ( 
.A(n_686),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_701),
.Y(n_871)
);

AND2x6_ASAP7_75t_L g872 ( 
.A(n_710),
.B(n_573),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_771),
.B(n_456),
.Y(n_873)
);

OAI22xp33_ASAP7_75t_L g874 ( 
.A1(n_768),
.A2(n_452),
.B1(n_458),
.B2(n_457),
.Y(n_874)
);

BUFx10_ASAP7_75t_L g875 ( 
.A(n_748),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_734),
.B(n_485),
.Y(n_876)
);

AND2x6_ASAP7_75t_L g877 ( 
.A(n_710),
.B(n_600),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_747),
.B(n_458),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_771),
.Y(n_879)
);

INVxp67_ASAP7_75t_SL g880 ( 
.A(n_714),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_774),
.B(n_507),
.Y(n_881)
);

BUFx10_ASAP7_75t_L g882 ( 
.A(n_765),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_778),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_775),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_775),
.Y(n_885)
);

NAND2xp33_ASAP7_75t_SL g886 ( 
.A(n_758),
.B(n_441),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_751),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_701),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_701),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_722),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_751),
.Y(n_891)
);

NAND3xp33_ASAP7_75t_L g892 ( 
.A(n_686),
.B(n_463),
.C(n_461),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_734),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_773),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_711),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_711),
.Y(n_896)
);

OAI21xp33_ASAP7_75t_SL g897 ( 
.A1(n_737),
.A2(n_476),
.B(n_475),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_773),
.B(n_565),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_735),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_770),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_735),
.A2(n_488),
.B1(n_489),
.B2(n_483),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_736),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_736),
.A2(n_495),
.B1(n_500),
.B2(n_493),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_762),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_742),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_742),
.Y(n_906)
);

AND3x2_ASAP7_75t_L g907 ( 
.A(n_709),
.B(n_506),
.C(n_505),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_722),
.B(n_523),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_754),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_754),
.B(n_463),
.Y(n_910)
);

AND3x2_ASAP7_75t_L g911 ( 
.A(n_709),
.B(n_518),
.C(n_513),
.Y(n_911)
);

NAND3xp33_ASAP7_75t_L g912 ( 
.A(n_686),
.B(n_471),
.C(n_466),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_762),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_770),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_722),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_711),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_755),
.A2(n_530),
.B1(n_534),
.B2(n_528),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_711),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_755),
.B(n_466),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_716),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_711),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_757),
.B(n_471),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_763),
.B(n_666),
.Y(n_923)
);

INVxp33_ASAP7_75t_L g924 ( 
.A(n_766),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_769),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_713),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_769),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_702),
.Y(n_928)
);

OAI22xp33_ASAP7_75t_L g929 ( 
.A1(n_776),
.A2(n_532),
.B1(n_626),
.B2(n_526),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_713),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_805),
.B(n_524),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_880),
.B(n_469),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_852),
.Y(n_933)
);

INVx8_ASAP7_75t_L g934 ( 
.A(n_779),
.Y(n_934)
);

NOR3xp33_ASAP7_75t_L g935 ( 
.A(n_847),
.B(n_731),
.C(n_586),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_822),
.A2(n_549),
.B1(n_550),
.B2(n_538),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_779),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_854),
.B(n_531),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_844),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_782),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_924),
.B(n_923),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_789),
.B(n_502),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_789),
.B(n_502),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_801),
.B(n_502),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_832),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_809),
.B(n_666),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_835),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_783),
.A2(n_737),
.B(n_553),
.C(n_557),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_811),
.B(n_612),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_SL g950 ( 
.A(n_853),
.B(n_473),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_898),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_882),
.B(n_658),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_782),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_887),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_882),
.B(n_824),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_893),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_839),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_824),
.B(n_658),
.Y(n_958)
);

OAI21xp33_ASAP7_75t_L g959 ( 
.A1(n_833),
.A2(n_919),
.B(n_910),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_817),
.B(n_632),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_780),
.A2(n_568),
.B1(n_572),
.B2(n_552),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_839),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_922),
.B(n_867),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_899),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_902),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_905),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_878),
.B(n_660),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_787),
.B(n_482),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_906),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_804),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_SL g971 ( 
.A1(n_920),
.A2(n_472),
.B1(n_479),
.B2(n_477),
.Y(n_971)
);

AND2x4_ASAP7_75t_SL g972 ( 
.A(n_875),
.B(n_482),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_814),
.B(n_487),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_794),
.A2(n_809),
.B1(n_825),
.B2(n_874),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_909),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_815),
.B(n_491),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_800),
.B(n_499),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_784),
.B(n_526),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_875),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_856),
.B(n_532),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_819),
.B(n_511),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_SL g982 ( 
.A(n_806),
.B(n_564),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_925),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_807),
.B(n_533),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_834),
.B(n_522),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_840),
.B(n_626),
.Y(n_986)
);

AND2x6_ASAP7_75t_SL g987 ( 
.A(n_900),
.B(n_574),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_927),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_875),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_798),
.B(n_628),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_838),
.B(n_547),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_863),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_843),
.B(n_559),
.Y(n_993)
);

AND2x6_ASAP7_75t_SL g994 ( 
.A(n_914),
.B(n_575),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_860),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_857),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_781),
.B(n_589),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_865),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_812),
.B(n_535),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_796),
.B(n_596),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_827),
.B(n_831),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_812),
.B(n_536),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_820),
.B(n_539),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_901),
.B(n_671),
.Y(n_1004)
);

AND2x6_ASAP7_75t_L g1005 ( 
.A(n_876),
.B(n_640),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_879),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_849),
.B(n_628),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_891),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_901),
.B(n_673),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_792),
.B(n_551),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_903),
.A2(n_577),
.B1(n_564),
.B2(n_639),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_861),
.B(n_639),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_792),
.B(n_554),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_872),
.B(n_641),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_797),
.Y(n_1015)
);

NOR2xp67_ASAP7_75t_L g1016 ( 
.A(n_894),
.B(n_645),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_862),
.B(n_556),
.Y(n_1017)
);

NOR3xp33_ASAP7_75t_L g1018 ( 
.A(n_864),
.B(n_929),
.C(n_886),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_869),
.B(n_561),
.Y(n_1019)
);

AND2x2_ASAP7_75t_SL g1020 ( 
.A(n_785),
.B(n_702),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_883),
.B(n_562),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_884),
.B(n_569),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_885),
.B(n_571),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_873),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_876),
.B(n_828),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_903),
.B(n_481),
.Y(n_1026)
);

NAND2xp33_ASAP7_75t_L g1027 ( 
.A(n_892),
.B(n_576),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_877),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_917),
.B(n_651),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_877),
.B(n_651),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_877),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_826),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_873),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_830),
.Y(n_1034)
);

CKINVDCx8_ASAP7_75t_R g1035 ( 
.A(n_904),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_897),
.B(n_599),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_886),
.A2(n_577),
.B1(n_659),
.B2(n_654),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_868),
.B(n_605),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_881),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_868),
.B(n_870),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_870),
.B(n_606),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_850),
.B(n_654),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_881),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_785),
.A2(n_712),
.B(n_702),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_866),
.B(n_662),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_917),
.B(n_520),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_829),
.B(n_610),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_866),
.B(n_829),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_841),
.B(n_667),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_913),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_786),
.A2(n_580),
.B1(n_581),
.B2(n_579),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_836),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_795),
.A2(n_584),
.B1(n_587),
.B2(n_583),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_907),
.B(n_490),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_855),
.B(n_497),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_837),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_858),
.B(n_498),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_859),
.B(n_501),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_842),
.B(n_504),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_837),
.Y(n_1060)
);

NOR2xp67_ASAP7_75t_SL g1061 ( 
.A(n_795),
.B(n_712),
.Y(n_1061)
);

BUFx5_ASAP7_75t_L g1062 ( 
.A(n_890),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_842),
.B(n_623),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_911),
.B(n_563),
.Y(n_1064)
);

NOR2xp67_ASAP7_75t_SL g1065 ( 
.A(n_816),
.B(n_712),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_846),
.B(n_627),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_851),
.B(n_510),
.Y(n_1067)
);

INVx5_ASAP7_75t_L g1068 ( 
.A(n_890),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_851),
.A2(n_592),
.B(n_593),
.C(n_591),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_908),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_908),
.B(n_646),
.Y(n_1071)
);

INVx8_ASAP7_75t_L g1072 ( 
.A(n_816),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_788),
.B(n_648),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_920),
.A2(n_517),
.B1(n_519),
.B2(n_515),
.Y(n_1074)
);

O2A1O1Ixp5_ASAP7_75t_L g1075 ( 
.A1(n_790),
.A2(n_661),
.B(n_669),
.C(n_657),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_791),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_791),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_793),
.B(n_525),
.Y(n_1078)
);

OAI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_799),
.A2(n_479),
.B1(n_509),
.B2(n_477),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_802),
.B(n_555),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_808),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_808),
.B(n_677),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_810),
.Y(n_1083)
);

AND2x6_ASAP7_75t_SL g1084 ( 
.A(n_845),
.B(n_598),
.Y(n_1084)
);

AND2x6_ASAP7_75t_SL g1085 ( 
.A(n_845),
.B(n_601),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_813),
.B(n_566),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_818),
.B(n_821),
.Y(n_1087)
);

NOR2x1p5_ASAP7_75t_L g1088 ( 
.A(n_915),
.B(n_582),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_821),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_823),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_871),
.B(n_604),
.Y(n_1091)
);

BUFx8_ASAP7_75t_L g1092 ( 
.A(n_845),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_888),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_845),
.B(n_640),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_895),
.A2(n_615),
.B1(n_616),
.B2(n_613),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_895),
.B(n_621),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_896),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_918),
.B(n_588),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_918),
.B(n_622),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_930),
.B(n_635),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_921),
.B(n_602),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_926),
.B(n_607),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_957),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_1025),
.A2(n_636),
.B(n_643),
.C(n_638),
.Y(n_1104)
);

OAI321xp33_ASAP7_75t_L g1105 ( 
.A1(n_959),
.A2(n_655),
.A3(n_650),
.B1(n_668),
.B2(n_652),
.C(n_644),
.Y(n_1105)
);

AOI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1061),
.A2(n_760),
.B(n_744),
.Y(n_1106)
);

AOI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1065),
.A2(n_760),
.B(n_744),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1040),
.A2(n_760),
.B(n_744),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_996),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_970),
.B(n_608),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1090),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_941),
.B(n_672),
.Y(n_1112)
);

NOR3xp33_ASAP7_75t_L g1113 ( 
.A(n_1079),
.B(n_971),
.C(n_1011),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_974),
.A2(n_527),
.B1(n_546),
.B2(n_509),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1069),
.A2(n_664),
.B(n_675),
.C(n_595),
.Y(n_1115)
);

CKINVDCx10_ASAP7_75t_R g1116 ( 
.A(n_1035),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1038),
.A2(n_772),
.B(n_647),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_951),
.B(n_674),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1041),
.A2(n_451),
.B(n_480),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_978),
.B(n_527),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_968),
.B(n_546),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_962),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1041),
.A2(n_1020),
.B(n_1036),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_955),
.B(n_603),
.Y(n_1124)
);

CKINVDCx16_ASAP7_75t_R g1125 ( 
.A(n_950),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1020),
.A2(n_665),
.B(n_653),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1036),
.A2(n_679),
.B(n_665),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_1025),
.A2(n_679),
.B(n_680),
.C(n_663),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1001),
.A2(n_680),
.B(n_663),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_932),
.B(n_676),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_955),
.B(n_603),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_963),
.A2(n_889),
.B(n_848),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_SL g1133 ( 
.A(n_934),
.B(n_609),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_934),
.Y(n_1134)
);

AO32x2_ASAP7_75t_L g1135 ( 
.A1(n_1028),
.A2(n_723),
.A3(n_749),
.B1(n_720),
.B2(n_717),
.Y(n_1135)
);

NOR3xp33_ASAP7_75t_L g1136 ( 
.A(n_1079),
.B(n_614),
.C(n_609),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1048),
.A2(n_634),
.B(n_614),
.C(n_558),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_945),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_947),
.Y(n_1139)
);

OR2x6_ASAP7_75t_SL g1140 ( 
.A(n_1050),
.B(n_634),
.Y(n_1140)
);

NAND2x1p5_ASAP7_75t_L g1141 ( 
.A(n_979),
.B(n_558),
.Y(n_1141)
);

NAND2x1p5_ASAP7_75t_L g1142 ( 
.A(n_989),
.B(n_649),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1027),
.A2(n_733),
.B(n_728),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_1092),
.Y(n_1144)
);

NOR2x1_ASAP7_75t_R g1145 ( 
.A(n_968),
.B(n_670),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_964),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_936),
.B(n_1029),
.Y(n_1147)
);

NAND3xp33_ASAP7_75t_L g1148 ( 
.A(n_1018),
.B(n_670),
.C(n_733),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_980),
.B(n_29),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_931),
.A2(n_733),
.B(n_889),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_934),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1018),
.A2(n_720),
.B1(n_723),
.B2(n_717),
.Y(n_1152)
);

AO21x1_ASAP7_75t_L g1153 ( 
.A1(n_1066),
.A2(n_720),
.B(n_717),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_SL g1154 ( 
.A(n_935),
.B(n_30),
.C(n_31),
.Y(n_1154)
);

INVxp67_ASAP7_75t_SL g1155 ( 
.A(n_982),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_966),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_969),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_972),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_960),
.B(n_32),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1068),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1075),
.A2(n_916),
.B(n_749),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_946),
.B(n_33),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_975),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1037),
.B(n_34),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_938),
.B(n_952),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_SL g1166 ( 
.A1(n_1094),
.A2(n_295),
.B(n_297),
.C(n_294),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_1084),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1087),
.A2(n_750),
.B(n_723),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_995),
.B(n_750),
.Y(n_1169)
);

O2A1O1Ixp5_ASAP7_75t_L g1170 ( 
.A1(n_958),
.A2(n_299),
.B(n_303),
.C(n_298),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_SL g1171 ( 
.A(n_937),
.B(n_750),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1010),
.A2(n_756),
.B(n_36),
.C(n_35),
.Y(n_1172)
);

BUFx4f_ASAP7_75t_L g1173 ( 
.A(n_940),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1051),
.A2(n_756),
.B1(n_42),
.B2(n_37),
.Y(n_1174)
);

AO21x1_ASAP7_75t_L g1175 ( 
.A1(n_1066),
.A2(n_756),
.B(n_41),
.Y(n_1175)
);

BUFx12f_ASAP7_75t_L g1176 ( 
.A(n_953),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1059),
.A2(n_1067),
.B(n_1057),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_986),
.Y(n_1178)
);

AOI221xp5_ASAP7_75t_L g1179 ( 
.A1(n_961),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.C(n_44),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_958),
.B(n_43),
.Y(n_1180)
);

AOI221xp5_ASAP7_75t_L g1181 ( 
.A1(n_935),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.C(n_50),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_990),
.Y(n_1182)
);

OAI22x1_ASAP7_75t_L g1183 ( 
.A1(n_1015),
.A2(n_54),
.B1(n_51),
.B2(n_52),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1042),
.A2(n_55),
.B(n_52),
.C(n_54),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_1074),
.B(n_56),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1012),
.B(n_942),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_988),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_944),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_942),
.B(n_59),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_1088),
.Y(n_1190)
);

INVx1_ASAP7_75t_SL g1191 ( 
.A(n_1085),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_997),
.A2(n_311),
.B(n_309),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_943),
.B(n_60),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1053),
.A2(n_63),
.B1(n_60),
.B2(n_62),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1007),
.B(n_65),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1015),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1013),
.A2(n_70),
.B(n_67),
.C(n_69),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1068),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_SL g1199 ( 
.A(n_1092),
.B(n_71),
.Y(n_1199)
);

OAI22x1_ASAP7_75t_L g1200 ( 
.A1(n_1064),
.A2(n_1054),
.B1(n_1046),
.B2(n_1026),
.Y(n_1200)
);

CKINVDCx10_ASAP7_75t_R g1201 ( 
.A(n_987),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1053),
.A2(n_75),
.B1(n_72),
.B2(n_73),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1068),
.Y(n_1203)
);

INVxp67_ASAP7_75t_L g1204 ( 
.A(n_967),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1016),
.B(n_77),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1068),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1045),
.A2(n_80),
.B1(n_77),
.B2(n_78),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_933),
.A2(n_84),
.B1(n_81),
.B2(n_83),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1091),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_SL g1210 ( 
.A(n_1031),
.B(n_83),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1000),
.A2(n_322),
.B(n_321),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_984),
.B(n_84),
.Y(n_1212)
);

BUFx8_ASAP7_75t_L g1213 ( 
.A(n_1008),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1055),
.A2(n_411),
.B(n_325),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1058),
.A2(n_326),
.B(n_324),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_991),
.B(n_86),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1078),
.A2(n_336),
.B(n_333),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1004),
.A2(n_91),
.B(n_87),
.C(n_90),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_949),
.B(n_92),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1009),
.A2(n_98),
.B(n_93),
.C(n_95),
.Y(n_1220)
);

OR2x6_ASAP7_75t_L g1221 ( 
.A(n_1072),
.B(n_101),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1091),
.Y(n_1222)
);

O2A1O1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1049),
.A2(n_105),
.B(n_102),
.C(n_104),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_999),
.B(n_105),
.Y(n_1224)
);

OR2x6_ASAP7_75t_SL g1225 ( 
.A(n_1014),
.B(n_106),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1080),
.A2(n_409),
.B(n_339),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_956),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_965),
.A2(n_112),
.B1(n_107),
.B2(n_108),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1002),
.B(n_112),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_985),
.A2(n_345),
.B(n_344),
.Y(n_1230)
);

INVx6_ASAP7_75t_SL g1231 ( 
.A(n_994),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1002),
.B(n_113),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_983),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1003),
.B(n_114),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_939),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1003),
.B(n_116),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1086),
.Y(n_1237)
);

BUFx12f_ASAP7_75t_L g1238 ( 
.A(n_1005),
.Y(n_1238)
);

AO22x1_ASAP7_75t_L g1239 ( 
.A1(n_1005),
.A2(n_1030),
.B1(n_1033),
.B2(n_1024),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_992),
.B(n_121),
.Y(n_1240)
);

BUFx4f_ASAP7_75t_L g1241 ( 
.A(n_1005),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_998),
.B(n_125),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1005),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_1243)
);

AOI33xp33_ASAP7_75t_L g1244 ( 
.A1(n_1095),
.A2(n_126),
.A3(n_128),
.B1(n_129),
.B2(n_130),
.B3(n_131),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1047),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1006),
.B(n_132),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1017),
.B(n_133),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1062),
.Y(n_1248)
);

AND2x4_ASAP7_75t_SL g1249 ( 
.A(n_954),
.B(n_134),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1076),
.A2(n_405),
.B(n_358),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1077),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1017),
.B(n_139),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1019),
.B(n_140),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_993),
.A2(n_359),
.B(n_355),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1072),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1083),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_973),
.A2(n_361),
.B(n_360),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1021),
.B(n_141),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_976),
.A2(n_141),
.B(n_142),
.C(n_143),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1021),
.B(n_144),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_981),
.A2(n_401),
.B(n_370),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1022),
.B(n_144),
.Y(n_1262)
);

AOI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1022),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1023),
.B(n_146),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1063),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1073),
.A2(n_148),
.B(n_149),
.C(n_150),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1081),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1062),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1039),
.B(n_151),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1043),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1089),
.A2(n_375),
.B(n_369),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1062),
.B(n_153),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1071),
.B(n_155),
.Y(n_1273)
);

O2A1O1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1082),
.A2(n_155),
.B(n_156),
.C(n_157),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_R g1275 ( 
.A(n_1070),
.B(n_1071),
.Y(n_1275)
);

OR2x6_ASAP7_75t_L g1276 ( 
.A(n_977),
.B(n_159),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1056),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1096),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1099),
.B(n_161),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1098),
.B(n_163),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1099),
.B(n_164),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1101),
.B(n_165),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1102),
.A2(n_400),
.B(n_399),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1100),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1106),
.A2(n_1032),
.B(n_1034),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1107),
.A2(n_1060),
.B(n_1052),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1138),
.Y(n_1287)
);

BUFx12f_ASAP7_75t_L g1288 ( 
.A(n_1158),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1153),
.A2(n_1097),
.A3(n_1093),
.B(n_175),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_1116),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1139),
.Y(n_1291)
);

OR2x2_ASAP7_75t_L g1292 ( 
.A(n_1109),
.B(n_174),
.Y(n_1292)
);

NOR2xp67_ASAP7_75t_L g1293 ( 
.A(n_1144),
.B(n_174),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1113),
.B(n_175),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1146),
.B(n_176),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_SL g1296 ( 
.A(n_1133),
.B(n_1199),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1156),
.B(n_1157),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1120),
.B(n_180),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1151),
.Y(n_1299)
);

CKINVDCx20_ASAP7_75t_R g1300 ( 
.A(n_1125),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1163),
.Y(n_1301)
);

A2O1A1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1177),
.A2(n_181),
.B(n_182),
.C(n_184),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1175),
.A2(n_184),
.A3(n_186),
.B(n_187),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1164),
.A2(n_186),
.B1(n_187),
.B2(n_190),
.Y(n_1304)
);

INVx8_ASAP7_75t_L g1305 ( 
.A(n_1176),
.Y(n_1305)
);

AO32x2_ASAP7_75t_L g1306 ( 
.A1(n_1207),
.A2(n_191),
.A3(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_1306)
);

AOI21xp33_ASAP7_75t_L g1307 ( 
.A1(n_1145),
.A2(n_194),
.B(n_197),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1241),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1123),
.A2(n_378),
.B(n_376),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1140),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1126),
.A2(n_198),
.B(n_201),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1187),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1132),
.A2(n_205),
.B(n_207),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1231),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1240),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1237),
.B(n_208),
.Y(n_1316)
);

AO31x2_ASAP7_75t_L g1317 ( 
.A1(n_1129),
.A2(n_209),
.A3(n_210),
.B(n_211),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1241),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_1318)
);

NAND3xp33_ASAP7_75t_SL g1319 ( 
.A(n_1181),
.B(n_217),
.C(n_218),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1251),
.Y(n_1320)
);

INVxp67_ASAP7_75t_L g1321 ( 
.A(n_1178),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1165),
.B(n_219),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1117),
.A2(n_222),
.B(n_223),
.Y(n_1323)
);

INVx4_ASAP7_75t_L g1324 ( 
.A(n_1221),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1231),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_1191),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1235),
.B(n_224),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1104),
.B(n_226),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1221),
.Y(n_1329)
);

NOR2x1_ASAP7_75t_SL g1330 ( 
.A(n_1221),
.B(n_227),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1127),
.A2(n_228),
.B(n_229),
.C(n_232),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1173),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_1160),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1167),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1129),
.A2(n_233),
.B(n_235),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1195),
.B(n_237),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_1249),
.Y(n_1337)
);

AO21x2_ASAP7_75t_L g1338 ( 
.A1(n_1161),
.A2(n_1152),
.B(n_1168),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1255),
.B(n_238),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1173),
.Y(n_1340)
);

OA21x2_ASAP7_75t_L g1341 ( 
.A1(n_1271),
.A2(n_240),
.B(n_241),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1209),
.A2(n_241),
.B1(n_242),
.B2(n_244),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1114),
.B(n_242),
.Y(n_1343)
);

OAI22x1_ASAP7_75t_L g1344 ( 
.A1(n_1121),
.A2(n_1205),
.B1(n_1124),
.B2(n_1131),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1248),
.B(n_244),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1136),
.B(n_246),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1182),
.B(n_250),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1222),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1112),
.B(n_251),
.Y(n_1349)
);

BUFx4f_ASAP7_75t_L g1350 ( 
.A(n_1276),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1149),
.B(n_1196),
.Y(n_1351)
);

AO21x2_ASAP7_75t_L g1352 ( 
.A1(n_1119),
.A2(n_255),
.B(n_256),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1227),
.Y(n_1353)
);

O2A1O1Ixp33_ASAP7_75t_L g1354 ( 
.A1(n_1128),
.A2(n_259),
.B(n_260),
.C(n_262),
.Y(n_1354)
);

A2O1A1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1127),
.A2(n_262),
.B(n_263),
.C(n_264),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1233),
.Y(n_1356)
);

A2O1A1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1184),
.A2(n_263),
.B(n_264),
.C(n_265),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1256),
.Y(n_1358)
);

O2A1O1Ixp5_ASAP7_75t_L g1359 ( 
.A1(n_1170),
.A2(n_1239),
.B(n_1261),
.C(n_1257),
.Y(n_1359)
);

BUFx4_ASAP7_75t_SL g1360 ( 
.A(n_1276),
.Y(n_1360)
);

BUFx10_ASAP7_75t_L g1361 ( 
.A(n_1205),
.Y(n_1361)
);

A2O1A1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1223),
.A2(n_1259),
.B(n_1218),
.C(n_1220),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1201),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1198),
.Y(n_1364)
);

NOR3xp33_ASAP7_75t_SL g1365 ( 
.A(n_1154),
.B(n_1181),
.C(n_1194),
.Y(n_1365)
);

OR2x6_ASAP7_75t_L g1366 ( 
.A(n_1238),
.B(n_1190),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1118),
.B(n_1162),
.Y(n_1367)
);

OA21x2_ASAP7_75t_L g1368 ( 
.A1(n_1283),
.A2(n_1226),
.B(n_1217),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1213),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_1213),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1130),
.B(n_1185),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1253),
.B(n_1200),
.Y(n_1372)
);

NOR2x1_ASAP7_75t_SL g1373 ( 
.A(n_1255),
.B(n_1276),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_SL g1374 ( 
.A1(n_1137),
.A2(n_1179),
.B(n_1263),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1214),
.A2(n_1215),
.B(n_1250),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1250),
.A2(n_1215),
.B(n_1214),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1103),
.B(n_1122),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1219),
.A2(n_1266),
.B(n_1274),
.C(n_1179),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_SL g1379 ( 
.A1(n_1141),
.A2(n_1142),
.B(n_1155),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1150),
.A2(n_1159),
.B(n_1273),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1242),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1150),
.A2(n_1189),
.B(n_1193),
.Y(n_1382)
);

AOI221xp5_ASAP7_75t_L g1383 ( 
.A1(n_1115),
.A2(n_1105),
.B1(n_1110),
.B2(n_1202),
.C(n_1216),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1246),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1277),
.A2(n_1192),
.B(n_1211),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1277),
.A2(n_1254),
.B(n_1230),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1268),
.B(n_1210),
.Y(n_1387)
);

NOR2xp67_ASAP7_75t_SL g1388 ( 
.A(n_1255),
.B(n_1203),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1141),
.Y(n_1389)
);

INVx5_ASAP7_75t_L g1390 ( 
.A(n_1203),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1143),
.A2(n_1269),
.B(n_1169),
.Y(n_1391)
);

BUFx6f_ASAP7_75t_L g1392 ( 
.A(n_1203),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1206),
.Y(n_1393)
);

A2O1A1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1172),
.A2(n_1197),
.B(n_1282),
.C(n_1280),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1247),
.A2(n_1260),
.B(n_1262),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1265),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1252),
.A2(n_1258),
.B(n_1264),
.Y(n_1397)
);

OR2x6_ASAP7_75t_SL g1398 ( 
.A(n_1208),
.B(n_1270),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1206),
.Y(n_1399)
);

OAI21xp33_ASAP7_75t_SL g1400 ( 
.A1(n_1279),
.A2(n_1281),
.B(n_1243),
.Y(n_1400)
);

AO31x2_ASAP7_75t_L g1401 ( 
.A1(n_1183),
.A2(n_1284),
.A3(n_1228),
.B(n_1174),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1212),
.A2(n_1236),
.B(n_1234),
.Y(n_1402)
);

CKINVDCx11_ASAP7_75t_R g1403 ( 
.A(n_1225),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1224),
.A2(n_1229),
.B(n_1232),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1135),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1111),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1135),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1135),
.Y(n_1408)
);

AO31x2_ASAP7_75t_L g1409 ( 
.A1(n_1166),
.A2(n_1278),
.A3(n_1188),
.B(n_1245),
.Y(n_1409)
);

BUFx10_ASAP7_75t_L g1410 ( 
.A(n_1171),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1275),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1204),
.B(n_941),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1204),
.B(n_941),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1251),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1221),
.A2(n_1145),
.B(n_948),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1138),
.Y(n_1416)
);

NAND3xp33_ASAP7_75t_L g1417 ( 
.A(n_1148),
.B(n_955),
.C(n_1180),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1204),
.B(n_941),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1133),
.A2(n_784),
.B1(n_1011),
.B2(n_1109),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1204),
.B(n_941),
.Y(n_1420)
);

AOI211x1_ASAP7_75t_L g1421 ( 
.A1(n_1154),
.A2(n_822),
.B(n_1147),
.C(n_959),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1109),
.Y(n_1422)
);

INVx3_ASAP7_75t_SL g1423 ( 
.A(n_1158),
.Y(n_1423)
);

O2A1O1Ixp5_ASAP7_75t_L g1424 ( 
.A1(n_1175),
.A2(n_1153),
.B(n_1036),
.C(n_1272),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1204),
.B(n_941),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1109),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1204),
.B(n_941),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1138),
.Y(n_1428)
);

CKINVDCx6p67_ASAP7_75t_R g1429 ( 
.A(n_1116),
.Y(n_1429)
);

CKINVDCx11_ASAP7_75t_R g1430 ( 
.A(n_1140),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1109),
.Y(n_1431)
);

NOR2xp67_ASAP7_75t_SL g1432 ( 
.A(n_1134),
.B(n_1151),
.Y(n_1432)
);

NOR2x1_ASAP7_75t_SL g1433 ( 
.A(n_1221),
.B(n_1238),
.Y(n_1433)
);

AO31x2_ASAP7_75t_L g1434 ( 
.A1(n_1153),
.A2(n_1175),
.A3(n_1126),
.B(n_948),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1204),
.B(n_974),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1251),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1177),
.A2(n_1040),
.B(n_912),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_SL g1438 ( 
.A(n_1248),
.B(n_1267),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1116),
.Y(n_1439)
);

NAND3xp33_ASAP7_75t_L g1440 ( 
.A(n_1148),
.B(n_955),
.C(n_1180),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1204),
.B(n_941),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1108),
.A2(n_1040),
.B(n_1044),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1177),
.A2(n_1040),
.B(n_912),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1204),
.B(n_941),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1109),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1248),
.B(n_1267),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1251),
.Y(n_1447)
);

BUFx10_ASAP7_75t_L g1448 ( 
.A(n_1158),
.Y(n_1448)
);

AO31x2_ASAP7_75t_L g1449 ( 
.A1(n_1153),
.A2(n_1175),
.A3(n_1126),
.B(n_948),
.Y(n_1449)
);

OAI22x1_ASAP7_75t_L g1450 ( 
.A1(n_1167),
.A2(n_968),
.B1(n_1109),
.B2(n_1191),
.Y(n_1450)
);

A2O1A1Ixp33_ASAP7_75t_L g1451 ( 
.A1(n_1177),
.A2(n_1126),
.B(n_783),
.C(n_1244),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1116),
.Y(n_1452)
);

AOI21xp33_ASAP7_75t_L g1453 ( 
.A1(n_1145),
.A2(n_797),
.B(n_1124),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_SL g1454 ( 
.A(n_1248),
.B(n_1267),
.Y(n_1454)
);

A2O1A1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1177),
.A2(n_1126),
.B(n_783),
.C(n_1244),
.Y(n_1455)
);

AO31x2_ASAP7_75t_L g1456 ( 
.A1(n_1153),
.A2(n_1175),
.A3(n_1126),
.B(n_948),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1109),
.B(n_803),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1251),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1204),
.B(n_941),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1204),
.B(n_941),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1109),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1133),
.A2(n_784),
.B1(n_1011),
.B2(n_1109),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1248),
.B(n_1267),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1138),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1138),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1138),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_SL g1467 ( 
.A(n_1133),
.B(n_934),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1221),
.A2(n_1145),
.B(n_948),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1109),
.B(n_803),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1204),
.B(n_941),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1204),
.B(n_974),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1204),
.B(n_974),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1109),
.B(n_803),
.Y(n_1473)
);

AOI221xp5_ASAP7_75t_L g1474 ( 
.A1(n_1113),
.A2(n_1018),
.B1(n_847),
.B2(n_1114),
.C(n_1079),
.Y(n_1474)
);

NOR2x1_ASAP7_75t_L g1475 ( 
.A(n_1134),
.B(n_1144),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1138),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_1134),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1147),
.A2(n_822),
.B1(n_794),
.B2(n_1241),
.Y(n_1478)
);

AO32x2_ASAP7_75t_L g1479 ( 
.A1(n_1207),
.A2(n_868),
.A3(n_870),
.B1(n_928),
.B2(n_1284),
.Y(n_1479)
);

AND2x6_ASAP7_75t_L g1480 ( 
.A(n_1255),
.B(n_1144),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1109),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1138),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1109),
.B(n_803),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1109),
.B(n_803),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1147),
.A2(n_822),
.B1(n_794),
.B2(n_1241),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1177),
.A2(n_1126),
.B(n_783),
.C(n_1244),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1116),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1138),
.Y(n_1488)
);

NOR2xp67_ASAP7_75t_L g1489 ( 
.A(n_1144),
.B(n_784),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1109),
.B(n_803),
.Y(n_1490)
);

OAI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1177),
.A2(n_1040),
.B(n_912),
.Y(n_1491)
);

INVx6_ASAP7_75t_SL g1492 ( 
.A(n_1221),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1138),
.Y(n_1493)
);

AO31x2_ASAP7_75t_L g1494 ( 
.A1(n_1153),
.A2(n_1175),
.A3(n_1126),
.B(n_948),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1435),
.B(n_1471),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_SL g1496 ( 
.A1(n_1373),
.A2(n_1433),
.B(n_1330),
.Y(n_1496)
);

BUFx12f_ASAP7_75t_L g1497 ( 
.A(n_1290),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1287),
.Y(n_1498)
);

AO31x2_ASAP7_75t_L g1499 ( 
.A1(n_1451),
.A2(n_1486),
.A3(n_1455),
.B(n_1442),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_SL g1500 ( 
.A(n_1290),
.B(n_1452),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1291),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1320),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1416),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1402),
.A2(n_1404),
.B(n_1397),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1324),
.B(n_1390),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1435),
.B(n_1471),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1390),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1324),
.B(n_1390),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1390),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1472),
.B(n_1371),
.Y(n_1510)
);

NAND2x1_ASAP7_75t_L g1511 ( 
.A(n_1388),
.B(n_1379),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1472),
.B(n_1474),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1376),
.A2(n_1285),
.B(n_1286),
.Y(n_1513)
);

CKINVDCx11_ASAP7_75t_R g1514 ( 
.A(n_1305),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1371),
.B(n_1419),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1414),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1412),
.B(n_1413),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1378),
.A2(n_1394),
.B(n_1362),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1385),
.A2(n_1386),
.B(n_1359),
.Y(n_1519)
);

NAND2x1p5_ASAP7_75t_L g1520 ( 
.A(n_1350),
.B(n_1432),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1378),
.A2(n_1394),
.B(n_1362),
.Y(n_1521)
);

INVx2_ASAP7_75t_SL g1522 ( 
.A(n_1305),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1411),
.B(n_1301),
.Y(n_1523)
);

OAI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1367),
.A2(n_1322),
.B(n_1424),
.Y(n_1524)
);

OA21x2_ASAP7_75t_L g1525 ( 
.A1(n_1405),
.A2(n_1408),
.B(n_1407),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1428),
.Y(n_1526)
);

OR2x6_ASAP7_75t_L g1527 ( 
.A(n_1305),
.B(n_1369),
.Y(n_1527)
);

NAND3xp33_ASAP7_75t_L g1528 ( 
.A(n_1421),
.B(n_1302),
.C(n_1357),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1464),
.Y(n_1529)
);

INVx6_ASAP7_75t_L g1530 ( 
.A(n_1448),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1465),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1312),
.B(n_1466),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1418),
.B(n_1420),
.Y(n_1533)
);

AOI22x1_ASAP7_75t_L g1534 ( 
.A1(n_1344),
.A2(n_1389),
.B1(n_1309),
.B2(n_1313),
.Y(n_1534)
);

O2A1O1Ixp5_ASAP7_75t_L g1535 ( 
.A1(n_1387),
.A2(n_1350),
.B(n_1443),
.C(n_1437),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1462),
.B(n_1425),
.Y(n_1536)
);

CKINVDCx16_ASAP7_75t_R g1537 ( 
.A(n_1467),
.Y(n_1537)
);

NAND2x1p5_ASAP7_75t_L g1538 ( 
.A(n_1399),
.B(n_1431),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1476),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1482),
.B(n_1488),
.Y(n_1540)
);

BUFx8_ASAP7_75t_L g1541 ( 
.A(n_1288),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_SL g1542 ( 
.A1(n_1296),
.A2(n_1329),
.B1(n_1310),
.B2(n_1316),
.Y(n_1542)
);

AO21x2_ASAP7_75t_L g1543 ( 
.A1(n_1311),
.A2(n_1338),
.B(n_1491),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1427),
.B(n_1441),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1493),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1368),
.A2(n_1375),
.B(n_1391),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1353),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1445),
.Y(n_1548)
);

INVx4_ASAP7_75t_L g1549 ( 
.A(n_1370),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1473),
.B(n_1484),
.Y(n_1550)
);

BUFx2_ASAP7_75t_SL g1551 ( 
.A(n_1448),
.Y(n_1551)
);

OAI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1367),
.A2(n_1322),
.B(n_1417),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1329),
.B(n_1381),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1356),
.Y(n_1554)
);

NAND2x1p5_ASAP7_75t_L g1555 ( 
.A(n_1422),
.B(n_1426),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1490),
.B(n_1444),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1297),
.Y(n_1557)
);

AO21x2_ASAP7_75t_L g1558 ( 
.A1(n_1338),
.A2(n_1335),
.B(n_1372),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1459),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1460),
.B(n_1470),
.Y(n_1560)
);

BUFx2_ASAP7_75t_R g1561 ( 
.A(n_1452),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1384),
.B(n_1436),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1457),
.B(n_1469),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1480),
.Y(n_1564)
);

INVx8_ASAP7_75t_L g1565 ( 
.A(n_1480),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1445),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1447),
.B(n_1458),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1440),
.A2(n_1374),
.B(n_1400),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1447),
.B(n_1458),
.Y(n_1569)
);

OR2x6_ASAP7_75t_L g1570 ( 
.A(n_1461),
.B(n_1481),
.Y(n_1570)
);

AND2x4_ASAP7_75t_SL g1571 ( 
.A(n_1361),
.B(n_1483),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1377),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1321),
.B(n_1299),
.Y(n_1573)
);

BUFx4f_ASAP7_75t_SL g1574 ( 
.A(n_1429),
.Y(n_1574)
);

OAI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1438),
.A2(n_1454),
.B(n_1446),
.Y(n_1575)
);

OAI21x1_ASAP7_75t_L g1576 ( 
.A1(n_1454),
.A2(n_1463),
.B(n_1341),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1319),
.A2(n_1294),
.B1(n_1343),
.B2(n_1403),
.Y(n_1577)
);

A2O1A1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1354),
.A2(n_1365),
.B(n_1319),
.C(n_1331),
.Y(n_1578)
);

BUFx12f_ASAP7_75t_L g1579 ( 
.A(n_1439),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1321),
.B(n_1453),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1360),
.Y(n_1581)
);

AO21x2_ASAP7_75t_L g1582 ( 
.A1(n_1352),
.A2(n_1365),
.B(n_1355),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1358),
.Y(n_1583)
);

INVx8_ASAP7_75t_L g1584 ( 
.A(n_1480),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1298),
.B(n_1346),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1316),
.B(n_1347),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1360),
.Y(n_1587)
);

OAI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1349),
.A2(n_1478),
.B(n_1485),
.Y(n_1588)
);

OR2x6_ASAP7_75t_L g1589 ( 
.A(n_1415),
.B(n_1468),
.Y(n_1589)
);

OR2x6_ASAP7_75t_L g1590 ( 
.A(n_1288),
.B(n_1366),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1295),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1327),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1315),
.B(n_1347),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1334),
.B(n_1292),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1396),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1489),
.B(n_1349),
.Y(n_1596)
);

A2O1A1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1383),
.A2(n_1328),
.B(n_1304),
.C(n_1307),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1406),
.Y(n_1598)
);

AO21x2_ASAP7_75t_L g1599 ( 
.A1(n_1352),
.A2(n_1336),
.B(n_1351),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1337),
.Y(n_1600)
);

OAI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1406),
.A2(n_1293),
.B(n_1342),
.Y(n_1601)
);

OAI21x1_ASAP7_75t_L g1602 ( 
.A1(n_1308),
.A2(n_1318),
.B(n_1393),
.Y(n_1602)
);

NOR2xp67_ASAP7_75t_L g1603 ( 
.A(n_1314),
.B(n_1325),
.Y(n_1603)
);

NOR2x1_ASAP7_75t_R g1604 ( 
.A(n_1430),
.B(n_1487),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_SL g1605 ( 
.A1(n_1492),
.A2(n_1304),
.B(n_1348),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1333),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1317),
.Y(n_1607)
);

OR2x6_ASAP7_75t_L g1608 ( 
.A(n_1366),
.B(n_1340),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1317),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1434),
.A2(n_1494),
.B(n_1456),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1475),
.A2(n_1332),
.B(n_1477),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1317),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1434),
.A2(n_1494),
.B(n_1456),
.Y(n_1613)
);

OA21x2_ASAP7_75t_L g1614 ( 
.A1(n_1289),
.A2(n_1494),
.B(n_1449),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1434),
.A2(n_1494),
.B(n_1456),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1434),
.Y(n_1616)
);

OA21x2_ASAP7_75t_L g1617 ( 
.A1(n_1289),
.A2(n_1449),
.B(n_1456),
.Y(n_1617)
);

BUFx8_ASAP7_75t_L g1618 ( 
.A(n_1306),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1317),
.Y(n_1619)
);

OAI21x1_ASAP7_75t_L g1620 ( 
.A1(n_1449),
.A2(n_1289),
.B(n_1479),
.Y(n_1620)
);

AO21x2_ASAP7_75t_L g1621 ( 
.A1(n_1289),
.A2(n_1449),
.B(n_1479),
.Y(n_1621)
);

OAI21x1_ASAP7_75t_L g1622 ( 
.A1(n_1479),
.A2(n_1410),
.B(n_1303),
.Y(n_1622)
);

OA21x2_ASAP7_75t_L g1623 ( 
.A1(n_1479),
.A2(n_1303),
.B(n_1409),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_SL g1624 ( 
.A1(n_1492),
.A2(n_1398),
.B(n_1361),
.Y(n_1624)
);

BUFx4_ASAP7_75t_R g1625 ( 
.A(n_1492),
.Y(n_1625)
);

OA21x2_ASAP7_75t_L g1626 ( 
.A1(n_1409),
.A2(n_1306),
.B(n_1401),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1306),
.Y(n_1627)
);

AO21x2_ASAP7_75t_L g1628 ( 
.A1(n_1409),
.A2(n_1401),
.B(n_1306),
.Y(n_1628)
);

OAI21x1_ASAP7_75t_L g1629 ( 
.A1(n_1364),
.A2(n_1392),
.B(n_1401),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1450),
.B(n_1326),
.Y(n_1630)
);

OAI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1392),
.A2(n_1403),
.B(n_1423),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1392),
.A2(n_1310),
.B(n_1300),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1430),
.Y(n_1633)
);

INVx3_ASAP7_75t_L g1634 ( 
.A(n_1423),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1300),
.Y(n_1635)
);

INVx4_ASAP7_75t_SL g1636 ( 
.A(n_1363),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1305),
.Y(n_1637)
);

OAI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1378),
.A2(n_783),
.B(n_1186),
.Y(n_1638)
);

OAI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1378),
.A2(n_783),
.B(n_1186),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1435),
.B(n_1471),
.Y(n_1640)
);

NAND2x1p5_ASAP7_75t_L g1641 ( 
.A(n_1390),
.B(n_1144),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1390),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1402),
.A2(n_1404),
.B(n_1397),
.Y(n_1643)
);

AOI22x1_ASAP7_75t_L g1644 ( 
.A1(n_1382),
.A2(n_1200),
.B1(n_1380),
.B2(n_1395),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1435),
.B(n_1471),
.Y(n_1645)
);

AO21x1_ASAP7_75t_L g1646 ( 
.A1(n_1345),
.A2(n_1323),
.B(n_1339),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1287),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1287),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1474),
.A2(n_1113),
.B1(n_1471),
.B2(n_1435),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1390),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1287),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1435),
.B(n_1471),
.Y(n_1652)
);

INVx5_ASAP7_75t_L g1653 ( 
.A(n_1480),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1350),
.A2(n_1419),
.B1(n_1462),
.B2(n_1221),
.Y(n_1654)
);

OAI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1378),
.A2(n_783),
.B(n_1186),
.Y(n_1655)
);

NAND3xp33_ASAP7_75t_L g1656 ( 
.A(n_1421),
.B(n_1302),
.C(n_1357),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1431),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_SL g1658 ( 
.A1(n_1373),
.A2(n_1433),
.B(n_1330),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1435),
.B(n_1471),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_SL g1660 ( 
.A1(n_1373),
.A2(n_1433),
.B(n_1330),
.Y(n_1660)
);

OAI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1378),
.A2(n_783),
.B(n_1186),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1324),
.B(n_1433),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1287),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_SL g1664 ( 
.A(n_1350),
.B(n_1387),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1287),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_1565),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1589),
.B(n_1567),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1583),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1502),
.Y(n_1669)
);

AO21x1_ASAP7_75t_SL g1670 ( 
.A1(n_1606),
.A2(n_1568),
.B(n_1521),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1567),
.B(n_1569),
.Y(n_1671)
);

CKINVDCx20_ASAP7_75t_R g1672 ( 
.A(n_1514),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1567),
.B(n_1569),
.Y(n_1673)
);

INVxp67_ASAP7_75t_L g1674 ( 
.A(n_1560),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1559),
.Y(n_1675)
);

INVx2_ASAP7_75t_SL g1676 ( 
.A(n_1565),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1595),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1569),
.B(n_1516),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1560),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_1653),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1498),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1583),
.B(n_1550),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1659),
.B(n_1517),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1606),
.Y(n_1684)
);

BUFx3_ASAP7_75t_L g1685 ( 
.A(n_1514),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1501),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1503),
.Y(n_1687)
);

BUFx3_ASAP7_75t_L g1688 ( 
.A(n_1509),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1570),
.Y(n_1689)
);

INVx2_ASAP7_75t_SL g1690 ( 
.A(n_1565),
.Y(n_1690)
);

INVx6_ASAP7_75t_L g1691 ( 
.A(n_1653),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1570),
.Y(n_1692)
);

INVxp67_ASAP7_75t_SL g1693 ( 
.A(n_1548),
.Y(n_1693)
);

INVx2_ASAP7_75t_SL g1694 ( 
.A(n_1584),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_SL g1695 ( 
.A1(n_1578),
.A2(n_1589),
.B(n_1654),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1556),
.B(n_1512),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1570),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1548),
.B(n_1566),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1566),
.B(n_1495),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1664),
.B(n_1505),
.Y(n_1700)
);

INVx4_ASAP7_75t_L g1701 ( 
.A(n_1584),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1563),
.Y(n_1702)
);

BUFx8_ASAP7_75t_L g1703 ( 
.A(n_1497),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1525),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1562),
.B(n_1557),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1562),
.B(n_1572),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1526),
.Y(n_1707)
);

OR2x6_ASAP7_75t_L g1708 ( 
.A(n_1584),
.B(n_1624),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1529),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1531),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1562),
.B(n_1649),
.Y(n_1711)
);

BUFx3_ASAP7_75t_L g1712 ( 
.A(n_1509),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1539),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1659),
.B(n_1533),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1573),
.Y(n_1715)
);

INVx3_ASAP7_75t_L g1716 ( 
.A(n_1650),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1657),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1545),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1649),
.B(n_1532),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1607),
.Y(n_1720)
);

BUFx4f_ASAP7_75t_SL g1721 ( 
.A(n_1541),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1544),
.B(n_1506),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1647),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1640),
.B(n_1645),
.Y(n_1724)
);

CKINVDCx12_ASAP7_75t_R g1725 ( 
.A(n_1527),
.Y(n_1725)
);

AO21x2_ASAP7_75t_L g1726 ( 
.A1(n_1504),
.A2(n_1643),
.B(n_1546),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1652),
.B(n_1510),
.Y(n_1727)
);

CKINVDCx20_ASAP7_75t_R g1728 ( 
.A(n_1541),
.Y(n_1728)
);

AO21x2_ASAP7_75t_L g1729 ( 
.A1(n_1518),
.A2(n_1519),
.B(n_1622),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1532),
.B(n_1540),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1510),
.B(n_1536),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1515),
.B(n_1577),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1648),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1651),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1532),
.B(n_1540),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1540),
.B(n_1515),
.Y(n_1736)
);

BUFx12f_ASAP7_75t_L g1737 ( 
.A(n_1541),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1638),
.B(n_1639),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1663),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1551),
.Y(n_1740)
);

INVx1_ASAP7_75t_SL g1741 ( 
.A(n_1571),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1665),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1547),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1555),
.Y(n_1744)
);

OR2x6_ASAP7_75t_L g1745 ( 
.A(n_1496),
.B(n_1658),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1554),
.Y(n_1746)
);

AO21x2_ASAP7_75t_L g1747 ( 
.A1(n_1513),
.A2(n_1620),
.B(n_1612),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1598),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1628),
.B(n_1626),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1555),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1577),
.B(n_1585),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_SL g1752 ( 
.A(n_1561),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_SL g1753 ( 
.A(n_1604),
.B(n_1500),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1523),
.Y(n_1754)
);

AO21x2_ASAP7_75t_L g1755 ( 
.A1(n_1620),
.A2(n_1619),
.B(n_1609),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_1530),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1655),
.B(n_1661),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1553),
.Y(n_1758)
);

OAI21xp33_ASAP7_75t_SL g1759 ( 
.A1(n_1664),
.A2(n_1602),
.B(n_1524),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1552),
.B(n_1553),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1626),
.B(n_1591),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1520),
.Y(n_1762)
);

BUFx2_ASAP7_75t_L g1763 ( 
.A(n_1629),
.Y(n_1763)
);

BUFx4f_ASAP7_75t_SL g1764 ( 
.A(n_1497),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1586),
.B(n_1593),
.Y(n_1765)
);

AO31x2_ASAP7_75t_L g1766 ( 
.A1(n_1616),
.A2(n_1646),
.A3(n_1627),
.B(n_1578),
.Y(n_1766)
);

BUFx2_ASAP7_75t_L g1767 ( 
.A(n_1618),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1626),
.B(n_1610),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1592),
.B(n_1582),
.Y(n_1769)
);

AO21x1_ASAP7_75t_SL g1770 ( 
.A1(n_1588),
.A2(n_1601),
.B(n_1511),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1520),
.Y(n_1771)
);

INVx2_ASAP7_75t_SL g1772 ( 
.A(n_1745),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1704),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1720),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1667),
.B(n_1575),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1698),
.B(n_1610),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1675),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_1745),
.Y(n_1778)
);

INVxp67_ASAP7_75t_SL g1779 ( 
.A(n_1693),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1731),
.B(n_1580),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1732),
.A2(n_1605),
.B1(n_1618),
.B2(n_1580),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1761),
.B(n_1613),
.Y(n_1782)
);

NOR2x1_ASAP7_75t_L g1783 ( 
.A(n_1728),
.B(n_1590),
.Y(n_1783)
);

BUFx3_ASAP7_75t_L g1784 ( 
.A(n_1688),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1696),
.B(n_1542),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1769),
.B(n_1615),
.Y(n_1786)
);

INVxp67_ASAP7_75t_L g1787 ( 
.A(n_1702),
.Y(n_1787)
);

BUFx2_ASAP7_75t_L g1788 ( 
.A(n_1684),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1769),
.B(n_1615),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1678),
.B(n_1623),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1698),
.B(n_1614),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1677),
.Y(n_1792)
);

NOR2x1_ASAP7_75t_SL g1793 ( 
.A(n_1745),
.B(n_1564),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1682),
.B(n_1614),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1682),
.B(n_1614),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1696),
.B(n_1635),
.Y(n_1796)
);

OR2x6_ASAP7_75t_L g1797 ( 
.A(n_1695),
.B(n_1631),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1681),
.Y(n_1798)
);

INVx1_ASAP7_75t_SL g1799 ( 
.A(n_1672),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1668),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1738),
.B(n_1623),
.Y(n_1801)
);

BUFx3_ASAP7_75t_L g1802 ( 
.A(n_1688),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1683),
.B(n_1635),
.Y(n_1803)
);

AOI21xp33_ASAP7_75t_L g1804 ( 
.A1(n_1759),
.A2(n_1596),
.B(n_1599),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1686),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1699),
.B(n_1617),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1738),
.B(n_1757),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1714),
.B(n_1594),
.Y(n_1808)
);

INVx2_ASAP7_75t_SL g1809 ( 
.A(n_1745),
.Y(n_1809)
);

BUFx3_ASAP7_75t_L g1810 ( 
.A(n_1712),
.Y(n_1810)
);

BUFx3_ASAP7_75t_L g1811 ( 
.A(n_1712),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1687),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1757),
.B(n_1617),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1671),
.B(n_1617),
.Y(n_1814)
);

OAI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1727),
.A2(n_1674),
.B1(n_1679),
.B2(n_1630),
.C(n_1722),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1719),
.A2(n_1618),
.B1(n_1633),
.B2(n_1581),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1724),
.B(n_1662),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1673),
.B(n_1621),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1724),
.B(n_1662),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1707),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1699),
.B(n_1662),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1736),
.B(n_1621),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_1737),
.Y(n_1823)
);

INVxp67_ASAP7_75t_L g1824 ( 
.A(n_1717),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1751),
.B(n_1600),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1705),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1736),
.B(n_1558),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1709),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1710),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1719),
.B(n_1582),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1713),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1718),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1711),
.B(n_1706),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1723),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1711),
.B(n_1543),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1715),
.Y(n_1836)
);

AND2x4_ASAP7_75t_L g1837 ( 
.A(n_1667),
.B(n_1575),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1765),
.B(n_1538),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1733),
.B(n_1597),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1734),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1739),
.B(n_1742),
.Y(n_1841)
);

NOR2x1_ASAP7_75t_SL g1842 ( 
.A(n_1708),
.B(n_1770),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1743),
.B(n_1537),
.Y(n_1843)
);

HB1xp67_ASAP7_75t_L g1844 ( 
.A(n_1744),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1746),
.B(n_1599),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1762),
.B(n_1522),
.Y(n_1846)
);

INVx2_ASAP7_75t_SL g1847 ( 
.A(n_1691),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1669),
.B(n_1499),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1748),
.Y(n_1849)
);

BUFx2_ASAP7_75t_L g1850 ( 
.A(n_1767),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1771),
.B(n_1637),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1760),
.B(n_1499),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1708),
.B(n_1576),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1814),
.B(n_1766),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1774),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1774),
.Y(n_1856)
);

INVx1_ASAP7_75t_SL g1857 ( 
.A(n_1799),
.Y(n_1857)
);

AOI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1785),
.A2(n_1760),
.B1(n_1753),
.B2(n_1735),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1773),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1779),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1807),
.B(n_1730),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1814),
.B(n_1766),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1806),
.B(n_1768),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1777),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1792),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1806),
.B(n_1794),
.Y(n_1866)
);

HB1xp67_ASAP7_75t_L g1867 ( 
.A(n_1800),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1822),
.B(n_1766),
.Y(n_1868)
);

BUFx2_ASAP7_75t_L g1869 ( 
.A(n_1850),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1822),
.B(n_1766),
.Y(n_1870)
);

INVx3_ASAP7_75t_L g1871 ( 
.A(n_1778),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1807),
.B(n_1766),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1796),
.B(n_1689),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1813),
.B(n_1768),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1787),
.B(n_1692),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1813),
.B(n_1755),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1788),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1818),
.B(n_1755),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1836),
.B(n_1697),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1780),
.B(n_1758),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1794),
.B(n_1749),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1818),
.B(n_1755),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1823),
.B(n_1549),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1795),
.B(n_1749),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1849),
.B(n_1826),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1782),
.B(n_1729),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1782),
.B(n_1729),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1798),
.Y(n_1888)
);

INVxp67_ASAP7_75t_L g1889 ( 
.A(n_1844),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1786),
.B(n_1789),
.Y(n_1890)
);

NAND2x1p5_ASAP7_75t_L g1891 ( 
.A(n_1784),
.B(n_1680),
.Y(n_1891)
);

AOI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1825),
.A2(n_1725),
.B1(n_1737),
.B2(n_1700),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1805),
.B(n_1812),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1788),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1786),
.B(n_1729),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1789),
.B(n_1747),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_1823),
.B(n_1549),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1827),
.B(n_1747),
.Y(n_1898)
);

AND2x4_ASAP7_75t_L g1899 ( 
.A(n_1775),
.B(n_1837),
.Y(n_1899)
);

BUFx4_ASAP7_75t_SL g1900 ( 
.A(n_1784),
.Y(n_1900)
);

INVx1_ASAP7_75t_SL g1901 ( 
.A(n_1802),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1820),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1795),
.B(n_1726),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1827),
.B(n_1747),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1830),
.B(n_1670),
.Y(n_1905)
);

INVxp33_ASAP7_75t_L g1906 ( 
.A(n_1783),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1830),
.B(n_1835),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1775),
.B(n_1763),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1866),
.B(n_1791),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1859),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1866),
.B(n_1791),
.Y(n_1911)
);

OAI21xp5_ASAP7_75t_SL g1912 ( 
.A1(n_1906),
.A2(n_1850),
.B(n_1740),
.Y(n_1912)
);

INVx2_ASAP7_75t_SL g1913 ( 
.A(n_1900),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1899),
.B(n_1853),
.Y(n_1914)
);

NAND2x1p5_ASAP7_75t_L g1915 ( 
.A(n_1901),
.B(n_1802),
.Y(n_1915)
);

NOR2x1p5_ASAP7_75t_L g1916 ( 
.A(n_1871),
.B(n_1810),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1855),
.Y(n_1917)
);

INVx1_ASAP7_75t_SL g1918 ( 
.A(n_1869),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1855),
.Y(n_1919)
);

AND2x4_ASAP7_75t_L g1920 ( 
.A(n_1899),
.B(n_1853),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1860),
.Y(n_1921)
);

NAND2x1p5_ASAP7_75t_L g1922 ( 
.A(n_1869),
.B(n_1810),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1890),
.B(n_1801),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1856),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1863),
.B(n_1776),
.Y(n_1925)
);

OR3x2_ASAP7_75t_L g1926 ( 
.A(n_1863),
.B(n_1721),
.C(n_1752),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1857),
.B(n_1685),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1872),
.B(n_1801),
.Y(n_1928)
);

INVx1_ASAP7_75t_SL g1929 ( 
.A(n_1877),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1890),
.B(n_1835),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1856),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1874),
.B(n_1896),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1874),
.B(n_1790),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1872),
.B(n_1848),
.Y(n_1934)
);

INVxp67_ASAP7_75t_SL g1935 ( 
.A(n_1894),
.Y(n_1935)
);

NOR3x1_ASAP7_75t_L g1936 ( 
.A(n_1879),
.B(n_1587),
.C(n_1631),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1896),
.B(n_1790),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1867),
.B(n_1833),
.Y(n_1938)
);

INVx2_ASAP7_75t_SL g1939 ( 
.A(n_1891),
.Y(n_1939)
);

AOI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1926),
.A2(n_1858),
.B1(n_1815),
.B2(n_1781),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1921),
.Y(n_1941)
);

INVx1_ASAP7_75t_SL g1942 ( 
.A(n_1913),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1925),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1910),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1910),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1925),
.Y(n_1946)
);

INVx2_ASAP7_75t_SL g1947 ( 
.A(n_1916),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1909),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1932),
.B(n_1886),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1909),
.B(n_1881),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1911),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1930),
.B(n_1907),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1911),
.B(n_1881),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1917),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1917),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1919),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1932),
.B(n_1886),
.Y(n_1957)
);

OAI22xp33_ASAP7_75t_L g1958 ( 
.A1(n_1912),
.A2(n_1797),
.B1(n_1892),
.B2(n_1891),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1930),
.B(n_1907),
.Y(n_1959)
);

OR2x2_ASAP7_75t_SL g1960 ( 
.A(n_1926),
.B(n_1884),
.Y(n_1960)
);

OR2x2_ASAP7_75t_L g1961 ( 
.A(n_1928),
.B(n_1884),
.Y(n_1961)
);

NAND2x1p5_ASAP7_75t_L g1962 ( 
.A(n_1916),
.B(n_1685),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_L g1963 ( 
.A(n_1912),
.B(n_1889),
.Y(n_1963)
);

AOI21xp33_ASAP7_75t_SL g1964 ( 
.A1(n_1913),
.A2(n_1897),
.B(n_1883),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1923),
.B(n_1887),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1919),
.Y(n_1966)
);

NOR2x1p5_ASAP7_75t_L g1967 ( 
.A(n_1935),
.B(n_1811),
.Y(n_1967)
);

NAND2x1_ASAP7_75t_SL g1968 ( 
.A(n_1914),
.B(n_1920),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1923),
.B(n_1887),
.Y(n_1969)
);

INVxp67_ASAP7_75t_L g1970 ( 
.A(n_1927),
.Y(n_1970)
);

NOR2xp33_ASAP7_75t_L g1971 ( 
.A(n_1929),
.B(n_1824),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1924),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1950),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1950),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1965),
.B(n_1969),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1953),
.Y(n_1976)
);

AOI21xp33_ASAP7_75t_L g1977 ( 
.A1(n_1963),
.A2(n_1958),
.B(n_1942),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1953),
.Y(n_1978)
);

AND2x4_ASAP7_75t_L g1979 ( 
.A(n_1947),
.B(n_1914),
.Y(n_1979)
);

O2A1O1Ixp33_ASAP7_75t_L g1980 ( 
.A1(n_1963),
.A2(n_1875),
.B(n_1843),
.C(n_1839),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1948),
.B(n_1929),
.Y(n_1981)
);

INVxp33_ASAP7_75t_L g1982 ( 
.A(n_1962),
.Y(n_1982)
);

OAI221xp5_ASAP7_75t_L g1983 ( 
.A1(n_1940),
.A2(n_1816),
.B1(n_1938),
.B2(n_1918),
.C(n_1922),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1951),
.B(n_1934),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1943),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1965),
.B(n_1933),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1946),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1969),
.B(n_1933),
.Y(n_1988)
);

AOI221xp5_ASAP7_75t_L g1989 ( 
.A1(n_1941),
.A2(n_1928),
.B1(n_1934),
.B2(n_1885),
.C(n_1918),
.Y(n_1989)
);

OR4x1_ASAP7_75t_L g1990 ( 
.A(n_1947),
.B(n_1939),
.C(n_1772),
.D(n_1809),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1944),
.Y(n_1991)
);

AOI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1962),
.A2(n_1842),
.B(n_1939),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1961),
.B(n_1937),
.Y(n_1993)
);

O2A1O1Ixp33_ASAP7_75t_L g1994 ( 
.A1(n_1964),
.A2(n_1590),
.B(n_1808),
.C(n_1803),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1961),
.B(n_1937),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1954),
.Y(n_1996)
);

AOI22xp5_ASAP7_75t_L g1997 ( 
.A1(n_1971),
.A2(n_1914),
.B1(n_1920),
.B2(n_1905),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1971),
.A2(n_1842),
.B(n_1793),
.Y(n_1998)
);

AOI211x1_ASAP7_75t_L g1999 ( 
.A1(n_1952),
.A2(n_1632),
.B(n_1893),
.C(n_1861),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1949),
.B(n_1868),
.Y(n_2000)
);

AOI222xp33_ASAP7_75t_L g2001 ( 
.A1(n_1970),
.A2(n_1854),
.B1(n_1862),
.B2(n_1902),
.C1(n_1864),
.C2(n_1865),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1944),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1955),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1996),
.Y(n_2004)
);

AOI221xp5_ASAP7_75t_L g2005 ( 
.A1(n_1977),
.A2(n_1888),
.B1(n_1880),
.B2(n_1959),
.C(n_1956),
.Y(n_2005)
);

NAND3xp33_ASAP7_75t_SL g2006 ( 
.A(n_1994),
.B(n_1672),
.C(n_1728),
.Y(n_2006)
);

OAI21xp33_ASAP7_75t_L g2007 ( 
.A1(n_2001),
.A2(n_1968),
.B(n_1957),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1983),
.B(n_1960),
.Y(n_2008)
);

OAI22xp33_ASAP7_75t_SL g2009 ( 
.A1(n_1997),
.A2(n_1915),
.B1(n_1922),
.B2(n_1891),
.Y(n_2009)
);

AOI21xp33_ASAP7_75t_SL g2010 ( 
.A1(n_1982),
.A2(n_1915),
.B(n_1922),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_2003),
.Y(n_2011)
);

AOI21xp5_ASAP7_75t_L g2012 ( 
.A1(n_1982),
.A2(n_1915),
.B(n_1914),
.Y(n_2012)
);

OAI21xp33_ASAP7_75t_L g2013 ( 
.A1(n_1989),
.A2(n_1957),
.B(n_1949),
.Y(n_2013)
);

OAI21xp33_ASAP7_75t_L g2014 ( 
.A1(n_1981),
.A2(n_1905),
.B(n_1920),
.Y(n_2014)
);

AOI322xp5_ASAP7_75t_L g2015 ( 
.A1(n_1973),
.A2(n_1862),
.A3(n_1854),
.B1(n_1870),
.B2(n_1868),
.C1(n_1920),
.C2(n_1833),
.Y(n_2015)
);

AOI221xp5_ASAP7_75t_L g2016 ( 
.A1(n_1999),
.A2(n_1966),
.B1(n_1972),
.B2(n_1873),
.C(n_1695),
.Y(n_2016)
);

NAND3xp33_ASAP7_75t_SL g2017 ( 
.A(n_1992),
.B(n_1936),
.C(n_1741),
.Y(n_2017)
);

AOI322xp5_ASAP7_75t_L g2018 ( 
.A1(n_1974),
.A2(n_1870),
.A3(n_1895),
.B1(n_1882),
.B2(n_1878),
.C1(n_1898),
.C2(n_1904),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1976),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1978),
.Y(n_2020)
);

AOI22xp33_ASAP7_75t_L g2021 ( 
.A1(n_1979),
.A2(n_1899),
.B1(n_1908),
.B2(n_1967),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1993),
.Y(n_2022)
);

OAI21xp33_ASAP7_75t_L g2023 ( 
.A1(n_2007),
.A2(n_1980),
.B(n_1985),
.Y(n_2023)
);

INVxp67_ASAP7_75t_SL g2024 ( 
.A(n_2012),
.Y(n_2024)
);

NAND3xp33_ASAP7_75t_L g2025 ( 
.A(n_2008),
.B(n_1703),
.C(n_1987),
.Y(n_2025)
);

AOI21xp33_ASAP7_75t_L g2026 ( 
.A1(n_2009),
.A2(n_2005),
.B(n_1703),
.Y(n_2026)
);

AOI22xp5_ASAP7_75t_L g2027 ( 
.A1(n_2006),
.A2(n_1979),
.B1(n_1984),
.B2(n_1975),
.Y(n_2027)
);

OAI211xp5_ASAP7_75t_L g2028 ( 
.A1(n_2017),
.A2(n_1998),
.B(n_1603),
.C(n_1634),
.Y(n_2028)
);

OAI32xp33_ASAP7_75t_L g2029 ( 
.A1(n_2013),
.A2(n_1995),
.A3(n_1990),
.B1(n_2000),
.B2(n_1988),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_2004),
.Y(n_2030)
);

AOI211xp5_ASAP7_75t_SL g2031 ( 
.A1(n_2005),
.A2(n_1574),
.B(n_1764),
.C(n_1979),
.Y(n_2031)
);

OAI22xp33_ASAP7_75t_SL g2032 ( 
.A1(n_2019),
.A2(n_1990),
.B1(n_2002),
.B2(n_1797),
.Y(n_2032)
);

NOR3x1_ASAP7_75t_L g2033 ( 
.A(n_2020),
.B(n_1703),
.C(n_1772),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2011),
.Y(n_2034)
);

AOI211xp5_ASAP7_75t_L g2035 ( 
.A1(n_2010),
.A2(n_1634),
.B(n_1809),
.C(n_1975),
.Y(n_2035)
);

NOR3xp33_ASAP7_75t_L g2036 ( 
.A(n_2016),
.B(n_1756),
.C(n_1846),
.Y(n_2036)
);

OAI322xp33_ASAP7_75t_L g2037 ( 
.A1(n_2022),
.A2(n_1991),
.A3(n_2002),
.B1(n_1988),
.B2(n_1903),
.C1(n_1852),
.C2(n_1986),
.Y(n_2037)
);

XNOR2xp5_ASAP7_75t_L g2038 ( 
.A(n_2021),
.B(n_1590),
.Y(n_2038)
);

NOR3xp33_ASAP7_75t_L g2039 ( 
.A(n_2014),
.B(n_1756),
.C(n_1851),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_2015),
.B(n_1991),
.Y(n_2040)
);

OAI221xp5_ASAP7_75t_L g2041 ( 
.A1(n_2018),
.A2(n_1797),
.B1(n_1527),
.B2(n_1608),
.C(n_1871),
.Y(n_2041)
);

INVxp67_ASAP7_75t_SL g2042 ( 
.A(n_2012),
.Y(n_2042)
);

NAND3xp33_ASAP7_75t_L g2043 ( 
.A(n_2008),
.B(n_1804),
.C(n_1656),
.Y(n_2043)
);

AOI211x1_ASAP7_75t_L g2044 ( 
.A1(n_2029),
.A2(n_1611),
.B(n_1936),
.C(n_1841),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_2026),
.B(n_1574),
.Y(n_2045)
);

AOI221xp5_ASAP7_75t_L g2046 ( 
.A1(n_2026),
.A2(n_1831),
.B1(n_1832),
.B2(n_1829),
.C(n_1828),
.Y(n_2046)
);

NAND3xp33_ASAP7_75t_L g2047 ( 
.A(n_2024),
.B(n_1527),
.C(n_1534),
.Y(n_2047)
);

AOI21xp5_ASAP7_75t_L g2048 ( 
.A1(n_2031),
.A2(n_1793),
.B(n_1708),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_2042),
.B(n_1945),
.Y(n_2049)
);

NOR3xp33_ASAP7_75t_L g2050 ( 
.A(n_2028),
.B(n_1535),
.C(n_1507),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_SL g2051 ( 
.A(n_2032),
.B(n_1636),
.Y(n_2051)
);

NAND3xp33_ASAP7_75t_L g2052 ( 
.A(n_2023),
.B(n_1750),
.C(n_1644),
.Y(n_2052)
);

OAI21xp5_ASAP7_75t_L g2053 ( 
.A1(n_2025),
.A2(n_1528),
.B(n_1797),
.Y(n_2053)
);

NOR2x1_ASAP7_75t_L g2054 ( 
.A(n_2038),
.B(n_1608),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_2043),
.B(n_1945),
.Y(n_2055)
);

NOR2xp67_ASAP7_75t_L g2056 ( 
.A(n_2027),
.B(n_1579),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_2030),
.B(n_1924),
.Y(n_2057)
);

NOR3xp33_ASAP7_75t_SL g2058 ( 
.A(n_2041),
.B(n_1636),
.C(n_1579),
.Y(n_2058)
);

HB1xp67_ASAP7_75t_L g2059 ( 
.A(n_2049),
.Y(n_2059)
);

NOR2xp67_ASAP7_75t_SL g2060 ( 
.A(n_2045),
.B(n_1530),
.Y(n_2060)
);

OAI22xp33_ASAP7_75t_L g2061 ( 
.A1(n_2051),
.A2(n_2040),
.B1(n_2035),
.B2(n_2034),
.Y(n_2061)
);

AOI211xp5_ASAP7_75t_L g2062 ( 
.A1(n_2056),
.A2(n_2036),
.B(n_2037),
.C(n_2039),
.Y(n_2062)
);

AOI221xp5_ASAP7_75t_L g2063 ( 
.A1(n_2044),
.A2(n_2046),
.B1(n_2055),
.B2(n_2052),
.C(n_2047),
.Y(n_2063)
);

NAND4xp25_ASAP7_75t_SL g2064 ( 
.A(n_2054),
.B(n_2033),
.C(n_1636),
.D(n_1625),
.Y(n_2064)
);

NOR4xp25_ASAP7_75t_L g2065 ( 
.A(n_2057),
.B(n_1834),
.C(n_1840),
.D(n_1725),
.Y(n_2065)
);

NOR2xp67_ASAP7_75t_SL g2066 ( 
.A(n_2048),
.B(n_1530),
.Y(n_2066)
);

NAND4xp25_ASAP7_75t_SL g2067 ( 
.A(n_2058),
.B(n_1625),
.C(n_1819),
.D(n_1817),
.Y(n_2067)
);

NOR3xp33_ASAP7_75t_SL g2068 ( 
.A(n_2053),
.B(n_1838),
.C(n_1821),
.Y(n_2068)
);

OAI211xp5_ASAP7_75t_SL g2069 ( 
.A1(n_2050),
.A2(n_1676),
.B(n_1690),
.C(n_1666),
.Y(n_2069)
);

OR2x2_ASAP7_75t_L g2070 ( 
.A(n_2055),
.B(n_1903),
.Y(n_2070)
);

NAND3xp33_ASAP7_75t_L g2071 ( 
.A(n_2044),
.B(n_1608),
.C(n_1845),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2049),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_SL g2073 ( 
.A(n_2061),
.B(n_1811),
.Y(n_2073)
);

NAND4xp75_ASAP7_75t_L g2074 ( 
.A(n_2063),
.B(n_1666),
.C(n_1690),
.D(n_1676),
.Y(n_2074)
);

AOI211xp5_ASAP7_75t_L g2075 ( 
.A1(n_2064),
.A2(n_1505),
.B(n_1508),
.C(n_1694),
.Y(n_2075)
);

NAND3xp33_ASAP7_75t_SL g2076 ( 
.A(n_2062),
.B(n_1641),
.C(n_1701),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2059),
.B(n_2072),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_2070),
.Y(n_2078)
);

OR2x2_ASAP7_75t_L g2079 ( 
.A(n_2071),
.B(n_1931),
.Y(n_2079)
);

OR2x2_ASAP7_75t_L g2080 ( 
.A(n_2065),
.B(n_1931),
.Y(n_2080)
);

AND3x4_ASAP7_75t_L g2081 ( 
.A(n_2068),
.B(n_1508),
.C(n_1700),
.Y(n_2081)
);

NAND2x1p5_ASAP7_75t_L g2082 ( 
.A(n_2060),
.B(n_2066),
.Y(n_2082)
);

XNOR2xp5_ASAP7_75t_L g2083 ( 
.A(n_2082),
.B(n_2067),
.Y(n_2083)
);

NAND2x1p5_ASAP7_75t_L g2084 ( 
.A(n_2073),
.B(n_1508),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2077),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_2078),
.Y(n_2086)
);

INVx3_ASAP7_75t_L g2087 ( 
.A(n_2074),
.Y(n_2087)
);

NAND2x1p5_ASAP7_75t_L g2088 ( 
.A(n_2080),
.B(n_1701),
.Y(n_2088)
);

XOR2xp5_ASAP7_75t_L g2089 ( 
.A(n_2074),
.B(n_1641),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2079),
.B(n_1876),
.Y(n_2090)
);

NOR2x1_ASAP7_75t_L g2091 ( 
.A(n_2076),
.B(n_2069),
.Y(n_2091)
);

BUFx2_ASAP7_75t_L g2092 ( 
.A(n_2091),
.Y(n_2092)
);

OAI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_2087),
.A2(n_2081),
.B1(n_2075),
.B2(n_1708),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2086),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2085),
.Y(n_2095)
);

XNOR2xp5_ASAP7_75t_L g2096 ( 
.A(n_2083),
.B(n_1694),
.Y(n_2096)
);

AOI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_2091),
.A2(n_1700),
.B1(n_1847),
.B2(n_1754),
.Y(n_2097)
);

XNOR2x1_ASAP7_75t_L g2098 ( 
.A(n_2087),
.B(n_1564),
.Y(n_2098)
);

AO211x2_ASAP7_75t_L g2099 ( 
.A1(n_2094),
.A2(n_2085),
.B(n_2089),
.C(n_2088),
.Y(n_2099)
);

OAI22xp5_ASAP7_75t_L g2100 ( 
.A1(n_2096),
.A2(n_2084),
.B1(n_2090),
.B2(n_1701),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2095),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_SL g2102 ( 
.A(n_2101),
.B(n_2092),
.Y(n_2102)
);

AOI21xp5_ASAP7_75t_L g2103 ( 
.A1(n_2102),
.A2(n_2099),
.B(n_2098),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2103),
.B(n_2093),
.Y(n_2104)
);

OR2x2_ASAP7_75t_L g2105 ( 
.A(n_2104),
.B(n_2100),
.Y(n_2105)
);

AOI222xp33_ASAP7_75t_L g2106 ( 
.A1(n_2105),
.A2(n_1660),
.B1(n_2097),
.B2(n_1642),
.C1(n_1507),
.C2(n_1716),
.Y(n_2106)
);


endmodule