module real_aes_15649_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_397;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_0), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g621 ( .A(n_1), .Y(n_621) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_2), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_3), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g581 ( .A(n_3), .Y(n_581) );
BUFx3_ASAP7_75t_L g224 ( .A(n_4), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_5), .Y(n_524) );
OAI22xp33_ASAP7_75t_L g588 ( .A1(n_6), .A2(n_73), .B1(n_589), .B2(n_593), .Y(n_588) );
OAI22xp33_ASAP7_75t_L g634 ( .A1(n_6), .A2(n_73), .B1(n_635), .B2(n_638), .Y(n_634) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_7), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_8), .B(n_187), .Y(n_186) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_8), .Y(n_689) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_9), .Y(n_92) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_10), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_11), .B(n_116), .Y(n_211) );
XNOR2xp5_ASAP7_75t_L g482 ( .A(n_12), .B(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_13), .B(n_125), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g115 ( .A1(n_14), .A2(n_64), .B1(n_113), .B2(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g712 ( .A(n_14), .Y(n_712) );
INVx1_ASAP7_75t_L g501 ( .A(n_15), .Y(n_501) );
INVx1_ASAP7_75t_L g508 ( .A(n_15), .Y(n_508) );
INVx2_ASAP7_75t_L g494 ( .A(n_16), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_17), .Y(n_528) );
OAI21x1_ASAP7_75t_L g107 ( .A1(n_18), .A2(n_31), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g681 ( .A(n_19), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_20), .B(n_132), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_21), .A2(n_69), .B1(n_600), .B2(n_603), .Y(n_599) );
OAI22xp33_ASAP7_75t_L g659 ( .A1(n_21), .A2(n_69), .B1(n_660), .B2(n_662), .Y(n_659) );
AO32x1_ASAP7_75t_L g105 ( .A1(n_22), .A2(n_106), .A3(n_109), .B1(n_117), .B2(n_119), .Y(n_105) );
AO32x2_ASAP7_75t_L g232 ( .A1(n_22), .A2(n_106), .A3(n_109), .B1(n_117), .B2(n_119), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_23), .A2(n_34), .B1(n_132), .B2(n_133), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_24), .B(n_157), .Y(n_156) );
AOI22xp5_ASAP7_75t_L g112 ( .A1(n_25), .A2(n_70), .B1(n_113), .B2(n_114), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_26), .B(n_155), .Y(n_160) );
INVx2_ASAP7_75t_L g493 ( .A(n_27), .Y(n_493) );
INVx1_ASAP7_75t_L g537 ( .A(n_27), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_28), .A2(n_48), .B1(n_114), .B2(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g704 ( .A(n_29), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_30), .B(n_162), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_32), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_33), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_35), .A2(n_59), .B1(n_141), .B2(n_155), .Y(n_171) );
BUFx3_ASAP7_75t_L g499 ( .A(n_36), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_37), .A2(n_61), .B1(n_113), .B2(n_116), .Y(n_220) );
AND2x4_ASAP7_75t_L g84 ( .A(n_38), .B(n_85), .Y(n_84) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_38), .Y(n_674) );
INVx1_ASAP7_75t_L g108 ( .A(n_39), .Y(n_108) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_40), .Y(n_557) );
INVx1_ASAP7_75t_L g627 ( .A(n_41), .Y(n_627) );
OAI211xp5_ASAP7_75t_L g641 ( .A1(n_41), .A2(n_642), .B(n_645), .C(n_649), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_42), .B(n_113), .Y(n_185) );
INVx1_ASAP7_75t_L g85 ( .A(n_43), .Y(n_85) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_44), .B(n_119), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_45), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g137 ( .A1(n_46), .A2(n_138), .B(n_139), .C(n_142), .Y(n_137) );
NAND3xp33_ASAP7_75t_L g191 ( .A(n_47), .B(n_113), .C(n_190), .Y(n_191) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_49), .Y(n_556) );
OAI211xp5_ASAP7_75t_L g609 ( .A1(n_50), .A2(n_610), .B(n_613), .C(n_618), .Y(n_609) );
INVx1_ASAP7_75t_L g658 ( .A(n_50), .Y(n_658) );
BUFx2_ASAP7_75t_L g683 ( .A(n_51), .Y(n_683) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_52), .Y(n_542) );
AND2x2_ASAP7_75t_L g145 ( .A(n_53), .B(n_146), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_54), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_55), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_56), .A2(n_74), .B1(n_116), .B2(n_141), .Y(n_173) );
INVx2_ASAP7_75t_L g94 ( .A(n_57), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_58), .B(n_208), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_60), .Y(n_131) );
BUFx3_ASAP7_75t_L g549 ( .A(n_62), .Y(n_549) );
INVx1_ASAP7_75t_L g596 ( .A(n_62), .Y(n_596) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_63), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_65), .B(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g491 ( .A(n_66), .Y(n_491) );
INVx1_ASAP7_75t_L g536 ( .A(n_66), .Y(n_536) );
INVx2_ASAP7_75t_L g547 ( .A(n_66), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_67), .A2(n_76), .B1(n_114), .B2(n_133), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_68), .B(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g723 ( .A(n_70), .Y(n_723) );
BUFx2_ASAP7_75t_L g691 ( .A(n_71), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_72), .B(n_125), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_75), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_95), .B(n_481), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
BUFx3_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NOR2xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_86), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
BUFx10_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx1_ASAP7_75t_L g118 ( .A(n_84), .Y(n_118) );
INVx1_ASAP7_75t_L g144 ( .A(n_84), .Y(n_144) );
BUFx10_ASAP7_75t_L g192 ( .A(n_84), .Y(n_192) );
AO31x2_ASAP7_75t_L g244 ( .A1(n_84), .A2(n_169), .A3(n_245), .B(n_249), .Y(n_244) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_85), .Y(n_676) );
AOI21xp5_ASAP7_75t_SL g725 ( .A1(n_86), .A2(n_675), .B(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g86 ( .A(n_87), .B(n_93), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx2_ASAP7_75t_L g113 ( .A(n_92), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_92), .Y(n_114) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_92), .Y(n_116) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_92), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_92), .Y(n_133) );
INVx1_ASAP7_75t_L g138 ( .A(n_92), .Y(n_138) );
INVx1_ASAP7_75t_L g141 ( .A(n_92), .Y(n_141) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_92), .Y(n_187) );
INVx1_ASAP7_75t_L g204 ( .A(n_92), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g109 ( .A1(n_93), .A2(n_110), .B1(n_112), .B2(n_115), .Y(n_109) );
INVx6_ASAP7_75t_L g163 ( .A(n_93), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_93), .A2(n_185), .B(n_186), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_93), .A2(n_163), .B1(n_220), .B2(n_221), .Y(n_219) );
BUFx8_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g111 ( .A(n_94), .Y(n_111) );
INVx1_ASAP7_75t_L g136 ( .A(n_94), .Y(n_136) );
INVx2_ASAP7_75t_L g143 ( .A(n_94), .Y(n_143) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
NOR2x1p5_ASAP7_75t_L g96 ( .A(n_97), .B(n_401), .Y(n_96) );
NAND4xp75_ASAP7_75t_L g97 ( .A(n_98), .B(n_280), .C(n_333), .D(n_378), .Y(n_97) );
NOR2x1_ASAP7_75t_L g98 ( .A(n_99), .B(n_237), .Y(n_98) );
OAI21xp33_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_165), .B(n_194), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_120), .Y(n_101) );
AND2x4_ASAP7_75t_L g369 ( .A(n_102), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_102), .B(n_243), .Y(n_397) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_103), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g362 ( .A(n_104), .Y(n_362) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_104), .Y(n_384) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_L g268 ( .A(n_105), .B(n_244), .Y(n_268) );
INVx1_ASAP7_75t_L g290 ( .A(n_105), .Y(n_290) );
AND2x2_ASAP7_75t_L g324 ( .A(n_105), .B(n_244), .Y(n_324) );
INVx4_ASAP7_75t_L g119 ( .A(n_106), .Y(n_119) );
INVx2_ASAP7_75t_SL g151 ( .A(n_106), .Y(n_151) );
BUFx3_ASAP7_75t_L g169 ( .A(n_106), .Y(n_169) );
INVx2_ASAP7_75t_L g199 ( .A(n_106), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_106), .B(n_223), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_106), .B(n_250), .Y(n_249) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g127 ( .A(n_107), .Y(n_127) );
O2A1O1Ixp5_ASAP7_75t_L g201 ( .A1(n_110), .A2(n_202), .B(n_203), .C(n_205), .Y(n_201) );
BUFx4f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g190 ( .A(n_111), .Y(n_190) );
INVx2_ASAP7_75t_SL g155 ( .A(n_113), .Y(n_155) );
INVx2_ASAP7_75t_L g157 ( .A(n_114), .Y(n_157) );
INVx3_ASAP7_75t_L g162 ( .A(n_116), .Y(n_162) );
OAI21x1_ASAP7_75t_L g152 ( .A1(n_117), .A2(n_153), .B(n_159), .Y(n_152) );
INVx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g174 ( .A(n_118), .Y(n_174) );
INVx2_ASAP7_75t_L g218 ( .A(n_119), .Y(n_218) );
INVxp33_ASAP7_75t_L g319 ( .A(n_120), .Y(n_319) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g431 ( .A(n_121), .B(n_268), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_148), .Y(n_121) );
OR2x2_ASAP7_75t_L g311 ( .A(n_122), .B(n_149), .Y(n_311) );
INVx1_ASAP7_75t_L g344 ( .A(n_122), .Y(n_344) );
INVx1_ASAP7_75t_L g348 ( .A(n_122), .Y(n_348) );
AND2x2_ASAP7_75t_L g464 ( .A(n_122), .B(n_279), .Y(n_464) );
OR2x2_ASAP7_75t_L g470 ( .A(n_122), .B(n_290), .Y(n_470) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g229 ( .A(n_123), .Y(n_229) );
AOI21x1_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_128), .B(n_145), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g147 ( .A(n_127), .Y(n_147) );
INVx2_ASAP7_75t_L g182 ( .A(n_127), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_137), .B(n_144), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g129 ( .A(n_130), .B(n_135), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_132), .B1(n_133), .B2(n_134), .Y(n_130) );
INVx2_ASAP7_75t_L g247 ( .A(n_132), .Y(n_247) );
INVx1_ASAP7_75t_L g210 ( .A(n_133), .Y(n_210) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_SL g172 ( .A(n_136), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
INVx2_ASAP7_75t_L g158 ( .A(n_142), .Y(n_158) );
BUFx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g209 ( .A(n_143), .Y(n_209) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_147), .B(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g364 ( .A(n_148), .B(n_314), .Y(n_364) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g230 ( .A(n_149), .B(n_231), .Y(n_230) );
OR2x2_ASAP7_75t_L g234 ( .A(n_149), .B(n_231), .Y(n_234) );
AND2x2_ASAP7_75t_L g241 ( .A(n_149), .B(n_232), .Y(n_241) );
INVx2_ASAP7_75t_L g265 ( .A(n_149), .Y(n_265) );
INVx1_ASAP7_75t_L g288 ( .A(n_149), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_149), .B(n_244), .Y(n_361) );
AND2x2_ASAP7_75t_L g370 ( .A(n_149), .B(n_228), .Y(n_370) );
INVxp67_ASAP7_75t_L g440 ( .A(n_149), .Y(n_440) );
BUFx2_ASAP7_75t_L g448 ( .A(n_149), .Y(n_448) );
INVx1_ASAP7_75t_L g478 ( .A(n_149), .Y(n_478) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OAI21x1_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_164), .Y(n_150) );
AOI21x1_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_156), .B(n_158), .Y(n_153) );
OAI21xp5_ASAP7_75t_L g188 ( .A1(n_157), .A2(n_189), .B(n_191), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_158), .A2(n_163), .B1(n_246), .B2(n_248), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_163), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g170 ( .A1(n_163), .A2(n_171), .B1(n_172), .B2(n_173), .Y(n_170) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_167), .B(n_177), .Y(n_166) );
OR2x2_ASAP7_75t_L g236 ( .A(n_167), .B(n_197), .Y(n_236) );
AND2x2_ASAP7_75t_L g386 ( .A(n_167), .B(n_270), .Y(n_386) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OR2x2_ASAP7_75t_L g214 ( .A(n_168), .B(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g262 ( .A(n_168), .Y(n_262) );
AND2x2_ASAP7_75t_L g285 ( .A(n_168), .B(n_256), .Y(n_285) );
INVx1_ASAP7_75t_L g318 ( .A(n_168), .Y(n_318) );
AND2x2_ASAP7_75t_L g354 ( .A(n_168), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g359 ( .A(n_168), .B(n_215), .Y(n_359) );
AND2x2_ASAP7_75t_L g417 ( .A(n_168), .B(n_259), .Y(n_417) );
OR2x2_ASAP7_75t_L g426 ( .A(n_168), .B(n_198), .Y(n_426) );
AO31x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .A3(n_174), .B(n_175), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_177), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g302 ( .A(n_178), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_178), .B(n_255), .Y(n_343) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g272 ( .A(n_179), .Y(n_272) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
OR2x2_ASAP7_75t_L g296 ( .A(n_180), .B(n_216), .Y(n_296) );
OAI21x1_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_183), .B(n_193), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_181), .A2(n_183), .B(n_193), .Y(n_213) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
OAI21x1_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_188), .B(n_192), .Y(n_183) );
OAI21x1_ASAP7_75t_L g200 ( .A1(n_192), .A2(n_201), .B(n_206), .Y(n_200) );
AOI31xp67_ASAP7_75t_L g217 ( .A1(n_192), .A2(n_218), .A3(n_219), .B(n_222), .Y(n_217) );
AOI22xp33_ASAP7_75t_SL g194 ( .A1(n_195), .A2(n_225), .B1(n_233), .B2(n_235), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_196), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_214), .Y(n_196) );
INVx1_ASAP7_75t_L g367 ( .A(n_197), .Y(n_367) );
OR2x2_ASAP7_75t_L g480 ( .A(n_197), .B(n_376), .Y(n_480) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_213), .Y(n_197) );
INVx2_ASAP7_75t_SL g252 ( .A(n_198), .Y(n_252) );
BUFx2_ASAP7_75t_L g293 ( .A(n_198), .Y(n_293) );
AND2x2_ASAP7_75t_L g317 ( .A(n_198), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g355 ( .A(n_198), .Y(n_355) );
OA21x2_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_212), .Y(n_198) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_199), .A2(n_200), .B(n_212), .Y(n_259) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_209), .B1(n_210), .B2(n_211), .Y(n_206) );
INVx2_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g258 ( .A(n_213), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g418 ( .A(n_213), .B(n_256), .Y(n_418) );
INVx1_ASAP7_75t_L g275 ( .A(n_214), .Y(n_275) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g256 ( .A(n_217), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_230), .Y(n_226) );
AND2x2_ASAP7_75t_L g474 ( .A(n_227), .B(n_241), .Y(n_474) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g243 ( .A(n_229), .B(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g278 ( .A(n_229), .Y(n_278) );
INVx1_ASAP7_75t_L g291 ( .A(n_229), .Y(n_291) );
INVx1_ASAP7_75t_L g383 ( .A(n_229), .Y(n_383) );
NAND2x1p5_ASAP7_75t_L g276 ( .A(n_230), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g282 ( .A(n_230), .B(n_243), .Y(n_282) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x4_ASAP7_75t_L g314 ( .A(n_232), .B(n_279), .Y(n_314) );
INVx1_ASAP7_75t_L g332 ( .A(n_232), .Y(n_332) );
INVx2_ASAP7_75t_L g427 ( .A(n_233), .Y(n_427) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AOI321xp33_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_251), .A3(n_253), .B1(n_257), .B2(n_263), .C(n_266), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g263 ( .A(n_243), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g304 ( .A(n_243), .B(n_305), .Y(n_304) );
INVx3_ASAP7_75t_L g279 ( .A(n_244), .Y(n_279) );
AND2x2_ASAP7_75t_L g382 ( .A(n_244), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_252), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_254), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g327 ( .A(n_255), .Y(n_327) );
AND2x2_ASAP7_75t_L g389 ( .A(n_255), .B(n_318), .Y(n_389) );
AND2x2_ASAP7_75t_L g409 ( .A(n_255), .B(n_272), .Y(n_409) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g303 ( .A(n_256), .B(n_259), .Y(n_303) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
AND2x2_ASAP7_75t_L g388 ( .A(n_258), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g428 ( .A(n_258), .Y(n_428) );
INVx1_ASAP7_75t_L g273 ( .A(n_259), .Y(n_273) );
OAI32xp33_ASAP7_75t_L g266 ( .A1(n_260), .A2(n_267), .A3(n_269), .B1(n_274), .B2(n_276), .Y(n_266) );
OR2x2_ASAP7_75t_L g300 ( .A(n_260), .B(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g294 ( .A(n_261), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_261), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g461 ( .A(n_261), .B(n_296), .Y(n_461) );
INVx2_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g308 ( .A(n_262), .B(n_272), .Y(n_308) );
OR2x2_ASAP7_75t_L g477 ( .A(n_262), .B(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_264), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g267 ( .A(n_265), .B(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_265), .Y(n_305) );
OR2x2_ASAP7_75t_L g322 ( .A(n_265), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g455 ( .A(n_265), .B(n_382), .Y(n_455) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_265), .Y(n_469) );
INVx2_ASAP7_75t_L g406 ( .A(n_268), .Y(n_406) );
OR2x2_ASAP7_75t_L g447 ( .A(n_268), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g451 ( .A(n_269), .Y(n_451) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g465 ( .A(n_270), .B(n_285), .Y(n_465) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g326 ( .A(n_271), .B(n_327), .Y(n_326) );
NAND2x1p5_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx2_ASAP7_75t_L g422 ( .A(n_277), .Y(n_422) );
AND2x4_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g338 ( .A(n_279), .Y(n_338) );
INVx1_ASAP7_75t_L g374 ( .A(n_279), .Y(n_374) );
NOR2x1_ASAP7_75t_L g280 ( .A(n_281), .B(n_297), .Y(n_280) );
AO22x1_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B1(n_286), .B2(n_292), .Y(n_281) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g376 ( .A(n_285), .Y(n_376) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_287), .A2(n_380), .B1(n_385), .B2(n_387), .Y(n_379) );
NAND2x1p5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g330 ( .A(n_291), .Y(n_330) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
AND2x2_ASAP7_75t_L g358 ( .A(n_293), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g395 ( .A(n_293), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_294), .A2(n_400), .B1(n_433), .B2(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g316 ( .A(n_296), .Y(n_316) );
OR2x2_ASAP7_75t_L g441 ( .A(n_296), .B(n_426), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_298), .B(n_320), .Y(n_297) );
AOI21xp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_304), .B(n_306), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_299), .A2(n_321), .B1(n_325), .B2(n_328), .Y(n_320) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g351 ( .A(n_301), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx2_ASAP7_75t_L g377 ( .A(n_302), .Y(n_377) );
AND2x2_ASAP7_75t_L g434 ( .A(n_302), .B(n_317), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_303), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g336 ( .A(n_305), .B(n_337), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_309), .B1(n_315), .B2(n_319), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_311), .B(n_323), .Y(n_433) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp33_ASAP7_75t_R g328 ( .A(n_313), .B(n_329), .Y(n_328) );
INVx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g346 ( .A(n_314), .B(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g400 ( .A(n_314), .B(n_344), .Y(n_400) );
BUFx2_ASAP7_75t_L g463 ( .A(n_314), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x2_ASAP7_75t_L g394 ( .A(n_316), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g438 ( .A(n_316), .B(n_354), .Y(n_438) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_323), .Y(n_393) );
INVx2_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g411 ( .A(n_324), .B(n_348), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g459 ( .A(n_330), .Y(n_459) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g454 ( .A(n_332), .Y(n_454) );
NOR2x1_ASAP7_75t_L g333 ( .A(n_334), .B(n_356), .Y(n_333) );
OAI21xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_339), .B(n_345), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g435 ( .A1(n_335), .A2(n_436), .B(n_444), .Y(n_435) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_343), .B(n_344), .Y(n_342) );
AND2x2_ASAP7_75t_L g405 ( .A(n_344), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_349), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g408 ( .A(n_354), .B(n_409), .Y(n_408) );
OAI211xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_360), .B(n_363), .C(n_368), .Y(n_356) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI21xp5_ASAP7_75t_SL g444 ( .A1(n_360), .A2(n_441), .B(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI211xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_371), .B(n_375), .C(n_377), .Y(n_368) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_370), .Y(n_443) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g472 ( .A(n_377), .Y(n_472) );
NOR3x1_ASAP7_75t_L g378 ( .A(n_379), .B(n_390), .C(n_398), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_388), .A2(n_392), .B1(n_394), .B2(n_396), .Y(n_391) );
INVx2_ASAP7_75t_L g473 ( .A(n_389), .Y(n_473) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_394), .B(n_400), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_394), .A2(n_468), .B1(n_471), .B2(n_474), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_394), .A2(n_411), .B1(n_476), .B2(n_479), .Y(n_475) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND4xp75_ASAP7_75t_L g401 ( .A(n_402), .B(n_435), .C(n_449), .D(n_466), .Y(n_401) );
NOR2xp67_ASAP7_75t_L g402 ( .A(n_403), .B(n_419), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_407), .B1(n_410), .B2(n_412), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g414 ( .A(n_408), .Y(n_414) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
AND2x2_ASAP7_75t_L g424 ( .A(n_418), .B(n_425), .Y(n_424) );
OAI321xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_423), .A3(n_427), .B1(n_428), .B2(n_429), .C(n_432), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_422), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_424), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_439), .B1(n_441), .B2(n_442), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVxp67_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_447), .Y(n_460) );
NOR2x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_456), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_455), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_460), .B(n_461), .C(n_462), .Y(n_456) );
INVxp33_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI21xp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .B(n_465), .Y(n_462) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_475), .Y(n_466) );
NOR2x1p5_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
NOR2xp67_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
INVx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OAI221xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B1(n_670), .B2(n_677), .C(n_718), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_483), .A2(n_719), .B1(n_722), .B2(n_724), .Y(n_718) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND3x1_ASAP7_75t_L g484 ( .A(n_485), .B(n_587), .C(n_633), .Y(n_484) );
NOR2xp33_ASAP7_75t_SL g485 ( .A(n_486), .B(n_543), .Y(n_485) );
OAI33xp33_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_495), .A3(n_510), .B1(n_523), .B2(n_531), .B3(n_538), .Y(n_486) );
BUFx8_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_492), .Y(n_488) );
INVx1_ASAP7_75t_L g583 ( .A(n_489), .Y(n_583) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_489), .Y(n_669) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx2_ASAP7_75t_L g632 ( .A(n_490), .Y(n_632) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g709 ( .A(n_492), .Y(n_709) );
NAND2xp33_ASAP7_75t_SL g492 ( .A(n_493), .B(n_494), .Y(n_492) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_493), .Y(n_667) );
INVx1_ASAP7_75t_L g703 ( .A(n_493), .Y(n_703) );
INVx3_ASAP7_75t_L g534 ( .A(n_494), .Y(n_534) );
BUFx3_ASAP7_75t_L g653 ( .A(n_494), .Y(n_653) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B1(n_502), .B2(n_503), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_496), .A2(n_539), .B1(n_551), .B2(n_558), .Y(n_550) );
OAI22xp33_ASAP7_75t_L g538 ( .A1(n_497), .A2(n_539), .B1(n_540), .B2(n_542), .Y(n_538) );
BUFx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OR2x4_ASAP7_75t_L g637 ( .A(n_498), .B(n_534), .Y(n_637) );
OR2x4_ASAP7_75t_L g661 ( .A(n_498), .B(n_640), .Y(n_661) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_499), .Y(n_509) );
INVx2_ASAP7_75t_L g517 ( .A(n_499), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_499), .B(n_508), .Y(n_522) );
AND2x4_ASAP7_75t_L g647 ( .A(n_499), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVxp67_ASAP7_75t_L g516 ( .A(n_501), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_502), .A2(n_542), .B1(n_573), .B2(n_575), .Y(n_572) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_506), .Y(n_541) );
BUFx2_ASAP7_75t_L g644 ( .A(n_506), .Y(n_644) );
NAND2x1p5_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
BUFx2_ASAP7_75t_L g657 ( .A(n_507), .Y(n_657) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g648 ( .A(n_508), .Y(n_648) );
BUFx2_ASAP7_75t_L g654 ( .A(n_509), .Y(n_654) );
INVx2_ASAP7_75t_L g701 ( .A(n_509), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_518), .B2(n_519), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_511), .A2(n_524), .B1(n_565), .B2(n_569), .Y(n_564) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x4_ASAP7_75t_L g639 ( .A(n_514), .B(n_640), .Y(n_639) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g527 ( .A(n_515), .Y(n_527) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_518), .A2(n_528), .B1(n_551), .B2(n_585), .Y(n_584) );
CKINVDCx8_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
BUFx2_ASAP7_75t_L g530 ( .A(n_522), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B1(n_528), .B2(n_529), .Y(n_523) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OR2x6_ASAP7_75t_L g664 ( .A(n_530), .B(n_534), .Y(n_664) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND3x1_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .C(n_537), .Y(n_533) );
INVx1_ASAP7_75t_L g640 ( .A(n_534), .Y(n_640) );
AND2x4_ASAP7_75t_L g646 ( .A(n_534), .B(n_647), .Y(n_646) );
AND2x4_ASAP7_75t_L g702 ( .A(n_534), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OAI33xp33_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_550), .A3(n_564), .B1(n_572), .B2(n_578), .B3(n_584), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x4_ASAP7_75t_L g545 ( .A(n_546), .B(n_548), .Y(n_545) );
BUFx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x4_ASAP7_75t_L g580 ( .A(n_549), .B(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g592 ( .A(n_549), .Y(n_592) );
BUFx2_ASAP7_75t_L g608 ( .A(n_549), .Y(n_608) );
AND2x4_ASAP7_75t_L g624 ( .A(n_549), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx4f_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g590 ( .A(n_554), .Y(n_590) );
INVx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
INVx2_ASAP7_75t_L g563 ( .A(n_556), .Y(n_563) );
INVx2_ASAP7_75t_L g568 ( .A(n_556), .Y(n_568) );
NAND2x1_ASAP7_75t_L g571 ( .A(n_556), .B(n_557), .Y(n_571) );
AND2x2_ASAP7_75t_L g597 ( .A(n_556), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g617 ( .A(n_556), .B(n_557), .Y(n_617) );
INVx1_ASAP7_75t_L g626 ( .A(n_556), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_557), .B(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g567 ( .A(n_557), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g598 ( .A(n_557), .Y(n_598) );
BUFx2_ASAP7_75t_L g620 ( .A(n_557), .Y(n_620) );
INVx6_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g586 ( .A(n_560), .Y(n_586) );
INVx8_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g607 ( .A(n_561), .B(n_608), .Y(n_607) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g574 ( .A(n_565), .Y(n_574) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
BUFx4f_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx4f_ASAP7_75t_L g612 ( .A(n_570), .Y(n_612) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
BUFx3_ASAP7_75t_L g577 ( .A(n_571), .Y(n_577) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx5_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
INVx1_ASAP7_75t_L g630 ( .A(n_581), .Y(n_630) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
BUFx3_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OAI31xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_599), .A3(n_609), .B(n_628), .Y(n_587) );
OR2x6_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
OR2x6_ASAP7_75t_L g602 ( .A(n_590), .B(n_595), .Y(n_602) );
INVxp67_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g615 ( .A(n_592), .Y(n_615) );
INVx4_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g619 ( .A(n_608), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_621), .B1(n_622), .B2(n_627), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_621), .A2(n_650), .B1(n_655), .B2(n_658), .Y(n_649) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
BUFx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x4_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI31xp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_641), .A3(n_659), .B(n_665), .Y(n_633) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVxp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
CKINVDCx8_ASAP7_75t_R g645 ( .A(n_646), .Y(n_645) );
BUFx3_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
AND2x4_ASAP7_75t_L g656 ( .A(n_652), .B(n_657), .Y(n_656) );
INVx3_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
BUFx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_SL g665 ( .A(n_666), .B(n_668), .Y(n_665) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_671), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g671 ( .A(n_672), .Y(n_671) );
BUFx6f_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g711 ( .A(n_674), .Y(n_711) );
BUFx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_676), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g726 ( .A(n_676), .B(n_711), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_694), .B1(n_712), .B2(n_713), .Y(n_677) );
OAI22xp33_ASAP7_75t_L g719 ( .A1(n_678), .A2(n_712), .B1(n_720), .B2(n_721), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B1(n_684), .B2(n_693), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
XNOR2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g693 ( .A(n_684), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_686), .B1(n_687), .B2(n_688), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_690), .B1(n_691), .B2(n_692), .Y(n_688) );
INVx1_ASAP7_75t_L g692 ( .A(n_689), .Y(n_692) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx3_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
BUFx12f_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
BUFx4f_ASAP7_75t_SL g720 ( .A(n_696), .Y(n_720) );
BUFx8_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI211xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_704), .B(n_705), .C(n_710), .Y(n_697) );
AND2x2_ASAP7_75t_L g717 ( .A(n_698), .B(n_705), .Y(n_717) );
INVx4_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AND2x6_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
NAND3xp33_ASAP7_75t_L g705 ( .A(n_700), .B(n_706), .C(n_709), .Y(n_705) );
INVx3_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx3_ASAP7_75t_L g708 ( .A(n_704), .Y(n_708) );
INVx2_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
BUFx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g716 ( .A(n_710), .Y(n_716) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
BUFx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
BUFx3_ASAP7_75t_L g721 ( .A(n_715), .Y(n_721) );
OR2x6_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
endmodule