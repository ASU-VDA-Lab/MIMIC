module fake_jpeg_25876_n_33 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_33);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_33;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

AOI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_5),
.A2(n_1),
.B1(n_2),
.B2(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_7),
.C(n_1),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

NOR4xp25_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_17),
.C(n_15),
.D(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_25),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_20),
.A2(n_16),
.B1(n_9),
.B2(n_10),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_26),
.A2(n_3),
.B(n_5),
.Y(n_28)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_22),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_26),
.C(n_24),
.Y(n_30)
);

AOI322xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.A3(n_29),
.B1(n_28),
.B2(n_6),
.C1(n_27),
.C2(n_12),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_29),
.C(n_6),
.Y(n_33)
);


endmodule