module fake_jpeg_20253_n_168 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_27),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_0),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_21),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_85),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_51),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_80),
.A2(n_53),
.B1(n_61),
.B2(n_76),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_87),
.B(n_60),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_85),
.A2(n_69),
.B1(n_77),
.B2(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_92),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_57),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_66),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_70),
.C(n_58),
.Y(n_125)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_74),
.B1(n_64),
.B2(n_62),
.Y(n_120)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_60),
.B(n_75),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_82),
.B1(n_48),
.B2(n_49),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_56),
.B1(n_59),
.B2(n_67),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_115),
.B1(n_119),
.B2(n_5),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_50),
.B1(n_68),
.B2(n_71),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_66),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_116),
.A2(n_1),
.B(n_2),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_64),
.B1(n_62),
.B2(n_66),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_125),
.Y(n_133)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_1),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_127),
.Y(n_140)
);

AO22x2_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_78),
.B1(n_22),
.B2(n_23),
.Y(n_127)
);

OR2x6_ASAP7_75t_SL g128 ( 
.A(n_113),
.B(n_18),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_128),
.A2(n_135),
.B(n_127),
.Y(n_147)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_130),
.A2(n_131),
.B(n_141),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_127),
.A2(n_2),
.B(n_3),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_117),
.B(n_4),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_136),
.Y(n_149)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_134),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_119),
.B1(n_8),
.B2(n_9),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_7),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_150),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_128),
.A2(n_111),
.B(n_8),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_148),
.A2(n_131),
.B1(n_137),
.B2(n_140),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_150)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_151),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_143),
.B1(n_152),
.B2(n_155),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_155),
.C(n_150),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_153),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_133),
.B(n_149),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_145),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_162),
.A2(n_144),
.B(n_29),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

AOI31xp67_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_17),
.A3(n_30),
.B(n_32),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_165),
.A2(n_34),
.B(n_37),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_43),
.C(n_45),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_46),
.Y(n_168)
);


endmodule