module fake_netlist_6_984_n_761 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_761);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_761;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_685;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_746;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_683;
wire n_420;
wire n_620;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

BUFx3_ASAP7_75t_L g154 ( 
.A(n_14),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_14),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_37),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_45),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_55),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_93),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_31),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_127),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_26),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_32),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_79),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_113),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_0),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_48),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_57),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_44),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_73),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_74),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_96),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_63),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_101),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_8),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_28),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_1),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_19),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_82),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_65),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_114),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_78),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_77),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_51),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_53),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_13),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_68),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_49),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_39),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_59),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_106),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_60),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_105),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_102),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_104),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_163),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_171),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_156),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_165),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_0),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_166),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_167),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_169),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_174),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_161),
.B(n_172),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_174),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_174),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_181),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_170),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_193),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_172),
.B(n_1),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_155),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_158),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_175),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_164),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_157),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_157),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_177),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_178),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_179),
.B(n_2),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_176),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_180),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

OAI21x1_ASAP7_75t_L g255 ( 
.A1(n_222),
.A2(n_199),
.B(n_179),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_212),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_206),
.B(n_186),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_207),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_224),
.B(n_159),
.Y(n_261)
);

OA21x2_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_199),
.B(n_186),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_208),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_210),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_162),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_221),
.A2(n_162),
.B1(n_204),
.B2(n_187),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_213),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_215),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_223),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_223),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_211),
.B(n_189),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_220),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_214),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_208),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_230),
.B(n_190),
.Y(n_278)
);

AND2x4_ASAP7_75t_L g279 ( 
.A(n_229),
.B(n_191),
.Y(n_279)
);

AND2x6_ASAP7_75t_L g280 ( 
.A(n_227),
.B(n_192),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_233),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_216),
.Y(n_282)
);

CKINVDCx6p67_ASAP7_75t_R g283 ( 
.A(n_221),
.Y(n_283)
);

AND2x4_ASAP7_75t_L g284 ( 
.A(n_217),
.B(n_194),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_228),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_235),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_240),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_241),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_218),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_239),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_225),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_250),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_247),
.Y(n_294)
);

NAND2x1p5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_197),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_247),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_250),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_253),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_198),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_225),
.Y(n_301)
);

OR2x6_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_201),
.Y(n_302)
);

CKINVDCx8_ASAP7_75t_R g303 ( 
.A(n_289),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_248),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_279),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_284),
.B(n_202),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_283),
.Y(n_307)
);

OR2x6_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_203),
.Y(n_308)
);

BUFx10_ASAP7_75t_L g309 ( 
.A(n_279),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_276),
.B(n_183),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_275),
.B(n_226),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_253),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_247),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_280),
.A2(n_226),
.B1(n_204),
.B2(n_200),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_258),
.B(n_187),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_254),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_248),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_247),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_284),
.B(n_205),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_247),
.Y(n_320)
);

AND2x6_ASAP7_75t_L g321 ( 
.A(n_278),
.B(n_286),
.Y(n_321)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_248),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_284),
.B(n_188),
.Y(n_323)
);

AND2x6_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_273),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_252),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_274),
.B(n_188),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_272),
.B(n_270),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_264),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_273),
.B(n_195),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_254),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_256),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_272),
.B(n_195),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_246),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_252),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_262),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_275),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_246),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_261),
.B(n_200),
.Y(n_338)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_252),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_L g340 ( 
.A1(n_265),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_277),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_256),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_265),
.Y(n_343)
);

INVx6_ASAP7_75t_L g344 ( 
.A(n_284),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_260),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_280),
.B(n_3),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_280),
.B(n_4),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g348 ( 
.A1(n_278),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_260),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_263),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_283),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_270),
.B(n_20),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_271),
.B(n_153),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_263),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_262),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_343),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_336),
.B(n_268),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_304),
.Y(n_358)
);

BUFx6f_ASAP7_75t_SL g359 ( 
.A(n_302),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_293),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_261),
.Y(n_361)
);

BUFx8_ASAP7_75t_L g362 ( 
.A(n_301),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_298),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_316),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_317),
.B(n_278),
.Y(n_365)
);

A2O1A1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_326),
.A2(n_255),
.B(n_266),
.C(n_285),
.Y(n_366)
);

AO22x2_ASAP7_75t_L g367 ( 
.A1(n_323),
.A2(n_279),
.B1(n_291),
.B2(n_306),
.Y(n_367)
);

BUFx8_ASAP7_75t_L g368 ( 
.A(n_311),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_326),
.B(n_282),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_330),
.B(n_268),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_331),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_342),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_296),
.Y(n_373)
);

AO22x2_ASAP7_75t_L g374 ( 
.A1(n_323),
.A2(n_279),
.B1(n_291),
.B2(n_290),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_345),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_327),
.Y(n_376)
);

AO22x2_ASAP7_75t_L g377 ( 
.A1(n_306),
.A2(n_290),
.B1(n_292),
.B2(n_288),
.Y(n_377)
);

NAND2x1p5_ASAP7_75t_L g378 ( 
.A(n_325),
.B(n_282),
.Y(n_378)
);

NAND2xp33_ASAP7_75t_SL g379 ( 
.A(n_348),
.B(n_267),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_317),
.B(n_280),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_322),
.B(n_280),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_327),
.Y(n_382)
);

AO22x2_ASAP7_75t_L g383 ( 
.A1(n_299),
.A2(n_290),
.B1(n_292),
.B2(n_288),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_329),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_329),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_312),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_322),
.B(n_280),
.Y(n_387)
);

AO22x2_ASAP7_75t_L g388 ( 
.A1(n_340),
.A2(n_292),
.B1(n_287),
.B2(n_285),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_349),
.Y(n_389)
);

AO22x2_ASAP7_75t_L g390 ( 
.A1(n_340),
.A2(n_287),
.B1(n_266),
.B2(n_269),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_350),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_345),
.Y(n_393)
);

AO22x2_ASAP7_75t_L g394 ( 
.A1(n_348),
.A2(n_269),
.B1(n_259),
.B2(n_271),
.Y(n_394)
);

OR2x6_ASAP7_75t_L g395 ( 
.A(n_302),
.B(n_289),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_354),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_307),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_333),
.Y(n_398)
);

NOR2xp67_ASAP7_75t_L g399 ( 
.A(n_315),
.B(n_257),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_337),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_318),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_339),
.B(n_280),
.Y(n_402)
);

AO22x2_ASAP7_75t_L g403 ( 
.A1(n_319),
.A2(n_249),
.B1(n_6),
.B2(n_7),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_318),
.Y(n_404)
);

A2O1A1Ixp33_ASAP7_75t_L g405 ( 
.A1(n_310),
.A2(n_255),
.B(n_251),
.C(n_249),
.Y(n_405)
);

AO22x2_ASAP7_75t_L g406 ( 
.A1(n_319),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_406)
);

AO22x2_ASAP7_75t_L g407 ( 
.A1(n_346),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_334),
.B(n_289),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_294),
.Y(n_409)
);

AO22x2_ASAP7_75t_L g410 ( 
.A1(n_347),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_410)
);

OAI221xp5_ASAP7_75t_L g411 ( 
.A1(n_300),
.A2(n_310),
.B1(n_332),
.B2(n_295),
.C(n_344),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_332),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_295),
.B(n_314),
.Y(n_413)
);

AO22x2_ASAP7_75t_L g414 ( 
.A1(n_328),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_352),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_352),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_353),
.Y(n_417)
);

NAND2x1p5_ASAP7_75t_L g418 ( 
.A(n_339),
.B(n_262),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_353),
.Y(n_419)
);

BUFx8_ASAP7_75t_L g420 ( 
.A(n_303),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_344),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_344),
.A2(n_262),
.B1(n_88),
.B2(n_89),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_392),
.B(n_305),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_369),
.B(n_305),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_384),
.B(n_309),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_376),
.B(n_321),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_385),
.B(n_309),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_399),
.B(n_300),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_361),
.B(n_341),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_412),
.B(n_379),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_408),
.B(n_335),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_382),
.B(n_335),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_357),
.B(n_335),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_373),
.B(n_335),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_321),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_416),
.B(n_321),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_370),
.B(n_355),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_413),
.B(n_386),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_358),
.B(n_355),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_358),
.B(n_355),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_356),
.B(n_355),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_360),
.B(n_351),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_363),
.B(n_297),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_364),
.B(n_313),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_417),
.B(n_321),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_371),
.B(n_372),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_378),
.B(n_419),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_421),
.B(n_320),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_365),
.B(n_321),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_389),
.B(n_324),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_391),
.B(n_324),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_395),
.B(n_302),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_375),
.B(n_324),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_393),
.B(n_324),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_396),
.B(n_324),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_380),
.B(n_308),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_394),
.B(n_308),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_381),
.B(n_308),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_387),
.B(n_21),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_395),
.B(n_15),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_402),
.B(n_22),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_398),
.B(n_23),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_400),
.B(n_24),
.Y(n_463)
);

NAND2xp33_ASAP7_75t_SL g464 ( 
.A(n_359),
.B(n_16),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_394),
.B(n_16),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_397),
.B(n_25),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_SL g467 ( 
.A(n_420),
.B(n_17),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_411),
.B(n_17),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_422),
.B(n_27),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_368),
.B(n_29),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_362),
.B(n_18),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_409),
.B(n_30),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_401),
.B(n_33),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_404),
.B(n_34),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_366),
.B(n_35),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_405),
.B(n_36),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_418),
.B(n_38),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_367),
.B(n_40),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_367),
.B(n_41),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_446),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_430),
.A2(n_390),
.B(n_388),
.Y(n_481)
);

AOI21x1_ASAP7_75t_SL g482 ( 
.A1(n_468),
.A2(n_403),
.B(n_406),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_449),
.A2(n_374),
.B(n_377),
.Y(n_483)
);

AO31x2_ASAP7_75t_L g484 ( 
.A1(n_457),
.A2(n_374),
.A3(n_377),
.B(n_403),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_465),
.A2(n_410),
.B1(n_407),
.B2(n_390),
.Y(n_485)
);

OA21x2_ASAP7_75t_L g486 ( 
.A1(n_475),
.A2(n_406),
.B(n_410),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_428),
.B(n_388),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_472),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_450),
.A2(n_407),
.B(n_42),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_472),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_429),
.B(n_383),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_452),
.B(n_383),
.Y(n_492)
);

BUFx6f_ASAP7_75t_SL g493 ( 
.A(n_452),
.Y(n_493)
);

AOI31xp67_ASAP7_75t_L g494 ( 
.A1(n_476),
.A2(n_414),
.A3(n_43),
.B(n_46),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_435),
.A2(n_414),
.B(n_47),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_436),
.A2(n_103),
.B(n_50),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_460),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_438),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_426),
.A2(n_18),
.B1(n_52),
.B2(n_54),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_445),
.A2(n_56),
.B(n_58),
.Y(n_500)
);

AOI21x1_ASAP7_75t_SL g501 ( 
.A1(n_474),
.A2(n_61),
.B(n_62),
.Y(n_501)
);

A2O1A1Ixp33_ASAP7_75t_L g502 ( 
.A1(n_447),
.A2(n_64),
.B(n_66),
.C(n_67),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_433),
.B(n_69),
.Y(n_503)
);

AOI221x1_ASAP7_75t_L g504 ( 
.A1(n_474),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.C(n_75),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_443),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_437),
.A2(n_76),
.B(n_80),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_431),
.A2(n_81),
.B(n_83),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_432),
.A2(n_84),
.B(n_85),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_471),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_466),
.Y(n_510)
);

AO31x2_ASAP7_75t_L g511 ( 
.A1(n_478),
.A2(n_86),
.A3(n_87),
.B(n_90),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_441),
.B(n_91),
.Y(n_512)
);

AO21x1_ASAP7_75t_L g513 ( 
.A1(n_479),
.A2(n_92),
.B(n_94),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_455),
.A2(n_95),
.B(n_97),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_453),
.A2(n_98),
.B(n_99),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_444),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_442),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_424),
.B(n_100),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_454),
.A2(n_107),
.B(n_108),
.Y(n_519)
);

CKINVDCx14_ASAP7_75t_R g520 ( 
.A(n_467),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_451),
.A2(n_110),
.B(n_111),
.Y(n_521)
);

OAI21x1_ASAP7_75t_L g522 ( 
.A1(n_448),
.A2(n_112),
.B(n_115),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_423),
.B(n_116),
.Y(n_523)
);

AO31x2_ASAP7_75t_L g524 ( 
.A1(n_456),
.A2(n_118),
.A3(n_119),
.B(n_120),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_425),
.B(n_121),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_480),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_521),
.A2(n_461),
.B(n_459),
.Y(n_527)
);

NAND2x1p5_ASAP7_75t_L g528 ( 
.A(n_488),
.B(n_439),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_483),
.A2(n_458),
.B(n_469),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_509),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_505),
.Y(n_531)
);

NAND3xp33_ASAP7_75t_L g532 ( 
.A(n_517),
.B(n_464),
.C(n_427),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_485),
.A2(n_477),
.B1(n_434),
.B2(n_470),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_501),
.A2(n_473),
.B(n_463),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_512),
.A2(n_440),
.B(n_462),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g536 ( 
.A1(n_500),
.A2(n_515),
.B(n_519),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_516),
.Y(n_537)
);

AO31x2_ASAP7_75t_L g538 ( 
.A1(n_485),
.A2(n_122),
.A3(n_123),
.B(n_124),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_497),
.Y(n_539)
);

CKINVDCx11_ASAP7_75t_R g540 ( 
.A(n_510),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_512),
.A2(n_125),
.B(n_126),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_486),
.A2(n_129),
.B1(n_130),
.B2(n_132),
.Y(n_542)
);

AO21x2_ASAP7_75t_L g543 ( 
.A1(n_508),
.A2(n_134),
.B(n_135),
.Y(n_543)
);

OAI22xp33_ASAP7_75t_L g544 ( 
.A1(n_498),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_490),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_487),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_484),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_484),
.Y(n_548)
);

OA21x2_ASAP7_75t_L g549 ( 
.A1(n_504),
.A2(n_141),
.B(n_142),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_523),
.B(n_143),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_503),
.A2(n_144),
.B(n_145),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_520),
.Y(n_552)
);

AOI21x1_ASAP7_75t_L g553 ( 
.A1(n_518),
.A2(n_149),
.B(n_150),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_493),
.Y(n_554)
);

OAI21x1_ASAP7_75t_L g555 ( 
.A1(n_522),
.A2(n_151),
.B(n_152),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_486),
.A2(n_495),
.B1(n_499),
.B2(n_523),
.Y(n_556)
);

NOR2xp67_ASAP7_75t_L g557 ( 
.A(n_518),
.B(n_525),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_481),
.B(n_491),
.Y(n_558)
);

NOR4xp25_ASAP7_75t_L g559 ( 
.A(n_492),
.B(n_499),
.C(n_481),
.D(n_502),
.Y(n_559)
);

OAI21x1_ASAP7_75t_L g560 ( 
.A1(n_489),
.A2(n_514),
.B(n_496),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_484),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_513),
.A2(n_508),
.B1(n_503),
.B2(n_507),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_494),
.A2(n_506),
.B(n_482),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_493),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_511),
.A2(n_411),
.B(n_449),
.Y(n_565)
);

BUFx12f_ASAP7_75t_L g566 ( 
.A(n_511),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_555),
.Y(n_567)
);

OAI21x1_ASAP7_75t_L g568 ( 
.A1(n_536),
.A2(n_524),
.B(n_511),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_531),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_547),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_548),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_561),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_540),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_546),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_550),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_530),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_558),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_537),
.Y(n_578)
);

BUFx10_ASAP7_75t_L g579 ( 
.A(n_550),
.Y(n_579)
);

BUFx2_ASAP7_75t_SL g580 ( 
.A(n_530),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_558),
.B(n_524),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_558),
.Y(n_582)
);

BUFx2_ASAP7_75t_SL g583 ( 
.A(n_557),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_538),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_526),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_545),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_532),
.B(n_540),
.Y(n_587)
);

BUFx4f_ASAP7_75t_SL g588 ( 
.A(n_552),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_550),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_545),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_538),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_543),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_528),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_528),
.Y(n_594)
);

CKINVDCx16_ASAP7_75t_R g595 ( 
.A(n_552),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_538),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_543),
.Y(n_597)
);

INVx8_ASAP7_75t_L g598 ( 
.A(n_566),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_549),
.Y(n_599)
);

AO21x2_ASAP7_75t_L g600 ( 
.A1(n_565),
.A2(n_529),
.B(n_563),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_538),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_566),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_560),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_549),
.Y(n_604)
);

OAI22xp33_ASAP7_75t_L g605 ( 
.A1(n_551),
.A2(n_541),
.B1(n_564),
.B2(n_539),
.Y(n_605)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_527),
.A2(n_534),
.B(n_553),
.Y(n_606)
);

AND2x2_ASAP7_75t_SL g607 ( 
.A(n_549),
.B(n_559),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_556),
.B(n_542),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_574),
.B(n_533),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_574),
.B(n_533),
.Y(n_610)
);

INVx8_ASAP7_75t_L g611 ( 
.A(n_573),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_580),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_R g613 ( 
.A(n_573),
.B(n_564),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_569),
.B(n_556),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_580),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_569),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_589),
.B(n_554),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_578),
.Y(n_618)
);

NAND2xp33_ASAP7_75t_R g619 ( 
.A(n_587),
.B(n_535),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_R g620 ( 
.A(n_589),
.B(n_534),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_577),
.B(n_542),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_575),
.Y(n_622)
);

NAND2xp33_ASAP7_75t_R g623 ( 
.A(n_589),
.B(n_544),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_578),
.B(n_562),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_577),
.B(n_562),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_570),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_582),
.B(n_575),
.Y(n_627)
);

CKINVDCx16_ASAP7_75t_R g628 ( 
.A(n_595),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_582),
.B(n_575),
.Y(n_629)
);

NAND2x1p5_ASAP7_75t_L g630 ( 
.A(n_576),
.B(n_575),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_575),
.B(n_602),
.Y(n_631)
);

XOR2x2_ASAP7_75t_L g632 ( 
.A(n_595),
.B(n_588),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_R g633 ( 
.A(n_602),
.B(n_579),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_570),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_585),
.B(n_590),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_585),
.B(n_605),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_586),
.B(n_590),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_R g638 ( 
.A(n_579),
.B(n_598),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_586),
.B(n_579),
.Y(n_639)
);

OR2x4_ASAP7_75t_L g640 ( 
.A(n_571),
.B(n_572),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_571),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_593),
.B(n_594),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_583),
.B(n_608),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_R g644 ( 
.A(n_579),
.B(n_598),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_598),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_625),
.B(n_581),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_643),
.B(n_608),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_626),
.B(n_634),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_645),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_626),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_641),
.B(n_581),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_634),
.B(n_584),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_640),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_616),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_618),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_636),
.B(n_583),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_635),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_621),
.B(n_596),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_637),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_627),
.B(n_596),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_614),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_624),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_613),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_642),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_642),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_609),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_610),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_627),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_629),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_617),
.B(n_607),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_631),
.B(n_572),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_617),
.B(n_607),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_648),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_650),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_658),
.B(n_591),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_648),
.Y(n_676)
);

AND2x4_ASAP7_75t_SL g677 ( 
.A(n_664),
.B(n_631),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_650),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_658),
.B(n_591),
.Y(n_679)
);

INVxp67_ASAP7_75t_SL g680 ( 
.A(n_654),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_646),
.B(n_601),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_655),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_653),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_653),
.B(n_629),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_647),
.B(n_670),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_666),
.B(n_607),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_682),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_685),
.B(n_667),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_681),
.B(n_660),
.Y(n_689)
);

NOR2x1p5_ASAP7_75t_L g690 ( 
.A(n_686),
.B(n_649),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_681),
.B(n_660),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_680),
.B(n_673),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_682),
.Y(n_693)
);

NAND2x1_ASAP7_75t_SL g694 ( 
.A(n_683),
.B(n_667),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_675),
.B(n_646),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_674),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_SL g697 ( 
.A(n_694),
.B(n_633),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_688),
.B(n_662),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_695),
.B(n_661),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_SL g700 ( 
.A(n_690),
.B(n_644),
.Y(n_700)
);

NOR4xp25_ASAP7_75t_SL g701 ( 
.A(n_687),
.B(n_619),
.C(n_620),
.D(n_623),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_697),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_699),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_698),
.B(n_695),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_700),
.B(n_692),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_701),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_699),
.Y(n_707)
);

NOR2x1_ASAP7_75t_L g708 ( 
.A(n_702),
.B(n_706),
.Y(n_708)
);

O2A1O1Ixp33_ASAP7_75t_SL g709 ( 
.A1(n_702),
.A2(n_663),
.B(n_615),
.C(n_612),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_703),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_705),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_708),
.B(n_707),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_710),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_711),
.B(n_628),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_713),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_712),
.Y(n_716)
);

INVxp33_ASAP7_75t_SL g717 ( 
.A(n_714),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_714),
.B(n_704),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_715),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_716),
.B(n_709),
.Y(n_720)
);

NOR2xp67_ASAP7_75t_L g721 ( 
.A(n_718),
.B(n_649),
.Y(n_721)
);

NAND3xp33_ASAP7_75t_L g722 ( 
.A(n_717),
.B(n_656),
.C(n_669),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_717),
.B(n_632),
.Y(n_723)
);

AOI211xp5_ASAP7_75t_L g724 ( 
.A1(n_716),
.A2(n_638),
.B(n_684),
.C(n_611),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_716),
.B(n_669),
.C(n_655),
.Y(n_725)
);

AOI211xp5_ASAP7_75t_L g726 ( 
.A1(n_721),
.A2(n_611),
.B(n_684),
.C(n_584),
.Y(n_726)
);

AOI222xp33_ASAP7_75t_L g727 ( 
.A1(n_723),
.A2(n_601),
.B1(n_684),
.B2(n_677),
.C1(n_696),
.C2(n_693),
.Y(n_727)
);

OAI31xp33_ASAP7_75t_L g728 ( 
.A1(n_720),
.A2(n_722),
.A3(n_719),
.B(n_725),
.Y(n_728)
);

OAI21xp5_ASAP7_75t_L g729 ( 
.A1(n_724),
.A2(n_630),
.B(n_676),
.Y(n_729)
);

AOI211x1_ASAP7_75t_SL g730 ( 
.A1(n_721),
.A2(n_593),
.B(n_594),
.C(n_674),
.Y(n_730)
);

NOR3xp33_ASAP7_75t_L g731 ( 
.A(n_723),
.B(n_672),
.C(n_668),
.Y(n_731)
);

NAND5xp2_ASAP7_75t_L g732 ( 
.A(n_724),
.B(n_691),
.C(n_689),
.D(n_639),
.E(n_651),
.Y(n_732)
);

AOI211xp5_ASAP7_75t_L g733 ( 
.A1(n_721),
.A2(n_622),
.B(n_671),
.C(n_659),
.Y(n_733)
);

XOR2x1_ASAP7_75t_L g734 ( 
.A(n_728),
.B(n_691),
.Y(n_734)
);

NOR2x1_ASAP7_75t_L g735 ( 
.A(n_732),
.B(n_689),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_731),
.Y(n_736)
);

NAND2x1p5_ASAP7_75t_L g737 ( 
.A(n_733),
.B(n_726),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_730),
.Y(n_738)
);

NOR2x1_ASAP7_75t_L g739 ( 
.A(n_729),
.B(n_678),
.Y(n_739)
);

XOR2xp5_ASAP7_75t_L g740 ( 
.A(n_727),
.B(n_622),
.Y(n_740)
);

NAND2x1p5_ASAP7_75t_L g741 ( 
.A(n_728),
.B(n_622),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_734),
.B(n_678),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_741),
.B(n_736),
.Y(n_743)
);

XNOR2x1_ASAP7_75t_L g744 ( 
.A(n_737),
.B(n_671),
.Y(n_744)
);

NOR3xp33_ASAP7_75t_SL g745 ( 
.A(n_738),
.B(n_659),
.C(n_598),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_SL g746 ( 
.A(n_740),
.B(n_679),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_R g747 ( 
.A(n_739),
.B(n_598),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_746),
.A2(n_735),
.B1(n_671),
.B2(n_677),
.Y(n_748)
);

AOI222xp33_ASAP7_75t_L g749 ( 
.A1(n_743),
.A2(n_742),
.B1(n_745),
.B2(n_744),
.C1(n_747),
.C2(n_597),
.Y(n_749)
);

NOR4xp25_ASAP7_75t_L g750 ( 
.A(n_743),
.B(n_679),
.C(n_675),
.D(n_652),
.Y(n_750)
);

AOI22x1_ASAP7_75t_L g751 ( 
.A1(n_743),
.A2(n_668),
.B1(n_657),
.B2(n_597),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_751),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_748),
.A2(n_657),
.B1(n_665),
.B2(n_592),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_752),
.Y(n_754)
);

XNOR2xp5_ASAP7_75t_L g755 ( 
.A(n_753),
.B(n_750),
.Y(n_755)
);

AOI31xp33_ASAP7_75t_L g756 ( 
.A1(n_754),
.A2(n_749),
.A3(n_665),
.B(n_651),
.Y(n_756)
);

NAND4xp25_ASAP7_75t_L g757 ( 
.A(n_756),
.B(n_755),
.C(n_597),
.D(n_592),
.Y(n_757)
);

OAI222xp33_ASAP7_75t_L g758 ( 
.A1(n_757),
.A2(n_652),
.B1(n_604),
.B2(n_592),
.C1(n_567),
.C2(n_599),
.Y(n_758)
);

INVxp67_ASAP7_75t_SL g759 ( 
.A(n_758),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_759),
.A2(n_567),
.B1(n_600),
.B2(n_603),
.Y(n_760)
);

AOI211xp5_ASAP7_75t_L g761 ( 
.A1(n_760),
.A2(n_606),
.B(n_604),
.C(n_568),
.Y(n_761)
);


endmodule