module fake_jpeg_137_n_216 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_216);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_35),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_10),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_2),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_30),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_84),
.B(n_57),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_86),
.Y(n_87)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_94),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_59),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_85),
.A2(n_86),
.B1(n_79),
.B2(n_74),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_77),
.B1(n_66),
.B2(n_65),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_81),
.A2(n_56),
.B1(n_69),
.B2(n_60),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_67),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_71),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_78),
.B1(n_68),
.B2(n_74),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_100),
.A2(n_113),
.B1(n_22),
.B2(n_46),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_65),
.C(n_75),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_76),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_98),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

AO22x1_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_60),
.B1(n_56),
.B2(n_68),
.Y(n_104)
);

OA21x2_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_55),
.B(n_1),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_81),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_78),
.B1(n_58),
.B2(n_77),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_112),
.B1(n_117),
.B2(n_106),
.Y(n_121)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_83),
.B(n_63),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_83),
.B(n_63),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_110),
.Y(n_131)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_66),
.B1(n_56),
.B2(n_76),
.Y(n_113)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_73),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_4),
.B(n_5),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_90),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_123),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_134),
.B1(n_136),
.B2(n_28),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_125),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_0),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_115),
.A2(n_72),
.B1(n_55),
.B2(n_3),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_140),
.B1(n_119),
.B2(n_126),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_132),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_112),
.A2(n_104),
.B1(n_115),
.B2(n_113),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_55),
.B1(n_1),
.B2(n_3),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_101),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_29),
.Y(n_162)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_146),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_21),
.C(n_44),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_150),
.C(n_33),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_143),
.A2(n_159),
.B1(n_131),
.B2(n_19),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_20),
.Y(n_173)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

AND2x4_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_152),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_23),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_124),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_156),
.B1(n_158),
.B2(n_18),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_120),
.B(n_24),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_6),
.B(n_7),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_8),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_163),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_140),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_128),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_12),
.B(n_15),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_160),
.A2(n_34),
.B(n_36),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_162),
.B(n_164),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_15),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_16),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g165 ( 
.A(n_145),
.B(n_17),
.CI(n_18),
.CON(n_165),
.SN(n_165)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_165),
.A2(n_182),
.B(n_151),
.Y(n_192)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_161),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_170),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_178),
.B1(n_179),
.B2(n_182),
.Y(n_184)
);

NOR2x1_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_19),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_173),
.B(n_179),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_25),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_142),
.C(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_177),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_154),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_192),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_150),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_186),
.B(n_190),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_153),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_166),
.C(n_181),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_SL g194 ( 
.A(n_183),
.B(n_181),
.C(n_165),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_199),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_196),
.C(n_191),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_174),
.C(n_180),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_172),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_198),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_185),
.A2(n_188),
.B1(n_176),
.B2(n_157),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_193),
.A2(n_176),
.B1(n_157),
.B2(n_158),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_176),
.B1(n_156),
.B2(n_186),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_204),
.Y(n_208)
);

NAND4xp25_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_207),
.C(n_194),
.D(n_203),
.Y(n_210)
);

BUFx24_ASAP7_75t_SL g207 ( 
.A(n_201),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_208),
.A2(n_205),
.B(n_187),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_SL g211 ( 
.A(n_209),
.B(n_210),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_204),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_202),
.B(n_200),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_200),
.C(n_39),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_214),
.A2(n_37),
.B(n_40),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_50),
.Y(n_216)
);


endmodule