module fake_jpeg_30312_n_86 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_86);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

AOI21xp33_ASAP7_75t_L g32 ( 
.A1(n_2),
.A2(n_28),
.B(n_31),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_3),
.B(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_27),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

HAxp5_ASAP7_75t_SL g44 ( 
.A(n_32),
.B(n_0),
.CON(n_44),
.SN(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_34),
.B(n_43),
.C(n_3),
.Y(n_56)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_49),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_32),
.B(n_40),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_56),
.B(n_59),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_52),
.B(n_54),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_42),
.C(n_38),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_55),
.C(n_56),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_45),
.A2(n_33),
.B1(n_36),
.B2(n_4),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_64)
);

OA21x2_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_43),
.B(n_2),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_1),
.B1(n_6),
.B2(n_7),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_64),
.B1(n_16),
.B2(n_17),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_66),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_8),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_67),
.A2(n_69),
.B(n_9),
.Y(n_72)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_68),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_73),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_68),
.A2(n_13),
.B(n_14),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_76),
.Y(n_78)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_18),
.C(n_21),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_81),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_77),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_75),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_84),
.A2(n_71),
.B1(n_81),
.B2(n_70),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_79),
.C(n_70),
.Y(n_86)
);


endmodule