module real_aes_10500_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1845;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1441;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1225;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1284;
wire n_1095;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_346;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1853;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_733;
wire n_402;
wire n_1404;
wire n_1856;
wire n_658;
wire n_676;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1855;
wire n_1056;
wire n_1802;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1790;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_1596;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1842;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_729;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
CKINVDCx5p33_ASAP7_75t_R g1207 ( .A(n_0), .Y(n_1207) );
AOI22xp5_ASAP7_75t_L g1593 ( .A1(n_1), .A2(n_333), .B1(n_1568), .B2(n_1572), .Y(n_1593) );
INVx1_ASAP7_75t_L g938 ( .A(n_2), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g1504 ( .A(n_3), .Y(n_1504) );
CKINVDCx5p33_ASAP7_75t_R g1530 ( .A(n_4), .Y(n_1530) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_5), .A2(n_92), .B1(n_432), .B2(n_440), .Y(n_431) );
INVx1_ASAP7_75t_L g533 ( .A(n_5), .Y(n_533) );
INVx1_ASAP7_75t_L g1443 ( .A(n_6), .Y(n_1443) );
AOI22xp33_ASAP7_75t_L g1458 ( .A1(n_6), .A2(n_102), .B1(n_857), .B2(n_1459), .Y(n_1458) );
OAI22xp33_ASAP7_75t_L g599 ( .A1(n_7), .A2(n_89), .B1(n_600), .B2(n_602), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_7), .A2(n_89), .B1(n_609), .B2(n_621), .C(n_623), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g917 ( .A1(n_8), .A2(n_257), .B1(n_574), .B2(n_577), .C(n_918), .Y(n_917) );
OAI22xp33_ASAP7_75t_L g926 ( .A1(n_8), .A2(n_99), .B1(n_751), .B2(n_753), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g1449 ( .A1(n_9), .A2(n_108), .B1(n_1006), .B2(n_1450), .Y(n_1449) );
AOI22xp33_ASAP7_75t_SL g1456 ( .A1(n_9), .A2(n_108), .B1(n_812), .B2(n_1246), .Y(n_1456) );
INVx1_ASAP7_75t_L g1110 ( .A(n_10), .Y(n_1110) );
OAI211xp5_ASAP7_75t_SL g1130 ( .A1(n_10), .A2(n_602), .B(n_1131), .C(n_1137), .Y(n_1130) );
AOI221xp5_ASAP7_75t_L g845 ( .A1(n_11), .A2(n_287), .B1(n_511), .B2(n_577), .C(n_738), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_11), .A2(n_287), .B1(n_857), .B2(n_858), .Y(n_856) );
INVx1_ASAP7_75t_L g789 ( .A(n_12), .Y(n_789) );
AOI22xp33_ASAP7_75t_SL g805 ( .A1(n_12), .A2(n_276), .B1(n_806), .B2(n_808), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g1104 ( .A(n_13), .Y(n_1104) );
OAI22xp33_ASAP7_75t_L g1054 ( .A1(n_14), .A2(n_65), .B1(n_432), .B2(n_440), .Y(n_1054) );
OAI22xp33_ASAP7_75t_L g1060 ( .A1(n_14), .A2(n_174), .B1(n_358), .B2(n_1040), .Y(n_1060) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_15), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g1594 ( .A1(n_16), .A2(n_293), .B1(n_1539), .B2(n_1585), .Y(n_1594) );
XNOR2xp5_ASAP7_75t_L g664 ( .A(n_17), .B(n_665), .Y(n_664) );
CKINVDCx16_ASAP7_75t_R g1610 ( .A(n_17), .Y(n_1610) );
INVx1_ASAP7_75t_L g1378 ( .A(n_18), .Y(n_1378) );
AOI22xp33_ASAP7_75t_L g1418 ( .A1(n_18), .A2(n_112), .B1(n_697), .B2(n_1080), .Y(n_1418) );
AOI22xp33_ASAP7_75t_SL g1451 ( .A1(n_19), .A2(n_84), .B1(n_1006), .B2(n_1452), .Y(n_1451) );
INVxp67_ASAP7_75t_SL g1471 ( .A(n_19), .Y(n_1471) );
INVx1_ASAP7_75t_L g1051 ( .A(n_20), .Y(n_1051) );
OAI222xp33_ASAP7_75t_L g1057 ( .A1(n_20), .A2(n_223), .B1(n_318), .B2(n_571), .C1(n_1058), .C2(n_1059), .Y(n_1057) );
OAI222xp33_ASAP7_75t_L g1199 ( .A1(n_21), .A2(n_63), .B1(n_134), .B2(n_989), .C1(n_1200), .C2(n_1203), .Y(n_1199) );
INVx1_ASAP7_75t_L g1220 ( .A(n_21), .Y(n_1220) );
CKINVDCx5p33_ASAP7_75t_R g1282 ( .A(n_22), .Y(n_1282) );
AOI22xp33_ASAP7_75t_SL g1002 ( .A1(n_23), .A2(n_123), .B1(n_803), .B2(n_1003), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_23), .A2(n_123), .B1(n_1013), .B2(n_1014), .Y(n_1012) );
AOI221xp5_ASAP7_75t_L g830 ( .A1(n_24), .A2(n_186), .B1(n_770), .B2(n_831), .C(n_832), .Y(n_830) );
INVx1_ASAP7_75t_L g865 ( .A(n_24), .Y(n_865) );
INVx1_ASAP7_75t_L g984 ( .A(n_25), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_25), .A2(n_321), .B1(n_736), .B2(n_738), .Y(n_1009) );
INVx1_ASAP7_75t_L g1483 ( .A(n_26), .Y(n_1483) );
AOI221xp5_ASAP7_75t_L g1511 ( .A1(n_26), .A2(n_147), .B1(n_1512), .B2(n_1513), .C(n_1514), .Y(n_1511) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_27), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g531 ( .A(n_27), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g1107 ( .A(n_28), .Y(n_1107) );
CKINVDCx5p33_ASAP7_75t_R g765 ( .A(n_29), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_30), .A2(n_141), .B1(n_1023), .B2(n_1024), .Y(n_1255) );
AOI22xp33_ASAP7_75t_SL g1272 ( .A1(n_30), .A2(n_141), .B1(n_776), .B2(n_1273), .Y(n_1272) );
INVx1_ASAP7_75t_L g349 ( .A(n_31), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_32), .A2(n_107), .B1(n_422), .B2(n_1053), .Y(n_1052) );
AOI22xp33_ASAP7_75t_SL g1071 ( .A1(n_32), .A2(n_107), .B1(n_1008), .B2(n_1013), .Y(n_1071) );
INVx1_ASAP7_75t_L g941 ( .A(n_33), .Y(n_941) );
OAI211xp5_ASAP7_75t_SL g963 ( .A1(n_33), .A2(n_602), .B(n_964), .C(n_969), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_34), .A2(n_146), .B1(n_828), .B2(n_829), .Y(n_827) );
INVx1_ASAP7_75t_L g866 ( .A(n_34), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g1589 ( .A1(n_35), .A2(n_144), .B1(n_1568), .B2(n_1572), .Y(n_1589) );
AOI22xp33_ASAP7_75t_L g1574 ( .A1(n_36), .A2(n_211), .B1(n_1537), .B2(n_1545), .Y(n_1574) );
INVxp67_ASAP7_75t_SL g1444 ( .A(n_37), .Y(n_1444) );
OAI22xp33_ASAP7_75t_L g1465 ( .A1(n_37), .A2(n_169), .B1(n_989), .B2(n_1200), .Y(n_1465) );
INVx1_ASAP7_75t_L g1849 ( .A(n_38), .Y(n_1849) );
AOI22xp33_ASAP7_75t_L g1877 ( .A1(n_38), .A2(n_205), .B1(n_736), .B2(n_1067), .Y(n_1877) );
INVx1_ASAP7_75t_L g1303 ( .A(n_39), .Y(n_1303) );
AOI22xp33_ASAP7_75t_L g1327 ( .A1(n_39), .A2(n_279), .B1(n_1328), .B2(n_1331), .Y(n_1327) );
INVx1_ASAP7_75t_L g1062 ( .A(n_40), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_40), .A2(n_220), .B1(n_682), .B2(n_1088), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g1874 ( .A1(n_41), .A2(n_135), .B1(n_1067), .B2(n_1229), .Y(n_1874) );
AOI22xp33_ASAP7_75t_L g1880 ( .A1(n_41), .A2(n_135), .B1(n_609), .B2(n_806), .Y(n_1880) );
INVx1_ASAP7_75t_L g1492 ( .A(n_42), .Y(n_1492) );
AOI22xp33_ASAP7_75t_L g1528 ( .A1(n_42), .A2(n_121), .B1(n_894), .B2(n_1080), .Y(n_1528) );
CKINVDCx5p33_ASAP7_75t_R g1386 ( .A(n_43), .Y(n_1386) );
AOI22x1_ASAP7_75t_SL g1042 ( .A1(n_44), .A2(n_1043), .B1(n_1089), .B2(n_1090), .Y(n_1042) );
INVx1_ASAP7_75t_L g1089 ( .A(n_44), .Y(n_1089) );
AO221x2_ASAP7_75t_L g1595 ( .A1(n_44), .A2(n_249), .B1(n_1539), .B2(n_1585), .C(n_1596), .Y(n_1595) );
AOI22xp5_ASAP7_75t_L g1583 ( .A1(n_45), .A2(n_125), .B1(n_1568), .B2(n_1572), .Y(n_1583) );
CKINVDCx16_ASAP7_75t_R g1611 ( .A(n_46), .Y(n_1611) );
XNOR2xp5_ASAP7_75t_L g1093 ( .A(n_47), .B(n_1094), .Y(n_1093) );
AOI22xp5_ASAP7_75t_SL g1578 ( .A1(n_47), .A2(n_228), .B1(n_1539), .B2(n_1545), .Y(n_1578) );
INVx1_ASAP7_75t_L g890 ( .A(n_48), .Y(n_890) );
OAI221xp5_ASAP7_75t_L g900 ( .A1(n_48), .A2(n_600), .B1(n_725), .B2(n_901), .C(n_907), .Y(n_900) );
INVx1_ASAP7_75t_L g1155 ( .A(n_49), .Y(n_1155) );
OAI221xp5_ASAP7_75t_L g1172 ( .A1(n_49), .A2(n_602), .B1(n_1173), .B2(n_1178), .C(n_1183), .Y(n_1172) );
OAI22xp33_ASAP7_75t_L g948 ( .A1(n_50), .A2(n_235), .B1(n_659), .B2(n_662), .Y(n_948) );
INVx1_ASAP7_75t_L g967 ( .A(n_50), .Y(n_967) );
INVx1_ASAP7_75t_L g996 ( .A(n_51), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_51), .A2(n_172), .B1(n_1006), .B2(n_1008), .Y(n_1005) );
INVx1_ASAP7_75t_L g734 ( .A(n_52), .Y(n_734) );
OAI22xp33_ASAP7_75t_L g748 ( .A1(n_52), .A2(n_122), .B1(n_662), .B2(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g1317 ( .A(n_53), .Y(n_1317) );
AOI22xp33_ASAP7_75t_L g1343 ( .A1(n_53), .A2(n_270), .B1(n_682), .B2(n_1088), .Y(n_1343) );
INVx1_ASAP7_75t_L g1319 ( .A(n_54), .Y(n_1319) );
AOI22xp33_ASAP7_75t_L g1342 ( .A1(n_54), .A2(n_302), .B1(n_1048), .B2(n_1080), .Y(n_1342) );
INVx1_ASAP7_75t_L g1224 ( .A(n_55), .Y(n_1224) );
AOI22xp33_ASAP7_75t_SL g1243 ( .A1(n_55), .A2(n_106), .B1(n_609), .B2(n_1244), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_56), .A2(n_343), .B1(n_682), .B2(n_684), .Y(n_681) );
INVx1_ASAP7_75t_L g715 ( .A(n_56), .Y(n_715) );
CKINVDCx14_ASAP7_75t_R g1555 ( .A(n_57), .Y(n_1555) );
INVx1_ASAP7_75t_L g560 ( .A(n_58), .Y(n_560) );
AOI221xp5_ASAP7_75t_L g608 ( .A1(n_58), .A2(n_242), .B1(n_609), .B2(n_611), .C(n_614), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_59), .B(n_824), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g1102 ( .A(n_60), .Y(n_1102) );
OAI22xp33_ASAP7_75t_L g761 ( .A1(n_61), .A2(n_306), .B1(n_708), .B2(n_709), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_61), .A2(n_306), .B1(n_482), .B2(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g1308 ( .A(n_62), .Y(n_1308) );
OAI22xp5_ASAP7_75t_L g1313 ( .A1(n_62), .A2(n_320), .B1(n_1032), .B2(n_1314), .Y(n_1313) );
AOI22xp33_ASAP7_75t_SL g1228 ( .A1(n_63), .A2(n_296), .B1(n_1016), .B2(n_1229), .Y(n_1228) );
AOI22xp33_ASAP7_75t_L g1873 ( .A1(n_64), .A2(n_182), .B1(n_1006), .B2(n_1182), .Y(n_1873) );
AOI22xp33_ASAP7_75t_L g1879 ( .A1(n_64), .A2(n_182), .B1(n_697), .B2(n_1246), .Y(n_1879) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_65), .A2(n_131), .B1(n_1067), .B2(n_1073), .Y(n_1072) );
CKINVDCx5p33_ASAP7_75t_R g1149 ( .A(n_66), .Y(n_1149) );
AOI21xp33_ASAP7_75t_L g1799 ( .A1(n_67), .A2(n_1084), .B(n_1411), .Y(n_1799) );
INVxp33_ASAP7_75t_L g1816 ( .A(n_67), .Y(n_1816) );
AOI22xp33_ASAP7_75t_L g1567 ( .A1(n_68), .A2(n_193), .B1(n_1568), .B2(n_1571), .Y(n_1567) );
AOI22xp33_ASAP7_75t_SL g1066 ( .A1(n_69), .A2(n_138), .B1(n_577), .B2(n_1067), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_69), .A2(n_138), .B1(n_1080), .B2(n_1081), .Y(n_1079) );
OAI22xp33_ASAP7_75t_L g1117 ( .A1(n_70), .A2(n_334), .B1(n_896), .B2(n_897), .Y(n_1117) );
INVx1_ASAP7_75t_L g1139 ( .A(n_70), .Y(n_1139) );
INVx1_ASAP7_75t_L g1174 ( .A(n_71), .Y(n_1174) );
OAI22xp33_ASAP7_75t_L g1187 ( .A1(n_71), .A2(n_160), .B1(n_659), .B2(n_662), .Y(n_1187) );
INVx1_ASAP7_75t_L g945 ( .A(n_72), .Y(n_945) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_72), .A2(n_218), .B1(n_589), .B2(n_595), .Y(n_953) );
CKINVDCx5p33_ASAP7_75t_R g1396 ( .A(n_73), .Y(n_1396) );
INVx1_ASAP7_75t_L g1850 ( .A(n_74), .Y(n_1850) );
AOI22xp33_ASAP7_75t_L g1876 ( .A1(n_74), .A2(n_159), .B1(n_905), .B2(n_1006), .Y(n_1876) );
INVx1_ASAP7_75t_L g1481 ( .A(n_75), .Y(n_1481) );
AOI22xp33_ASAP7_75t_L g1516 ( .A1(n_75), .A2(n_210), .B1(n_1517), .B2(n_1518), .Y(n_1516) );
CKINVDCx20_ASAP7_75t_R g1790 ( .A(n_76), .Y(n_1790) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_77), .Y(n_677) );
INVx1_ASAP7_75t_L g1116 ( .A(n_78), .Y(n_1116) );
OAI22xp5_ASAP7_75t_L g1121 ( .A1(n_78), .A2(n_288), .B1(n_589), .B2(n_595), .Y(n_1121) );
CKINVDCx14_ASAP7_75t_R g1597 ( .A(n_79), .Y(n_1597) );
XNOR2x2_ASAP7_75t_L g548 ( .A(n_80), .B(n_549), .Y(n_548) );
INVxp67_ASAP7_75t_SL g1438 ( .A(n_81), .Y(n_1438) );
AOI22xp33_ASAP7_75t_L g1461 ( .A1(n_81), .A2(n_248), .B1(n_894), .B2(n_1246), .Y(n_1461) );
OAI221xp5_ASAP7_75t_L g1488 ( .A1(n_82), .A2(n_111), .B1(n_1363), .B2(n_1368), .C(n_1489), .Y(n_1488) );
OAI22xp5_ASAP7_75t_L g1519 ( .A1(n_82), .A2(n_111), .B1(n_1405), .B2(n_1520), .Y(n_1519) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_83), .Y(n_576) );
INVxp33_ASAP7_75t_L g1470 ( .A(n_84), .Y(n_1470) );
BUFx2_ASAP7_75t_L g374 ( .A(n_85), .Y(n_374) );
BUFx2_ASAP7_75t_L g472 ( .A(n_85), .Y(n_472) );
INVx1_ASAP7_75t_L g543 ( .A(n_85), .Y(n_543) );
OR2x2_ASAP7_75t_L g1367 ( .A(n_85), .B(n_587), .Y(n_1367) );
AOI22xp33_ASAP7_75t_SL g1069 ( .A1(n_86), .A2(n_231), .B1(n_1008), .B2(n_1070), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_86), .A2(n_231), .B1(n_1077), .B2(n_1078), .Y(n_1076) );
CKINVDCx5p33_ASAP7_75t_R g1389 ( .A(n_87), .Y(n_1389) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_88), .A2(n_329), .B1(n_609), .B2(n_806), .Y(n_1001) );
AOI22xp33_ASAP7_75t_SL g1015 ( .A1(n_88), .A2(n_329), .B1(n_736), .B2(n_1016), .Y(n_1015) );
CKINVDCx5p33_ASAP7_75t_R g1355 ( .A(n_90), .Y(n_1355) );
CKINVDCx5p33_ASAP7_75t_R g1787 ( .A(n_91), .Y(n_1787) );
INVx1_ASAP7_75t_L g411 ( .A(n_92), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g1325 ( .A1(n_93), .A2(n_340), .B1(n_1070), .B2(n_1326), .Y(n_1325) );
AOI22xp33_ASAP7_75t_SL g1336 ( .A1(n_93), .A2(n_340), .B1(n_1337), .B2(n_1338), .Y(n_1336) );
AOI221xp5_ASAP7_75t_L g1802 ( .A1(n_94), .A2(n_219), .B1(n_1525), .B2(n_1803), .C(n_1804), .Y(n_1802) );
INVxp67_ASAP7_75t_SL g1826 ( .A(n_94), .Y(n_1826) );
INVx1_ASAP7_75t_L g1179 ( .A(n_95), .Y(n_1179) );
OAI22xp33_ASAP7_75t_L g1188 ( .A1(n_95), .A2(n_183), .B1(n_751), .B2(n_753), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_96), .A2(n_149), .B1(n_987), .B2(n_989), .Y(n_986) );
OAI22xp33_ASAP7_75t_L g1030 ( .A1(n_96), .A2(n_149), .B1(n_1031), .B2(n_1032), .Y(n_1030) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_97), .Y(n_558) );
INVx1_ASAP7_75t_L g1158 ( .A(n_98), .Y(n_1158) );
OAI22xp5_ASAP7_75t_L g1163 ( .A1(n_98), .A2(n_103), .B1(n_589), .B2(n_595), .Y(n_1163) );
INVx1_ASAP7_75t_L g914 ( .A(n_99), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g1453 ( .A1(n_100), .A2(n_190), .B1(n_736), .B2(n_1454), .Y(n_1453) );
INVxp67_ASAP7_75t_SL g1464 ( .A(n_100), .Y(n_1464) );
INVx1_ASAP7_75t_L g1305 ( .A(n_101), .Y(n_1305) );
AOI22xp33_ASAP7_75t_L g1332 ( .A1(n_101), .A2(n_119), .B1(n_1219), .B2(n_1333), .Y(n_1332) );
INVxp33_ASAP7_75t_L g1440 ( .A(n_102), .Y(n_1440) );
INVx1_ASAP7_75t_L g1157 ( .A(n_103), .Y(n_1157) );
AO221x1_ASAP7_75t_L g1277 ( .A1(n_104), .A2(n_185), .B1(n_573), .B2(n_574), .C(n_1017), .Y(n_1277) );
INVx1_ASAP7_75t_L g1286 ( .A(n_104), .Y(n_1286) );
INVx1_ASAP7_75t_L g1215 ( .A(n_105), .Y(n_1215) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_105), .A2(n_207), .B1(n_1024), .B2(n_1246), .Y(n_1245) );
INVx1_ASAP7_75t_L g1218 ( .A(n_106), .Y(n_1218) );
XNOR2x2_ASAP7_75t_L g1295 ( .A(n_109), .B(n_1296), .Y(n_1295) );
AO22x2_ASAP7_75t_L g1194 ( .A1(n_110), .A2(n_1195), .B1(n_1196), .B2(n_1247), .Y(n_1194) );
INVxp67_ASAP7_75t_SL g1195 ( .A(n_110), .Y(n_1195) );
INVx1_ASAP7_75t_L g1382 ( .A(n_112), .Y(n_1382) );
INVx1_ASAP7_75t_L g940 ( .A(n_113), .Y(n_940) );
OAI221xp5_ASAP7_75t_L g954 ( .A1(n_113), .A2(n_600), .B1(n_955), .B2(n_958), .C(n_962), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g1256 ( .A1(n_114), .A2(n_273), .B1(n_806), .B2(n_1257), .Y(n_1256) );
AOI221xp5_ASAP7_75t_L g1274 ( .A1(n_114), .A2(n_273), .B1(n_511), .B2(n_577), .C(n_918), .Y(n_1274) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_115), .A2(n_188), .B1(n_1229), .B2(n_1237), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g1239 ( .A1(n_115), .A2(n_188), .B1(n_609), .B2(n_806), .Y(n_1239) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_116), .A2(n_181), .B1(n_638), .B2(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g743 ( .A(n_116), .Y(n_743) );
INVx1_ASAP7_75t_L g1152 ( .A(n_117), .Y(n_1152) );
CKINVDCx5p33_ASAP7_75t_R g884 ( .A(n_118), .Y(n_884) );
INVx1_ASAP7_75t_L g1299 ( .A(n_119), .Y(n_1299) );
OA22x2_ASAP7_75t_L g371 ( .A1(n_120), .A2(n_372), .B1(n_546), .B2(n_547), .Y(n_371) );
INVxp67_ASAP7_75t_SL g547 ( .A(n_120), .Y(n_547) );
INVx1_ASAP7_75t_L g1501 ( .A(n_121), .Y(n_1501) );
AOI221xp5_ASAP7_75t_L g735 ( .A1(n_122), .A2(n_294), .B1(n_574), .B2(n_736), .C(n_737), .Y(n_735) );
CKINVDCx5p33_ASAP7_75t_R g777 ( .A(n_124), .Y(n_777) );
INVx1_ASAP7_75t_L g1865 ( .A(n_126), .Y(n_1865) );
AOI22xp33_ASAP7_75t_SL g1882 ( .A1(n_126), .A2(n_303), .B1(n_609), .B2(n_1244), .Y(n_1882) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_127), .A2(n_151), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
INVx1_ASAP7_75t_L g1035 ( .A(n_127), .Y(n_1035) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_128), .Y(n_568) );
INVx1_ASAP7_75t_L g787 ( .A(n_129), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_129), .A2(n_280), .B1(n_803), .B2(n_804), .Y(n_802) );
INVx1_ASAP7_75t_L g729 ( .A(n_130), .Y(n_729) );
OAI22xp33_ASAP7_75t_L g750 ( .A1(n_130), .A2(n_294), .B1(n_751), .B2(n_753), .Y(n_750) );
INVx1_ASAP7_75t_L g1047 ( .A(n_131), .Y(n_1047) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_132), .Y(n_412) );
AOI22xp5_ASAP7_75t_SL g1577 ( .A1(n_133), .A2(n_155), .B1(n_1568), .B2(n_1572), .Y(n_1577) );
INVx1_ASAP7_75t_L g1222 ( .A(n_134), .Y(n_1222) );
INVx1_ASAP7_75t_L g1543 ( .A(n_136), .Y(n_1543) );
OAI22xp33_ASAP7_75t_L g895 ( .A1(n_137), .A2(n_322), .B1(n_896), .B2(n_897), .Y(n_895) );
INVx1_ASAP7_75t_L g920 ( .A(n_137), .Y(n_920) );
INVx1_ASAP7_75t_L g1860 ( .A(n_139), .Y(n_1860) );
AOI22xp33_ASAP7_75t_L g1883 ( .A1(n_139), .A2(n_180), .B1(n_654), .B2(n_697), .Y(n_1883) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_140), .A2(n_339), .B1(n_696), .B2(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g903 ( .A(n_140), .Y(n_903) );
CKINVDCx16_ASAP7_75t_R g1607 ( .A(n_142), .Y(n_1607) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_143), .A2(n_297), .B1(n_733), .B2(n_828), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_143), .A2(n_297), .B1(n_616), .B2(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g794 ( .A(n_145), .Y(n_794) );
INVx1_ASAP7_75t_L g862 ( .A(n_146), .Y(n_862) );
INVx1_ASAP7_75t_L g1485 ( .A(n_147), .Y(n_1485) );
INVx1_ASAP7_75t_L g1441 ( .A(n_148), .Y(n_1441) );
INVx1_ASAP7_75t_L g1379 ( .A(n_150), .Y(n_1379) );
AOI221xp5_ASAP7_75t_L g1413 ( .A1(n_150), .A2(n_195), .B1(n_616), .B2(n_1414), .C(n_1416), .Y(n_1413) );
INVx1_ASAP7_75t_L g1036 ( .A(n_151), .Y(n_1036) );
INVx1_ASAP7_75t_L g935 ( .A(n_152), .Y(n_935) );
INVx1_ASAP7_75t_L g1541 ( .A(n_153), .Y(n_1541) );
NAND2xp5_ASAP7_75t_L g1560 ( .A(n_153), .B(n_1554), .Y(n_1560) );
INVx1_ASAP7_75t_L g891 ( .A(n_154), .Y(n_891) );
OAI211xp5_ASAP7_75t_SL g911 ( .A1(n_154), .A2(n_602), .B(n_912), .C(n_919), .Y(n_911) );
INVx1_ASAP7_75t_L g1358 ( .A(n_156), .Y(n_1358) );
AOI21xp33_ASAP7_75t_L g1410 ( .A1(n_156), .A2(n_1261), .B(n_1411), .Y(n_1410) );
INVx2_ASAP7_75t_L g361 ( .A(n_157), .Y(n_361) );
INVx1_ASAP7_75t_L g1360 ( .A(n_158), .Y(n_1360) );
AOI22xp33_ASAP7_75t_L g1409 ( .A1(n_158), .A2(n_215), .B1(n_686), .B2(n_696), .Y(n_1409) );
INVx1_ASAP7_75t_L g1853 ( .A(n_159), .Y(n_1853) );
INVx1_ASAP7_75t_L g1180 ( .A(n_160), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1232 ( .A1(n_161), .A2(n_261), .B1(n_1013), .B2(n_1233), .Y(n_1232) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_161), .A2(n_261), .B1(n_1024), .B2(n_1241), .Y(n_1240) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_162), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_163), .A2(n_335), .B1(n_694), .B2(n_697), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_163), .A2(n_335), .B1(n_708), .B2(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g430 ( .A(n_164), .Y(n_430) );
BUFx3_ASAP7_75t_L g446 ( .A(n_164), .Y(n_446) );
INVx1_ASAP7_75t_L g916 ( .A(n_165), .Y(n_916) );
OAI22xp33_ASAP7_75t_L g925 ( .A1(n_165), .A2(n_257), .B1(n_662), .B2(n_749), .Y(n_925) );
INVx1_ASAP7_75t_L g844 ( .A(n_166), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_166), .A2(n_251), .B1(n_642), .B2(n_647), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_167), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g1280 ( .A(n_168), .Y(n_1280) );
INVx1_ASAP7_75t_L g1445 ( .A(n_169), .Y(n_1445) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_170), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_171), .A2(n_309), .B1(n_589), .B2(n_595), .Y(n_588) );
INVx1_ASAP7_75t_L g627 ( .A(n_171), .Y(n_627) );
INVx1_ASAP7_75t_L g998 ( .A(n_172), .Y(n_998) );
OAI221xp5_ASAP7_75t_L g1854 ( .A1(n_173), .A2(n_241), .B1(n_989), .B2(n_1855), .C(n_1856), .Y(n_1854) );
INVx1_ASAP7_75t_L g1863 ( .A(n_173), .Y(n_1863) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_174), .A2(n_223), .B1(n_1083), .B2(n_1085), .Y(n_1082) );
CKINVDCx5p33_ASAP7_75t_R g1265 ( .A(n_175), .Y(n_1265) );
OAI221xp5_ASAP7_75t_SL g1791 ( .A1(n_176), .A2(n_330), .B1(n_1792), .B2(n_1793), .C(n_1795), .Y(n_1791) );
OAI221xp5_ASAP7_75t_L g1818 ( .A1(n_176), .A2(n_330), .B1(n_1369), .B2(n_1489), .C(n_1819), .Y(n_1818) );
AOI22xp33_ASAP7_75t_SL g1262 ( .A1(n_177), .A2(n_341), .B1(n_654), .B2(n_812), .Y(n_1262) );
INVx1_ASAP7_75t_L g1269 ( .A(n_177), .Y(n_1269) );
CKINVDCx5p33_ASAP7_75t_R g1506 ( .A(n_178), .Y(n_1506) );
AOI221xp5_ASAP7_75t_L g1136 ( .A1(n_179), .A2(n_342), .B1(n_577), .B2(n_738), .C(n_770), .Y(n_1136) );
OAI22xp33_ASAP7_75t_L g1142 ( .A1(n_179), .A2(n_281), .B1(n_751), .B2(n_753), .Y(n_1142) );
INVx1_ASAP7_75t_L g1861 ( .A(n_180), .Y(n_1861) );
INVx1_ASAP7_75t_L g740 ( .A(n_181), .Y(n_740) );
INVx1_ASAP7_75t_L g1177 ( .A(n_183), .Y(n_1177) );
CKINVDCx5p33_ASAP7_75t_R g768 ( .A(n_184), .Y(n_768) );
INVx1_ASAP7_75t_L g1288 ( .A(n_185), .Y(n_1288) );
INVx1_ASAP7_75t_L g863 ( .A(n_186), .Y(n_863) );
INVx1_ASAP7_75t_L g1808 ( .A(n_187), .Y(n_1808) );
INVx1_ASAP7_75t_L g470 ( .A(n_189), .Y(n_470) );
INVx1_ASAP7_75t_L g636 ( .A(n_189), .Y(n_636) );
INVxp33_ASAP7_75t_L g1467 ( .A(n_190), .Y(n_1467) );
OAI22xp33_ASAP7_75t_L g949 ( .A1(n_191), .A2(n_267), .B1(n_751), .B2(n_753), .Y(n_949) );
AOI221xp5_ASAP7_75t_L g968 ( .A1(n_191), .A2(n_235), .B1(n_574), .B2(n_910), .C(n_918), .Y(n_968) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_192), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g1548 ( .A(n_194), .Y(n_1548) );
INVx1_ASAP7_75t_L g1381 ( .A(n_195), .Y(n_1381) );
CKINVDCx5p33_ASAP7_75t_R g1503 ( .A(n_196), .Y(n_1503) );
INVx1_ASAP7_75t_L g841 ( .A(n_197), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_197), .A2(n_246), .B1(n_616), .B2(n_686), .Y(n_860) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_198), .Y(n_779) );
XOR2x2_ASAP7_75t_L g758 ( .A(n_199), .B(n_759), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g1258 ( .A1(n_200), .A2(n_317), .B1(n_609), .B2(n_1259), .Y(n_1258) );
OAI221xp5_ASAP7_75t_L g1276 ( .A1(n_200), .A2(n_602), .B1(n_1277), .B2(n_1278), .C(n_1281), .Y(n_1276) );
INVx1_ASAP7_75t_L g1109 ( .A(n_201), .Y(n_1109) );
OAI221xp5_ASAP7_75t_L g1122 ( .A1(n_201), .A2(n_600), .B1(n_725), .B2(n_1123), .C(n_1129), .Y(n_1122) );
CKINVDCx5p33_ASAP7_75t_R g1507 ( .A(n_202), .Y(n_1507) );
CKINVDCx5p33_ASAP7_75t_R g994 ( .A(n_203), .Y(n_994) );
XOR2xp5_ASAP7_75t_L g1476 ( .A(n_204), .B(n_1477), .Y(n_1476) );
INVx1_ASAP7_75t_L g1857 ( .A(n_205), .Y(n_1857) );
INVx1_ASAP7_75t_L g1494 ( .A(n_206), .Y(n_1494) );
AOI221xp5_ASAP7_75t_L g1523 ( .A1(n_206), .A2(n_224), .B1(n_1337), .B2(n_1524), .C(n_1525), .Y(n_1523) );
INVx1_ASAP7_75t_L g1214 ( .A(n_207), .Y(n_1214) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_208), .Y(n_581) );
OAI221xp5_ASAP7_75t_L g628 ( .A1(n_208), .A2(n_629), .B1(n_637), .B2(n_638), .C(n_641), .Y(n_628) );
CKINVDCx5p33_ASAP7_75t_R g1384 ( .A(n_209), .Y(n_1384) );
INVx1_ASAP7_75t_L g1486 ( .A(n_210), .Y(n_1486) );
CKINVDCx14_ASAP7_75t_R g1598 ( .A(n_212), .Y(n_1598) );
OAI22xp5_ASAP7_75t_L g835 ( .A1(n_213), .A2(n_237), .B1(n_745), .B2(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g870 ( .A(n_213), .Y(n_870) );
INVx1_ASAP7_75t_L g1161 ( .A(n_214), .Y(n_1161) );
INVx1_ASAP7_75t_L g1351 ( .A(n_215), .Y(n_1351) );
INVx1_ASAP7_75t_L g871 ( .A(n_216), .Y(n_871) );
CKINVDCx5p33_ASAP7_75t_R g937 ( .A(n_217), .Y(n_937) );
INVx1_ASAP7_75t_L g943 ( .A(n_218), .Y(n_943) );
INVx1_ASAP7_75t_L g1824 ( .A(n_219), .Y(n_1824) );
INVx1_ASAP7_75t_L g1063 ( .A(n_220), .Y(n_1063) );
CKINVDCx5p33_ASAP7_75t_R g774 ( .A(n_221), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g1805 ( .A1(n_222), .A2(n_299), .B1(n_886), .B2(n_1341), .Y(n_1805) );
INVx1_ASAP7_75t_L g1823 ( .A(n_222), .Y(n_1823) );
INVx1_ASAP7_75t_L g1498 ( .A(n_224), .Y(n_1498) );
CKINVDCx5p33_ASAP7_75t_R g1852 ( .A(n_225), .Y(n_1852) );
OAI22xp33_ASAP7_75t_L g1159 ( .A1(n_226), .A2(n_315), .B1(n_896), .B2(n_897), .Y(n_1159) );
INVx1_ASAP7_75t_L g1185 ( .A(n_226), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g1324 ( .A1(n_227), .A2(n_307), .B1(n_1028), .B2(n_1073), .Y(n_1324) );
AOI22xp33_ASAP7_75t_SL g1340 ( .A1(n_227), .A2(n_307), .B1(n_1048), .B2(n_1341), .Y(n_1340) );
INVx1_ASAP7_75t_L g692 ( .A(n_229), .Y(n_692) );
OAI211xp5_ASAP7_75t_SL g726 ( .A1(n_229), .A2(n_602), .B(n_727), .C(n_739), .Y(n_726) );
CKINVDCx16_ASAP7_75t_R g1433 ( .A(n_230), .Y(n_1433) );
INVx1_ASAP7_75t_L g877 ( .A(n_232), .Y(n_877) );
INVx1_ASAP7_75t_L g689 ( .A(n_233), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g710 ( .A1(n_233), .A2(n_600), .B1(n_711), .B2(n_720), .C(n_725), .Y(n_710) );
INVx1_ASAP7_75t_L g1154 ( .A(n_234), .Y(n_1154) );
OAI221xp5_ASAP7_75t_L g1164 ( .A1(n_234), .A2(n_600), .B1(n_725), .B2(n_1165), .C(n_1169), .Y(n_1164) );
INVx1_ASAP7_75t_L g933 ( .A(n_236), .Y(n_933) );
INVx1_ASAP7_75t_L g868 ( .A(n_237), .Y(n_868) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_238), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_239), .A2(n_263), .B1(n_379), .B2(n_387), .Y(n_378) );
INVx1_ASAP7_75t_L g503 ( .A(n_239), .Y(n_503) );
INVx1_ASAP7_75t_L g882 ( .A(n_240), .Y(n_882) );
AOI21xp33_ASAP7_75t_L g909 ( .A1(n_240), .A2(n_511), .B(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g1864 ( .A(n_241), .Y(n_1864) );
AOI21xp33_ASAP7_75t_L g562 ( .A1(n_242), .A2(n_511), .B(n_563), .Y(n_562) );
CKINVDCx5p33_ASAP7_75t_R g676 ( .A(n_243), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g1798 ( .A1(n_244), .A2(n_260), .B1(n_686), .B2(n_696), .Y(n_1798) );
INVxp33_ASAP7_75t_L g1817 ( .A(n_244), .Y(n_1817) );
OAI221xp5_ASAP7_75t_L g762 ( .A1(n_245), .A2(n_602), .B1(n_763), .B2(n_772), .C(n_778), .Y(n_762) );
AOI22xp33_ASAP7_75t_SL g810 ( .A1(n_245), .A2(n_316), .B1(n_621), .B2(n_808), .Y(n_810) );
INVx1_ASAP7_75t_L g842 ( .A(n_246), .Y(n_842) );
OAI211xp5_ASAP7_75t_L g393 ( .A1(n_247), .A2(n_394), .B(n_399), .C(n_406), .Y(n_393) );
INVx1_ASAP7_75t_L g499 ( .A(n_247), .Y(n_499) );
INVx1_ASAP7_75t_L g1437 ( .A(n_248), .Y(n_1437) );
XNOR2xp5_ASAP7_75t_L g874 ( .A(n_250), .B(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g834 ( .A(n_251), .Y(n_834) );
INVx1_ASAP7_75t_L g1148 ( .A(n_252), .Y(n_1148) );
AOI22xp33_ASAP7_75t_SL g892 ( .A1(n_253), .A2(n_282), .B1(n_893), .B2(n_894), .Y(n_892) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_253), .A2(n_282), .B1(n_708), .B2(n_709), .Y(n_899) );
CKINVDCx20_ASAP7_75t_R g1606 ( .A(n_254), .Y(n_1606) );
BUFx3_ASAP7_75t_L g429 ( .A(n_255), .Y(n_429) );
INVx1_ASAP7_75t_L g439 ( .A(n_255), .Y(n_439) );
AO221x2_ASAP7_75t_L g1536 ( .A1(n_256), .A2(n_323), .B1(n_1537), .B2(n_1544), .C(n_1547), .Y(n_1536) );
INVx1_ASAP7_75t_L g951 ( .A(n_258), .Y(n_951) );
CKINVDCx5p33_ASAP7_75t_R g1264 ( .A(n_259), .Y(n_1264) );
INVxp33_ASAP7_75t_L g1814 ( .A(n_260), .Y(n_1814) );
AOI22xp5_ASAP7_75t_L g1584 ( .A1(n_262), .A2(n_265), .B1(n_1539), .B2(n_1585), .Y(n_1584) );
INVx1_ASAP7_75t_L g501 ( .A(n_263), .Y(n_501) );
XNOR2xp5_ASAP7_75t_L g928 ( .A(n_264), .B(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g1832 ( .A(n_265), .Y(n_1832) );
AOI22xp33_ASAP7_75t_L g1838 ( .A1(n_265), .A2(n_1839), .B1(n_1843), .B2(n_1884), .Y(n_1838) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_266), .Y(n_357) );
INVx1_ASAP7_75t_L g545 ( .A(n_266), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_266), .B(n_325), .Y(n_587) );
AND2x2_ASAP7_75t_L g591 ( .A(n_266), .B(n_383), .Y(n_591) );
INVx1_ASAP7_75t_L g966 ( .A(n_267), .Y(n_966) );
CKINVDCx5p33_ASAP7_75t_R g1279 ( .A(n_268), .Y(n_1279) );
AOI21xp33_ASAP7_75t_L g572 ( .A1(n_269), .A2(n_573), .B(n_574), .Y(n_572) );
INVx1_ASAP7_75t_L g652 ( .A(n_269), .Y(n_652) );
INVx1_ASAP7_75t_L g1316 ( .A(n_270), .Y(n_1316) );
XNOR2xp5_ASAP7_75t_L g979 ( .A(n_271), .B(n_980), .Y(n_979) );
INVx2_ASAP7_75t_L g426 ( .A(n_272), .Y(n_426) );
OR2x2_ASAP7_75t_L g651 ( .A(n_272), .B(n_636), .Y(n_651) );
XNOR2xp5_ASAP7_75t_L g1844 ( .A(n_274), .B(n_1845), .Y(n_1844) );
CKINVDCx5p33_ASAP7_75t_R g1100 ( .A(n_275), .Y(n_1100) );
INVx1_ASAP7_75t_L g792 ( .A(n_276), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_277), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_278), .Y(n_480) );
INVx1_ASAP7_75t_L g1300 ( .A(n_279), .Y(n_1300) );
INVx1_ASAP7_75t_L g784 ( .A(n_280), .Y(n_784) );
INVx1_ASAP7_75t_L g1132 ( .A(n_281), .Y(n_1132) );
INVx1_ASAP7_75t_L g1801 ( .A(n_283), .Y(n_1801) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_284), .Y(n_566) );
INVx1_ASAP7_75t_L g1135 ( .A(n_285), .Y(n_1135) );
OAI22xp33_ASAP7_75t_L g1141 ( .A1(n_285), .A2(n_342), .B1(n_659), .B2(n_662), .Y(n_1141) );
INVx1_ASAP7_75t_L g1346 ( .A(n_286), .Y(n_1346) );
AOI22xp5_ASAP7_75t_SL g1590 ( .A1(n_286), .A2(n_290), .B1(n_1539), .B2(n_1545), .Y(n_1590) );
INVx1_ASAP7_75t_L g1113 ( .A(n_288), .Y(n_1113) );
INVx1_ASAP7_75t_L g1210 ( .A(n_289), .Y(n_1210) );
AOI22xp33_ASAP7_75t_L g1230 ( .A1(n_289), .A2(n_300), .B1(n_1006), .B2(n_1127), .Y(n_1230) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_291), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_292), .A2(n_308), .B1(n_609), .B2(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g1038 ( .A(n_292), .Y(n_1038) );
AOI22x1_ASAP7_75t_L g1249 ( .A1(n_295), .A2(n_1250), .B1(n_1251), .B2(n_1289), .Y(n_1249) );
INVxp67_ASAP7_75t_SL g1289 ( .A(n_295), .Y(n_1289) );
INVx1_ASAP7_75t_L g1206 ( .A(n_296), .Y(n_1206) );
AOI22xp33_ASAP7_75t_L g1448 ( .A1(n_298), .A2(n_337), .B1(n_736), .B2(n_737), .Y(n_1448) );
AOI22xp33_ASAP7_75t_L g1457 ( .A1(n_298), .A2(n_337), .B1(n_451), .B2(n_806), .Y(n_1457) );
INVx1_ASAP7_75t_L g1827 ( .A(n_299), .Y(n_1827) );
INVx1_ASAP7_75t_L g1209 ( .A(n_300), .Y(n_1209) );
CKINVDCx5p33_ASAP7_75t_R g1388 ( .A(n_301), .Y(n_1388) );
INVx1_ASAP7_75t_L g1312 ( .A(n_302), .Y(n_1312) );
INVx1_ASAP7_75t_L g1870 ( .A(n_303), .Y(n_1870) );
CKINVDCx5p33_ASAP7_75t_R g1302 ( .A(n_304), .Y(n_1302) );
OAI22xp33_ASAP7_75t_L g946 ( .A1(n_305), .A2(n_328), .B1(n_896), .B2(n_897), .Y(n_946) );
INVx1_ASAP7_75t_L g972 ( .A(n_305), .Y(n_972) );
INVx1_ASAP7_75t_L g1027 ( .A(n_308), .Y(n_1027) );
INVx1_ASAP7_75t_L g624 ( .A(n_309), .Y(n_624) );
INVx1_ASAP7_75t_L g1796 ( .A(n_310), .Y(n_1796) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_311), .Y(n_351) );
AND3x2_ASAP7_75t_L g1542 ( .A(n_311), .B(n_349), .C(n_1543), .Y(n_1542) );
NAND2xp5_ASAP7_75t_L g1552 ( .A(n_311), .B(n_349), .Y(n_1552) );
CKINVDCx5p33_ASAP7_75t_R g1119 ( .A(n_312), .Y(n_1119) );
INVx2_ASAP7_75t_L g362 ( .A(n_313), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g1151 ( .A(n_314), .Y(n_1151) );
INVx1_ASAP7_75t_L g1184 ( .A(n_315), .Y(n_1184) );
OAI221xp5_ASAP7_75t_L g781 ( .A1(n_316), .A2(n_600), .B1(n_725), .B2(n_782), .C(n_788), .Y(n_781) );
INVx1_ASAP7_75t_L g1275 ( .A(n_317), .Y(n_1275) );
CKINVDCx5p33_ASAP7_75t_R g1050 ( .A(n_318), .Y(n_1050) );
XNOR2xp5_ASAP7_75t_L g1143 ( .A(n_319), .B(n_1144), .Y(n_1143) );
INVx1_ASAP7_75t_L g1306 ( .A(n_320), .Y(n_1306) );
INVx1_ASAP7_75t_L g991 ( .A(n_321), .Y(n_991) );
INVx1_ASAP7_75t_L g921 ( .A(n_322), .Y(n_921) );
OAI221xp5_ASAP7_75t_L g1362 ( .A1(n_324), .A2(n_326), .B1(n_1363), .B2(n_1368), .C(n_1370), .Y(n_1362) );
OAI221xp5_ASAP7_75t_L g1401 ( .A1(n_324), .A2(n_326), .B1(n_1402), .B2(n_1405), .C(n_1407), .Y(n_1401) );
INVx1_ASAP7_75t_L g364 ( .A(n_325), .Y(n_364) );
INVx2_ASAP7_75t_L g383 ( .A(n_325), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_327), .Y(n_377) );
INVx1_ASAP7_75t_L g970 ( .A(n_328), .Y(n_970) );
INVx1_ASAP7_75t_L g580 ( .A(n_331), .Y(n_580) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_331), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g448 ( .A1(n_332), .A2(n_449), .B(n_454), .C(n_465), .Y(n_448) );
INVx1_ASAP7_75t_L g538 ( .A(n_332), .Y(n_538) );
INVx1_ASAP7_75t_L g1138 ( .A(n_334), .Y(n_1138) );
INVx1_ASAP7_75t_L g1807 ( .A(n_336), .Y(n_1807) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_338), .Y(n_780) );
INVx1_ASAP7_75t_L g906 ( .A(n_339), .Y(n_906) );
INVx1_ASAP7_75t_L g1270 ( .A(n_341), .Y(n_1270) );
INVx1_ASAP7_75t_L g719 ( .A(n_343), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_365), .B(n_1533), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_347), .B(n_352), .Y(n_346) );
AND2x4_ASAP7_75t_L g1837 ( .A(n_347), .B(n_353), .Y(n_1837) );
NOR2xp33_ASAP7_75t_SL g347 ( .A(n_348), .B(n_350), .Y(n_347) );
INVx1_ASAP7_75t_SL g1842 ( .A(n_348), .Y(n_1842) );
NAND2xp5_ASAP7_75t_L g1890 ( .A(n_348), .B(n_350), .Y(n_1890) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g1841 ( .A(n_350), .B(n_1842), .Y(n_1841) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_354), .B(n_358), .Y(n_353) );
INVxp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g373 ( .A(n_355), .B(n_374), .Y(n_373) );
OR2x6_ASAP7_75t_L g1041 ( .A(n_355), .B(n_374), .Y(n_1041) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g724 ( .A(n_356), .B(n_364), .Y(n_724) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g511 ( .A(n_357), .B(n_382), .Y(n_511) );
INVx8_ASAP7_75t_L g376 ( .A(n_358), .Y(n_376) );
OR2x6_ASAP7_75t_L g358 ( .A(n_359), .B(n_363), .Y(n_358) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_359), .Y(n_513) );
BUFx2_ASAP7_75t_L g961 ( .A(n_359), .Y(n_961) );
OR2x6_ASAP7_75t_L g1040 ( .A(n_359), .B(n_381), .Y(n_1040) );
INVx2_ASAP7_75t_SL g1171 ( .A(n_359), .Y(n_1171) );
INVx1_ASAP7_75t_L g1176 ( .A(n_359), .Y(n_1176) );
INVx2_ASAP7_75t_SL g1377 ( .A(n_359), .Y(n_1377) );
OR2x2_ASAP7_75t_L g1394 ( .A(n_359), .B(n_1367), .Y(n_1394) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx2_ASAP7_75t_L g386 ( .A(n_361), .Y(n_386) );
AND2x4_ASAP7_75t_L g391 ( .A(n_361), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g398 ( .A(n_361), .Y(n_398) );
INVx1_ASAP7_75t_L g405 ( .A(n_361), .Y(n_405) );
AND2x2_ASAP7_75t_L g410 ( .A(n_361), .B(n_362), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_362), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g392 ( .A(n_362), .Y(n_392) );
INVx1_ASAP7_75t_L g397 ( .A(n_362), .Y(n_397) );
INVx1_ASAP7_75t_L g414 ( .A(n_362), .Y(n_414) );
INVx1_ASAP7_75t_L g594 ( .A(n_362), .Y(n_594) );
AND2x4_ASAP7_75t_L g413 ( .A(n_363), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_364), .B(n_417), .Y(n_1032) );
OR2x2_ASAP7_75t_L g1059 ( .A(n_364), .B(n_417), .Y(n_1059) );
OAI22xp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_1290), .B1(n_1291), .B2(n_1532), .Y(n_365) );
INVx1_ASAP7_75t_L g1532 ( .A(n_366), .Y(n_1532) );
XNOR2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_976), .Y(n_366) );
XOR2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_755), .Y(n_367) );
XNOR2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_663), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
XNOR2x1_ASAP7_75t_L g370 ( .A(n_371), .B(n_548), .Y(n_370) );
INVx1_ASAP7_75t_L g546 ( .A(n_372), .Y(n_546) );
OAI211xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_375), .B(n_420), .C(n_473), .Y(n_372) );
AND2x4_ASAP7_75t_L g506 ( .A(n_374), .B(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_L g655 ( .A(n_374), .B(n_656), .Y(n_655) );
AND2x4_ASAP7_75t_L g815 ( .A(n_374), .B(n_507), .Y(n_815) );
AOI211xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B(n_378), .C(n_393), .Y(n_375) );
AOI22xp33_ASAP7_75t_SL g1037 ( .A1(n_376), .A2(n_994), .B1(n_1038), .B2(n_1039), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_376), .A2(n_1039), .B1(n_1207), .B2(n_1224), .Y(n_1223) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_376), .A2(n_1302), .B1(n_1319), .B2(n_1320), .Y(n_1318) );
AOI22xp33_ASAP7_75t_L g1439 ( .A1(n_376), .A2(n_1320), .B1(n_1440), .B2(n_1441), .Y(n_1439) );
AOI22xp33_ASAP7_75t_L g1869 ( .A1(n_376), .A2(n_1320), .B1(n_1852), .B2(n_1870), .Y(n_1869) );
OAI22xp33_ASAP7_75t_L g496 ( .A1(n_377), .A2(n_490), .B1(n_497), .B2(n_499), .Y(n_496) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_384), .Y(n_379) );
AOI322xp5_ASAP7_75t_L g406 ( .A1(n_380), .A2(n_407), .A3(n_411), .B1(n_412), .B2(n_413), .C1(n_415), .C2(n_419), .Y(n_406) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x4_ASAP7_75t_L g388 ( .A(n_381), .B(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g1034 ( .A(n_381), .B(n_592), .Y(n_1034) );
AND2x4_ASAP7_75t_L g1216 ( .A(n_381), .B(n_389), .Y(n_1216) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g403 ( .A(n_383), .Y(n_403) );
INVx2_ASAP7_75t_L g519 ( .A(n_384), .Y(n_519) );
BUFx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g526 ( .A(n_385), .Y(n_526) );
INVx1_ASAP7_75t_L g554 ( .A(n_385), .Y(n_554) );
INVx1_ASAP7_75t_L g583 ( .A(n_386), .Y(n_583) );
AND2x4_ASAP7_75t_L g592 ( .A(n_386), .B(n_593), .Y(n_592) );
INVx5_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
AOI22xp33_ASAP7_75t_SL g1033 ( .A1(n_388), .A2(n_1034), .B1(n_1035), .B2(n_1036), .Y(n_1033) );
AOI22xp5_ASAP7_75t_L g1061 ( .A1(n_388), .A2(n_1034), .B1(n_1062), .B2(n_1063), .Y(n_1061) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g1168 ( .A(n_390), .Y(n_1168) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g522 ( .A(n_391), .Y(n_522) );
INVx3_ASAP7_75t_L g530 ( .A(n_391), .Y(n_530) );
BUFx6f_ASAP7_75t_L g776 ( .A(n_391), .Y(n_776) );
AND2x4_ASAP7_75t_L g404 ( .A(n_392), .B(n_405), .Y(n_404) );
OAI22xp33_ASAP7_75t_L g1375 ( .A1(n_394), .A2(n_1376), .B1(n_1378), .B2(n_1379), .Y(n_1375) );
OAI22xp33_ASAP7_75t_L g1387 ( .A1(n_394), .A2(n_721), .B1(n_1388), .B2(n_1389), .Y(n_1387) );
OAI22xp33_ASAP7_75t_L g1821 ( .A1(n_394), .A2(n_1822), .B1(n_1823), .B2(n_1824), .Y(n_1821) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g516 ( .A(n_396), .Y(n_516) );
INVx3_ASAP7_75t_L g561 ( .A(n_396), .Y(n_561) );
INVx2_ASAP7_75t_L g571 ( .A(n_396), .Y(n_571) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_397), .B(n_398), .Y(n_537) );
INVx1_ASAP7_75t_L g417 ( .A(n_398), .Y(n_417) );
NAND4xp25_ASAP7_75t_SL g1212 ( .A(n_399), .B(n_1213), .C(n_1217), .D(n_1223), .Y(n_1212) );
NAND4xp25_ASAP7_75t_SL g1435 ( .A(n_399), .B(n_1436), .C(n_1439), .D(n_1442), .Y(n_1435) );
NAND4xp25_ASAP7_75t_SL g1858 ( .A(n_399), .B(n_1859), .C(n_1862), .D(n_1869), .Y(n_1858) );
CKINVDCx11_ASAP7_75t_R g399 ( .A(n_400), .Y(n_399) );
AOI211xp5_ASAP7_75t_L g1026 ( .A1(n_400), .A2(n_1027), .B(n_1028), .C(n_1030), .Y(n_1026) );
NOR3xp33_ASAP7_75t_L g1056 ( .A(n_400), .B(n_1057), .C(n_1060), .Y(n_1056) );
AOI211xp5_ASAP7_75t_L g1311 ( .A1(n_400), .A2(n_1067), .B(n_1312), .C(n_1313), .Y(n_1311) );
AND2x4_ASAP7_75t_L g400 ( .A(n_401), .B(n_404), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g418 ( .A(n_402), .Y(n_418) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2x1p5_ASAP7_75t_L g544 ( .A(n_403), .B(n_545), .Y(n_544) );
BUFx3_ASAP7_75t_L g604 ( .A(n_404), .Y(n_604) );
BUFx6f_ASAP7_75t_L g738 ( .A(n_404), .Y(n_738) );
BUFx3_ASAP7_75t_L g918 ( .A(n_404), .Y(n_918) );
BUFx6f_ASAP7_75t_L g1017 ( .A(n_404), .Y(n_1017) );
BUFx2_ASAP7_75t_L g1868 ( .A(n_404), .Y(n_1868) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g1229 ( .A(n_408), .Y(n_1229) );
INVx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_409), .Y(n_577) );
AND2x4_ASAP7_75t_L g601 ( .A(n_409), .B(n_591), .Y(n_601) );
BUFx2_ASAP7_75t_L g831 ( .A(n_409), .Y(n_831) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g564 ( .A(n_410), .Y(n_564) );
AOI322xp5_ASAP7_75t_L g454 ( .A1(n_412), .A2(n_419), .A3(n_455), .B1(n_457), .B2(n_458), .C1(n_459), .C2(n_463), .Y(n_454) );
INVx2_ASAP7_75t_L g1031 ( .A(n_413), .Y(n_1031) );
INVx2_ASAP7_75t_L g1058 ( .A(n_413), .Y(n_1058) );
INVx2_ASAP7_75t_L g1314 ( .A(n_413), .Y(n_1314) );
AOI222xp33_ASAP7_75t_L g1862 ( .A1(n_413), .A2(n_415), .B1(n_1863), .B2(n_1864), .C1(n_1865), .C2(n_1866), .Y(n_1862) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_414), .A2(n_580), .B1(n_581), .B2(n_582), .Y(n_579) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_414), .Y(n_742) );
INVx1_ASAP7_75t_L g838 ( .A(n_414), .Y(n_838) );
AOI222xp33_ASAP7_75t_L g1217 ( .A1(n_415), .A2(n_1218), .B1(n_1219), .B2(n_1220), .C1(n_1221), .C2(n_1222), .Y(n_1217) );
AOI222xp33_ASAP7_75t_L g1442 ( .A1(n_415), .A2(n_1219), .B1(n_1221), .B2(n_1443), .C1(n_1444), .C2(n_1445), .Y(n_1442) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g1284 ( .A1(n_416), .A2(n_837), .B1(n_1264), .B2(n_1265), .Y(n_1284) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI31xp33_ASAP7_75t_SL g420 ( .A1(n_421), .A2(n_431), .A3(n_448), .B(n_468), .Y(n_420) );
INVx4_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_423), .A2(n_996), .B1(n_997), .B2(n_998), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_423), .A2(n_997), .B1(n_1209), .B2(n_1210), .Y(n_1208) );
AOI22xp33_ASAP7_75t_L g1301 ( .A1(n_423), .A2(n_441), .B1(n_1302), .B2(n_1303), .Y(n_1301) );
AOI22xp33_ASAP7_75t_L g1469 ( .A1(n_423), .A2(n_997), .B1(n_1470), .B2(n_1471), .Y(n_1469) );
AOI22xp33_ASAP7_75t_L g1848 ( .A1(n_423), .A2(n_992), .B1(n_1849), .B2(n_1850), .Y(n_1848) );
AND2x6_ASAP7_75t_L g423 ( .A(n_424), .B(n_427), .Y(n_423) );
AND2x4_ASAP7_75t_L g992 ( .A(n_424), .B(n_993), .Y(n_992) );
AND2x4_ASAP7_75t_L g1468 ( .A(n_424), .B(n_993), .Y(n_1468) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_425), .B(n_1202), .Y(n_1201) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g435 ( .A(n_426), .Y(n_435) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_426), .Y(n_443) );
AND2x2_ASAP7_75t_L g477 ( .A(n_426), .B(n_470), .Y(n_477) );
INVx2_ASAP7_75t_L g508 ( .A(n_426), .Y(n_508) );
INVx1_ASAP7_75t_L g504 ( .A(n_427), .Y(n_504) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_427), .Y(n_812) );
BUFx6f_ASAP7_75t_L g886 ( .A(n_427), .Y(n_886) );
BUFx6f_ASAP7_75t_L g894 ( .A(n_427), .Y(n_894) );
INVx2_ASAP7_75t_L g1339 ( .A(n_427), .Y(n_1339) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g487 ( .A(n_428), .Y(n_487) );
INVx1_ASAP7_75t_L g617 ( .A(n_428), .Y(n_617) );
INVx1_ASAP7_75t_L g660 ( .A(n_428), .Y(n_660) );
BUFx6f_ASAP7_75t_L g686 ( .A(n_428), .Y(n_686) );
AND2x4_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx2_ASAP7_75t_L g447 ( .A(n_429), .Y(n_447) );
AND2x2_ASAP7_75t_L g453 ( .A(n_429), .B(n_446), .Y(n_453) );
INVx1_ASAP7_75t_L g437 ( .A(n_430), .Y(n_437) );
OR2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g457 ( .A(n_433), .Y(n_457) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g450 ( .A(n_434), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g467 ( .A(n_434), .Y(n_467) );
AND2x6_ASAP7_75t_L g997 ( .A(n_434), .B(n_456), .Y(n_997) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AND2x6_ASAP7_75t_L g463 ( .A(n_435), .B(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g491 ( .A(n_436), .Y(n_491) );
INVx1_ASAP7_75t_L g675 ( .A(n_436), .Y(n_675) );
BUFx2_ASAP7_75t_L g881 ( .A(n_436), .Y(n_881) );
OR2x2_ASAP7_75t_L g1426 ( .A(n_436), .B(n_651), .Y(n_1426) );
OR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
AND2x2_ASAP7_75t_L g495 ( .A(n_437), .B(n_438), .Y(n_495) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g456 ( .A(n_439), .B(n_446), .Y(n_456) );
INVx4_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_441), .A2(n_991), .B1(n_992), .B2(n_994), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g1205 ( .A1(n_441), .A2(n_992), .B1(n_1206), .B2(n_1207), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g1466 ( .A1(n_441), .A2(n_1441), .B1(n_1467), .B2(n_1468), .Y(n_1466) );
AOI221xp5_ASAP7_75t_L g1851 ( .A1(n_441), .A2(n_997), .B1(n_1852), .B2(n_1853), .C(n_1854), .Y(n_1851) );
AND2x4_ASAP7_75t_L g441 ( .A(n_442), .B(n_444), .Y(n_441) );
AND2x2_ASAP7_75t_SL g459 ( .A(n_442), .B(n_460), .Y(n_459) );
AND2x4_ASAP7_75t_L g988 ( .A(n_442), .B(n_460), .Y(n_988) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx6_ASAP7_75t_L g613 ( .A(n_444), .Y(n_613) );
INVx2_ASAP7_75t_L g648 ( .A(n_444), .Y(n_648) );
AND2x2_ASAP7_75t_L g656 ( .A(n_444), .B(n_634), .Y(n_656) );
BUFx2_ASAP7_75t_L g857 ( .A(n_444), .Y(n_857) );
AND2x4_ASAP7_75t_L g444 ( .A(n_445), .B(n_447), .Y(n_444) );
INVx1_ASAP7_75t_L g464 ( .A(n_445), .Y(n_464) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g462 ( .A(n_447), .Y(n_462) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI211xp5_ASAP7_75t_L g1463 ( .A1(n_450), .A2(n_466), .B(n_1464), .C(n_1465), .Y(n_1463) );
HB1xp67_ASAP7_75t_L g985 ( .A(n_451), .Y(n_985) );
HB1xp67_ASAP7_75t_L g1513 ( .A(n_451), .Y(n_1513) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g466 ( .A(n_452), .B(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g610 ( .A(n_452), .Y(n_610) );
INVx1_ASAP7_75t_L g670 ( .A(n_452), .Y(n_670) );
BUFx6f_ASAP7_75t_L g1086 ( .A(n_452), .Y(n_1086) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_453), .Y(n_643) );
INVx2_ASAP7_75t_L g483 ( .A(n_455), .Y(n_483) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_SL g502 ( .A(n_456), .Y(n_502) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_456), .Y(n_616) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_456), .Y(n_683) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_456), .Y(n_696) );
BUFx3_ASAP7_75t_L g893 ( .A(n_456), .Y(n_893) );
BUFx2_ASAP7_75t_L g1241 ( .A(n_456), .Y(n_1241) );
BUFx2_ASAP7_75t_L g1246 ( .A(n_456), .Y(n_1246) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_458), .A2(n_524), .B1(n_527), .B2(n_531), .Y(n_523) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g1202 ( .A(n_461), .Y(n_1202) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g631 ( .A(n_462), .Y(n_631) );
INVx3_ASAP7_75t_L g989 ( .A(n_463), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_463), .A2(n_988), .B1(n_1050), .B2(n_1051), .Y(n_1049) );
AOI222xp33_ASAP7_75t_L g1304 ( .A1(n_463), .A2(n_1257), .B1(n_1305), .B2(n_1306), .C1(n_1307), .C2(n_1308), .Y(n_1304) );
BUFx3_ASAP7_75t_L g640 ( .A(n_464), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g1045 ( .A(n_465), .B(n_1046), .C(n_1049), .Y(n_1045) );
CKINVDCx8_ASAP7_75t_R g465 ( .A(n_466), .Y(n_465) );
AOI211xp5_ASAP7_75t_L g983 ( .A1(n_466), .A2(n_984), .B(n_985), .C(n_986), .Y(n_983) );
NOR2xp33_ASAP7_75t_L g1198 ( .A(n_466), .B(n_1199), .Y(n_1198) );
INVx5_ASAP7_75t_L g1309 ( .A(n_466), .Y(n_1309) );
OAI21xp33_ASAP7_75t_L g1856 ( .A1(n_467), .A2(n_1086), .B(n_1857), .Y(n_1856) );
OAI31xp33_ASAP7_75t_L g1044 ( .A1(n_468), .A2(n_1045), .A3(n_1052), .B(n_1054), .Y(n_1044) );
INVx1_ASAP7_75t_SL g1472 ( .A(n_468), .Y(n_1472) );
AND2x4_ASAP7_75t_L g468 ( .A(n_469), .B(n_471), .Y(n_468) );
AND2x4_ASAP7_75t_L g981 ( .A(n_469), .B(n_471), .Y(n_981) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x4_ASAP7_75t_L g507 ( .A(n_470), .B(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g923 ( .A(n_471), .Y(n_923) );
BUFx2_ASAP7_75t_L g1810 ( .A(n_471), .Y(n_1810) );
BUFx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g478 ( .A(n_472), .Y(n_478) );
OR2x6_ASAP7_75t_L g510 ( .A(n_472), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_509), .Y(n_473) );
OAI33xp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_479), .A3(n_488), .B1(n_496), .B2(n_500), .B3(n_505), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_475), .A2(n_880), .B1(n_887), .B2(n_889), .Y(n_879) );
OAI33xp33_ASAP7_75t_L g931 ( .A1(n_475), .A2(n_505), .A3(n_932), .B1(n_936), .B2(n_939), .B3(n_942), .Y(n_931) );
OAI33xp33_ASAP7_75t_L g1097 ( .A1(n_475), .A2(n_505), .A3(n_1098), .B1(n_1103), .B2(n_1108), .B3(n_1111), .Y(n_1097) );
OAI33xp33_ASAP7_75t_L g1146 ( .A1(n_475), .A2(n_505), .A3(n_1147), .B1(n_1150), .B2(n_1153), .B3(n_1156), .Y(n_1146) );
INVx1_ASAP7_75t_SL g1254 ( .A(n_475), .Y(n_1254) );
OR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_478), .Y(n_475) );
OR2x6_ASAP7_75t_L g619 ( .A(n_476), .B(n_478), .Y(n_619) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g853 ( .A(n_477), .Y(n_853) );
BUFx3_ASAP7_75t_L g1417 ( .A(n_477), .Y(n_1417) );
INVx2_ASAP7_75t_SL g1527 ( .A(n_477), .Y(n_1527) );
INVx2_ASAP7_75t_L g606 ( .A(n_478), .Y(n_606) );
BUFx2_ASAP7_75t_L g746 ( .A(n_478), .Y(n_746) );
OAI31xp33_ASAP7_75t_L g760 ( .A1(n_478), .A2(n_761), .A3(n_762), .B(n_781), .Y(n_760) );
OR2x2_ASAP7_75t_L g852 ( .A(n_478), .B(n_853), .Y(n_852) );
AND2x4_ASAP7_75t_L g1018 ( .A(n_478), .B(n_724), .Y(n_1018) );
AND2x4_ASAP7_75t_L g1065 ( .A(n_478), .B(n_724), .Y(n_1065) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_484), .B2(n_485), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_480), .A2(n_484), .B1(n_518), .B2(n_520), .Y(n_517) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_483), .A2(n_624), .B1(n_625), .B2(n_627), .Y(n_623) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g626 ( .A(n_487), .Y(n_626) );
OR2x2_ASAP7_75t_L g1428 ( .A(n_487), .B(n_651), .Y(n_1428) );
OAI22xp33_ASAP7_75t_SL g488 ( .A1(n_489), .A2(n_490), .B1(n_492), .B2(n_493), .Y(n_488) );
OAI22xp33_ASAP7_75t_L g512 ( .A1(n_489), .A2(n_492), .B1(n_513), .B2(n_514), .Y(n_512) );
OAI22xp33_ASAP7_75t_L g936 ( .A1(n_490), .A2(n_690), .B1(n_937), .B2(n_938), .Y(n_936) );
OAI22xp33_ASAP7_75t_L g939 ( .A1(n_490), .A2(n_883), .B1(n_940), .B2(n_941), .Y(n_939) );
OAI22xp33_ASAP7_75t_L g1153 ( .A1(n_490), .A2(n_497), .B1(n_1154), .B2(n_1155), .Y(n_1153) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g688 ( .A(n_491), .Y(n_688) );
INVx1_ASAP7_75t_L g752 ( .A(n_491), .Y(n_752) );
OAI221xp5_ASAP7_75t_L g889 ( .A1(n_493), .A2(n_881), .B1(n_890), .B2(n_891), .C(n_892), .Y(n_889) );
BUFx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g691 ( .A(n_494), .Y(n_691) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g498 ( .A(n_495), .Y(n_498) );
BUFx4f_ASAP7_75t_L g680 ( .A(n_495), .Y(n_680) );
INVx1_ASAP7_75t_L g1106 ( .A(n_495), .Y(n_1106) );
OAI22xp33_ASAP7_75t_L g1150 ( .A1(n_497), .A2(n_881), .B1(n_1151), .B2(n_1152), .Y(n_1150) );
BUFx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OR2x6_ASAP7_75t_L g662 ( .A(n_498), .B(n_650), .Y(n_662) );
OAI22xp33_ASAP7_75t_L g1108 ( .A1(n_498), .A2(n_674), .B1(n_1109), .B2(n_1110), .Y(n_1108) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B1(n_503), .B2(n_504), .Y(n_500) );
INVx2_ASAP7_75t_L g654 ( .A(n_502), .Y(n_654) );
INVx1_ASAP7_75t_L g1023 ( .A(n_502), .Y(n_1023) );
OAI22xp5_ASAP7_75t_SL g671 ( .A1(n_505), .A2(n_619), .B1(n_672), .B2(n_687), .Y(n_671) );
INVx4_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AOI221xp5_ASAP7_75t_L g607 ( .A1(n_506), .A2(n_608), .B1(n_618), .B2(n_620), .C(n_628), .Y(n_607) );
BUFx4f_ASAP7_75t_L g888 ( .A(n_506), .Y(n_888) );
AOI33xp33_ASAP7_75t_L g1074 ( .A1(n_506), .A2(n_1075), .A3(n_1076), .B1(n_1079), .B2(n_1082), .B3(n_1087), .Y(n_1074) );
BUFx4f_ASAP7_75t_L g1344 ( .A(n_506), .Y(n_1344) );
CKINVDCx5p33_ASAP7_75t_R g1411 ( .A(n_507), .Y(n_1411) );
INVx2_ASAP7_75t_L g1515 ( .A(n_507), .Y(n_1515) );
AND2x4_ASAP7_75t_L g634 ( .A(n_508), .B(n_635), .Y(n_634) );
OAI33xp33_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_512), .A3(n_517), .B1(n_523), .B2(n_532), .B3(n_539), .Y(n_509) );
INVx1_ASAP7_75t_L g1374 ( .A(n_510), .Y(n_1374) );
OAI33xp33_ASAP7_75t_L g1490 ( .A1(n_510), .A2(n_1390), .A3(n_1491), .B1(n_1497), .B2(n_1502), .B3(n_1505), .Y(n_1490) );
OAI33xp33_ASAP7_75t_L g1820 ( .A1(n_510), .A2(n_1390), .A3(n_1821), .B1(n_1825), .B2(n_1828), .B3(n_1830), .Y(n_1820) );
OAI22xp33_ASAP7_75t_L g532 ( .A1(n_513), .A2(n_533), .B1(n_534), .B2(n_538), .Y(n_532) );
BUFx2_ASAP7_75t_L g721 ( .A(n_513), .Y(n_721) );
INVx1_ASAP7_75t_L g767 ( .A(n_513), .Y(n_767) );
INVx1_ASAP7_75t_L g791 ( .A(n_513), .Y(n_791) );
OAI221xp5_ASAP7_75t_L g1129 ( .A1(n_513), .A2(n_536), .B1(n_722), .B2(n_1104), .C(n_1107), .Y(n_1129) );
OAI221xp5_ASAP7_75t_L g788 ( .A1(n_514), .A2(n_722), .B1(n_789), .B2(n_790), .C(n_792), .Y(n_788) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_516), .B(n_579), .Y(n_578) );
OR2x6_ASAP7_75t_L g725 ( .A(n_516), .B(n_585), .Y(n_725) );
OR2x2_ASAP7_75t_L g962 ( .A(n_516), .B(n_585), .Y(n_962) );
OAI221xp5_ASAP7_75t_L g1131 ( .A1(n_518), .A2(n_1132), .B1(n_1133), .B2(n_1135), .C(n_1136), .Y(n_1131) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g1014 ( .A(n_520), .Y(n_1014) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x4_ASAP7_75t_L g596 ( .A(n_521), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g733 ( .A(n_522), .Y(n_733) );
INVx2_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g902 ( .A(n_525), .Y(n_902) );
INVx2_ASAP7_75t_L g913 ( .A(n_525), .Y(n_913) );
INVx2_ASAP7_75t_L g965 ( .A(n_525), .Y(n_965) );
BUFx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g714 ( .A(n_526), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g1380 ( .A1(n_527), .A2(n_712), .B1(n_1381), .B2(n_1382), .Y(n_1380) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g786 ( .A(n_529), .Y(n_786) );
INVx2_ASAP7_75t_L g905 ( .A(n_529), .Y(n_905) );
INVx2_ASAP7_75t_L g1134 ( .A(n_529), .Y(n_1134) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx3_ASAP7_75t_L g557 ( .A(n_530), .Y(n_557) );
INVx3_ASAP7_75t_L g1235 ( .A(n_530), .Y(n_1235) );
OAI221xp5_ASAP7_75t_L g1173 ( .A1(n_534), .A2(n_769), .B1(n_1174), .B2(n_1175), .C(n_1177), .Y(n_1173) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g764 ( .A(n_535), .Y(n_764) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx3_ASAP7_75t_L g908 ( .A(n_536), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g1283 ( .A(n_536), .B(n_1284), .Y(n_1283) );
BUFx3_ASAP7_75t_L g1496 ( .A(n_536), .Y(n_1496) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AOI33xp33_ASAP7_75t_L g1064 ( .A1(n_540), .A2(n_1065), .A3(n_1066), .B1(n_1069), .B2(n_1071), .B3(n_1072), .Y(n_1064) );
AOI33xp33_ASAP7_75t_L g1322 ( .A1(n_540), .A2(n_1323), .A3(n_1324), .B1(n_1325), .B2(n_1327), .B3(n_1332), .Y(n_1322) );
AOI33xp33_ASAP7_75t_L g1447 ( .A1(n_540), .A2(n_1065), .A3(n_1448), .B1(n_1449), .B2(n_1451), .B3(n_1453), .Y(n_1447) );
INVx6_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx5_ASAP7_75t_L g1010 ( .A(n_541), .Y(n_1010) );
OR2x6_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .Y(n_541) );
NAND2x1p5_ASAP7_75t_L g633 ( .A(n_542), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g650 ( .A(n_543), .B(n_651), .Y(n_650) );
AND2x4_ASAP7_75t_L g1354 ( .A(n_543), .B(n_591), .Y(n_1354) );
BUFx2_ASAP7_75t_L g574 ( .A(n_544), .Y(n_574) );
INVx2_ASAP7_75t_L g771 ( .A(n_544), .Y(n_771) );
NAND4xp25_ASAP7_75t_L g549 ( .A(n_550), .B(n_607), .C(n_645), .D(n_657), .Y(n_549) );
OAI31xp33_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_588), .A3(n_599), .B(n_605), .Y(n_550) );
OAI221xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_559), .B1(n_565), .B2(n_569), .C(n_575), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_555), .B1(n_556), .B2(n_558), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_553), .A2(n_566), .B1(n_567), .B2(n_568), .Y(n_565) );
BUFx2_ASAP7_75t_L g773 ( .A(n_553), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g1278 ( .A1(n_553), .A2(n_567), .B1(n_1279), .B2(n_1280), .Y(n_1278) );
OAI22xp5_ASAP7_75t_L g1825 ( .A1(n_553), .A2(n_1385), .B1(n_1826), .B2(n_1827), .Y(n_1825) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
HB1xp67_ASAP7_75t_L g1125 ( .A(n_554), .Y(n_1125) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_555), .A2(n_558), .B1(n_615), .B2(n_617), .Y(n_614) );
INVx2_ASAP7_75t_SL g1182 ( .A(n_556), .Y(n_1182) );
INVx2_ASAP7_75t_L g1452 ( .A(n_556), .Y(n_1452) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g567 ( .A(n_557), .Y(n_567) );
INVx1_ASAP7_75t_L g718 ( .A(n_557), .Y(n_718) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_557), .Y(n_829) );
INVx2_ASAP7_75t_L g1128 ( .A(n_557), .Y(n_1128) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B(n_562), .Y(n_559) );
OAI221xp5_ASAP7_75t_L g958 ( .A1(n_561), .A2(n_722), .B1(n_937), .B2(n_938), .C(n_959), .Y(n_958) );
OAI221xp5_ASAP7_75t_L g1169 ( .A1(n_561), .A2(n_722), .B1(n_1151), .B2(n_1152), .C(n_1170), .Y(n_1169) );
BUFx2_ASAP7_75t_L g1831 ( .A(n_561), .Y(n_1831) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_563), .B(n_705), .Y(n_704) );
BUFx2_ASAP7_75t_L g736 ( .A(n_563), .Y(n_736) );
INVx2_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g573 ( .A(n_564), .Y(n_573) );
INVx2_ASAP7_75t_SL g910 ( .A(n_564), .Y(n_910) );
AOI222xp33_ASAP7_75t_L g645 ( .A1(n_566), .A2(n_576), .B1(n_646), .B2(n_652), .C1(n_653), .C2(n_655), .Y(n_645) );
INVx1_ASAP7_75t_L g957 ( .A(n_567), .Y(n_957) );
INVx2_ASAP7_75t_L g1008 ( .A(n_567), .Y(n_1008) );
INVx1_ASAP7_75t_L g1450 ( .A(n_567), .Y(n_1450) );
HB1xp67_ASAP7_75t_L g1829 ( .A(n_567), .Y(n_1829) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_568), .A2(n_570), .B1(n_658), .B2(n_661), .Y(n_657) );
OAI21xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_571), .B(n_572), .Y(n_569) );
OAI221xp5_ASAP7_75t_L g720 ( .A1(n_571), .A2(n_676), .B1(n_677), .B2(n_721), .C(n_722), .Y(n_720) );
OAI22xp33_ASAP7_75t_L g1505 ( .A1(n_571), .A2(n_1175), .B1(n_1506), .B2(n_1507), .Y(n_1505) );
BUFx3_ASAP7_75t_L g1073 ( .A(n_573), .Y(n_1073) );
A2O1A1Ixp33_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B(n_578), .C(n_584), .Y(n_575) );
INVx1_ASAP7_75t_L g1334 ( .A(n_577), .Y(n_1334) );
NAND2x1p5_ASAP7_75t_L g1369 ( .A(n_582), .B(n_1366), .Y(n_1369) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x6_ASAP7_75t_L g745 ( .A(n_583), .B(n_585), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g1281 ( .A1(n_584), .A2(n_1229), .B(n_1282), .C(n_1283), .Y(n_1281) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g705 ( .A(n_585), .Y(n_705) );
INVx1_ASAP7_75t_L g839 ( .A(n_585), .Y(n_839) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx3_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx3_ASAP7_75t_L g708 ( .A(n_590), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_590), .A2(n_596), .B1(n_841), .B2(n_842), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g1268 ( .A1(n_590), .A2(n_596), .B1(n_1269), .B2(n_1270), .Y(n_1268) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx2_ASAP7_75t_L g598 ( .A(n_591), .Y(n_598) );
BUFx6f_ASAP7_75t_L g828 ( .A(n_592), .Y(n_828) );
INVx1_ASAP7_75t_L g1007 ( .A(n_592), .Y(n_1007) );
BUFx2_ASAP7_75t_L g1013 ( .A(n_592), .Y(n_1013) );
BUFx2_ASAP7_75t_L g1070 ( .A(n_592), .Y(n_1070) );
BUFx6f_ASAP7_75t_L g1273 ( .A(n_592), .Y(n_1273) );
BUFx6f_ASAP7_75t_L g1330 ( .A(n_592), .Y(n_1330) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx3_ASAP7_75t_L g709 ( .A(n_596), .Y(n_709) );
AND2x4_ASAP7_75t_L g603 ( .A(n_597), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
CKINVDCx6p67_ASAP7_75t_R g600 ( .A(n_601), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g843 ( .A1(n_601), .A2(n_844), .B1(n_845), .B2(n_846), .C(n_847), .Y(n_843) );
AOI22xp5_ASAP7_75t_L g1271 ( .A1(n_601), .A2(n_1272), .B1(n_1274), .B2(n_1275), .Y(n_1271) );
INVx8_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AOI221xp5_ASAP7_75t_SL g826 ( .A1(n_603), .A2(n_827), .B1(n_830), .B2(n_834), .C(n_835), .Y(n_826) );
INVx1_ASAP7_75t_L g833 ( .A(n_604), .Y(n_833) );
INVx1_ASAP7_75t_L g848 ( .A(n_605), .Y(n_848) );
OAI31xp33_ASAP7_75t_L g1120 ( .A1(n_605), .A2(n_1121), .A3(n_1122), .B(n_1130), .Y(n_1120) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NOR2xp67_ASAP7_75t_L g703 ( .A(n_606), .B(n_704), .Y(n_703) );
INVx3_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g858 ( .A(n_610), .Y(n_858) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_613), .Y(n_622) );
INVx2_ASAP7_75t_L g807 ( .A(n_613), .Y(n_807) );
INVx2_ASAP7_75t_L g993 ( .A(n_613), .Y(n_993) );
INVx2_ASAP7_75t_L g1084 ( .A(n_613), .Y(n_1084) );
INVx1_ASAP7_75t_L g1244 ( .A(n_613), .Y(n_1244) );
INVx2_ASAP7_75t_SL g1261 ( .A(n_613), .Y(n_1261) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_615), .A2(n_943), .B1(n_944), .B2(n_945), .Y(n_942) );
INVx1_ASAP7_75t_L g1077 ( .A(n_615), .Y(n_1077) );
INVx2_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
AND2x4_ASAP7_75t_L g1399 ( .A(n_616), .B(n_1400), .Y(n_1399) );
BUFx3_ASAP7_75t_L g1517 ( .A(n_616), .Y(n_1517) );
INVx1_ASAP7_75t_L g1078 ( .A(n_617), .Y(n_1078) );
INVx1_ASAP7_75t_L g1088 ( .A(n_617), .Y(n_1088) );
INVx1_ASAP7_75t_L g1115 ( .A(n_617), .Y(n_1115) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g801 ( .A(n_619), .Y(n_801) );
CKINVDCx5p33_ASAP7_75t_R g1075 ( .A(n_619), .Y(n_1075) );
INVx4_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g1021 ( .A(n_622), .Y(n_1021) );
INVx1_ASAP7_75t_L g1512 ( .A(n_622), .Y(n_1512) );
INVx2_ASAP7_75t_SL g804 ( .A(n_625), .Y(n_804) );
INVx1_ASAP7_75t_L g1003 ( .A(n_625), .Y(n_1003) );
INVx1_ASAP7_75t_L g1024 ( .A(n_625), .Y(n_1024) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_629), .Y(n_699) );
INVx1_ASAP7_75t_L g798 ( .A(n_629), .Y(n_798) );
INVx2_ASAP7_75t_L g869 ( .A(n_629), .Y(n_869) );
NAND2x1p5_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g1404 ( .A(n_631), .Y(n_1404) );
INVx2_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
OR2x6_ASAP7_75t_L g638 ( .A(n_633), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g644 ( .A(n_633), .Y(n_644) );
OR2x2_ASAP7_75t_L g897 ( .A(n_633), .B(n_639), .Y(n_897) );
AND2x4_ASAP7_75t_L g1403 ( .A(n_634), .B(n_1404), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_634), .B(n_640), .Y(n_1406) );
INVx1_ASAP7_75t_L g1423 ( .A(n_634), .Y(n_1423) );
AND2x4_ASAP7_75t_L g1521 ( .A(n_634), .B(n_1404), .Y(n_1521) );
AND2x2_ASAP7_75t_L g1794 ( .A(n_634), .B(n_640), .Y(n_1794) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g799 ( .A(n_638), .Y(n_799) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g817 ( .A(n_641), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_SL g809 ( .A(n_643), .Y(n_809) );
BUFx3_ASAP7_75t_L g1081 ( .A(n_643), .Y(n_1081) );
BUFx4f_ASAP7_75t_L g1257 ( .A(n_643), .Y(n_1257) );
AND2x4_ASAP7_75t_L g1420 ( .A(n_643), .B(n_1400), .Y(n_1420) );
INVx1_ASAP7_75t_L g1460 ( .A(n_643), .Y(n_1460) );
AND2x2_ASAP7_75t_L g668 ( .A(n_644), .B(n_669), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_646), .A2(n_653), .B1(n_768), .B2(n_774), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g864 ( .A1(n_646), .A2(n_653), .B1(n_865), .B2(n_866), .Y(n_864) );
AOI222xp33_ASAP7_75t_L g1285 ( .A1(n_646), .A2(n_655), .B1(n_658), .B2(n_1279), .C1(n_1282), .C2(n_1286), .Y(n_1285) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g1080 ( .A(n_648), .Y(n_1080) );
AND2x2_ASAP7_75t_L g653 ( .A(n_649), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OR2x6_ASAP7_75t_L g659 ( .A(n_650), .B(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g749 ( .A(n_650), .B(n_660), .Y(n_749) );
OR2x2_ASAP7_75t_L g751 ( .A(n_650), .B(n_752), .Y(n_751) );
OR2x2_ASAP7_75t_L g753 ( .A(n_650), .B(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g1400 ( .A(n_651), .Y(n_1400) );
AOI22xp5_ASAP7_75t_L g1287 ( .A1(n_653), .A2(n_661), .B1(n_1280), .B2(n_1288), .Y(n_1287) );
OR2x6_ASAP7_75t_L g702 ( .A(n_655), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g1395 ( .A(n_655), .Y(n_1395) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_658), .A2(n_661), .B1(n_765), .B2(n_777), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g861 ( .A1(n_658), .A2(n_661), .B1(n_862), .B2(n_863), .Y(n_861) );
CKINVDCx6p67_ASAP7_75t_R g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g855 ( .A(n_660), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g1156 ( .A1(n_660), .A2(n_1099), .B1(n_1157), .B2(n_1158), .Y(n_1156) );
CKINVDCx6p67_ASAP7_75t_R g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND4x1_ASAP7_75t_L g665 ( .A(n_666), .B(n_700), .C(n_706), .D(n_747), .Y(n_665) );
NOR3xp33_ASAP7_75t_SL g666 ( .A(n_667), .B(n_671), .C(n_698), .Y(n_666) );
BUFx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g867 ( .A1(n_668), .A2(n_799), .B1(n_868), .B2(n_869), .C(n_870), .Y(n_867) );
NOR3xp33_ASAP7_75t_SL g878 ( .A(n_668), .B(n_879), .C(n_895), .Y(n_878) );
NOR3xp33_ASAP7_75t_SL g930 ( .A(n_668), .B(n_931), .C(n_946), .Y(n_930) );
HB1xp67_ASAP7_75t_L g1096 ( .A(n_668), .Y(n_1096) );
AOI221xp5_ASAP7_75t_L g1263 ( .A1(n_668), .A2(n_799), .B1(n_869), .B2(n_1264), .C(n_1265), .Y(n_1263) );
HB1xp67_ASAP7_75t_L g1804 ( .A(n_669), .Y(n_1804) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g1524 ( .A(n_670), .Y(n_1524) );
OAI221xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_676), .B1(n_677), .B2(n_678), .C(n_681), .Y(n_672) );
BUFx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
BUFx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g883 ( .A(n_680), .Y(n_883) );
INVx2_ASAP7_75t_SL g1408 ( .A(n_680), .Y(n_1408) );
INVx2_ASAP7_75t_L g1797 ( .A(n_680), .Y(n_1797) );
BUFx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g754 ( .A(n_683), .Y(n_754) );
BUFx4f_ASAP7_75t_L g803 ( .A(n_683), .Y(n_803) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OAI22xp33_ASAP7_75t_L g1147 ( .A1(n_685), .A2(n_695), .B1(n_1148), .B2(n_1149), .Y(n_1147) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_686), .Y(n_697) );
INVx1_ASAP7_75t_L g934 ( .A(n_686), .Y(n_934) );
OAI221xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .B1(n_690), .B2(n_692), .C(n_693), .Y(n_687) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI22xp33_ASAP7_75t_L g932 ( .A1(n_695), .A2(n_933), .B1(n_934), .B2(n_935), .Y(n_932) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g1112 ( .A(n_696), .Y(n_1112) );
BUFx3_ASAP7_75t_L g1337 ( .A(n_696), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_702), .B(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g824 ( .A(n_702), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_702), .B(n_877), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_702), .B(n_951), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_702), .B(n_1119), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_702), .B(n_1161), .Y(n_1160) );
AND2x2_ASAP7_75t_L g741 ( .A(n_705), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g971 ( .A(n_705), .B(n_742), .Y(n_971) );
OAI31xp33_ASAP7_75t_SL g706 ( .A1(n_707), .A2(n_710), .A3(n_726), .B(n_746), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_715), .B1(n_716), .B2(n_719), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g1383 ( .A1(n_712), .A2(n_1384), .B1(n_1385), .B2(n_1386), .Y(n_1383) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g728 ( .A(n_713), .Y(n_728) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
BUFx2_ASAP7_75t_L g783 ( .A(n_714), .Y(n_783) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g847 ( .A(n_725), .Y(n_847) );
OAI221xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B1(n_730), .B2(n_734), .C(n_735), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_SL g1029 ( .A(n_738), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B1(n_743), .B2(n_744), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_741), .A2(n_744), .B1(n_779), .B2(n_780), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_741), .A2(n_744), .B1(n_920), .B2(n_921), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_741), .A2(n_744), .B1(n_1138), .B2(n_1139), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_744), .A2(n_970), .B1(n_971), .B2(n_972), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_744), .A2(n_971), .B1(n_1184), .B2(n_1185), .Y(n_1183) );
CKINVDCx11_ASAP7_75t_R g744 ( .A(n_745), .Y(n_744) );
CKINVDCx8_ASAP7_75t_R g974 ( .A(n_746), .Y(n_974) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_750), .Y(n_747) );
INVx1_ASAP7_75t_L g1803 ( .A(n_754), .Y(n_1803) );
XNOR2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_873), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B1(n_821), .B2(n_872), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NAND3xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_793), .C(n_795), .Y(n_759) );
OAI221xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B1(n_766), .B2(n_768), .C(n_769), .Y(n_763) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx2_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_774), .B1(n_775), .B2(n_777), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g1502 ( .A1(n_775), .A2(n_1499), .B1(n_1503), .B2(n_1504), .Y(n_1502) );
INVx2_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
INVx4_ASAP7_75t_L g915 ( .A(n_776), .Y(n_915) );
BUFx3_ASAP7_75t_L g1331 ( .A(n_776), .Y(n_1331) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_779), .A2(n_780), .B1(n_798), .B2(n_799), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_784), .B1(n_785), .B2(n_787), .Y(n_782) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
OAI22xp33_ASAP7_75t_L g1830 ( .A1(n_790), .A2(n_1801), .B1(n_1807), .B2(n_1831), .Y(n_1830) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NOR2xp33_ASAP7_75t_SL g795 ( .A(n_796), .B(n_818), .Y(n_795) );
NAND3xp33_ASAP7_75t_SL g796 ( .A(n_797), .B(n_800), .C(n_816), .Y(n_796) );
AOI33xp33_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_802), .A3(n_805), .B1(n_810), .B2(n_811), .B3(n_813), .Y(n_800) );
INVx1_ASAP7_75t_L g1101 ( .A(n_804), .Y(n_1101) );
BUFx6f_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g1048 ( .A(n_809), .Y(n_1048) );
NAND3xp33_ASAP7_75t_L g1242 ( .A(n_813), .B(n_1243), .C(n_1245), .Y(n_1242) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
AOI33xp33_ASAP7_75t_L g850 ( .A1(n_815), .A2(n_851), .A3(n_854), .B1(n_856), .B2(n_859), .B3(n_860), .Y(n_850) );
NAND3xp33_ASAP7_75t_L g1019 ( .A(n_815), .B(n_1020), .C(n_1022), .Y(n_1019) );
AOI33xp33_ASAP7_75t_L g1253 ( .A1(n_815), .A2(n_1254), .A3(n_1255), .B1(n_1256), .B2(n_1258), .B3(n_1262), .Y(n_1253) );
AOI33xp33_ASAP7_75t_L g1455 ( .A1(n_815), .A2(n_1254), .A3(n_1456), .B1(n_1457), .B2(n_1458), .B3(n_1461), .Y(n_1455) );
NAND3xp33_ASAP7_75t_L g1881 ( .A(n_815), .B(n_1882), .C(n_1883), .Y(n_1881) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
INVx2_ASAP7_75t_L g872 ( .A(n_821), .Y(n_872) );
XOR2x2_ASAP7_75t_L g821 ( .A(n_822), .B(n_871), .Y(n_821) );
NOR3xp33_ASAP7_75t_L g822 ( .A(n_823), .B(n_825), .C(n_849), .Y(n_822) );
AOI31xp33_ASAP7_75t_L g825 ( .A1(n_826), .A2(n_840), .A3(n_843), .B(n_848), .Y(n_825) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g1237 ( .A(n_833), .Y(n_1237) );
NAND2x1p5_ASAP7_75t_L g836 ( .A(n_837), .B(n_839), .Y(n_836) );
NAND2x1_ASAP7_75t_SL g1365 ( .A(n_837), .B(n_1366), .Y(n_1365) );
INVx2_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g1508 ( .A1(n_848), .A2(n_1392), .B1(n_1509), .B2(n_1530), .Y(n_1508) );
NAND4xp25_ASAP7_75t_L g849 ( .A(n_850), .B(n_861), .C(n_864), .D(n_867), .Y(n_849) );
NAND3xp33_ASAP7_75t_L g1000 ( .A(n_851), .B(n_1001), .C(n_1002), .Y(n_1000) );
NAND3xp33_ASAP7_75t_L g1238 ( .A(n_851), .B(n_1239), .C(n_1240), .Y(n_1238) );
NAND3xp33_ASAP7_75t_L g1878 ( .A(n_851), .B(n_1879), .C(n_1880), .Y(n_1878) );
INVx3_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
BUFx2_ASAP7_75t_L g1518 ( .A(n_855), .Y(n_1518) );
INVx2_ASAP7_75t_L g896 ( .A(n_869), .Y(n_896) );
AO22x2_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_927), .B1(n_928), .B2(n_975), .Y(n_873) );
INVx1_ASAP7_75t_L g975 ( .A(n_874), .Y(n_975) );
AND4x1_ASAP7_75t_L g875 ( .A(n_876), .B(n_878), .C(n_898), .D(n_924), .Y(n_875) );
OAI221xp5_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_882), .B1(n_883), .B2(n_884), .C(n_885), .Y(n_880) );
OAI22xp33_ASAP7_75t_L g1103 ( .A1(n_881), .A2(n_1104), .B1(n_1105), .B2(n_1107), .Y(n_1103) );
OAI21xp33_ASAP7_75t_L g907 ( .A1(n_884), .A2(n_908), .B(n_909), .Y(n_907) );
INVx2_ASAP7_75t_SL g944 ( .A(n_886), .Y(n_944) );
CKINVDCx5p33_ASAP7_75t_R g887 ( .A(n_888), .Y(n_887) );
INVx2_ASAP7_75t_SL g1099 ( .A(n_893), .Y(n_1099) );
OAI31xp33_ASAP7_75t_L g898 ( .A1(n_899), .A2(n_900), .A3(n_911), .B(n_922), .Y(n_898) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_902), .A2(n_903), .B1(n_904), .B2(n_906), .Y(n_901) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_902), .A2(n_933), .B1(n_935), .B2(n_956), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g1165 ( .A1(n_902), .A2(n_1148), .B1(n_1149), .B2(n_1166), .Y(n_1165) );
OAI22xp5_ASAP7_75t_SL g1178 ( .A1(n_902), .A2(n_1179), .B1(n_1180), .B2(n_1181), .Y(n_1178) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
AND2x4_ASAP7_75t_L g1359 ( .A(n_910), .B(n_1354), .Y(n_1359) );
OAI221xp5_ASAP7_75t_L g912 ( .A1(n_913), .A2(n_914), .B1(n_915), .B2(n_916), .C(n_917), .Y(n_912) );
INVx2_ASAP7_75t_L g1500 ( .A(n_913), .Y(n_1500) );
OAI22xp5_ASAP7_75t_L g1828 ( .A1(n_913), .A2(n_1790), .B1(n_1808), .B2(n_1829), .Y(n_1828) );
OAI221xp5_ASAP7_75t_L g964 ( .A1(n_915), .A2(n_965), .B1(n_966), .B2(n_967), .C(n_968), .Y(n_964) );
INVx2_ASAP7_75t_SL g1326 ( .A(n_915), .Y(n_1326) );
AND2x6_ASAP7_75t_L g1356 ( .A(n_918), .B(n_1354), .Y(n_1356) );
NAND2x1p5_ASAP7_75t_L g1371 ( .A(n_918), .B(n_1366), .Y(n_1371) );
OAI21xp5_ASAP7_75t_L g1266 ( .A1(n_922), .A2(n_1267), .B(n_1276), .Y(n_1266) );
BUFx8_ASAP7_75t_SL g922 ( .A(n_923), .Y(n_922) );
NOR2xp33_ASAP7_75t_L g924 ( .A(n_925), .B(n_926), .Y(n_924) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
AND4x1_ASAP7_75t_L g929 ( .A(n_930), .B(n_947), .C(n_950), .D(n_952), .Y(n_929) );
NOR2xp33_ASAP7_75t_L g947 ( .A(n_948), .B(n_949), .Y(n_947) );
OAI31xp33_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_954), .A3(n_963), .B(n_973), .Y(n_952) );
INVx1_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
INVx2_ASAP7_75t_SL g959 ( .A(n_960), .Y(n_959) );
INVx2_ASAP7_75t_SL g960 ( .A(n_961), .Y(n_960) );
OAI31xp33_ASAP7_75t_L g1162 ( .A1(n_973), .A2(n_1163), .A3(n_1164), .B(n_1172), .Y(n_1162) );
AOI31xp33_ASAP7_75t_L g1397 ( .A1(n_973), .A2(n_1398), .A3(n_1412), .B(n_1424), .Y(n_1397) );
INVx2_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
XNOR2x1_ASAP7_75t_L g976 ( .A(n_977), .B(n_1190), .Y(n_976) );
XNOR2xp5_ASAP7_75t_L g977 ( .A(n_978), .B(n_1091), .Y(n_977) );
XNOR2x1_ASAP7_75t_L g978 ( .A(n_979), .B(n_1042), .Y(n_978) );
AO211x2_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_982), .B(n_999), .C(n_1025), .Y(n_980) );
BUFx6f_ASAP7_75t_L g1211 ( .A(n_981), .Y(n_1211) );
NAND3xp33_ASAP7_75t_L g982 ( .A(n_983), .B(n_990), .C(n_995), .Y(n_982) );
INVx1_ASAP7_75t_L g1307 ( .A(n_987), .Y(n_1307) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g1298 ( .A1(n_992), .A2(n_997), .B1(n_1299), .B2(n_1300), .Y(n_1298) );
CKINVDCx6p67_ASAP7_75t_R g1053 ( .A(n_997), .Y(n_1053) );
NAND4xp25_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1004), .C(n_1011), .D(n_1019), .Y(n_999) );
NAND3xp33_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1009), .C(n_1010), .Y(n_1004) );
INVx2_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
NAND3xp33_ASAP7_75t_L g1227 ( .A(n_1010), .B(n_1228), .C(n_1230), .Y(n_1227) );
CKINVDCx8_ASAP7_75t_R g1390 ( .A(n_1010), .Y(n_1390) );
NAND3xp33_ASAP7_75t_L g1875 ( .A(n_1010), .B(n_1876), .C(n_1877), .Y(n_1875) );
NAND3xp33_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1015), .C(n_1018), .Y(n_1011) );
HB1xp67_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
INVx2_ASAP7_75t_SL g1068 ( .A(n_1017), .Y(n_1068) );
BUFx2_ASAP7_75t_L g1454 ( .A(n_1017), .Y(n_1454) );
BUFx3_ASAP7_75t_L g1323 ( .A(n_1018), .Y(n_1323) );
AOI31xp33_ASAP7_75t_L g1025 ( .A1(n_1026), .A2(n_1033), .A3(n_1037), .B(n_1041), .Y(n_1025) );
INVx2_ASAP7_75t_SL g1028 ( .A(n_1029), .Y(n_1028) );
INVx2_ASAP7_75t_L g1219 ( .A(n_1029), .Y(n_1219) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1031), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g1213 ( .A1(n_1034), .A2(n_1214), .B1(n_1215), .B2(n_1216), .Y(n_1213) );
AOI22xp33_ASAP7_75t_L g1315 ( .A1(n_1034), .A2(n_1216), .B1(n_1316), .B2(n_1317), .Y(n_1315) );
AOI22xp5_ASAP7_75t_L g1436 ( .A1(n_1034), .A2(n_1216), .B1(n_1437), .B2(n_1438), .Y(n_1436) );
AOI22xp33_ASAP7_75t_L g1859 ( .A1(n_1034), .A2(n_1216), .B1(n_1860), .B2(n_1861), .Y(n_1859) );
INVx5_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
INVx4_ASAP7_75t_L g1320 ( .A(n_1040), .Y(n_1320) );
AO21x1_ASAP7_75t_SL g1055 ( .A1(n_1041), .A2(n_1056), .B(n_1061), .Y(n_1055) );
CKINVDCx16_ASAP7_75t_R g1225 ( .A(n_1041), .Y(n_1225) );
AOI31xp33_ASAP7_75t_L g1310 ( .A1(n_1041), .A2(n_1311), .A3(n_1315), .B(n_1318), .Y(n_1310) );
AND4x1_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1055), .C(n_1064), .D(n_1074), .Y(n_1043) );
NAND4xp25_ASAP7_75t_L g1090 ( .A(n_1044), .B(n_1055), .C(n_1064), .D(n_1074), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1048), .Y(n_1046) );
NAND3xp33_ASAP7_75t_L g1231 ( .A(n_1065), .B(n_1232), .C(n_1236), .Y(n_1231) );
NAND3xp33_ASAP7_75t_L g1872 ( .A(n_1065), .B(n_1873), .C(n_1874), .Y(n_1872) );
INVx2_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
AOI33xp33_ASAP7_75t_L g1335 ( .A1(n_1075), .A2(n_1336), .A3(n_1340), .B1(n_1342), .B2(n_1343), .B3(n_1344), .Y(n_1335) );
HB1xp67_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
BUFx3_ASAP7_75t_L g1341 ( .A(n_1084), .Y(n_1341) );
BUFx6f_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1086), .Y(n_1415) );
AND2x4_ASAP7_75t_L g1421 ( .A(n_1086), .B(n_1422), .Y(n_1421) );
AOI22xp5_ASAP7_75t_L g1091 ( .A1(n_1092), .A2(n_1093), .B1(n_1143), .B2(n_1189), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
AND4x1_ASAP7_75t_L g1094 ( .A(n_1095), .B(n_1118), .C(n_1120), .D(n_1140), .Y(n_1094) );
NOR3xp33_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1097), .C(n_1117), .Y(n_1095) );
NOR3xp33_ASAP7_75t_SL g1145 ( .A(n_1096), .B(n_1146), .C(n_1159), .Y(n_1145) );
OAI22xp33_ASAP7_75t_L g1098 ( .A1(n_1099), .A2(n_1100), .B1(n_1101), .B2(n_1102), .Y(n_1098) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_1100), .A2(n_1102), .B1(n_1124), .B2(n_1126), .Y(n_1123) );
HB1xp67_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1106), .Y(n_1204) );
OAI22xp5_ASAP7_75t_L g1111 ( .A1(n_1112), .A2(n_1113), .B1(n_1114), .B2(n_1116), .Y(n_1111) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
NOR2xp33_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1142), .Y(n_1140) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1143), .Y(n_1189) );
AND4x1_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1160), .C(n_1162), .D(n_1186), .Y(n_1144) );
OAI22xp5_ASAP7_75t_L g1497 ( .A1(n_1166), .A2(n_1498), .B1(n_1499), .B2(n_1501), .Y(n_1497) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
INVx2_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1176), .Y(n_1493) );
INVx1_ASAP7_75t_L g1822 ( .A(n_1176), .Y(n_1822) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
NOR2xp33_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1188), .Y(n_1186) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
OAI22x1_ASAP7_75t_L g1192 ( .A1(n_1193), .A2(n_1194), .B1(n_1248), .B2(n_1249), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1196), .Y(n_1247) );
AOI221x1_ASAP7_75t_L g1196 ( .A1(n_1197), .A2(n_1211), .B1(n_1212), .B2(n_1225), .C(n_1226), .Y(n_1196) );
NAND3xp33_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1205), .C(n_1208), .Y(n_1197) );
INVx2_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
INVx1_ASAP7_75t_L g1855 ( .A(n_1201), .Y(n_1855) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
AOI211x1_ASAP7_75t_L g1296 ( .A1(n_1211), .A2(n_1297), .B(n_1310), .C(n_1321), .Y(n_1296) );
AOI221x1_ASAP7_75t_L g1846 ( .A1(n_1211), .A2(n_1225), .B1(n_1847), .B2(n_1858), .C(n_1871), .Y(n_1846) );
AOI211xp5_ASAP7_75t_L g1434 ( .A1(n_1225), .A2(n_1435), .B(n_1446), .C(n_1462), .Y(n_1434) );
NAND4xp25_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1231), .C(n_1238), .D(n_1242), .Y(n_1226) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
INVx2_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
AND2x4_ASAP7_75t_L g1353 ( .A(n_1235), .B(n_1354), .Y(n_1353) );
INVx2_ASAP7_75t_SL g1248 ( .A(n_1249), .Y(n_1248) );
INVx2_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
NAND4xp75_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1266), .C(n_1285), .D(n_1287), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1263), .Y(n_1252) );
INVx2_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1261), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1271), .Y(n_1267) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
XOR2xp5_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1429), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
XNOR2xp5_ASAP7_75t_L g1294 ( .A(n_1295), .B(n_1345), .Y(n_1294) );
NAND4xp25_ASAP7_75t_SL g1297 ( .A(n_1298), .B(n_1301), .C(n_1304), .D(n_1309), .Y(n_1297) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1335), .Y(n_1321) );
INVx3_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
INVx2_ASAP7_75t_SL g1329 ( .A(n_1330), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_1330), .B(n_1354), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_1330), .B(n_1354), .Y(n_1487) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1331), .Y(n_1385) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
XNOR2x1_ASAP7_75t_L g1345 ( .A(n_1346), .B(n_1347), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1348), .B(n_1391), .Y(n_1347) );
NOR3xp33_ASAP7_75t_SL g1348 ( .A(n_1349), .B(n_1362), .C(n_1372), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1350), .B(n_1357), .Y(n_1349) );
AOI22xp33_ASAP7_75t_L g1350 ( .A1(n_1351), .A2(n_1352), .B1(n_1355), .B2(n_1356), .Y(n_1350) );
BUFx2_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
BUFx2_ASAP7_75t_L g1482 ( .A(n_1353), .Y(n_1482) );
OAI211xp5_ASAP7_75t_L g1407 ( .A1(n_1355), .A2(n_1408), .B(n_1409), .C(n_1410), .Y(n_1407) );
AOI22xp33_ASAP7_75t_L g1480 ( .A1(n_1356), .A2(n_1481), .B1(n_1482), .B2(n_1483), .Y(n_1480) );
AOI22xp33_ASAP7_75t_L g1813 ( .A1(n_1356), .A2(n_1482), .B1(n_1796), .B2(n_1814), .Y(n_1813) );
AOI22xp33_ASAP7_75t_L g1357 ( .A1(n_1358), .A2(n_1359), .B1(n_1360), .B2(n_1361), .Y(n_1357) );
AOI22xp33_ASAP7_75t_L g1484 ( .A1(n_1359), .A2(n_1485), .B1(n_1486), .B2(n_1487), .Y(n_1484) );
AOI22xp33_ASAP7_75t_L g1815 ( .A1(n_1359), .A2(n_1487), .B1(n_1816), .B2(n_1817), .Y(n_1815) );
INVx2_ASAP7_75t_SL g1363 ( .A(n_1364), .Y(n_1363) );
INVx2_ASAP7_75t_L g1819 ( .A(n_1364), .Y(n_1819) );
INVx2_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
INVx3_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
BUFx4f_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
BUFx2_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
BUFx2_ASAP7_75t_L g1489 ( .A(n_1371), .Y(n_1489) );
OAI33xp33_ASAP7_75t_L g1372 ( .A1(n_1373), .A2(n_1375), .A3(n_1380), .B1(n_1383), .B2(n_1387), .B3(n_1390), .Y(n_1372) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVx3_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
AOI21xp5_ASAP7_75t_L g1398 ( .A1(n_1384), .A2(n_1399), .B(n_1401), .Y(n_1398) );
AOI22xp33_ASAP7_75t_L g1424 ( .A1(n_1386), .A2(n_1388), .B1(n_1425), .B2(n_1427), .Y(n_1424) );
AOI221xp5_ASAP7_75t_L g1412 ( .A1(n_1389), .A2(n_1413), .B1(n_1418), .B2(n_1419), .C(n_1421), .Y(n_1412) );
AOI21xp33_ASAP7_75t_L g1391 ( .A1(n_1392), .A2(n_1396), .B(n_1397), .Y(n_1391) );
AOI21xp33_ASAP7_75t_SL g1786 ( .A1(n_1392), .A2(n_1787), .B(n_1788), .Y(n_1786) );
INVx5_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
AND2x4_ASAP7_75t_L g1393 ( .A(n_1394), .B(n_1395), .Y(n_1393) );
AOI221xp5_ASAP7_75t_L g1510 ( .A1(n_1399), .A2(n_1503), .B1(n_1511), .B2(n_1516), .C(n_1519), .Y(n_1510) );
AOI21xp5_ASAP7_75t_L g1789 ( .A1(n_1399), .A2(n_1790), .B(n_1791), .Y(n_1789) );
INVx1_ASAP7_75t_SL g1402 ( .A(n_1403), .Y(n_1402) );
INVx2_ASAP7_75t_L g1792 ( .A(n_1403), .Y(n_1792) );
INVx2_ASAP7_75t_SL g1405 ( .A(n_1406), .Y(n_1405) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1415), .Y(n_1414) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
AOI221xp5_ASAP7_75t_L g1522 ( .A1(n_1419), .A2(n_1421), .B1(n_1507), .B2(n_1523), .C(n_1528), .Y(n_1522) );
AOI221xp5_ASAP7_75t_L g1800 ( .A1(n_1419), .A2(n_1421), .B1(n_1801), .B2(n_1802), .C(n_1805), .Y(n_1800) );
BUFx6f_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
INVx1_ASAP7_75t_SL g1422 ( .A(n_1423), .Y(n_1422) );
AOI22xp33_ASAP7_75t_L g1529 ( .A1(n_1425), .A2(n_1427), .B1(n_1504), .B2(n_1506), .Y(n_1529) );
AOI22xp33_ASAP7_75t_L g1806 ( .A1(n_1425), .A2(n_1427), .B1(n_1807), .B2(n_1808), .Y(n_1806) );
INVx6_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
INVx4_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
AOI22xp5_ASAP7_75t_L g1429 ( .A1(n_1430), .A2(n_1473), .B1(n_1474), .B2(n_1531), .Y(n_1429) );
INVxp67_ASAP7_75t_SL g1531 ( .A(n_1430), .Y(n_1531) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
XNOR2xp5_ASAP7_75t_L g1432 ( .A(n_1433), .B(n_1434), .Y(n_1432) );
NAND2xp5_ASAP7_75t_SL g1446 ( .A(n_1447), .B(n_1455), .Y(n_1446) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
AOI31xp33_ASAP7_75t_SL g1462 ( .A1(n_1463), .A2(n_1466), .A3(n_1469), .B(n_1472), .Y(n_1462) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
HB1xp67_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
NAND2xp5_ASAP7_75t_L g1477 ( .A(n_1478), .B(n_1508), .Y(n_1477) );
NOR3xp33_ASAP7_75t_L g1478 ( .A(n_1479), .B(n_1488), .C(n_1490), .Y(n_1478) );
NAND2xp5_ASAP7_75t_L g1479 ( .A(n_1480), .B(n_1484), .Y(n_1479) );
OAI22xp33_ASAP7_75t_L g1491 ( .A1(n_1492), .A2(n_1493), .B1(n_1494), .B2(n_1495), .Y(n_1491) );
BUFx3_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
INVx2_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
NAND3xp33_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1522), .C(n_1529), .Y(n_1509) );
BUFx2_ASAP7_75t_L g1514 ( .A(n_1515), .Y(n_1514) );
INVx2_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
OAI221xp5_ASAP7_75t_L g1533 ( .A1(n_1534), .A2(n_1779), .B1(n_1783), .B2(n_1833), .C(n_1838), .Y(n_1533) );
AOI211xp5_ASAP7_75t_L g1534 ( .A1(n_1535), .A2(n_1561), .B(n_1692), .C(n_1746), .Y(n_1534) );
OAI321xp33_ASAP7_75t_L g1692 ( .A1(n_1535), .A2(n_1624), .A3(n_1693), .B1(n_1699), .B2(n_1703), .C(n_1718), .Y(n_1692) );
INVx3_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
AOI211xp5_ASAP7_75t_L g1718 ( .A1(n_1536), .A2(n_1719), .B(n_1733), .C(n_1742), .Y(n_1718) );
NAND2xp5_ASAP7_75t_L g1739 ( .A(n_1536), .B(n_1740), .Y(n_1739) );
INVx3_ASAP7_75t_L g1754 ( .A(n_1536), .Y(n_1754) );
NAND3xp33_ASAP7_75t_L g1760 ( .A(n_1536), .B(n_1595), .C(n_1654), .Y(n_1760) );
AND2x2_ASAP7_75t_L g1772 ( .A(n_1536), .B(n_1773), .Y(n_1772) );
INVx2_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
OAI22xp5_ASAP7_75t_L g1608 ( .A1(n_1538), .A2(n_1609), .B1(n_1610), .B2(n_1611), .Y(n_1608) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1538), .Y(n_1782) );
INVx2_ASAP7_75t_L g1538 ( .A(n_1539), .Y(n_1538) );
AND2x4_ASAP7_75t_L g1539 ( .A(n_1540), .B(n_1542), .Y(n_1539) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1540), .Y(n_1546) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
NAND2xp5_ASAP7_75t_L g1553 ( .A(n_1541), .B(n_1554), .Y(n_1553) );
AND2x4_ASAP7_75t_L g1545 ( .A(n_1542), .B(n_1546), .Y(n_1545) );
AND2x2_ASAP7_75t_L g1585 ( .A(n_1542), .B(n_1546), .Y(n_1585) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1543), .Y(n_1554) );
BUFx3_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1545), .Y(n_1609) );
HB1xp67_ASAP7_75t_L g1887 ( .A(n_1546), .Y(n_1887) );
OAI22xp33_ASAP7_75t_L g1547 ( .A1(n_1548), .A2(n_1549), .B1(n_1555), .B2(n_1556), .Y(n_1547) );
BUFx3_ASAP7_75t_L g1549 ( .A(n_1550), .Y(n_1549) );
OAI22xp5_ASAP7_75t_L g1605 ( .A1(n_1550), .A2(n_1557), .B1(n_1606), .B2(n_1607), .Y(n_1605) );
BUFx6f_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
OAI22xp5_ASAP7_75t_L g1596 ( .A1(n_1551), .A2(n_1559), .B1(n_1597), .B2(n_1598), .Y(n_1596) );
OR2x2_ASAP7_75t_L g1551 ( .A(n_1552), .B(n_1553), .Y(n_1551) );
OR2x2_ASAP7_75t_L g1559 ( .A(n_1552), .B(n_1560), .Y(n_1559) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1552), .Y(n_1570) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1553), .Y(n_1569) );
HB1xp67_ASAP7_75t_L g1889 ( .A(n_1554), .Y(n_1889) );
HB1xp67_ASAP7_75t_L g1556 ( .A(n_1557), .Y(n_1556) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1560), .Y(n_1573) );
NAND4xp25_ASAP7_75t_L g1561 ( .A(n_1562), .B(n_1642), .C(n_1655), .D(n_1677), .Y(n_1561) );
NOR3xp33_ASAP7_75t_L g1562 ( .A(n_1563), .B(n_1629), .C(n_1634), .Y(n_1562) );
OAI211xp5_ASAP7_75t_L g1563 ( .A1(n_1564), .A2(n_1579), .B(n_1599), .C(n_1621), .Y(n_1563) );
OAI221xp5_ASAP7_75t_L g1719 ( .A1(n_1564), .A2(n_1697), .B1(n_1720), .B2(n_1728), .C(n_1729), .Y(n_1719) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
NAND2xp5_ASAP7_75t_L g1657 ( .A(n_1565), .B(n_1658), .Y(n_1657) );
AND2x2_ASAP7_75t_L g1565 ( .A(n_1566), .B(n_1575), .Y(n_1565) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1566), .Y(n_1601) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1566), .Y(n_1620) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1566), .Y(n_1639) );
OR2x2_ASAP7_75t_L g1652 ( .A(n_1566), .B(n_1576), .Y(n_1652) );
AND2x2_ASAP7_75t_L g1566 ( .A(n_1567), .B(n_1574), .Y(n_1566) );
AND2x4_ASAP7_75t_L g1568 ( .A(n_1569), .B(n_1570), .Y(n_1568) );
AND2x4_ASAP7_75t_L g1572 ( .A(n_1570), .B(n_1573), .Y(n_1572) );
BUFx2_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
OR2x2_ASAP7_75t_L g1619 ( .A(n_1575), .B(n_1620), .Y(n_1619) );
AND2x4_ASAP7_75t_L g1624 ( .A(n_1575), .B(n_1603), .Y(n_1624) );
AND2x2_ASAP7_75t_L g1687 ( .A(n_1575), .B(n_1604), .Y(n_1687) );
INVx1_ASAP7_75t_L g1706 ( .A(n_1575), .Y(n_1706) );
NOR2xp33_ASAP7_75t_L g1713 ( .A(n_1575), .B(n_1714), .Y(n_1713) );
AOI221xp5_ASAP7_75t_L g1762 ( .A1(n_1575), .A2(n_1763), .B1(n_1765), .B2(n_1767), .C(n_1768), .Y(n_1762) );
INVx3_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1602 ( .A(n_1576), .B(n_1603), .Y(n_1602) );
AND2x2_ASAP7_75t_L g1641 ( .A(n_1576), .B(n_1604), .Y(n_1641) );
AND2x2_ASAP7_75t_L g1668 ( .A(n_1576), .B(n_1639), .Y(n_1668) );
AOI322xp5_ASAP7_75t_L g1677 ( .A1(n_1576), .A2(n_1581), .A3(n_1678), .B1(n_1680), .B2(n_1683), .C1(n_1686), .C2(n_1688), .Y(n_1677) );
AND2x2_ASAP7_75t_L g1576 ( .A(n_1577), .B(n_1578), .Y(n_1576) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1581), .B(n_1586), .Y(n_1580) );
AND2x2_ASAP7_75t_L g1649 ( .A(n_1581), .B(n_1627), .Y(n_1649) );
OR2x2_ASAP7_75t_L g1663 ( .A(n_1581), .B(n_1588), .Y(n_1663) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1581), .B(n_1595), .Y(n_1685) );
AND2x2_ASAP7_75t_L g1704 ( .A(n_1581), .B(n_1705), .Y(n_1704) );
NOR2xp33_ASAP7_75t_L g1723 ( .A(n_1581), .B(n_1592), .Y(n_1723) );
AND2x2_ASAP7_75t_L g1726 ( .A(n_1581), .B(n_1592), .Y(n_1726) );
AND2x2_ASAP7_75t_L g1740 ( .A(n_1581), .B(n_1628), .Y(n_1740) );
BUFx3_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
BUFx2_ASAP7_75t_L g1616 ( .A(n_1582), .Y(n_1616) );
INVxp67_ASAP7_75t_L g1626 ( .A(n_1582), .Y(n_1626) );
OR2x2_ASAP7_75t_L g1712 ( .A(n_1582), .B(n_1595), .Y(n_1712) );
AND2x2_ASAP7_75t_L g1750 ( .A(n_1582), .B(n_1613), .Y(n_1750) );
AND2x2_ASAP7_75t_L g1582 ( .A(n_1583), .B(n_1584), .Y(n_1582) );
AND2x2_ASAP7_75t_L g1586 ( .A(n_1587), .B(n_1591), .Y(n_1586) );
NOR2xp33_ASAP7_75t_L g1633 ( .A(n_1587), .B(n_1614), .Y(n_1633) );
NAND2xp5_ASAP7_75t_L g1679 ( .A(n_1587), .B(n_1624), .Y(n_1679) );
AND2x2_ASAP7_75t_L g1705 ( .A(n_1587), .B(n_1613), .Y(n_1705) );
OAI21xp5_ASAP7_75t_SL g1733 ( .A1(n_1587), .A2(n_1734), .B(n_1741), .Y(n_1733) );
AND2x2_ASAP7_75t_L g1757 ( .A(n_1587), .B(n_1672), .Y(n_1757) );
INVx2_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
AND2x2_ASAP7_75t_L g1600 ( .A(n_1588), .B(n_1601), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1615 ( .A(n_1588), .B(n_1616), .Y(n_1615) );
BUFx2_ASAP7_75t_L g1645 ( .A(n_1588), .Y(n_1645) );
INVx2_ASAP7_75t_L g1654 ( .A(n_1588), .Y(n_1654) );
NAND2xp5_ASAP7_75t_L g1684 ( .A(n_1588), .B(n_1685), .Y(n_1684) );
AND2x2_ASAP7_75t_L g1695 ( .A(n_1588), .B(n_1591), .Y(n_1695) );
A2O1A1Ixp33_ASAP7_75t_L g1707 ( .A1(n_1588), .A2(n_1640), .B(n_1708), .C(n_1710), .Y(n_1707) );
NAND2xp5_ASAP7_75t_L g1714 ( .A(n_1588), .B(n_1603), .Y(n_1714) );
NAND2xp5_ASAP7_75t_L g1752 ( .A(n_1588), .B(n_1687), .Y(n_1752) );
NAND2xp5_ASAP7_75t_L g1764 ( .A(n_1588), .B(n_1709), .Y(n_1764) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1589), .B(n_1590), .Y(n_1588) );
NAND2xp5_ASAP7_75t_L g1702 ( .A(n_1591), .B(n_1615), .Y(n_1702) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_1592), .B(n_1595), .Y(n_1591) );
OR2x2_ASAP7_75t_L g1614 ( .A(n_1592), .B(n_1595), .Y(n_1614) );
AND2x2_ASAP7_75t_L g1627 ( .A(n_1592), .B(n_1628), .Y(n_1627) );
INVx2_ASAP7_75t_L g1666 ( .A(n_1592), .Y(n_1666) );
AND2x2_ASAP7_75t_L g1592 ( .A(n_1593), .B(n_1594), .Y(n_1592) );
AOI32xp33_ASAP7_75t_L g1599 ( .A1(n_1595), .A2(n_1600), .A3(n_1602), .B1(n_1612), .B2(n_1617), .Y(n_1599) );
INVx2_ASAP7_75t_SL g1628 ( .A(n_1595), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1672 ( .A(n_1595), .B(n_1666), .Y(n_1672) );
NAND2xp5_ASAP7_75t_L g1647 ( .A(n_1601), .B(n_1648), .Y(n_1647) );
AND2x2_ASAP7_75t_L g1686 ( .A(n_1601), .B(n_1687), .Y(n_1686) );
O2A1O1Ixp33_ASAP7_75t_L g1751 ( .A1(n_1601), .A2(n_1666), .B(n_1702), .C(n_1752), .Y(n_1751) );
INVx1_ASAP7_75t_L g1661 ( .A(n_1602), .Y(n_1661) );
NAND2xp5_ASAP7_75t_L g1716 ( .A(n_1602), .B(n_1717), .Y(n_1716) );
INVx2_ASAP7_75t_SL g1618 ( .A(n_1603), .Y(n_1618) );
HB1xp67_ASAP7_75t_L g1630 ( .A(n_1603), .Y(n_1630) );
INVx1_ASAP7_75t_L g1658 ( .A(n_1603), .Y(n_1658) );
AOI21xp5_ASAP7_75t_L g1720 ( .A1(n_1603), .A2(n_1721), .B(n_1724), .Y(n_1720) );
AND2x2_ASAP7_75t_L g1727 ( .A(n_1603), .B(n_1654), .Y(n_1727) );
NAND2xp5_ASAP7_75t_L g1766 ( .A(n_1603), .B(n_1676), .Y(n_1766) );
OAI32xp33_ASAP7_75t_L g1770 ( .A1(n_1603), .A2(n_1618), .A3(n_1671), .B1(n_1705), .B2(n_1709), .Y(n_1770) );
CKINVDCx5p33_ASAP7_75t_R g1603 ( .A(n_1604), .Y(n_1603) );
OR2x2_ASAP7_75t_L g1604 ( .A(n_1605), .B(n_1608), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1767 ( .A(n_1612), .B(n_1618), .Y(n_1767) );
AND2x2_ASAP7_75t_L g1612 ( .A(n_1613), .B(n_1615), .Y(n_1612) );
AND2x2_ASAP7_75t_L g1659 ( .A(n_1613), .B(n_1626), .Y(n_1659) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1614), .Y(n_1613) );
OR2x2_ASAP7_75t_L g1662 ( .A(n_1614), .B(n_1663), .Y(n_1662) );
AND2x2_ASAP7_75t_L g1671 ( .A(n_1615), .B(n_1672), .Y(n_1671) );
NOR2xp33_ASAP7_75t_L g1665 ( .A(n_1616), .B(n_1666), .Y(n_1665) );
AND2x2_ASAP7_75t_L g1691 ( .A(n_1616), .B(n_1672), .Y(n_1691) );
NOR2x1_ASAP7_75t_L g1732 ( .A(n_1616), .B(n_1628), .Y(n_1732) );
NOR2xp33_ASAP7_75t_L g1617 ( .A(n_1618), .B(n_1619), .Y(n_1617) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1618), .Y(n_1648) );
INVx2_ASAP7_75t_L g1701 ( .A(n_1618), .Y(n_1701) );
NOR2xp33_ASAP7_75t_L g1730 ( .A(n_1619), .B(n_1731), .Y(n_1730) );
OAI22xp5_ASAP7_75t_L g1761 ( .A1(n_1619), .A2(n_1647), .B1(n_1673), .B2(n_1725), .Y(n_1761) );
INVxp67_ASAP7_75t_L g1621 ( .A(n_1622), .Y(n_1621) );
A2O1A1Ixp33_ASAP7_75t_L g1741 ( .A1(n_1622), .A2(n_1678), .B(n_1697), .C(n_1711), .Y(n_1741) );
NOR2xp33_ASAP7_75t_L g1622 ( .A(n_1623), .B(n_1625), .Y(n_1622) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
AOI22xp5_ASAP7_75t_L g1734 ( .A1(n_1624), .A2(n_1735), .B1(n_1737), .B2(n_1738), .Y(n_1734) );
AND2x2_ASAP7_75t_L g1744 ( .A(n_1624), .B(n_1676), .Y(n_1744) );
INVx2_ASAP7_75t_L g1717 ( .A(n_1625), .Y(n_1717) );
NAND2xp5_ASAP7_75t_L g1625 ( .A(n_1626), .B(n_1627), .Y(n_1625) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1626), .B(n_1633), .Y(n_1632) );
AND2x2_ASAP7_75t_L g1694 ( .A(n_1626), .B(n_1695), .Y(n_1694) );
AND2x2_ASAP7_75t_L g1709 ( .A(n_1626), .B(n_1672), .Y(n_1709) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1627), .Y(n_1635) );
NOR2xp33_ASAP7_75t_L g1629 ( .A(n_1630), .B(n_1631), .Y(n_1629) );
A2O1A1Ixp33_ASAP7_75t_L g1755 ( .A1(n_1631), .A2(n_1636), .B(n_1756), .C(n_1758), .Y(n_1755) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
NOR2xp33_ASAP7_75t_L g1634 ( .A(n_1635), .B(n_1636), .Y(n_1634) );
OR2x2_ASAP7_75t_L g1673 ( .A(n_1635), .B(n_1663), .Y(n_1673) );
NAND2xp5_ASAP7_75t_L g1681 ( .A(n_1635), .B(n_1682), .Y(n_1681) );
OR2x2_ASAP7_75t_L g1636 ( .A(n_1637), .B(n_1640), .Y(n_1636) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
INVx1_ASAP7_75t_L g1773 ( .A(n_1638), .Y(n_1773) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1639), .Y(n_1676) );
AOI21xp5_ASAP7_75t_L g1742 ( .A1(n_1640), .A2(n_1743), .B(n_1745), .Y(n_1742) );
CKINVDCx5p33_ASAP7_75t_R g1640 ( .A(n_1641), .Y(n_1640) );
NAND2xp5_ASAP7_75t_L g1644 ( .A(n_1641), .B(n_1645), .Y(n_1644) );
O2A1O1Ixp33_ASAP7_75t_L g1642 ( .A1(n_1643), .A2(n_1646), .B(n_1649), .C(n_1650), .Y(n_1642) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
INVx2_ASAP7_75t_L g1690 ( .A(n_1645), .Y(n_1690) );
NAND2xp5_ASAP7_75t_SL g1722 ( .A(n_1645), .B(n_1723), .Y(n_1722) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
OR2x2_ASAP7_75t_L g1776 ( .A(n_1648), .B(n_1764), .Y(n_1776) );
AND2x2_ASAP7_75t_L g1653 ( .A(n_1649), .B(n_1654), .Y(n_1653) );
NOR2xp33_ASAP7_75t_L g1736 ( .A(n_1649), .B(n_1709), .Y(n_1736) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_1651), .B(n_1653), .Y(n_1650) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1652), .Y(n_1651) );
NAND2xp5_ASAP7_75t_L g1664 ( .A(n_1654), .B(n_1665), .Y(n_1664) );
NAND2xp5_ASAP7_75t_L g1769 ( .A(n_1654), .B(n_1687), .Y(n_1769) );
AOI211xp5_ASAP7_75t_L g1655 ( .A1(n_1656), .A2(n_1659), .B(n_1660), .C(n_1669), .Y(n_1655) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1657), .Y(n_1656) );
NAND2xp5_ASAP7_75t_L g1667 ( .A(n_1658), .B(n_1668), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1675 ( .A(n_1658), .B(n_1676), .Y(n_1675) );
INVx1_ASAP7_75t_L g1698 ( .A(n_1658), .Y(n_1698) );
OAI22xp5_ASAP7_75t_L g1660 ( .A1(n_1661), .A2(n_1662), .B1(n_1664), .B2(n_1667), .Y(n_1660) );
OAI31xp33_ASAP7_75t_L g1774 ( .A1(n_1668), .A2(n_1704), .A3(n_1775), .B(n_1777), .Y(n_1774) );
AOI21xp33_ASAP7_75t_L g1669 ( .A1(n_1670), .A2(n_1673), .B(n_1674), .Y(n_1669) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1671), .Y(n_1670) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1672), .Y(n_1682) );
NOR2xp33_ASAP7_75t_L g1748 ( .A(n_1674), .B(n_1749), .Y(n_1748) );
INVx1_ASAP7_75t_L g1674 ( .A(n_1675), .Y(n_1674) );
INVx2_ASAP7_75t_L g1697 ( .A(n_1676), .Y(n_1697) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1684), .Y(n_1683) );
INVx1_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
NAND2xp5_ASAP7_75t_L g1689 ( .A(n_1690), .B(n_1691), .Y(n_1689) );
NAND2xp5_ASAP7_75t_L g1731 ( .A(n_1690), .B(n_1732), .Y(n_1731) );
NAND2xp5_ASAP7_75t_L g1778 ( .A(n_1691), .B(n_1701), .Y(n_1778) );
AOI21xp33_ASAP7_75t_SL g1693 ( .A1(n_1694), .A2(n_1696), .B(n_1698), .Y(n_1693) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1695), .Y(n_1728) );
INVx1_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
INVxp67_ASAP7_75t_SL g1699 ( .A(n_1700), .Y(n_1699) );
NAND2xp5_ASAP7_75t_L g1700 ( .A(n_1701), .B(n_1702), .Y(n_1700) );
AOI211xp5_ASAP7_75t_L g1703 ( .A1(n_1704), .A2(n_1706), .B(n_1707), .C(n_1715), .Y(n_1703) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1704), .Y(n_1745) );
INVx1_ASAP7_75t_L g1737 ( .A(n_1706), .Y(n_1737) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1709), .Y(n_1708) );
O2A1O1Ixp33_ASAP7_75t_L g1758 ( .A1(n_1709), .A2(n_1744), .B(n_1759), .C(n_1761), .Y(n_1758) );
NAND2xp5_ASAP7_75t_L g1710 ( .A(n_1711), .B(n_1713), .Y(n_1710) );
INVx1_ASAP7_75t_L g1711 ( .A(n_1712), .Y(n_1711) );
INVxp67_ASAP7_75t_L g1715 ( .A(n_1716), .Y(n_1715) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1724 ( .A(n_1725), .Y(n_1724) );
NAND2xp5_ASAP7_75t_L g1725 ( .A(n_1726), .B(n_1727), .Y(n_1725) );
O2A1O1Ixp33_ASAP7_75t_SL g1768 ( .A1(n_1726), .A2(n_1769), .B(n_1770), .C(n_1771), .Y(n_1768) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1730), .Y(n_1729) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1736), .Y(n_1735) );
INVx1_ASAP7_75t_L g1738 ( .A(n_1739), .Y(n_1738) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1744), .Y(n_1743) );
NAND3xp33_ASAP7_75t_L g1746 ( .A(n_1747), .B(n_1762), .C(n_1774), .Y(n_1746) );
O2A1O1Ixp33_ASAP7_75t_L g1747 ( .A1(n_1748), .A2(n_1751), .B(n_1753), .C(n_1755), .Y(n_1747) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1750), .Y(n_1749) );
INVx2_ASAP7_75t_L g1753 ( .A(n_1754), .Y(n_1753) );
INVx1_ASAP7_75t_L g1756 ( .A(n_1757), .Y(n_1756) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1760), .Y(n_1759) );
INVx1_ASAP7_75t_L g1763 ( .A(n_1764), .Y(n_1763) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1766), .Y(n_1765) );
INVx1_ASAP7_75t_L g1771 ( .A(n_1772), .Y(n_1771) );
INVxp67_ASAP7_75t_L g1775 ( .A(n_1776), .Y(n_1775) );
INVxp67_ASAP7_75t_L g1777 ( .A(n_1778), .Y(n_1777) );
CKINVDCx5p33_ASAP7_75t_R g1779 ( .A(n_1780), .Y(n_1779) );
INVx1_ASAP7_75t_L g1780 ( .A(n_1781), .Y(n_1780) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1782), .Y(n_1781) );
INVx1_ASAP7_75t_L g1783 ( .A(n_1784), .Y(n_1783) );
XNOR2x1_ASAP7_75t_L g1784 ( .A(n_1785), .B(n_1832), .Y(n_1784) );
AND2x2_ASAP7_75t_L g1785 ( .A(n_1786), .B(n_1811), .Y(n_1785) );
AOI31xp33_ASAP7_75t_L g1788 ( .A1(n_1789), .A2(n_1800), .A3(n_1806), .B(n_1809), .Y(n_1788) );
INVx3_ASAP7_75t_L g1793 ( .A(n_1794), .Y(n_1793) );
OAI211xp5_ASAP7_75t_L g1795 ( .A1(n_1796), .A2(n_1797), .B(n_1798), .C(n_1799), .Y(n_1795) );
INVx2_ASAP7_75t_L g1809 ( .A(n_1810), .Y(n_1809) );
NOR3xp33_ASAP7_75t_SL g1811 ( .A(n_1812), .B(n_1818), .C(n_1820), .Y(n_1811) );
NAND2xp5_ASAP7_75t_L g1812 ( .A(n_1813), .B(n_1815), .Y(n_1812) );
CKINVDCx14_ASAP7_75t_R g1833 ( .A(n_1834), .Y(n_1833) );
BUFx2_ASAP7_75t_L g1834 ( .A(n_1835), .Y(n_1834) );
INVx1_ASAP7_75t_L g1835 ( .A(n_1836), .Y(n_1835) );
INVx1_ASAP7_75t_L g1836 ( .A(n_1837), .Y(n_1836) );
INVx1_ASAP7_75t_L g1839 ( .A(n_1840), .Y(n_1839) );
CKINVDCx5p33_ASAP7_75t_R g1840 ( .A(n_1841), .Y(n_1840) );
A2O1A1Ixp33_ASAP7_75t_L g1885 ( .A1(n_1842), .A2(n_1886), .B(n_1888), .C(n_1890), .Y(n_1885) );
INVxp33_ASAP7_75t_SL g1843 ( .A(n_1844), .Y(n_1843) );
HB1xp67_ASAP7_75t_L g1845 ( .A(n_1846), .Y(n_1845) );
NAND2xp5_ASAP7_75t_L g1847 ( .A(n_1848), .B(n_1851), .Y(n_1847) );
INVx1_ASAP7_75t_L g1866 ( .A(n_1867), .Y(n_1866) );
INVx1_ASAP7_75t_L g1867 ( .A(n_1868), .Y(n_1867) );
NAND4xp25_ASAP7_75t_L g1871 ( .A(n_1872), .B(n_1875), .C(n_1878), .D(n_1881), .Y(n_1871) );
HB1xp67_ASAP7_75t_L g1884 ( .A(n_1885), .Y(n_1884) );
INVx1_ASAP7_75t_L g1886 ( .A(n_1887), .Y(n_1886) );
INVx1_ASAP7_75t_L g1888 ( .A(n_1889), .Y(n_1888) );
endmodule