module fake_jpeg_13986_n_362 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_362);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_362;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_6),
.B(n_3),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_28),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_54),
.Y(n_96)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_50),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_51),
.Y(n_146)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_52),
.Y(n_136)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_56),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_71),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_68),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_18),
.B(n_1),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_34),
.B(n_1),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_84),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_17),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_85),
.Y(n_105)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_83),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_35),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_42),
.B(n_4),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_86),
.B(n_89),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_88),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_42),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_91),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_25),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_41),
.B(n_5),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_92),
.B(n_9),
.Y(n_126)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_93),
.B(n_63),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_50),
.A2(n_23),
.B1(n_24),
.B2(n_47),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_95),
.A2(n_98),
.B1(n_100),
.B2(n_70),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_24),
.B1(n_43),
.B2(n_38),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_51),
.A2(n_22),
.B1(n_27),
.B2(n_21),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_60),
.B1(n_57),
.B2(n_55),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_101),
.A2(n_95),
.B1(n_100),
.B2(n_146),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_22),
.B1(n_27),
.B2(n_21),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_102),
.A2(n_127),
.B1(n_118),
.B2(n_129),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_20),
.C(n_43),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_108),
.B(n_128),
.C(n_107),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_62),
.A2(n_20),
.B1(n_38),
.B2(n_44),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_111),
.A2(n_116),
.B(n_88),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_67),
.A2(n_44),
.B1(n_25),
.B2(n_9),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_52),
.B(n_5),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_67),
.B(n_7),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_89),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_131),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_133),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_81),
.B(n_9),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_56),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_83),
.B(n_11),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_140),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_84),
.B(n_11),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_148),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_149),
.Y(n_219)
);

CKINVDCx12_ASAP7_75t_R g150 ( 
.A(n_136),
.Y(n_150)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_154),
.A2(n_155),
.B(n_169),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_111),
.A2(n_116),
.B(n_142),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_156),
.A2(n_180),
.B1(n_185),
.B2(n_162),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_112),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_165),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_105),
.Y(n_165)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_166),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_97),
.B(n_72),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_168),
.B(n_172),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_104),
.B(n_88),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_96),
.B(n_73),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_99),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_174),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_99),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_121),
.A2(n_137),
.B(n_113),
.C(n_134),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_175),
.A2(n_117),
.B(n_119),
.C(n_146),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_182),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_128),
.B(n_139),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_177),
.B(n_178),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_115),
.B(n_144),
.Y(n_178)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_181),
.A2(n_129),
.B1(n_135),
.B2(n_143),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_127),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_183),
.Y(n_204)
);

INVx2_ASAP7_75t_R g184 ( 
.A(n_101),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_186),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_94),
.A2(n_106),
.B1(n_117),
.B2(n_119),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_94),
.B(n_106),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_208),
.Y(n_223)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_122),
.B1(n_155),
.B2(n_154),
.Y(n_191)
);

AND2x4_ASAP7_75t_L g240 ( 
.A(n_191),
.B(n_202),
.Y(n_240)
);

AND2x6_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_122),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_206),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

MAJx2_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_160),
.C(n_158),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_166),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_148),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_186),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_157),
.A2(n_153),
.B(n_169),
.C(n_180),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_212),
.Y(n_225)
);

AO22x1_ASAP7_75t_SL g212 ( 
.A1(n_164),
.A2(n_147),
.B1(n_151),
.B2(n_171),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_169),
.A2(n_179),
.B(n_163),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_152),
.B(n_161),
.Y(n_230)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_212),
.Y(n_221)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_221),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_232),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_201),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_233),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_227),
.Y(n_265)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_230),
.A2(n_191),
.B(n_197),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_149),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_211),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_188),
.A2(n_149),
.B(n_183),
.C(n_170),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_234),
.A2(n_240),
.B(n_199),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_183),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_235),
.B(n_236),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_167),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_241),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_239),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_192),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_202),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_192),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_242),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_199),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_206),
.Y(n_252)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_189),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_189),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_246),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_251),
.A2(n_255),
.B(n_230),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_262),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_191),
.C(n_197),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_260),
.C(n_240),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_231),
.A2(n_200),
.B1(n_191),
.B2(n_196),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_263),
.B1(n_228),
.B2(n_225),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_242),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_266),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_220),
.B(n_193),
.C(n_204),
.Y(n_260)
);

XOR2x2_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_218),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_231),
.A2(n_221),
.B1(n_227),
.B2(n_240),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_225),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_247),
.B(n_224),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_269),
.B(n_276),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_261),
.Y(n_270)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_249),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_278),
.B1(n_284),
.B2(n_285),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_266),
.A2(n_231),
.B1(n_223),
.B2(n_228),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_277),
.Y(n_289)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_275),
.Y(n_303)
);

NOR4xp25_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_223),
.C(n_233),
.D(n_240),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_263),
.A2(n_265),
.B1(n_255),
.B2(n_250),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_281),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_240),
.C(n_245),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_260),
.C(n_267),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_282),
.A2(n_253),
.B(n_251),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_226),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_283),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_210),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_193),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_248),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_267),
.Y(n_295)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_287),
.Y(n_293)
);

NAND3xp33_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_276),
.C(n_280),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_262),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_257),
.Y(n_314)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_295),
.Y(n_318)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_297),
.Y(n_305)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_302),
.C(n_279),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_282),
.A2(n_246),
.B1(n_234),
.B2(n_261),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_301),
.A2(n_257),
.B1(n_270),
.B2(n_238),
.Y(n_316)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_275),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_304),
.Y(n_313)
);

OAI21xp33_ASAP7_75t_SL g322 ( 
.A1(n_306),
.A2(n_311),
.B(n_318),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_274),
.B1(n_286),
.B2(n_287),
.Y(n_307)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_295),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_315),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_291),
.B(n_302),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_309),
.B(n_312),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_304),
.C(n_297),
.Y(n_331)
);

OA21x2_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_273),
.B(n_278),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_298),
.B(n_274),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_301),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_294),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_292),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_238),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_319),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_290),
.B(n_244),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_288),
.C(n_289),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_324),
.C(n_331),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_L g338 ( 
.A(n_322),
.B(n_328),
.C(n_293),
.Y(n_338)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_311),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_299),
.C(n_303),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_327),
.B(n_314),
.Y(n_334)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_305),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_329),
.Y(n_336)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_332),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_325),
.B(n_293),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_338),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_334),
.B(n_337),
.Y(n_343)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_323),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_321),
.A2(n_313),
.B1(n_306),
.B2(n_237),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_339),
.A2(n_340),
.B(n_322),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_320),
.A2(n_313),
.B(n_229),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_330),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_341),
.B(n_344),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_326),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_345),
.B(n_195),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_338),
.A2(n_326),
.B1(n_194),
.B2(n_219),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_347),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_339),
.B(n_194),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_350),
.B(n_352),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_341),
.B(n_190),
.C(n_219),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_190),
.Y(n_353)
);

O2A1O1Ixp33_ASAP7_75t_L g355 ( 
.A1(n_353),
.A2(n_348),
.B(n_343),
.C(n_346),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_355),
.B(n_356),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_195),
.C(n_214),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_353),
.A2(n_214),
.B(n_218),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_357),
.A2(n_351),
.B(n_215),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_359),
.B(n_354),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_360),
.B(n_358),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_361),
.B(n_215),
.Y(n_362)
);


endmodule