module fake_jpeg_3254_n_94 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_94);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_94;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_17),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_3),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_24),
.B(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_10),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_0),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_16),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_29),
.A2(n_13),
.B1(n_15),
.B2(n_18),
.Y(n_42)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_10),
.B(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_13),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_21),
.B1(n_20),
.B2(n_19),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_43),
.B1(n_26),
.B2(n_32),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

OA22x2_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_45),
.B1(n_40),
.B2(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_5),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_15),
.B1(n_18),
.B2(n_4),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_22),
.A2(n_5),
.B1(n_30),
.B2(n_27),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_48),
.B1(n_40),
.B2(n_36),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_23),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_50),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_57),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_23),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_30),
.Y(n_57)
);

AOI21x1_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_44),
.B(n_35),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_57),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_63),
.B1(n_66),
.B2(n_68),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_52),
.Y(n_64)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_44),
.B1(n_34),
.B2(n_35),
.Y(n_66)
);

INVx2_ASAP7_75t_R g69 ( 
.A(n_68),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_54),
.C(n_55),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_60),
.C(n_65),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_54),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_62),
.B(n_51),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_48),
.B1(n_34),
.B2(n_51),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_67),
.B1(n_74),
.B2(n_69),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_74),
.A2(n_67),
.B(n_63),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_78),
.C(n_79),
.Y(n_84)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

AOI322xp5_ASAP7_75t_SL g82 ( 
.A1(n_76),
.A2(n_72),
.A3(n_71),
.B1(n_69),
.B2(n_70),
.C1(n_75),
.C2(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_82),
.B(n_69),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_79),
.C(n_76),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_86),
.B(n_87),
.Y(n_90)
);

NOR2xp67_ASAP7_75t_SL g88 ( 
.A(n_83),
.B(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_85),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_75),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_71),
.B(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_90),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_71),
.Y(n_94)
);


endmodule