module fake_jpeg_29800_n_177 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_26),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_30),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_25),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_0),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_72),
.Y(n_92)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_60),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_73),
.B(n_75),
.Y(n_80)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_44),
.Y(n_75)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_53),
.C(n_49),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_61),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_69),
.Y(n_90)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g112 ( 
.A(n_93),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_92),
.B(n_62),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_80),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_97),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_68),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_43),
.B1(n_45),
.B2(n_48),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_43),
.B1(n_54),
.B2(n_23),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_67),
.C(n_46),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_64),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_104),
.Y(n_133)
);

OA22x2_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_90),
.B1(n_85),
.B2(n_58),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

OR2x4_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_65),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_65),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_62),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_106),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_79),
.B(n_51),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_55),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_80),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_109),
.B(n_56),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_6),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_59),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_115),
.B(n_130),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_121),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_47),
.B(n_63),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_9),
.B(n_10),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_101),
.A2(n_54),
.B1(n_48),
.B2(n_45),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_1),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_128),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_106),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_112),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_131),
.Y(n_140)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_102),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_5),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_132),
.Y(n_148)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_136),
.Y(n_149)
);

NOR2x1_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_7),
.Y(n_141)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_27),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_143),
.A2(n_152),
.B(n_137),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

NAND2xp33_ASAP7_75t_SL g147 ( 
.A(n_134),
.B(n_7),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_SL g159 ( 
.A1(n_147),
.A2(n_15),
.B(n_16),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_150),
.A2(n_154),
.B(n_131),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_120),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_151),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_31),
.B(n_12),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_9),
.B1(n_13),
.B2(n_14),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_139),
.A2(n_135),
.B1(n_128),
.B2(n_129),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_156),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_159),
.Y(n_166)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_160),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_146),
.A2(n_19),
.B(n_21),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_142),
.B1(n_138),
.B2(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_SL g168 ( 
.A(n_166),
.B(n_140),
.C(n_157),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_167),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_170),
.B(n_169),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_SL g172 ( 
.A(n_171),
.B(n_165),
.C(n_163),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_172),
.B(n_163),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_162),
.B1(n_164),
.B2(n_147),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_149),
.C(n_148),
.Y(n_175)
);

AOI31xp67_ASAP7_75t_SL g176 ( 
.A1(n_175),
.A2(n_143),
.A3(n_153),
.B(n_141),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_153),
.Y(n_177)
);


endmodule