module fake_jpeg_27470_n_198 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_198);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

BUFx8_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_14),
.B(n_1),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_29),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_33),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_19),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_17),
.B1(n_23),
.B2(n_22),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_42),
.B1(n_31),
.B2(n_25),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_17),
.B1(n_24),
.B2(n_18),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_26),
.A2(n_13),
.B1(n_15),
.B2(n_22),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_15),
.B1(n_18),
.B2(n_25),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_34),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_47),
.B(n_31),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_20),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_57),
.Y(n_83)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_51),
.B(n_54),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_52),
.Y(n_84)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_12),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_34),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_32),
.Y(n_81)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_12),
.Y(n_58)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_62),
.B1(n_65),
.B2(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_64),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_30),
.B1(n_32),
.B2(n_13),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_20),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_21),
.B1(n_19),
.B2(n_16),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_30),
.B1(n_13),
.B2(n_20),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_41),
.B1(n_42),
.B2(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

AND2x6_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_86),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_82),
.B1(n_87),
.B2(n_65),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_46),
.B1(n_62),
.B2(n_48),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_79),
.A2(n_6),
.B1(n_7),
.B2(n_78),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_39),
.C(n_34),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_3),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_1),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_21),
.B1(n_19),
.B2(n_16),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_2),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_5),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_106),
.B1(n_78),
.B2(n_77),
.Y(n_134)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_108),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_59),
.B(n_68),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_100),
.A2(n_102),
.B(n_103),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_11),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_101),
.B(n_110),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_53),
.B(n_49),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_57),
.B(n_61),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_10),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_104),
.A2(n_105),
.B(n_107),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_64),
.B(n_70),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_16),
.B1(n_3),
.B2(n_4),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_71),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_72),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_89),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_111),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_112),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_113),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_86),
.B(n_8),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_116),
.A2(n_92),
.B1(n_100),
.B2(n_90),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_99),
.C(n_109),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_127),
.C(n_136),
.Y(n_150)
);

FAx1_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_72),
.CI(n_75),
.CON(n_120),
.SN(n_120)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_132),
.Y(n_147)
);

XNOR2x1_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_81),
.Y(n_122)
);

XNOR2x2_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_107),
.Y(n_144)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_92),
.B(n_88),
.Y(n_124)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_125),
.B(n_127),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_128),
.A2(n_134),
.B1(n_116),
.B2(n_90),
.Y(n_145)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_141),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_131),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_143),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_150),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_134),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_107),
.B1(n_91),
.B2(n_6),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_91),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_124),
.B(n_133),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_152),
.A2(n_145),
.B(n_146),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_142),
.A2(n_122),
.B1(n_125),
.B2(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_155),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_126),
.B1(n_120),
.B2(n_136),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_119),
.C(n_130),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_161),
.B(n_149),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_154),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_165),
.Y(n_177)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_170),
.B1(n_147),
.B2(n_151),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_161),
.C(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_169),
.Y(n_173)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_172),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_137),
.B(n_144),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_175),
.B(n_176),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_160),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_179),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_160),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_159),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_180),
.B(n_156),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_177),
.Y(n_183)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_185),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_166),
.B1(n_139),
.B2(n_143),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_140),
.B1(n_138),
.B2(n_141),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_174),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_188),
.B(n_190),
.Y(n_192)
);

NOR2xp67_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_120),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_183),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_189),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_193),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_192),
.A2(n_181),
.B(n_179),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_194),
.C(n_118),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_135),
.Y(n_198)
);


endmodule