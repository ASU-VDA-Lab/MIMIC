module fake_jpeg_32037_n_331 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_44),
.B(n_47),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_48),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_14),
.B(n_6),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_53),
.Y(n_81)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_23),
.Y(n_55)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_21),
.A2(n_27),
.B(n_31),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_35),
.B(n_33),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_61),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_95),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_29),
.B1(n_17),
.B2(n_38),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_77),
.A2(n_24),
.B1(n_15),
.B2(n_58),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_82),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_37),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g152 ( 
.A(n_84),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_35),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_87),
.B(n_0),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_57),
.B1(n_29),
.B2(n_17),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_94),
.A2(n_4),
.B1(n_12),
.B2(n_88),
.Y(n_157)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_37),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_104),
.Y(n_126)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_55),
.A2(n_29),
.B1(n_17),
.B2(n_32),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_105),
.B1(n_119),
.B2(n_48),
.Y(n_120)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_54),
.A2(n_32),
.B1(n_16),
.B2(n_19),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_63),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_109),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_53),
.B(n_25),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_53),
.B(n_25),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_116),
.Y(n_145)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_48),
.A2(n_19),
.B(n_33),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_0),
.C(n_2),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_63),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_43),
.B(n_14),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_117),
.B(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_67),
.A2(n_19),
.B1(n_36),
.B2(n_24),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_120),
.A2(n_123),
.B1(n_130),
.B2(n_134),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_122),
.B(n_127),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_68),
.B1(n_62),
.B2(n_69),
.Y(n_123)
);

NAND2x1p5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_63),
.Y(n_125)
);

NAND2x1_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_78),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_82),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_91),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_128),
.B(n_144),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_87),
.A2(n_114),
.B1(n_115),
.B2(n_76),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_81),
.B(n_36),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_136),
.B(n_154),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_137),
.A2(n_140),
.B(n_83),
.Y(n_181)
);

AO22x1_ASAP7_75t_SL g138 ( 
.A1(n_79),
.A2(n_46),
.B1(n_19),
.B2(n_3),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_113),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_139),
.B(n_112),
.Y(n_177)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_141),
.Y(n_171)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_73),
.B(n_8),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_71),
.B(n_2),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_153),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_71),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_147),
.A2(n_160),
.B1(n_161),
.B2(n_78),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_7),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_149),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_9),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_90),
.A2(n_11),
.B1(n_12),
.B2(n_5),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_150),
.A2(n_157),
.B1(n_89),
.B2(n_106),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_93),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_158),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_90),
.B(n_2),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_92),
.B(n_12),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_92),
.B(n_2),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_156),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_79),
.B(n_4),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_101),
.B(n_97),
.CI(n_74),
.CON(n_158),
.SN(n_158)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_97),
.A2(n_88),
.B1(n_110),
.B2(n_102),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_110),
.A2(n_72),
.B1(n_83),
.B2(n_118),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_113),
.B(n_72),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_158),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_93),
.B(n_86),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_163),
.A2(n_138),
.B(n_135),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_86),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_177),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_166),
.A2(n_172),
.B1(n_187),
.B2(n_193),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_167),
.A2(n_153),
.B(n_155),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_169),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_175),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_131),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_179),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_163),
.Y(n_222)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_133),
.Y(n_182)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_145),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_128),
.Y(n_212)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_89),
.B1(n_106),
.B2(n_96),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_127),
.B(n_78),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_191),
.B(n_126),
.Y(n_205)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_143),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_195),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_152),
.A2(n_75),
.B1(n_96),
.B2(n_157),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_137),
.A2(n_75),
.B(n_134),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_194),
.A2(n_167),
.B(n_187),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_139),
.B(n_146),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_135),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_141),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_197),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_152),
.A2(n_125),
.B1(n_156),
.B2(n_140),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_198),
.A2(n_154),
.B1(n_136),
.B2(n_121),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_200),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_211),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_193),
.A2(n_125),
.B1(n_130),
.B2(n_138),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_206),
.A2(n_207),
.B(n_224),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_165),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_219),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_209),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_179),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_214),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_222),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_190),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_183),
.A2(n_129),
.B1(n_132),
.B2(n_142),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_215),
.A2(n_218),
.B1(n_221),
.B2(n_226),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_166),
.A2(n_124),
.B1(n_151),
.B2(n_159),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_124),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_174),
.Y(n_220)
);

A2O1A1O1Ixp25_ASAP7_75t_L g255 ( 
.A1(n_220),
.A2(n_223),
.B(n_225),
.C(n_176),
.D(n_171),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_166),
.A2(n_194),
.B1(n_172),
.B2(n_198),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_174),
.B(n_195),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_190),
.A2(n_197),
.B(n_165),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_177),
.B(n_182),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_183),
.A2(n_167),
.B1(n_178),
.B2(n_181),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_230),
.A2(n_171),
.B(n_173),
.Y(n_248)
);

AOI22x1_ASAP7_75t_L g231 ( 
.A1(n_208),
.A2(n_164),
.B1(n_168),
.B2(n_192),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_231),
.Y(n_266)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_178),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_244),
.C(n_200),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_208),
.A2(n_186),
.B1(n_164),
.B2(n_175),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_255),
.Y(n_259)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_237),
.Y(n_268)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_241),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_196),
.C(n_185),
.Y(n_244)
);

AOI22x1_ASAP7_75t_SL g247 ( 
.A1(n_207),
.A2(n_173),
.B1(n_185),
.B2(n_188),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_247),
.A2(n_202),
.B(n_225),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_202),
.B(n_224),
.Y(n_257)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_250),
.Y(n_264)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_201),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_232),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_188),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_215),
.A2(n_176),
.B1(n_180),
.B2(n_230),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_256),
.A2(n_203),
.B1(n_218),
.B2(n_221),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_257),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_238),
.B(n_245),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_258),
.B(n_269),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_262),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_220),
.C(n_223),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_244),
.C(n_242),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_276),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_210),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_233),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_270),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_247),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_242),
.Y(n_280)
);

OAI322xp33_ASAP7_75t_L g272 ( 
.A1(n_255),
.A2(n_210),
.A3(n_219),
.B1(n_213),
.B2(n_211),
.C1(n_203),
.C2(n_206),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_261),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_246),
.A2(n_228),
.B(n_217),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_239),
.A2(n_209),
.B1(n_228),
.B2(n_256),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_277),
.A2(n_239),
.B1(n_248),
.B2(n_246),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_279),
.A2(n_282),
.B1(n_273),
.B2(n_274),
.Y(n_303)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_287),
.C(n_289),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_266),
.A2(n_243),
.B1(n_253),
.B2(n_231),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_285),
.B(n_288),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_253),
.C(n_243),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_231),
.C(n_252),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_259),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_274),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_286),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_297),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_292),
.B(n_267),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_271),
.C(n_270),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_302),
.C(n_290),
.Y(n_306)
);

NOR4xp25_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_275),
.C(n_264),
.D(n_272),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_299),
.B(n_303),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_284),
.A2(n_277),
.B1(n_265),
.B2(n_266),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_278),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_278),
.A2(n_259),
.B1(n_266),
.B2(n_264),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_301),
.A2(n_304),
.B1(n_260),
.B2(n_268),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_269),
.C(n_276),
.Y(n_302)
);

XOR2x1_ASAP7_75t_SL g304 ( 
.A(n_284),
.B(n_273),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_285),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_310),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_283),
.C(n_281),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_313),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_315),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_298),
.A2(n_289),
.B(n_268),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_311),
.A2(n_306),
.B(n_312),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_282),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_260),
.Y(n_314)
);

NAND2xp33_ASAP7_75t_SL g317 ( 
.A(n_314),
.B(n_308),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_314),
.A2(n_294),
.B(n_302),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_319),
.B(n_321),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_317),
.B(n_318),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_295),
.C(n_305),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_310),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_323),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_326),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_319),
.C(n_316),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_325),
.C(n_323),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_329),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_328),
.Y(n_331)
);


endmodule