module fake_jpeg_28950_n_401 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_401);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_401;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_48),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_49),
.B(n_21),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_53),
.Y(n_81)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_44),
.B1(n_38),
.B2(n_28),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_63),
.B1(n_38),
.B2(n_34),
.Y(n_79)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g104 ( 
.A(n_72),
.B(n_77),
.Y(n_104)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

BUFx4f_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_35),
.Y(n_108)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_21),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_43),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_79),
.A2(n_96),
.B1(n_100),
.B2(n_105),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_38),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_94),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_36),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_60),
.A2(n_30),
.B1(n_28),
.B2(n_42),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_21),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_54),
.A2(n_30),
.B1(n_22),
.B2(n_41),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_57),
.A2(n_30),
.B1(n_41),
.B2(n_23),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_110),
.B(n_116),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_51),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_34),
.B1(n_31),
.B2(n_45),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_59),
.B(n_65),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_115),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_27),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_47),
.B(n_40),
.C(n_22),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_21),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

NAND2xp33_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_73),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_140),
.Y(n_154)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_87),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_130),
.Y(n_160)
);

OA22x2_ASAP7_75t_SL g129 ( 
.A1(n_79),
.A2(n_76),
.B1(n_69),
.B2(n_53),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_129),
.A2(n_144),
.B(n_104),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_87),
.Y(n_130)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_145),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_81),
.A2(n_52),
.B1(n_39),
.B2(n_45),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_137),
.Y(n_156)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_139),
.Y(n_174)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_89),
.A2(n_39),
.B(n_34),
.C(n_23),
.Y(n_144)
);

BUFx4f_ASAP7_75t_SL g145 ( 
.A(n_118),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_108),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_81),
.A2(n_58),
.B1(n_72),
.B2(n_27),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_148),
.A2(n_69),
.B1(n_95),
.B2(n_103),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_111),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_96),
.Y(n_153)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_151),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_90),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_153),
.A2(n_155),
.B(n_140),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_113),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_161),
.A2(n_154),
.B(n_175),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_117),
.C(n_101),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_175),
.C(n_127),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_141),
.B(n_25),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_176),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_171),
.A2(n_131),
.B1(n_95),
.B2(n_129),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_132),
.A2(n_100),
.B1(n_108),
.B2(n_82),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_173),
.A2(n_179),
.B1(n_90),
.B2(n_151),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_121),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_132),
.A2(n_82),
.B1(n_56),
.B2(n_62),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_185),
.C(n_197),
.Y(n_216)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_124),
.C(n_131),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_160),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_186),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_187),
.A2(n_192),
.B1(n_201),
.B2(n_179),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_120),
.B(n_129),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_188),
.A2(n_161),
.B(n_153),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_168),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_189),
.Y(n_218)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_154),
.A2(n_144),
.B1(n_126),
.B2(n_135),
.Y(n_192)
);

NOR3xp33_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_25),
.C(n_149),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_194),
.Y(n_215)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_165),
.A2(n_103),
.B1(n_123),
.B2(n_122),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_106),
.C(n_104),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_158),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_198),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_199),
.A2(n_157),
.B1(n_177),
.B2(n_165),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_200),
.A2(n_171),
.B1(n_174),
.B2(n_151),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_66),
.B1(n_75),
.B2(n_55),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_202),
.A2(n_188),
.B(n_192),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_162),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_205),
.A2(n_213),
.B1(n_159),
.B2(n_157),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_208),
.A2(n_201),
.B1(n_190),
.B2(n_174),
.Y(n_238)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_174),
.B1(n_159),
.B2(n_142),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_220),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_185),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_232),
.C(n_236),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_225),
.A2(n_229),
.B(n_99),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_186),
.Y(n_226)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_203),
.B(n_181),
.CI(n_185),
.CON(n_228),
.SN(n_228)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_228),
.B(n_211),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_184),
.B(n_187),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_206),
.B(n_182),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_231),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_197),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_220),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_233),
.Y(n_252)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_189),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_235),
.B(n_243),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_177),
.C(n_195),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_191),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_214),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_238),
.A2(n_134),
.B1(n_125),
.B2(n_150),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_240),
.B1(n_222),
.B2(n_210),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_219),
.A2(n_218),
.B1(n_205),
.B2(n_215),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_145),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_245),
.C(n_249),
.Y(n_269)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_242),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_158),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_204),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_244),
.B(n_248),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_212),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_246),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_209),
.B(n_14),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_222),
.C(n_208),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_253),
.A2(n_255),
.B1(n_265),
.B2(n_272),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_217),
.B1(n_205),
.B2(n_213),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_237),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_256),
.B(n_261),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_214),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_257),
.B(n_267),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_237),
.Y(n_261)
);

OA22x2_ASAP7_75t_L g262 ( 
.A1(n_223),
.A2(n_230),
.B1(n_234),
.B2(n_229),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_262),
.B(n_266),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_264),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_213),
.B1(n_211),
.B2(n_210),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_233),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_270),
.A2(n_274),
.B1(n_275),
.B2(n_238),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_SL g271 ( 
.A1(n_245),
.A2(n_207),
.B(n_204),
.C(n_145),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_271),
.A2(n_246),
.B(n_109),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_223),
.A2(n_207),
.B1(n_178),
.B2(n_152),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_230),
.B(n_172),
.Y(n_273)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_273),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_239),
.A2(n_178),
.B1(n_152),
.B2(n_139),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_227),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_224),
.B(n_90),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_276),
.B(n_277),
.Y(n_292)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_278),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_236),
.C(n_228),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_291),
.C(n_296),
.Y(n_311)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_282),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_228),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_288),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_259),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_284),
.B(n_286),
.Y(n_309)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_260),
.A2(n_225),
.B1(n_242),
.B2(n_227),
.Y(n_287)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_287),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_241),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_250),
.Y(n_289)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_289),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_290),
.A2(n_264),
.B(n_272),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_172),
.C(n_163),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_269),
.B(n_21),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_295),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_269),
.B(n_21),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_277),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_262),
.B(n_138),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_301),
.C(n_302),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_266),
.B(n_133),
.C(n_83),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_262),
.B(n_83),
.C(n_99),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_303),
.B(n_307),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_297),
.A2(n_253),
.B1(n_252),
.B2(n_255),
.Y(n_305)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_323),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_294),
.Y(n_307)
);

MAJx2_ASAP7_75t_L g308 ( 
.A(n_279),
.B(n_264),
.C(n_263),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_308),
.B(n_314),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_302),
.A2(n_254),
.B(n_268),
.Y(n_310)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_310),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_300),
.A2(n_280),
.B1(n_265),
.B2(n_299),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_319),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_273),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_296),
.A2(n_271),
.B1(n_274),
.B2(n_298),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_283),
.B(n_251),
.C(n_271),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_281),
.C(n_86),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_292),
.A2(n_271),
.B1(n_278),
.B2(n_109),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_321),
.A2(n_322),
.B1(n_114),
.B2(n_70),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_292),
.A2(n_86),
.B1(n_71),
.B2(n_61),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_301),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_291),
.B(n_118),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_324),
.B(n_295),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_325),
.A2(n_337),
.B1(n_318),
.B2(n_12),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_331),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_315),
.A2(n_281),
.B1(n_293),
.B2(n_107),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_334),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_316),
.A2(n_321),
.B1(n_313),
.B2(n_320),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_333),
.B(n_305),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_114),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_322),
.A2(n_107),
.B1(n_48),
.B2(n_77),
.Y(n_336)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_336),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_319),
.A2(n_11),
.B1(n_20),
.B2(n_19),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_9),
.C(n_20),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_338),
.B(n_340),
.C(n_304),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_317),
.B(n_9),
.C(n_18),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_308),
.B(n_8),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_342),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_317),
.B(n_8),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_339),
.A2(n_313),
.B(n_324),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_343),
.A2(n_344),
.B(n_6),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_326),
.A2(n_312),
.B(n_314),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_349),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_330),
.B(n_304),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_351),
.B(n_7),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_337),
.B(n_309),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_352),
.B(n_353),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_328),
.A2(n_341),
.B1(n_335),
.B2(n_330),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_348),
.Y(n_369)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_329),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_355),
.B(n_356),
.Y(n_363)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_338),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_340),
.A2(n_8),
.B1(n_18),
.B2(n_17),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_12),
.B1(n_14),
.B2(n_18),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_358),
.B(n_360),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_334),
.C(n_332),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_353),
.B(n_342),
.Y(n_361)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_361),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_362),
.B(n_364),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_6),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_345),
.B(n_6),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_365),
.B(n_369),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_366),
.B(n_5),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_11),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_367),
.A2(n_347),
.B(n_14),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_359),
.A2(n_345),
.B(n_351),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_372),
.A2(n_0),
.B(n_1),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_SL g373 ( 
.A(n_369),
.B(n_347),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_373),
.Y(n_381)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_374),
.Y(n_388)
);

INVx11_ASAP7_75t_L g376 ( 
.A(n_368),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_377),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_363),
.B(n_29),
.C(n_5),
.Y(n_377)
);

BUFx24_ASAP7_75t_SL g379 ( 
.A(n_363),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_380),
.Y(n_385)
);

A2O1A1O1Ixp25_ASAP7_75t_L g382 ( 
.A1(n_370),
.A2(n_367),
.B(n_16),
.C(n_17),
.D(n_29),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_382),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_378),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_377),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_371),
.A2(n_0),
.B(n_1),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_386),
.B(n_383),
.C(n_388),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_387),
.A2(n_1),
.B(n_2),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_389),
.B(n_391),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_381),
.B(n_376),
.C(n_375),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_392),
.B(n_393),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_390),
.A2(n_385),
.B(n_2),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_396),
.A2(n_2),
.B(n_3),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_397),
.Y(n_399)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_394),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_399),
.B(n_398),
.C(n_395),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_400),
.B(n_3),
.Y(n_401)
);


endmodule