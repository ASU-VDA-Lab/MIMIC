module fake_jpeg_29436_n_207 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_207);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_207;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

NAND2x1_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_0),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_33),
.B1(n_21),
.B2(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_15),
.B(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_2),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_15),
.B(n_3),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_58),
.Y(n_64)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_3),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_4),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_34),
.C(n_27),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_26),
.B(n_4),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_59),
.Y(n_79)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_26),
.B(n_6),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_60),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_61),
.B(n_12),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

FAx1_ASAP7_75t_SL g115 ( 
.A(n_71),
.B(n_6),
.CI(n_8),
.CON(n_115),
.SN(n_115)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_34),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_73),
.B(n_82),
.Y(n_106)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_23),
.B1(n_29),
.B2(n_18),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_80),
.B1(n_36),
.B2(n_41),
.Y(n_105)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_50),
.A2(n_23),
.B1(n_40),
.B2(n_18),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_17),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_81),
.B(n_90),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_39),
.B(n_17),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_27),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_22),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_28),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_38),
.B(n_28),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_44),
.B(n_46),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_99),
.Y(n_127)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_46),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_103),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_37),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_89),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_109),
.B1(n_110),
.B2(n_70),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_33),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_107),
.B(n_106),
.Y(n_138)
);

INVx2_ASAP7_75t_R g108 ( 
.A(n_60),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_122),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_92),
.A2(n_29),
.B1(n_18),
.B2(n_13),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_75),
.A2(n_29),
.B1(n_13),
.B2(n_23),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

AND2x6_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_71),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_114),
.B(n_108),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_62),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_63),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_70),
.B1(n_89),
.B2(n_83),
.Y(n_129)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_123),
.B(n_138),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_129),
.B1(n_133),
.B2(n_116),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_SL g126 ( 
.A(n_108),
.B(n_64),
.C(n_88),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_126),
.B(n_137),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_142),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_77),
.C(n_78),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_107),
.C(n_109),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_65),
.B1(n_67),
.B2(n_63),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_136),
.B1(n_102),
.B2(n_112),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_104),
.A2(n_65),
.B1(n_74),
.B2(n_83),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_84),
.C(n_66),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_10),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_66),
.B(n_11),
.Y(n_145)
);

NAND2x1_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_115),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_103),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_153),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_152),
.C(n_130),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_150),
.A2(n_125),
.B1(n_144),
.B2(n_133),
.Y(n_169)
);

AO21x2_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_99),
.B(n_114),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_116),
.B1(n_119),
.B2(n_97),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_101),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_95),
.B(n_141),
.Y(n_173)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_135),
.B1(n_102),
.B2(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_137),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_134),
.C(n_97),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_163),
.B(n_164),
.Y(n_180)
);

AOI322xp5_ASAP7_75t_SL g164 ( 
.A1(n_162),
.A2(n_126),
.A3(n_123),
.B1(n_142),
.B2(n_144),
.C1(n_115),
.C2(n_128),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_174),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_161),
.A2(n_129),
.B1(n_135),
.B2(n_134),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_173),
.B1(n_169),
.B2(n_171),
.Y(n_183)
);

A2O1A1O1Ixp25_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_147),
.B(n_156),
.C(n_151),
.D(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_150),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_165),
.A2(n_153),
.B1(n_154),
.B2(n_160),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_181),
.A2(n_184),
.B(n_179),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_182),
.A2(n_183),
.B1(n_172),
.B2(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_168),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_188),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_163),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_149),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_180),
.B(n_152),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_189),
.A2(n_177),
.B(n_176),
.Y(n_195)
);

OAI321xp33_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_151),
.A3(n_156),
.B1(n_159),
.B2(n_155),
.C(n_175),
.Y(n_190)
);

AOI31xp67_ASAP7_75t_L g193 ( 
.A1(n_190),
.A2(n_178),
.A3(n_151),
.B(n_155),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_191),
.B(n_182),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_195),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_194),
.A2(n_185),
.B1(n_187),
.B2(n_191),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_194),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_197),
.B(n_198),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_192),
.A2(n_151),
.B(n_189),
.Y(n_198)
);

AOI322xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_170),
.A3(n_168),
.B1(n_148),
.B2(n_146),
.C1(n_140),
.C2(n_96),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

AOI322xp5_ASAP7_75t_L g203 ( 
.A1(n_199),
.A2(n_146),
.A3(n_112),
.B1(n_140),
.B2(n_124),
.C1(n_98),
.C2(n_12),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_SL g205 ( 
.A1(n_203),
.A2(n_140),
.B(n_12),
.C(n_197),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_202),
.C(n_124),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_204),
.Y(n_207)
);


endmodule