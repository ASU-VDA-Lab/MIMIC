module fake_jpeg_17602_n_146 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_26),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_18),
.B(n_21),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_65),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_0),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_1),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_1),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_51),
.Y(n_74)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_60),
.B1(n_44),
.B2(n_59),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_78),
.B1(n_84),
.B2(n_54),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_75),
.Y(n_91)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_44),
.B1(n_42),
.B2(n_46),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_81),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_2),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_55),
.B1(n_53),
.B2(n_50),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_87),
.B(n_99),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

BUFx4f_ASAP7_75t_SL g92 ( 
.A(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_92),
.Y(n_112)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_71),
.B(n_45),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_2),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_6),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_69),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_57),
.B1(n_56),
.B2(n_43),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_101),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_3),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_56),
.B1(n_52),
.B2(n_5),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_102),
.A2(n_3),
.B(n_4),
.Y(n_111)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_110),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_7),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_96),
.C(n_95),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_92),
.C(n_112),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_118),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_90),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_121),
.Y(n_127)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_116),
.A2(n_109),
.B(n_106),
.Y(n_123)
);

FAx1_ASAP7_75t_SL g128 ( 
.A(n_123),
.B(n_107),
.CI(n_52),
.CON(n_128),
.SN(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_89),
.C(n_86),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_109),
.B1(n_115),
.B2(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_125),
.B(n_126),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_100),
.B1(n_88),
.B2(n_105),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_129),
.C(n_126),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_7),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_133),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_128),
.C(n_10),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_8),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_29),
.Y(n_136)
);

FAx1_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_134),
.CI(n_13),
.CON(n_137),
.SN(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_31),
.C(n_15),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_32),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_130),
.C(n_16),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_27),
.Y(n_141)
);

AOI321xp33_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_33),
.A3(n_20),
.B1(n_22),
.B2(n_23),
.C(n_24),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_143),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_36),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_145),
.A2(n_38),
.B(n_25),
.Y(n_146)
);


endmodule