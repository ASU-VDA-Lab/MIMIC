module fake_aes_345_n_702 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_702);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_702;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_70), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_54), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_71), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_30), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_44), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_50), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_52), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_63), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_61), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_76), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_41), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_24), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_75), .Y(n_91) );
INVxp33_ASAP7_75t_SL g92 ( .A(n_42), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_60), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_48), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_43), .Y(n_95) );
CKINVDCx14_ASAP7_75t_R g96 ( .A(n_57), .Y(n_96) );
INVxp33_ASAP7_75t_L g97 ( .A(n_21), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_68), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_0), .Y(n_99) );
CKINVDCx14_ASAP7_75t_R g100 ( .A(n_40), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_62), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_26), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_5), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_11), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_58), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_36), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_49), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_47), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_6), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_19), .Y(n_110) );
INVxp33_ASAP7_75t_L g111 ( .A(n_9), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_25), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_15), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_34), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_66), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_18), .Y(n_116) );
INVx4_ASAP7_75t_R g117 ( .A(n_46), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_6), .Y(n_118) );
INVxp67_ASAP7_75t_SL g119 ( .A(n_13), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_0), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_33), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_2), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_16), .Y(n_123) );
INVxp33_ASAP7_75t_SL g124 ( .A(n_32), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_4), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_51), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_79), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_118), .B(n_1), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_90), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_90), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_81), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_81), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_82), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_82), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_106), .B(n_1), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_83), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
BUFx2_ASAP7_75t_L g139 ( .A(n_123), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_84), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g141 ( .A1(n_111), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_84), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_123), .B(n_3), .Y(n_143) );
OAI22xp5_ASAP7_75t_SL g144 ( .A1(n_99), .A2(n_5), .B1(n_7), .B2(n_8), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_85), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_85), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_86), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_118), .B(n_7), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_97), .B(n_8), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_122), .B(n_9), .Y(n_150) );
XOR2xp5_ASAP7_75t_L g151 ( .A(n_88), .B(n_10), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_86), .Y(n_152) );
AND3x2_ASAP7_75t_L g153 ( .A(n_122), .B(n_10), .C(n_11), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_89), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_89), .Y(n_155) );
AND2x4_ASAP7_75t_SL g156 ( .A(n_94), .B(n_38), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_93), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_93), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_95), .B(n_12), .Y(n_159) );
AOI22xp33_ASAP7_75t_SL g160 ( .A1(n_104), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_95), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_108), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_125), .B(n_14), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_103), .B(n_15), .Y(n_164) );
XNOR2xp5_ASAP7_75t_SL g165 ( .A(n_80), .B(n_16), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_108), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_121), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_121), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_101), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_107), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_131), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_131), .Y(n_172) );
NAND2x1p5_ASAP7_75t_L g173 ( .A(n_139), .B(n_125), .Y(n_173) );
NAND2x1p5_ASAP7_75t_L g174 ( .A(n_139), .B(n_109), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_131), .Y(n_175) );
INVx4_ASAP7_75t_L g176 ( .A(n_129), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_131), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_131), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_149), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_131), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_129), .Y(n_181) );
OAI21xp33_ASAP7_75t_L g182 ( .A1(n_127), .A2(n_116), .B(n_96), .Y(n_182) );
AND2x6_ASAP7_75t_L g183 ( .A(n_129), .B(n_110), .Y(n_183) );
NAND3xp33_ASAP7_75t_L g184 ( .A(n_149), .B(n_80), .C(n_87), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_129), .Y(n_185) );
OR2x2_ASAP7_75t_L g186 ( .A(n_136), .B(n_113), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_148), .B(n_120), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_127), .B(n_100), .Y(n_188) );
INVxp33_ASAP7_75t_L g189 ( .A(n_143), .Y(n_189) );
INVx2_ASAP7_75t_SL g190 ( .A(n_142), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_148), .B(n_119), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_142), .B(n_115), .Y(n_192) );
OR2x6_ASAP7_75t_L g193 ( .A(n_144), .B(n_112), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_148), .Y(n_194) );
INVx1_ASAP7_75t_SL g195 ( .A(n_156), .Y(n_195) );
BUFx10_ASAP7_75t_L g196 ( .A(n_148), .Y(n_196) );
INVxp67_ASAP7_75t_L g197 ( .A(n_128), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_128), .B(n_114), .Y(n_198) );
INVxp67_ASAP7_75t_L g199 ( .A(n_132), .Y(n_199) );
INVxp67_ASAP7_75t_L g200 ( .A(n_132), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_133), .B(n_124), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_150), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_150), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_133), .B(n_92), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_150), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_142), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_150), .B(n_105), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_163), .B(n_91), .Y(n_208) );
INVx4_ASAP7_75t_L g209 ( .A(n_163), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_135), .B(n_87), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_163), .A2(n_126), .B1(n_102), .B2(n_98), .Y(n_211) );
INVx5_ASAP7_75t_L g212 ( .A(n_163), .Y(n_212) );
OR2x2_ASAP7_75t_SL g213 ( .A(n_151), .B(n_17), .Y(n_213) );
BUFx3_ASAP7_75t_L g214 ( .A(n_169), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_142), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_155), .Y(n_216) );
INVx2_ASAP7_75t_SL g217 ( .A(n_155), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_135), .B(n_53), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_138), .B(n_55), .Y(n_219) );
INVx4_ASAP7_75t_L g220 ( .A(n_155), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_155), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_158), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_158), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_158), .Y(n_224) );
INVx1_ASAP7_75t_SL g225 ( .A(n_156), .Y(n_225) );
INVx1_ASAP7_75t_SL g226 ( .A(n_151), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_138), .B(n_17), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_220), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_220), .Y(n_229) );
BUFx4f_ASAP7_75t_SL g230 ( .A(n_195), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_215), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_216), .Y(n_232) );
BUFx8_ASAP7_75t_L g233 ( .A(n_188), .Y(n_233) );
BUFx2_ASAP7_75t_L g234 ( .A(n_173), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_176), .Y(n_235) );
NOR2x1_ASAP7_75t_R g236 ( .A(n_191), .B(n_165), .Y(n_236) );
BUFx3_ASAP7_75t_L g237 ( .A(n_183), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_179), .A2(n_141), .B1(n_144), .B2(n_140), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_197), .B(n_146), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_221), .Y(n_240) );
NOR2xp33_ASAP7_75t_R g241 ( .A(n_225), .B(n_168), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_181), .Y(n_242) );
BUFx2_ASAP7_75t_L g243 ( .A(n_173), .Y(n_243) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_174), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_222), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_172), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_222), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_185), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_223), .Y(n_249) );
BUFx4f_ASAP7_75t_L g250 ( .A(n_183), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_190), .Y(n_251) );
BUFx2_ASAP7_75t_L g252 ( .A(n_174), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_194), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_197), .B(n_146), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_196), .B(n_164), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_199), .B(n_166), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_187), .A2(n_166), .B1(n_140), .B2(n_161), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_206), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_191), .B(n_153), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_202), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_201), .A2(n_145), .B1(n_147), .B2(n_154), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_183), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_183), .Y(n_263) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_186), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_199), .B(n_147), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_176), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_196), .B(n_161), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_226), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_223), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_201), .A2(n_145), .B1(n_154), .B2(n_162), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_183), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_172), .Y(n_272) );
BUFx2_ASAP7_75t_L g273 ( .A(n_209), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_203), .Y(n_274) );
BUFx8_ASAP7_75t_L g275 ( .A(n_187), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_204), .A2(n_162), .B1(n_159), .B2(n_168), .Y(n_276) );
INVx2_ASAP7_75t_SL g277 ( .A(n_212), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_189), .B(n_170), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_200), .B(n_168), .Y(n_279) );
INVx5_ASAP7_75t_L g280 ( .A(n_209), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_171), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_205), .Y(n_282) );
INVx2_ASAP7_75t_SL g283 ( .A(n_212), .Y(n_283) );
INVx3_ASAP7_75t_L g284 ( .A(n_212), .Y(n_284) );
INVx2_ASAP7_75t_SL g285 ( .A(n_212), .Y(n_285) );
OAI21xp5_ASAP7_75t_L g286 ( .A1(n_200), .A2(n_168), .B(n_170), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_217), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_172), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_227), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_171), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_211), .Y(n_291) );
NAND3x1_ASAP7_75t_L g292 ( .A(n_238), .B(n_213), .C(n_165), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_264), .B(n_189), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_239), .A2(n_204), .B(n_192), .Y(n_294) );
INVx2_ASAP7_75t_SL g295 ( .A(n_275), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_280), .Y(n_296) );
AND2x2_ASAP7_75t_SL g297 ( .A(n_250), .B(n_208), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_232), .Y(n_298) );
O2A1O1Ixp5_ASAP7_75t_L g299 ( .A1(n_286), .A2(n_219), .B(n_218), .C(n_192), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_275), .Y(n_300) );
OR2x6_ASAP7_75t_L g301 ( .A(n_234), .B(n_193), .Y(n_301) );
BUFx12f_ASAP7_75t_L g302 ( .A(n_268), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_278), .B(n_187), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_231), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_231), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_240), .Y(n_306) );
NOR2xp33_ASAP7_75t_R g307 ( .A(n_275), .B(n_207), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_257), .B(n_210), .Y(n_308) );
INVx5_ASAP7_75t_L g309 ( .A(n_280), .Y(n_309) );
INVx5_ASAP7_75t_L g310 ( .A(n_280), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_234), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_240), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_237), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_254), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_242), .A2(n_193), .B1(n_207), .B2(n_208), .Y(n_315) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_237), .Y(n_316) );
NAND2x1p5_ASAP7_75t_L g317 ( .A(n_280), .B(n_137), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_235), .Y(n_318) );
BUFx2_ASAP7_75t_SL g319 ( .A(n_244), .Y(n_319) );
AND2x4_ASAP7_75t_L g320 ( .A(n_259), .B(n_184), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_280), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_261), .B(n_198), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_273), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_259), .B(n_198), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_243), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_228), .Y(n_326) );
OAI21xp33_ASAP7_75t_L g327 ( .A1(n_289), .A2(n_182), .B(n_193), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_256), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_259), .B(n_137), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_228), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_235), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_265), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_262), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_262), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_243), .A2(n_160), .B1(n_219), .B2(n_218), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_270), .B(n_134), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_289), .B(n_134), .Y(n_337) );
INVx4_ASAP7_75t_L g338 ( .A(n_230), .Y(n_338) );
BUFx2_ASAP7_75t_L g339 ( .A(n_233), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_279), .A2(n_175), .B(n_177), .Y(n_340) );
OR2x6_ASAP7_75t_L g341 ( .A(n_252), .B(n_152), .Y(n_341) );
NAND2xp33_ASAP7_75t_L g342 ( .A(n_241), .B(n_172), .Y(n_342) );
OR2x6_ASAP7_75t_L g343 ( .A(n_252), .B(n_152), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_229), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_263), .Y(n_345) );
NAND4xp25_ASAP7_75t_L g346 ( .A(n_315), .B(n_276), .C(n_236), .D(n_167), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_304), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_314), .B(n_233), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_309), .Y(n_349) );
CKINVDCx6p67_ASAP7_75t_R g350 ( .A(n_319), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_309), .B(n_263), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_324), .A2(n_291), .B1(n_233), .B2(n_268), .Y(n_352) );
OAI22xp33_ASAP7_75t_L g353 ( .A1(n_293), .A2(n_291), .B1(n_250), .B2(n_271), .Y(n_353) );
BUFx2_ASAP7_75t_L g354 ( .A(n_307), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_324), .A2(n_273), .B1(n_266), .B2(n_235), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_304), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_306), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_309), .B(n_271), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_328), .A2(n_250), .B1(n_260), .B2(n_248), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_315), .A2(n_266), .B1(n_253), .B2(n_260), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_332), .B(n_253), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_306), .Y(n_362) );
OAI22xp33_ASAP7_75t_L g363 ( .A1(n_301), .A2(n_242), .B1(n_282), .B2(n_274), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_307), .Y(n_364) );
OAI221xp5_ASAP7_75t_L g365 ( .A1(n_322), .A2(n_255), .B1(n_274), .B2(n_282), .C(n_248), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_320), .B(n_267), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_303), .B(n_229), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_305), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_312), .Y(n_369) );
AOI22xp33_ASAP7_75t_SL g370 ( .A1(n_300), .A2(n_266), .B1(n_287), .B2(n_284), .Y(n_370) );
AOI21xp33_ASAP7_75t_L g371 ( .A1(n_308), .A2(n_285), .B(n_283), .Y(n_371) );
O2A1O1Ixp33_ASAP7_75t_L g372 ( .A1(n_327), .A2(n_157), .B(n_167), .C(n_251), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_309), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_298), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_337), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_329), .B(n_287), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_302), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_326), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_326), .Y(n_379) );
NAND2x1p5_ASAP7_75t_L g380 ( .A(n_310), .B(n_284), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_347), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_347), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_374), .B(n_320), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g384 ( .A1(n_346), .A2(n_294), .B1(n_295), .B2(n_329), .C(n_336), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_375), .B(n_341), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_348), .Y(n_386) );
AOI22xp33_ASAP7_75t_SL g387 ( .A1(n_354), .A2(n_339), .B1(n_301), .B2(n_343), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_356), .B(n_341), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_375), .A2(n_343), .B1(n_341), .B2(n_335), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_346), .A2(n_292), .B1(n_301), .B2(n_343), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_356), .B(n_297), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_363), .A2(n_297), .B1(n_323), .B2(n_311), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_357), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_357), .Y(n_394) );
INVx4_ASAP7_75t_L g395 ( .A(n_350), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_359), .A2(n_299), .B(n_340), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_354), .A2(n_323), .B1(n_294), .B2(n_325), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g398 ( .A1(n_364), .A2(n_338), .B1(n_342), .B2(n_321), .Y(n_398) );
OR2x6_ASAP7_75t_L g399 ( .A(n_362), .B(n_313), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_362), .B(n_317), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_350), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_378), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_365), .A2(n_338), .B1(n_331), .B2(n_321), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_374), .A2(n_299), .B1(n_157), .B2(n_258), .C(n_130), .Y(n_404) );
OAI211xp5_ASAP7_75t_SL g405 ( .A1(n_352), .A2(n_130), .B(n_296), .C(n_287), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_364), .A2(n_317), .B1(n_310), .B2(n_296), .Y(n_406) );
INVx2_ASAP7_75t_SL g407 ( .A(n_351), .Y(n_407) );
BUFx4f_ASAP7_75t_SL g408 ( .A(n_349), .Y(n_408) );
INVx3_ASAP7_75t_L g409 ( .A(n_351), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_402), .B(n_378), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_402), .B(n_379), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_381), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_386), .B(n_353), .Y(n_413) );
OAI211xp5_ASAP7_75t_L g414 ( .A1(n_390), .A2(n_370), .B(n_366), .C(n_355), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_381), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_389), .A2(n_360), .B1(n_361), .B2(n_379), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_388), .Y(n_417) );
BUFx3_ASAP7_75t_L g418 ( .A(n_408), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_396), .A2(n_342), .B(n_371), .Y(n_419) );
NAND3xp33_ASAP7_75t_L g420 ( .A(n_384), .B(n_372), .C(n_368), .Y(n_420) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_399), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_402), .Y(n_422) );
AOI22xp33_ASAP7_75t_SL g423 ( .A1(n_389), .A2(n_373), .B1(n_349), .B2(n_369), .Y(n_423) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_399), .Y(n_424) );
AOI322xp5_ASAP7_75t_L g425 ( .A1(n_390), .A2(n_369), .A3(n_368), .B1(n_377), .B2(n_376), .C1(n_349), .C2(n_373), .Y(n_425) );
BUFx2_ASAP7_75t_L g426 ( .A(n_399), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_393), .Y(n_427) );
OAI21xp5_ASAP7_75t_L g428 ( .A1(n_405), .A2(n_367), .B(n_340), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_393), .B(n_373), .Y(n_429) );
NAND3xp33_ASAP7_75t_L g430 ( .A(n_404), .B(n_158), .C(n_169), .Y(n_430) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_387), .A2(n_392), .B1(n_397), .B2(n_403), .C(n_383), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_381), .Y(n_432) );
OAI211xp5_ASAP7_75t_SL g433 ( .A1(n_401), .A2(n_224), .B(n_175), .C(n_177), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_385), .A2(n_376), .B1(n_351), .B2(n_358), .Y(n_434) );
AO21x2_ASAP7_75t_L g435 ( .A1(n_382), .A2(n_180), .B(n_178), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_382), .Y(n_436) );
OAI211xp5_ASAP7_75t_SL g437 ( .A1(n_398), .A2(n_224), .B(n_180), .C(n_178), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_388), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_382), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_394), .Y(n_440) );
INVx2_ASAP7_75t_SL g441 ( .A(n_395), .Y(n_441) );
NAND4xp25_ASAP7_75t_L g442 ( .A(n_395), .B(n_214), .C(n_331), .D(n_318), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_385), .A2(n_358), .B1(n_351), .B2(n_169), .Y(n_443) );
NAND4xp25_ASAP7_75t_L g444 ( .A(n_425), .B(n_395), .C(n_391), .D(n_409), .Y(n_444) );
BUFx2_ASAP7_75t_L g445 ( .A(n_426), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_412), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_421), .B(n_394), .Y(n_447) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_425), .B(n_413), .C(n_420), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_410), .B(n_394), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_422), .Y(n_450) );
AND4x1_ASAP7_75t_L g451 ( .A(n_443), .B(n_395), .C(n_391), .D(n_400), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_412), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_426), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_415), .Y(n_454) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_422), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_415), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_427), .B(n_400), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_421), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_427), .Y(n_459) );
INVx2_ASAP7_75t_SL g460 ( .A(n_441), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_410), .B(n_409), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_421), .B(n_409), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_432), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_418), .B(n_377), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_439), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_411), .B(n_407), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_432), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_436), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_411), .B(n_409), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_436), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_440), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_429), .Y(n_472) );
OAI31xp33_ASAP7_75t_SL g473 ( .A1(n_423), .A2(n_406), .A3(n_358), .B(n_407), .Y(n_473) );
OAI22xp33_ASAP7_75t_L g474 ( .A1(n_431), .A2(n_399), .B1(n_310), .B2(n_380), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_440), .B(n_399), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_416), .A2(n_158), .B1(n_169), .B2(n_358), .Y(n_476) );
OAI221xp5_ASAP7_75t_SL g477 ( .A1(n_414), .A2(n_284), .B1(n_344), .B2(n_330), .C(n_285), .Y(n_477) );
BUFx3_ASAP7_75t_L g478 ( .A(n_441), .Y(n_478) );
INVx3_ASAP7_75t_L g479 ( .A(n_421), .Y(n_479) );
INVx3_ASAP7_75t_L g480 ( .A(n_421), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_439), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_429), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_424), .Y(n_483) );
AOI21x1_ASAP7_75t_L g484 ( .A1(n_419), .A2(n_344), .B(n_330), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_417), .B(n_158), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_438), .B(n_169), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_420), .A2(n_380), .B1(n_169), .B2(n_310), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_435), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_434), .B(n_380), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_434), .B(n_18), .Y(n_490) );
INVx1_ASAP7_75t_SL g491 ( .A(n_418), .Y(n_491) );
INVx3_ASAP7_75t_SL g492 ( .A(n_478), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_461), .B(n_424), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_459), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_491), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_472), .B(n_424), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_459), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_461), .B(n_424), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_446), .Y(n_499) );
NAND3xp33_ASAP7_75t_L g500 ( .A(n_448), .B(n_428), .C(n_442), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_469), .B(n_424), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_469), .B(n_435), .Y(n_502) );
BUFx3_ASAP7_75t_L g503 ( .A(n_478), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_455), .B(n_435), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_482), .B(n_430), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_450), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_475), .B(n_430), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_450), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_458), .B(n_20), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_475), .B(n_22), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_457), .B(n_23), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_464), .B(n_27), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_463), .Y(n_513) );
INVx3_ASAP7_75t_L g514 ( .A(n_478), .Y(n_514) );
NOR3xp33_ASAP7_75t_SL g515 ( .A(n_448), .B(n_437), .C(n_433), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_463), .B(n_467), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_446), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_467), .B(n_28), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_468), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_458), .B(n_29), .Y(n_520) );
OAI31xp33_ASAP7_75t_L g521 ( .A1(n_474), .A2(n_283), .A3(n_277), .B(n_214), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_468), .B(n_31), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_470), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_457), .B(n_35), .Y(n_524) );
OAI332xp33_ASAP7_75t_L g525 ( .A1(n_490), .A2(n_277), .A3(n_117), .B1(n_245), .B2(n_249), .B3(n_247), .C1(n_269), .C2(n_281), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_470), .B(n_37), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_460), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_471), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_471), .Y(n_529) );
INVx1_ASAP7_75t_SL g530 ( .A(n_460), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_481), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_446), .Y(n_532) );
NAND3xp33_ASAP7_75t_L g533 ( .A(n_477), .B(n_345), .C(n_334), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_483), .B(n_39), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_466), .B(n_45), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_481), .Y(n_536) );
NOR4xp75_ASAP7_75t_L g537 ( .A(n_489), .B(n_56), .C(n_59), .D(n_64), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_483), .B(n_65), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_449), .B(n_67), .Y(n_539) );
OAI21xp5_ASAP7_75t_SL g540 ( .A1(n_473), .A2(n_345), .B(n_334), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_452), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_445), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_452), .Y(n_543) );
OR2x6_ASAP7_75t_L g544 ( .A(n_445), .B(n_345), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_452), .B(n_69), .Y(n_545) );
OAI31xp33_ASAP7_75t_L g546 ( .A1(n_444), .A2(n_72), .A3(n_73), .B(n_74), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_454), .B(n_465), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_454), .B(n_77), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_499), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_493), .B(n_458), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_516), .B(n_485), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_495), .Y(n_552) );
NAND3xp33_ASAP7_75t_L g553 ( .A(n_500), .B(n_451), .C(n_485), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_527), .B(n_453), .Y(n_554) );
INVx3_ASAP7_75t_L g555 ( .A(n_514), .Y(n_555) );
AND3x1_ASAP7_75t_L g556 ( .A(n_546), .B(n_451), .C(n_487), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_494), .Y(n_557) );
AOI21xp33_ASAP7_75t_L g558 ( .A1(n_530), .A2(n_486), .B(n_458), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_499), .Y(n_559) );
NAND3xp33_ASAP7_75t_L g560 ( .A(n_515), .B(n_487), .C(n_476), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_493), .B(n_480), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_516), .B(n_453), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_494), .B(n_465), .Y(n_563) );
INVx1_ASAP7_75t_SL g564 ( .A(n_492), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_542), .B(n_465), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_498), .B(n_480), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_497), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_498), .B(n_480), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_501), .B(n_480), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_525), .B(n_479), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_501), .B(n_479), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_502), .B(n_479), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_497), .Y(n_573) );
NAND2x1p5_ASAP7_75t_L g574 ( .A(n_503), .B(n_447), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_502), .B(n_479), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_547), .B(n_447), .Y(n_576) );
OAI21xp5_ASAP7_75t_L g577 ( .A1(n_540), .A2(n_447), .B(n_488), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_547), .B(n_447), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_496), .B(n_456), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_503), .Y(n_580) );
NOR3xp33_ASAP7_75t_L g581 ( .A(n_535), .B(n_484), .C(n_488), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_507), .B(n_456), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_506), .B(n_456), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_492), .Y(n_584) );
OAI32xp33_ASAP7_75t_L g585 ( .A1(n_514), .A2(n_454), .A3(n_488), .B1(n_462), .B2(n_78), .Y(n_585) );
INVxp67_ASAP7_75t_L g586 ( .A(n_514), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_531), .B(n_462), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_531), .B(n_462), .Y(n_588) );
OAI211xp5_ASAP7_75t_SL g589 ( .A1(n_505), .A2(n_245), .B(n_269), .C(n_247), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_506), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_492), .B(n_462), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_536), .B(n_484), .Y(n_592) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_510), .B(n_345), .C(n_334), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_536), .B(n_334), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_507), .B(n_249), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_504), .B(n_333), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_517), .Y(n_597) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_504), .Y(n_598) );
INVx3_ASAP7_75t_L g599 ( .A(n_517), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_508), .B(n_333), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g601 ( .A1(n_521), .A2(n_333), .B(n_316), .C(n_313), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_512), .A2(n_333), .B1(n_316), .B2(n_313), .Y(n_602) );
XOR2x2_ASAP7_75t_SL g603 ( .A(n_574), .B(n_520), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_551), .B(n_541), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_598), .B(n_523), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_550), .B(n_523), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_556), .A2(n_533), .B(n_544), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_564), .B(n_543), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_582), .B(n_508), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_557), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_580), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_SL g612 ( .A1(n_584), .A2(n_511), .B(n_524), .C(n_519), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_550), .B(n_528), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_561), .B(n_528), .Y(n_614) );
INVx2_ASAP7_75t_SL g615 ( .A(n_555), .Y(n_615) );
OAI21xp5_ASAP7_75t_SL g616 ( .A1(n_553), .A2(n_510), .B(n_518), .Y(n_616) );
AOI21xp5_ASAP7_75t_SL g617 ( .A1(n_601), .A2(n_570), .B(n_593), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_582), .B(n_519), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_562), .B(n_513), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_561), .B(n_529), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_567), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_555), .B(n_543), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_573), .B(n_513), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_566), .B(n_529), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_590), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_599), .Y(n_626) );
INVx1_ASAP7_75t_SL g627 ( .A(n_552), .Y(n_627) );
AOI21xp33_ASAP7_75t_L g628 ( .A1(n_570), .A2(n_539), .B(n_518), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_579), .B(n_541), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_563), .Y(n_630) );
NAND3x1_ASAP7_75t_L g631 ( .A(n_555), .B(n_537), .C(n_522), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_554), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_583), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_586), .B(n_522), .Y(n_634) );
NAND4xp25_ASAP7_75t_L g635 ( .A(n_560), .B(n_526), .C(n_520), .D(n_509), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_565), .Y(n_636) );
XOR2x2_ASAP7_75t_L g637 ( .A(n_591), .B(n_520), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_572), .B(n_532), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_572), .B(n_532), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_587), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_575), .B(n_526), .Y(n_641) );
AOI211xp5_ASAP7_75t_SL g642 ( .A1(n_591), .A2(n_509), .B(n_534), .C(n_538), .Y(n_642) );
INVx2_ASAP7_75t_SL g643 ( .A(n_574), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_575), .B(n_538), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_588), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_566), .B(n_544), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_599), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_568), .B(n_509), .Y(n_648) );
AOI21xp5_ASAP7_75t_SL g649 ( .A1(n_601), .A2(n_548), .B(n_545), .Y(n_649) );
OAI21xp5_ASAP7_75t_SL g650 ( .A1(n_577), .A2(n_534), .B(n_548), .Y(n_650) );
NAND2x1p5_ASAP7_75t_L g651 ( .A(n_602), .B(n_545), .Y(n_651) );
XNOR2x1_ASAP7_75t_L g652 ( .A(n_568), .B(n_544), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g653 ( .A1(n_558), .A2(n_544), .B1(n_316), .B2(n_313), .C(n_288), .Y(n_653) );
AOI222xp33_ASAP7_75t_L g654 ( .A1(n_595), .A2(n_316), .B1(n_281), .B2(n_290), .C1(n_288), .C2(n_272), .Y(n_654) );
XOR2x2_ASAP7_75t_L g655 ( .A(n_576), .B(n_246), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_599), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_549), .Y(n_657) );
XOR2x2_ASAP7_75t_L g658 ( .A(n_576), .B(n_246), .Y(n_658) );
OA22x2_ASAP7_75t_L g659 ( .A1(n_569), .A2(n_290), .B1(n_272), .B2(n_288), .Y(n_659) );
NOR2xp67_ASAP7_75t_L g660 ( .A(n_549), .B(n_246), .Y(n_660) );
OAI211xp5_ASAP7_75t_L g661 ( .A1(n_589), .A2(n_246), .B(n_272), .C(n_288), .Y(n_661) );
XOR2x2_ASAP7_75t_L g662 ( .A(n_578), .B(n_246), .Y(n_662) );
NOR4xp25_ASAP7_75t_L g663 ( .A(n_595), .B(n_272), .C(n_288), .D(n_592), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_559), .Y(n_664) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_578), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_605), .Y(n_666) );
OAI221xp5_ASAP7_75t_L g667 ( .A1(n_616), .A2(n_635), .B1(n_617), .B2(n_607), .C(n_650), .Y(n_667) );
AOI221xp5_ASAP7_75t_SL g668 ( .A1(n_627), .A2(n_611), .B1(n_632), .B2(n_636), .C(n_640), .Y(n_668) );
INVx3_ASAP7_75t_L g669 ( .A(n_637), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_630), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_633), .Y(n_671) );
INVx2_ASAP7_75t_SL g672 ( .A(n_629), .Y(n_672) );
AOI21xp33_ASAP7_75t_SL g673 ( .A1(n_603), .A2(n_608), .B(n_659), .Y(n_673) );
NAND4xp25_ASAP7_75t_L g674 ( .A(n_628), .B(n_642), .C(n_612), .D(n_650), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_608), .A2(n_612), .B(n_637), .Y(n_675) );
OAI222xp33_ASAP7_75t_L g676 ( .A1(n_603), .A2(n_615), .B1(n_665), .B2(n_651), .C1(n_659), .C2(n_643), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_645), .B(n_619), .Y(n_677) );
NOR3xp33_ASAP7_75t_L g678 ( .A(n_661), .B(n_653), .C(n_615), .Y(n_678) );
OAI221xp5_ASAP7_75t_SL g679 ( .A1(n_649), .A2(n_648), .B1(n_641), .B2(n_663), .C(n_644), .Y(n_679) );
O2A1O1Ixp33_ASAP7_75t_L g680 ( .A1(n_675), .A2(n_585), .B(n_622), .C(n_663), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_667), .A2(n_652), .B1(n_631), .B2(n_651), .Y(n_681) );
OAI32xp33_ASAP7_75t_L g682 ( .A1(n_669), .A2(n_634), .A3(n_656), .B1(n_622), .B2(n_604), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_670), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_671), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_669), .B(n_620), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_667), .A2(n_610), .B1(n_621), .B2(n_625), .C(n_634), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_668), .A2(n_609), .B1(n_618), .B2(n_647), .C(n_624), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_681), .A2(n_674), .B1(n_666), .B2(n_678), .Y(n_688) );
OAI22x1_ASAP7_75t_L g689 ( .A1(n_683), .A2(n_676), .B1(n_673), .B2(n_672), .Y(n_689) );
XOR2xp5_ASAP7_75t_L g690 ( .A(n_685), .B(n_655), .Y(n_690) );
NOR3x1_ASAP7_75t_SL g691 ( .A(n_686), .B(n_679), .C(n_631), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_684), .A2(n_677), .B1(n_658), .B2(n_662), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_689), .A2(n_687), .B1(n_581), .B2(n_646), .Y(n_693) );
AND3x1_ASAP7_75t_L g694 ( .A(n_688), .B(n_680), .C(n_682), .Y(n_694) );
NOR4xp75_ASAP7_75t_L g695 ( .A(n_691), .B(n_639), .C(n_638), .D(n_614), .Y(n_695) );
OAI221xp5_ASAP7_75t_L g696 ( .A1(n_693), .A2(n_692), .B1(n_690), .B2(n_656), .C(n_626), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_694), .A2(n_626), .B1(n_657), .B2(n_664), .C(n_623), .Y(n_697) );
AO22x2_ASAP7_75t_L g698 ( .A1(n_696), .A2(n_695), .B1(n_613), .B2(n_606), .Y(n_698) );
OAI22x1_ASAP7_75t_L g699 ( .A1(n_697), .A2(n_569), .B1(n_571), .B2(n_559), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_698), .A2(n_660), .B1(n_596), .B2(n_597), .Y(n_700) );
AOI22x1_ASAP7_75t_L g701 ( .A1(n_700), .A2(n_699), .B1(n_654), .B2(n_571), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_701), .A2(n_600), .B1(n_597), .B2(n_594), .C(n_272), .Y(n_702) );
endmodule