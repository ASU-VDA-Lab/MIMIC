module fake_jpeg_25929_n_312 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_312);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_20),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_37),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_45),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_24),
.B(n_21),
.Y(n_45)
);

CKINVDCx12_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_47),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_46),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_49),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_22),
.B1(n_30),
.B2(n_24),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_55),
.B1(n_56),
.B2(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_58),
.B(n_63),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_51),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_30),
.B1(n_38),
.B2(n_44),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_22),
.B1(n_29),
.B2(n_28),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

OR2x2_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_22),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_26),
.Y(n_71)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_36),
.A2(n_14),
.B1(n_21),
.B2(n_28),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_72),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_44),
.B1(n_37),
.B2(n_43),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_55),
.B1(n_64),
.B2(n_49),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_54),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_71),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_39),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_78),
.Y(n_87)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_39),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_54),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_39),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_53),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_84),
.A2(n_55),
.B1(n_65),
.B2(n_63),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_88),
.B1(n_89),
.B2(n_77),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_84),
.A2(n_58),
.B1(n_61),
.B2(n_50),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_96),
.Y(n_139)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_44),
.Y(n_98)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_46),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_69),
.B(n_58),
.Y(n_100)
);

OAI32xp33_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_21),
.A3(n_19),
.B1(n_11),
.B2(n_13),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_56),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_101),
.A2(n_109),
.B(n_79),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_49),
.B1(n_64),
.B2(n_62),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_49),
.Y(n_106)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_31),
.C(n_25),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_33),
.C(n_17),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_62),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_108),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_32),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_110),
.A2(n_113),
.B(n_130),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_81),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_114),
.B(n_118),
.C(n_120),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_43),
.B1(n_36),
.B2(n_70),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_81),
.B1(n_73),
.B2(n_78),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_122),
.B1(n_124),
.B2(n_128),
.Y(n_149)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_90),
.C(n_97),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_93),
.A2(n_43),
.B1(n_76),
.B2(n_80),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_109),
.B(n_94),
.C(n_87),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_82),
.B1(n_27),
.B2(n_26),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_11),
.B(n_19),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_29),
.B1(n_27),
.B2(n_11),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_7),
.C(n_10),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_137),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_19),
.B1(n_40),
.B2(n_32),
.Y(n_134)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_33),
.B1(n_32),
.B2(n_31),
.Y(n_136)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_90),
.A2(n_13),
.B1(n_16),
.B2(n_15),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_95),
.A2(n_33),
.B1(n_31),
.B2(n_13),
.Y(n_138)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_95),
.Y(n_141)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_151),
.Y(n_178)
);

CKINVDCx12_ASAP7_75t_R g144 ( 
.A(n_116),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_144),
.Y(n_200)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_130),
.A2(n_91),
.B(n_106),
.C(n_108),
.D(n_109),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_145),
.B(n_12),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_125),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_146),
.Y(n_188)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_158),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_155),
.A2(n_12),
.B(n_15),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_87),
.Y(n_156)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

OAI31xp33_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_104),
.A3(n_94),
.B(n_18),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_157),
.A2(n_171),
.B(n_15),
.Y(n_196)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_16),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_161),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_121),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_132),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_164),
.Y(n_195)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_166),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_137),
.B(n_16),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_134),
.B(n_17),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_169),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_23),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_113),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_172),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_135),
.A2(n_18),
.B(n_8),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_121),
.B(n_18),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_114),
.B(n_120),
.Y(n_173)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_23),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_174),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_110),
.B(n_23),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_118),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_162),
.C(n_173),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_158),
.A2(n_135),
.B1(n_124),
.B2(n_128),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_SL g223 ( 
.A(n_180),
.B(n_183),
.C(n_193),
.Y(n_223)
);

AOI21x1_ASAP7_75t_SL g183 ( 
.A1(n_145),
.A2(n_123),
.B(n_140),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_17),
.B1(n_15),
.B2(n_23),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_184),
.A2(n_186),
.B1(n_150),
.B2(n_143),
.Y(n_221)
);

BUFx24_ASAP7_75t_SL g185 ( 
.A(n_141),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_191),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_152),
.A2(n_17),
.B1(n_15),
.B2(n_12),
.Y(n_186)
);

OA21x2_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_12),
.B(n_17),
.Y(n_187)
);

AO22x1_ASAP7_75t_SL g225 ( 
.A1(n_187),
.A2(n_153),
.B1(n_160),
.B2(n_151),
.Y(n_225)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g194 ( 
.A(n_147),
.B(n_10),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_202),
.Y(n_211)
);

AO22x1_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_157),
.B1(n_155),
.B2(n_167),
.Y(n_212)
);

AOI21x1_ASAP7_75t_SL g216 ( 
.A1(n_199),
.A2(n_169),
.B(n_154),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_170),
.A2(n_10),
.B(n_9),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_184),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_161),
.Y(n_206)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_201),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_210),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_212),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_148),
.C(n_147),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_219),
.C(n_193),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_195),
.A2(n_148),
.B1(n_165),
.B2(n_159),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

A2O1A1O1Ixp25_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_163),
.B(n_172),
.C(n_171),
.D(n_166),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_202),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_187),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_198),
.A2(n_159),
.B1(n_168),
.B2(n_164),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_221),
.B1(n_222),
.B2(n_224),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_178),
.B(n_149),
.C(n_168),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_220),
.B(n_225),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_192),
.B1(n_194),
.B2(n_196),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_149),
.B1(n_150),
.B2(n_153),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_181),
.A2(n_163),
.B1(n_9),
.B2(n_8),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_226),
.A2(n_203),
.B1(n_191),
.B2(n_9),
.Y(n_247)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_182),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_227),
.B(n_228),
.Y(n_238)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_240),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_241),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_189),
.C(n_197),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_233),
.C(n_239),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_188),
.C(n_190),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_204),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_236),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_211),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_190),
.C(n_186),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_223),
.B(n_200),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_200),
.B(n_187),
.Y(n_242)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_247),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_243),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_249),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_231),
.A2(n_224),
.B1(n_217),
.B2(n_214),
.Y(n_250)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_235),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_252),
.Y(n_267)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_238),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_208),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_225),
.C(n_206),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_259),
.C(n_241),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_225),
.C(n_223),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_221),
.B1(n_212),
.B2(n_216),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_262),
.A2(n_244),
.B1(n_246),
.B2(n_245),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_232),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_263),
.B(n_264),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_249),
.B1(n_250),
.B2(n_257),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_209),
.Y(n_268)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_268),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_229),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_270),
.B(n_272),
.Y(n_287)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_215),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_9),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_274),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_0),
.C(n_1),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_7),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_0),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_249),
.B(n_259),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_276),
.B(n_280),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_256),
.B(n_253),
.Y(n_277)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_284),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_260),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_265),
.A2(n_262),
.B(n_7),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_0),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_264),
.A2(n_7),
.B1(n_1),
.B2(n_2),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_286),
.A2(n_274),
.B1(n_1),
.B2(n_2),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_290),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_276),
.A2(n_263),
.B(n_270),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_292),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_0),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_2),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_294),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_287),
.A2(n_2),
.B(n_3),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_2),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_3),
.Y(n_303)
);

AOI32xp33_ASAP7_75t_L g298 ( 
.A1(n_291),
.A2(n_296),
.A3(n_297),
.B1(n_285),
.B2(n_280),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_298),
.B(n_303),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_SL g302 ( 
.A(n_296),
.B(n_279),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_302),
.A2(n_3),
.B(n_4),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_288),
.C(n_4),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_305),
.C(n_300),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_306),
.B(n_301),
.Y(n_308)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_3),
.B(n_4),
.Y(n_309)
);

NOR3xp33_ASAP7_75t_SL g310 ( 
.A(n_309),
.B(n_5),
.C(n_6),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_5),
.B(n_6),
.Y(n_311)
);

FAx1_ASAP7_75t_SL g312 ( 
.A(n_311),
.B(n_6),
.CI(n_211),
.CON(n_312),
.SN(n_312)
);


endmodule