module real_jpeg_22572_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_332, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_332;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_0),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_0),
.A2(n_9),
.B1(n_49),
.B2(n_61),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_0),
.A2(n_26),
.B1(n_33),
.B2(n_49),
.Y(n_284)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_2),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_2),
.A2(n_34),
.B1(n_46),
.B2(n_47),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_2),
.A2(n_9),
.B1(n_34),
.B2(n_61),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_3),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_3),
.B(n_29),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_3),
.A2(n_9),
.B(n_14),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_129),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_3),
.A2(n_103),
.B1(n_108),
.B2(n_189),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_3),
.B(n_85),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_3),
.B(n_31),
.Y(n_216)
);

AOI21xp33_ASAP7_75t_L g220 ( 
.A1(n_3),
.A2(n_31),
.B(n_216),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_4),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_4),
.A2(n_26),
.B1(n_33),
.B2(n_124),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_4),
.A2(n_9),
.B1(n_61),
.B2(n_124),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_124),
.Y(n_204)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_6),
.A2(n_26),
.B1(n_33),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_6),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_131),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_131),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_6),
.A2(n_9),
.B1(n_61),
.B2(n_131),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_7),
.B(n_61),
.Y(n_104)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_7),
.Y(n_108)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_7),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_8),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_8),
.A2(n_9),
.B1(n_61),
.B2(n_126),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_126),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_8),
.A2(n_26),
.B1(n_33),
.B2(n_126),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_9),
.A2(n_14),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_9),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_9),
.A2(n_13),
.B1(n_36),
.B2(n_61),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_9),
.A2(n_11),
.B1(n_56),
.B2(n_61),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_11),
.A2(n_26),
.B1(n_33),
.B2(n_56),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_56),
.Y(n_113)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_12),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_13),
.A2(n_26),
.B1(n_33),
.B2(n_36),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_13),
.A2(n_36),
.B1(n_46),
.B2(n_47),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_14),
.A2(n_46),
.B(n_59),
.C(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_14),
.B(n_46),
.Y(n_59)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_15),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_92),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_90),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_76),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_19),
.B(n_76),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_68),
.C(n_71),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_20),
.A2(n_21),
.B1(n_68),
.B2(n_318),
.Y(n_324)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_38),
.B1(n_39),
.B2(n_67),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_22),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_23),
.A2(n_37),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_23),
.A2(n_37),
.B1(n_142),
.B2(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_23),
.A2(n_264),
.B(n_283),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_23),
.A2(n_82),
.B(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_24),
.B(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_24),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_24),
.A2(n_29),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_25),
.B(n_31),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g128 ( 
.A(n_26),
.B(n_129),
.CON(n_128),
.SN(n_128)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_28),
.A2(n_30),
.B1(n_128),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_29),
.B(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_29),
.B(n_284),
.Y(n_283)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

AOI32xp33_ASAP7_75t_L g215 ( 
.A1(n_30),
.A2(n_45),
.A3(n_46),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_31),
.A2(n_43),
.B(n_44),
.C(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_44),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_32),
.A2(n_37),
.B(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_35),
.Y(n_80)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_57),
.B1(n_65),
.B2(n_66),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_50),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_42),
.A2(n_51),
.B(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_43),
.A2(n_52),
.B1(n_123),
.B2(n_125),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_43),
.A2(n_52),
.B1(n_162),
.B2(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_43),
.A2(n_50),
.B(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_43),
.A2(n_52),
.B1(n_74),
.B2(n_280),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g217 ( 
.A(n_44),
.B(n_47),
.Y(n_217)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_47),
.A2(n_62),
.B(n_129),
.C(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_73),
.B(n_75),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_51),
.A2(n_85),
.B(n_86),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_51),
.A2(n_85),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_51),
.A2(n_75),
.B(n_86),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_66),
.C(n_67),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_57),
.A2(n_65),
.B1(n_72),
.B2(n_321),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_60),
.B(n_63),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_58),
.A2(n_63),
.B(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_58),
.A2(n_60),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_58),
.A2(n_60),
.B1(n_184),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_58),
.A2(n_60),
.B1(n_204),
.B2(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_58),
.A2(n_223),
.B(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_58),
.A2(n_60),
.B1(n_111),
.B2(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_58),
.A2(n_119),
.B(n_256),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_60),
.A2(n_111),
.B(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_60),
.B(n_129),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_61),
.B(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_64),
.B(n_120),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_68),
.C(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_68),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_68),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_71),
.B(n_324),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_72),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_77),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_84),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI321xp33_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_315),
.A3(n_325),
.B1(n_328),
.B2(n_329),
.C(n_332),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_295),
.B(n_314),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_271),
.B(n_294),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_164),
.B(n_247),
.C(n_270),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_147),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_97),
.B(n_147),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_132),
.B2(n_146),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_116),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_100),
.B(n_116),
.C(n_146),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_110),
.B2(n_115),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_101),
.B(n_115),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_105),
.B(n_106),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_103),
.A2(n_105),
.B1(n_108),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_103),
.A2(n_156),
.B1(n_173),
.B2(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_103),
.A2(n_176),
.B(n_206),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_103),
.A2(n_156),
.B(n_290),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_104),
.B(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_104),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_104),
.A2(n_107),
.B(n_208),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_108),
.B(n_129),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_109),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_110),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_112),
.B(n_238),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_113),
.B(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_127),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_123),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_127),
.B(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_130),
.Y(n_141)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_133),
.B(n_139),
.C(n_144),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_136),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_137),
.A2(n_156),
.B(n_157),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_143),
.B2(n_144),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.C(n_152),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_148),
.B(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_159),
.C(n_160),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_154),
.A2(n_155),
.B1(n_159),
.B2(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_157),
.B(n_206),
.Y(n_254)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_159),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_160),
.B(n_233),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_246),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_241),
.B(n_245),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_228),
.B(n_240),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_210),
.B(n_227),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_196),
.B(n_209),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_185),
.B(n_195),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_177),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_179),
.B(n_181),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_190),
.B(n_194),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_188),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_197),
.B(n_198),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_205),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_203),
.C(n_205),
.Y(n_211)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_208),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_212),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_218),
.B1(n_225),
.B2(n_226),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_213),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_215),
.Y(n_239)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_218),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_221),
.B1(n_222),
.B2(n_224),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_219),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_224),
.C(n_225),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_229),
.B(n_230),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_235),
.B2(n_236),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_237),
.C(n_239),
.Y(n_242)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2x2_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_242),
.B(n_243),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_248),
.B(n_249),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_268),
.B2(n_269),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_257),
.B2(n_258),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_258),
.C(n_269),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_255),
.Y(n_277)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_267),
.Y(n_258)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_266),
.C(n_267),
.Y(n_293)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_268),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_272),
.B(n_273),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_293),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_286),
.B2(n_287),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_287),
.C(n_293),
.Y(n_296)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_281),
.C(n_285),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_281),
.B1(n_282),
.B2(n_285),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_279),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_284),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_288),
.A2(n_289),
.B1(n_309),
.B2(n_311),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_288),
.A2(n_305),
.B(n_309),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_291),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_291),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_296),
.B(n_297),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_312),
.B2(n_313),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_304),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_304),
.C(n_313),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B(n_303),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_302),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_317),
.C(n_322),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_303),
.B(n_317),
.CI(n_322),
.CON(n_327),
.SN(n_327)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_309),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_312),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_323),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_323),
.Y(n_329)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_326),
.B(n_327),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_327),
.Y(n_331)
);


endmodule