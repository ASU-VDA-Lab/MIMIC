module fake_jpeg_24434_n_28 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_28);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_28;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_26;
wire n_17;
wire n_25;
wire n_12;
wire n_15;

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

O2A1O1Ixp33_ASAP7_75t_SL g16 ( 
.A1(n_15),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_16),
.A2(n_17),
.B(n_18),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_21),
.B(n_22),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_11),
.B(n_4),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_3),
.Y(n_26)
);

OAI21x1_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_25),
.B(n_8),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_23),
.C(n_10),
.Y(n_28)
);


endmodule