module fake_netlist_6_4717_n_1974 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1974);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1974;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_92),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_101),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_146),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_73),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_132),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_2),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_137),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_23),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_40),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_12),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_43),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_56),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_176),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_63),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_9),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_62),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_102),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_160),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_93),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_138),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_38),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_55),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_25),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_63),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_163),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_57),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_84),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_41),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_53),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_152),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_40),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_70),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_185),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_100),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_107),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_8),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_140),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_23),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_113),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_51),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_32),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_85),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_38),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_10),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_47),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_18),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_42),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_72),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_5),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_168),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_166),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_90),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_5),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_36),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_11),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_162),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_78),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_151),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_6),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_12),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_161),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_17),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_139),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_115),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_118),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_52),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_30),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_51),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_42),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_175),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_10),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_29),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_31),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_28),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_171),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_69),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_44),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_69),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_94),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_89),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_135),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_33),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_41),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_164),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_157),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_20),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_18),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_2),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_31),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_9),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_75),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_99),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_32),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_26),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_123),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_15),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_36),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_116),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_104),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_179),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_33),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_67),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_59),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_130),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_0),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_6),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_77),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_61),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_24),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_110),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_3),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_1),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_180),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_27),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_169),
.Y(n_312)
);

BUFx10_ASAP7_75t_L g313 ( 
.A(n_142),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_43),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_88),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_167),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_55),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_25),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_17),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_172),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_136),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_122),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_96),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_143),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_49),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_74),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_39),
.Y(n_327)
);

BUFx10_ASAP7_75t_L g328 ( 
.A(n_46),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_28),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_57),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_183),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_45),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_8),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_21),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_82),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_37),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_124),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_24),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_109),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_11),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_103),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_150),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_35),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_64),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_66),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_16),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_27),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_29),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_121),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_67),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_1),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_61),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_34),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_76),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_4),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_173),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_13),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_125),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_106),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_21),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_87),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_97),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_13),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_81),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_79),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_66),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_112),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_0),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_165),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_62),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_129),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_188),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_134),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_39),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_189),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_154),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_174),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_133),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_156),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_178),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_251),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_210),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_299),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_299),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_235),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_193),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_202),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_282),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_204),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_208),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_234),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_209),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_219),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_235),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_222),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_193),
.Y(n_396)
);

BUFx10_ASAP7_75t_L g397 ( 
.A(n_303),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_192),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_237),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_254),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_240),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_241),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_248),
.B(n_3),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_320),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_192),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_372),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_373),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_380),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_196),
.Y(n_409)
);

BUFx6f_ASAP7_75t_SL g410 ( 
.A(n_301),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_250),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_248),
.B(n_4),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_196),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_256),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_265),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_227),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_268),
.Y(n_417)
);

INVxp33_ASAP7_75t_SL g418 ( 
.A(n_346),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_226),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_198),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_226),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_191),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_346),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_198),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_228),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_228),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_229),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_251),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_199),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_229),
.Y(n_430)
);

BUFx2_ASAP7_75t_SL g431 ( 
.A(n_207),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_230),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_199),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_230),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_269),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_231),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_205),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_194),
.Y(n_438)
);

BUFx2_ASAP7_75t_SL g439 ( 
.A(n_207),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_203),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_R g441 ( 
.A(n_195),
.B(n_71),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_231),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_255),
.Y(n_443)
);

BUFx6f_ASAP7_75t_SL g444 ( 
.A(n_301),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_255),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g446 ( 
.A(n_203),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_289),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_289),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_282),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_197),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_296),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_296),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_270),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_307),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_273),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_200),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_275),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_206),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_251),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_216),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_279),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_283),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_367),
.B(n_7),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_251),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_286),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_290),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_307),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_312),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_312),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_315),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_315),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_335),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_227),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_251),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_291),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_381),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_464),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_350),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_459),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_381),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_428),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_398),
.B(n_367),
.Y(n_483)
);

NAND2x1p5_ASAP7_75t_L g484 ( 
.A(n_412),
.B(n_367),
.Y(n_484)
);

BUFx8_ASAP7_75t_L g485 ( 
.A(n_410),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_388),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_405),
.B(n_302),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_459),
.B(n_350),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_388),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_416),
.B(n_302),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_428),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_474),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_384),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_474),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_464),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_388),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_461),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_388),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_449),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_449),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_449),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_418),
.A2(n_217),
.B1(n_214),
.B2(n_266),
.Y(n_502)
);

INVx6_ASAP7_75t_L g503 ( 
.A(n_449),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_449),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_386),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_396),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_409),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_413),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_420),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_424),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_425),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_426),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_427),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_430),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_432),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_434),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_436),
.B(n_350),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_442),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_443),
.B(n_350),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_445),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_447),
.B(n_448),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_451),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_422),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_473),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_452),
.B(n_233),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_454),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_403),
.B(n_277),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_467),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_468),
.B(n_350),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_469),
.B(n_379),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_470),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_471),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_472),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_473),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_431),
.B(n_211),
.Y(n_535)
);

AND3x2_ASAP7_75t_L g536 ( 
.A(n_385),
.B(n_253),
.C(n_233),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_463),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_418),
.A2(n_298),
.B1(n_370),
.B2(n_244),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_429),
.B(n_253),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_431),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_433),
.B(n_278),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_439),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_397),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_397),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_387),
.B(n_297),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_397),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_439),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_440),
.B(n_460),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_446),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_462),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_465),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_441),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_394),
.B(n_378),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_423),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_480),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_527),
.B(n_387),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_537),
.B(n_483),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_502),
.B(n_382),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_537),
.A2(n_242),
.B1(n_215),
.B2(n_263),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_478),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_524),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_549),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_480),
.Y(n_563)
);

BUFx6f_ASAP7_75t_SL g564 ( 
.A(n_543),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_523),
.Y(n_565)
);

BUFx8_ASAP7_75t_SL g566 ( 
.A(n_543),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_549),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_552),
.B(n_389),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_478),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_479),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_478),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_552),
.B(n_540),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_540),
.B(n_542),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_483),
.B(n_278),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_484),
.A2(n_450),
.B1(n_456),
.B2(n_438),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_495),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_484),
.B(n_389),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_495),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_543),
.B(n_437),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_538),
.A2(n_264),
.B1(n_306),
.B2(n_201),
.Y(n_580)
);

INVx5_ASAP7_75t_L g581 ( 
.A(n_477),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_484),
.A2(n_215),
.B1(n_242),
.B2(n_263),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_524),
.Y(n_583)
);

BUFx10_ASAP7_75t_L g584 ( 
.A(n_543),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_477),
.Y(n_585)
);

AO21x2_ASAP7_75t_L g586 ( 
.A1(n_535),
.A2(n_339),
.B(n_335),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_508),
.Y(n_587)
);

NAND3xp33_ASAP7_75t_L g588 ( 
.A(n_490),
.B(n_487),
.C(n_483),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_476),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_479),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_488),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_524),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_484),
.B(n_390),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_490),
.A2(n_284),
.B1(n_311),
.B2(n_271),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_534),
.B(n_339),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_490),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_488),
.Y(n_597)
);

NAND3xp33_ASAP7_75t_L g598 ( 
.A(n_487),
.B(n_359),
.C(n_349),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_476),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_481),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_551),
.A2(n_458),
.B1(n_384),
.B2(n_392),
.Y(n_601)
);

NOR3xp33_ASAP7_75t_L g602 ( 
.A(n_502),
.B(n_383),
.C(n_390),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_534),
.Y(n_603)
);

INVx5_ASAP7_75t_L g604 ( 
.A(n_477),
.Y(n_604)
);

BUFx6f_ASAP7_75t_SL g605 ( 
.A(n_543),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_543),
.B(n_544),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_542),
.B(n_392),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_534),
.B(n_349),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_506),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_525),
.A2(n_284),
.B1(n_311),
.B2(n_271),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_481),
.Y(n_611)
);

AND2x2_ASAP7_75t_SL g612 ( 
.A(n_545),
.B(n_304),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_547),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_482),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_506),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_482),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_507),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_535),
.B(n_393),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_547),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_477),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_507),
.Y(n_621)
);

OR2x6_ASAP7_75t_L g622 ( 
.A(n_551),
.B(n_359),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_554),
.B(n_393),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_525),
.B(n_362),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_509),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_508),
.Y(n_626)
);

INVx4_ASAP7_75t_SL g627 ( 
.A(n_503),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_551),
.B(n_544),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_544),
.B(n_395),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_491),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_491),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_508),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_492),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_509),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_544),
.B(n_395),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_492),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_494),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_485),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_525),
.A2(n_347),
.B1(n_302),
.B2(n_280),
.Y(n_639)
);

BUFx10_ASAP7_75t_L g640 ( 
.A(n_544),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_525),
.A2(n_541),
.B1(n_539),
.B2(n_554),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_554),
.Y(n_642)
);

INVx6_ASAP7_75t_L g643 ( 
.A(n_486),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_510),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_494),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_510),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_550),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_512),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_539),
.A2(n_347),
.B1(n_280),
.B2(n_353),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_512),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_498),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_477),
.Y(n_652)
);

INVx5_ASAP7_75t_L g653 ( 
.A(n_477),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_530),
.B(n_399),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_493),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_553),
.B(n_399),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_489),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_539),
.B(n_401),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_493),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_498),
.Y(n_660)
);

BUFx10_ASAP7_75t_L g661 ( 
.A(n_544),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_530),
.B(n_401),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_553),
.B(n_402),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_516),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_489),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_539),
.A2(n_353),
.B1(n_252),
.B2(n_232),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_498),
.Y(n_667)
);

INVxp67_ASAP7_75t_SL g668 ( 
.A(n_489),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_516),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_501),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_546),
.B(n_362),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_501),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_526),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_501),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_546),
.B(n_497),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_508),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_541),
.A2(n_246),
.B1(n_243),
.B2(n_252),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_526),
.Y(n_678)
);

AND2x6_ASAP7_75t_L g679 ( 
.A(n_541),
.B(n_304),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_508),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_497),
.B(n_402),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_504),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_533),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_SL g684 ( 
.A1(n_546),
.A2(n_421),
.B1(n_419),
.B2(n_410),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_504),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_508),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_511),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_496),
.B(n_411),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_504),
.Y(n_689)
);

XOR2x2_ASAP7_75t_L g690 ( 
.A(n_538),
.B(n_7),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_505),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_496),
.B(n_411),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_505),
.Y(n_693)
);

OR2x6_ASAP7_75t_L g694 ( 
.A(n_546),
.B(n_371),
.Y(n_694)
);

INVx1_ASAP7_75t_SL g695 ( 
.A(n_546),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_550),
.B(n_414),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_533),
.B(n_414),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_541),
.A2(n_505),
.B1(n_532),
.B2(n_531),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_546),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_499),
.B(n_415),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_513),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_511),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_513),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_511),
.Y(n_704)
);

INVx5_ASAP7_75t_L g705 ( 
.A(n_489),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_499),
.B(n_415),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_513),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_561),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_612),
.B(n_511),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_612),
.B(n_282),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_556),
.B(n_417),
.Y(n_711)
);

BUFx5_ASAP7_75t_L g712 ( 
.A(n_574),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_609),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_612),
.B(n_511),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_572),
.B(n_619),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_596),
.B(n_511),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_658),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_668),
.A2(n_486),
.B(n_521),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_596),
.B(n_515),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_588),
.A2(n_391),
.B1(n_400),
.B2(n_404),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_609),
.Y(n_721)
);

NAND2x1p5_ASAP7_75t_L g722 ( 
.A(n_695),
.B(n_371),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_588),
.B(n_282),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_642),
.B(n_548),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_570),
.B(n_515),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_656),
.B(n_485),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_561),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_570),
.B(n_515),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_590),
.B(n_515),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_577),
.B(n_282),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_603),
.Y(n_731)
);

NAND3xp33_ASAP7_75t_L g732 ( 
.A(n_697),
.B(n_435),
.C(n_417),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_590),
.B(n_515),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_591),
.B(n_515),
.Y(n_734)
);

A2O1A1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_573),
.A2(n_375),
.B(n_376),
.C(n_548),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_615),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_591),
.B(n_522),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_597),
.B(n_522),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_593),
.B(n_323),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_615),
.Y(n_740)
);

AND2x4_ASAP7_75t_SL g741 ( 
.A(n_584),
.B(n_406),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_589),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_597),
.B(n_522),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_589),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_555),
.B(n_522),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_642),
.B(n_435),
.Y(n_746)
);

AND2x4_ASAP7_75t_SL g747 ( 
.A(n_584),
.B(n_407),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_555),
.B(n_563),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_619),
.B(n_453),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_563),
.B(n_522),
.Y(n_750)
);

O2A1O1Ixp5_ASAP7_75t_L g751 ( 
.A1(n_617),
.A2(n_519),
.B(n_517),
.C(n_529),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_613),
.B(n_557),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_557),
.A2(n_285),
.B1(n_238),
.B2(n_224),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_613),
.B(n_522),
.Y(n_754)
);

O2A1O1Ixp5_ASAP7_75t_L g755 ( 
.A1(n_617),
.A2(n_519),
.B(n_517),
.C(n_529),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_621),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_621),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_663),
.B(n_453),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_599),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_623),
.B(n_455),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_658),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_599),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_623),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_696),
.B(n_457),
.C(n_455),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_600),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_562),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_600),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_565),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_625),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_592),
.B(n_536),
.Y(n_770)
);

INVxp67_ASAP7_75t_L g771 ( 
.A(n_681),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_603),
.B(n_457),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_586),
.A2(n_274),
.B1(n_224),
.B2(n_232),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_592),
.B(n_536),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_679),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_562),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_582),
.B(n_654),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_611),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_659),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_662),
.B(n_466),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_611),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_679),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_625),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_607),
.B(n_485),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_634),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_647),
.Y(n_786)
);

NAND2xp33_ASAP7_75t_L g787 ( 
.A(n_574),
.B(n_679),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_607),
.B(n_485),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_634),
.B(n_466),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_567),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_568),
.B(n_475),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_644),
.B(n_475),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_647),
.B(n_408),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_644),
.B(n_514),
.Y(n_794)
);

INVxp67_ASAP7_75t_L g795 ( 
.A(n_567),
.Y(n_795)
);

NOR2x1p5_ASAP7_75t_L g796 ( 
.A(n_638),
.B(n_293),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_584),
.B(n_323),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_646),
.B(n_514),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_618),
.B(n_410),
.Y(n_799)
);

OR2x6_ASAP7_75t_L g800 ( 
.A(n_628),
.B(n_216),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_565),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_614),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_583),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_640),
.B(n_212),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_601),
.B(n_521),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_614),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_646),
.B(n_514),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_648),
.B(n_518),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_586),
.A2(n_363),
.B1(n_221),
.B2(n_238),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_616),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_648),
.B(n_518),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_675),
.B(n_444),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_574),
.A2(n_500),
.B(n_310),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_616),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_650),
.B(n_518),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_650),
.Y(n_816)
);

NOR2xp67_ASAP7_75t_L g817 ( 
.A(n_575),
.B(n_638),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_664),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_566),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_664),
.B(n_669),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_669),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_630),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_630),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_SL g824 ( 
.A(n_564),
.B(n_444),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_673),
.B(n_520),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_673),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_631),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_640),
.B(n_213),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_640),
.B(n_323),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_661),
.B(n_218),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_678),
.B(n_520),
.Y(n_831)
);

NOR3xp33_ASAP7_75t_L g832 ( 
.A(n_602),
.B(n_305),
.C(n_300),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_558),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_655),
.Y(n_834)
);

NAND2x1p5_ASAP7_75t_L g835 ( 
.A(n_699),
.B(n_375),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_661),
.B(n_323),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_661),
.B(n_323),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_641),
.B(n_699),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_631),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_678),
.B(n_520),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_633),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_683),
.B(n_528),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_583),
.B(n_444),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_683),
.B(n_698),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_564),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_624),
.B(n_691),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_688),
.B(n_308),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_628),
.B(n_528),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_628),
.A2(n_376),
.B1(n_236),
.B2(n_225),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_574),
.B(n_586),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_574),
.B(n_528),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_624),
.B(n_342),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_558),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_692),
.B(n_309),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_579),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_633),
.Y(n_856)
);

INVx8_ASAP7_75t_L g857 ( 
.A(n_564),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_574),
.B(n_531),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_574),
.B(n_531),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_624),
.B(n_532),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_595),
.Y(n_861)
);

OAI221xp5_ASAP7_75t_L g862 ( 
.A1(n_594),
.A2(n_221),
.B1(n_243),
.B2(n_246),
.C(n_363),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_595),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_700),
.Y(n_864)
);

BUFx5_ASAP7_75t_L g865 ( 
.A(n_679),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_706),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_595),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_624),
.B(n_532),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_595),
.B(n_486),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_598),
.A2(n_259),
.B1(n_257),
.B2(n_285),
.Y(n_870)
);

INVx8_ASAP7_75t_L g871 ( 
.A(n_605),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_608),
.B(n_486),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_636),
.Y(n_873)
);

INVx4_ASAP7_75t_L g874 ( 
.A(n_605),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_608),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_629),
.B(n_314),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_608),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_608),
.B(n_257),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_636),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_715),
.B(n_606),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_715),
.B(n_628),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_866),
.B(n_684),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_803),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_771),
.B(n_635),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_710),
.A2(n_622),
.B(n_598),
.C(n_637),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_777),
.A2(n_580),
.B(n_637),
.C(n_645),
.Y(n_886)
);

NAND2x1_ASAP7_75t_L g887 ( 
.A(n_731),
.B(n_643),
.Y(n_887)
);

O2A1O1Ixp5_ASAP7_75t_L g888 ( 
.A1(n_710),
.A2(n_645),
.B(n_704),
.C(n_702),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_724),
.B(n_628),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_834),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_863),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_742),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_742),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_744),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_708),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_838),
.A2(n_626),
.B(n_587),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_709),
.A2(n_605),
.B1(n_694),
.B2(n_671),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_708),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_749),
.B(n_580),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_708),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_714),
.A2(n_626),
.B(n_587),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_723),
.A2(n_704),
.B(n_702),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_708),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_861),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_752),
.B(n_622),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_844),
.A2(n_626),
.B(n_587),
.Y(n_906)
);

O2A1O1Ixp5_ASAP7_75t_L g907 ( 
.A1(n_730),
.A2(n_651),
.B(n_660),
.C(n_667),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_844),
.A2(n_676),
.B(n_632),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_803),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_850),
.A2(n_694),
.B1(n_671),
.B2(n_622),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_760),
.B(n_622),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_748),
.B(n_622),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_867),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_711),
.B(n_671),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_875),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_768),
.Y(n_916)
);

O2A1O1Ixp5_ASAP7_75t_L g917 ( 
.A1(n_730),
.A2(n_651),
.B(n_660),
.C(n_667),
.Y(n_917)
);

AND3x2_ASAP7_75t_L g918 ( 
.A(n_824),
.B(n_274),
.C(n_259),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_863),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_864),
.B(n_666),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_766),
.B(n_677),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_723),
.A2(n_679),
.B(n_691),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_787),
.A2(n_676),
.B(n_632),
.Y(n_923)
);

NAND2x1p5_ASAP7_75t_L g924 ( 
.A(n_775),
.B(n_680),
.Y(n_924)
);

O2A1O1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_735),
.A2(n_671),
.B(n_694),
.C(n_701),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_869),
.A2(n_676),
.B(n_632),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_749),
.B(n_559),
.Y(n_927)
);

NAND3xp33_ASAP7_75t_L g928 ( 
.A(n_711),
.B(n_649),
.C(n_639),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_758),
.B(n_671),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_876),
.A2(n_707),
.B(n_703),
.C(n_701),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_780),
.B(n_694),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_847),
.B(n_694),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_790),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_872),
.A2(n_687),
.B(n_686),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_846),
.A2(n_687),
.B(n_686),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_846),
.A2(n_687),
.B(n_686),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_725),
.A2(n_680),
.B(n_652),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_847),
.B(n_854),
.Y(n_938)
);

AOI21x1_ASAP7_75t_L g939 ( 
.A1(n_739),
.A2(n_672),
.B(n_670),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_728),
.A2(n_652),
.B(n_585),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_763),
.B(n_690),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_791),
.B(n_643),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_854),
.B(n_713),
.Y(n_943)
);

O2A1O1Ixp5_ASAP7_75t_L g944 ( 
.A1(n_739),
.A2(n_829),
.B(n_836),
.C(n_797),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_716),
.A2(n_719),
.B(n_851),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_877),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_858),
.A2(n_703),
.B(n_693),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_859),
.A2(n_707),
.B(n_693),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_801),
.Y(n_949)
);

CKINVDCx10_ASAP7_75t_R g950 ( 
.A(n_833),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_717),
.A2(n_610),
.B1(n_643),
.B2(n_685),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_729),
.A2(n_672),
.B(n_670),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_759),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_761),
.A2(n_643),
.B1(n_689),
.B2(n_685),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_876),
.A2(n_576),
.B(n_578),
.C(n_689),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_795),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_721),
.B(n_679),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_791),
.A2(n_578),
.B(n_576),
.C(n_682),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_733),
.A2(n_679),
.B(n_674),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_727),
.B(n_786),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_779),
.B(n_317),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_762),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_805),
.A2(n_682),
.B(n_674),
.C(n_657),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_736),
.B(n_620),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_734),
.A2(n_569),
.B(n_560),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_764),
.B(n_319),
.Y(n_966)
);

CKINVDCx8_ASAP7_75t_R g967 ( 
.A(n_819),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_732),
.B(n_325),
.Y(n_968)
);

AO21x1_ASAP7_75t_L g969 ( 
.A1(n_722),
.A2(n_294),
.B(n_287),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_799),
.A2(n_620),
.B(n_657),
.C(n_560),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_855),
.A2(n_267),
.B1(n_261),
.B2(n_260),
.Y(n_971)
);

OAI321xp33_ASAP7_75t_L g972 ( 
.A1(n_870),
.A2(n_287),
.A3(n_294),
.B1(n_348),
.B2(n_351),
.C(n_318),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_848),
.A2(n_799),
.B1(n_772),
.B2(n_792),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_740),
.B(n_620),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_812),
.A2(n_657),
.B(n_569),
.C(n_571),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_727),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_746),
.B(n_690),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_756),
.B(n_571),
.Y(n_978)
);

NOR3xp33_ASAP7_75t_L g979 ( 
.A(n_853),
.B(n_333),
.C(n_344),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_737),
.A2(n_743),
.B(n_738),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_720),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_860),
.A2(n_665),
.B(n_585),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_868),
.A2(n_500),
.B(n_653),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_776),
.B(n_627),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_754),
.A2(n_665),
.B(n_585),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_757),
.B(n_585),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_741),
.B(n_205),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_769),
.B(n_585),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_765),
.Y(n_989)
);

NAND2xp33_ASAP7_75t_L g990 ( 
.A(n_712),
.B(n_652),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_765),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_789),
.B(n_327),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_783),
.B(n_652),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_741),
.B(n_205),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_731),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_857),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_745),
.A2(n_665),
.B(n_652),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_767),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_750),
.A2(n_665),
.B(n_489),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_820),
.A2(n_665),
.B(n_489),
.Y(n_1000)
);

NAND3xp33_ASAP7_75t_L g1001 ( 
.A(n_832),
.B(n_336),
.C(n_329),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_785),
.B(n_220),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_718),
.A2(n_705),
.B(n_653),
.Y(n_1003)
);

BUFx12f_ASAP7_75t_L g1004 ( 
.A(n_796),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_767),
.Y(n_1005)
);

BUFx4f_ASAP7_75t_L g1006 ( 
.A(n_747),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_816),
.B(n_223),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_773),
.A2(n_337),
.B1(n_331),
.B2(n_239),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_778),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_793),
.B(n_747),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_818),
.B(n_245),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_794),
.A2(n_705),
.B(n_653),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_821),
.B(n_247),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_798),
.A2(n_705),
.B(n_653),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_807),
.A2(n_705),
.B(n_653),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_826),
.B(n_249),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_770),
.B(n_330),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_843),
.B(n_205),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_778),
.B(n_258),
.Y(n_1019)
);

AO21x1_ASAP7_75t_L g1020 ( 
.A1(n_722),
.A2(n_318),
.B(n_348),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_812),
.A2(n_262),
.B1(n_272),
.B2(n_341),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_808),
.A2(n_705),
.B(n_653),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_781),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_857),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_811),
.A2(n_705),
.B(n_581),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_815),
.A2(n_581),
.B(n_604),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_825),
.A2(n_581),
.B(n_604),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_751),
.A2(n_351),
.B(n_321),
.C(n_316),
.Y(n_1028)
);

NAND3xp33_ASAP7_75t_L g1029 ( 
.A(n_753),
.B(n_374),
.C(n_368),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_802),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_802),
.B(n_276),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_784),
.B(n_332),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_755),
.A2(n_581),
.B(n_604),
.Y(n_1033)
);

INVx4_ASAP7_75t_L g1034 ( 
.A(n_857),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_806),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_878),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_831),
.A2(n_581),
.B(n_604),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_806),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_770),
.A2(n_774),
.B1(n_800),
.B2(n_817),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_810),
.B(n_281),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_843),
.B(n_328),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_788),
.B(n_334),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_813),
.A2(n_288),
.B(n_292),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_836),
.A2(n_342),
.B(n_322),
.Y(n_1044)
);

OAI21xp33_ASAP7_75t_L g1045 ( 
.A1(n_753),
.A2(n_360),
.B(n_357),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_840),
.A2(n_295),
.B(n_324),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_842),
.A2(n_354),
.B(n_326),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_814),
.A2(n_361),
.B(n_356),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_774),
.B(n_338),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_871),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_837),
.A2(n_364),
.B(n_377),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_837),
.A2(n_358),
.B(n_369),
.Y(n_1052)
);

AND2x6_ASAP7_75t_L g1053 ( 
.A(n_775),
.B(n_782),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_712),
.B(n_365),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_862),
.A2(n_301),
.B(n_313),
.C(n_328),
.Y(n_1055)
);

INVxp67_ASAP7_75t_L g1056 ( 
.A(n_878),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_773),
.A2(n_342),
.B1(n_355),
.B2(n_352),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_726),
.B(n_340),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_809),
.A2(n_343),
.B(n_345),
.C(n_342),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_852),
.A2(n_342),
.B(n_627),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_712),
.B(n_313),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_712),
.B(n_313),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_809),
.A2(n_301),
.B(n_313),
.C(n_328),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_852),
.A2(n_627),
.B(n_503),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_814),
.B(n_503),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_822),
.A2(n_503),
.B(n_83),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_990),
.A2(n_871),
.B(n_874),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_996),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_909),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_938),
.B(n_943),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_928),
.A2(n_870),
.B1(n_800),
.B2(n_782),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_996),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_904),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_913),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_945),
.A2(n_879),
.B(n_839),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_884),
.B(n_845),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_883),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_945),
.A2(n_871),
.B(n_874),
.Y(n_1078)
);

AND2x2_ASAP7_75t_SL g1079 ( 
.A(n_1006),
.B(n_899),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_942),
.B(n_822),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_915),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_946),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_939),
.A2(n_879),
.B(n_873),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_962),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_880),
.A2(n_800),
.B1(n_782),
.B2(n_775),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_933),
.B(n_849),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_941),
.B(n_823),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_889),
.B(n_873),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_992),
.B(n_804),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_890),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_923),
.A2(n_712),
.B(n_782),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_927),
.A2(n_823),
.B1(n_856),
.B2(n_841),
.Y(n_1092)
);

INVx5_ASAP7_75t_L g1093 ( 
.A(n_1053),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_977),
.B(n_827),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_892),
.Y(n_1095)
);

NAND3xp33_ASAP7_75t_SL g1096 ( 
.A(n_1058),
.B(n_835),
.C(n_830),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_956),
.Y(n_1097)
);

BUFx12f_ASAP7_75t_L g1098 ( 
.A(n_916),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_973),
.B(n_827),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_SL g1100 ( 
.A1(n_1059),
.A2(n_932),
.B(n_1028),
.C(n_914),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_882),
.A2(n_828),
.B(n_839),
.C(n_841),
.Y(n_1101)
);

BUFx8_ASAP7_75t_L g1102 ( 
.A(n_1004),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_893),
.Y(n_1103)
);

NOR3xp33_ASAP7_75t_SL g1104 ( 
.A(n_1010),
.B(n_328),
.C(n_366),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_881),
.A2(n_835),
.B1(n_856),
.B2(n_712),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_931),
.B(n_865),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_996),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_929),
.B(n_865),
.Y(n_1108)
);

INVx5_ASAP7_75t_L g1109 ( 
.A(n_1053),
.Y(n_1109)
);

OAI21xp33_ASAP7_75t_SL g1110 ( 
.A1(n_920),
.A2(n_865),
.B(n_366),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_960),
.Y(n_1111)
);

BUFx10_ASAP7_75t_L g1112 ( 
.A(n_1049),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_1050),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_SL g1114 ( 
.A1(n_1063),
.A2(n_865),
.B(n_86),
.C(n_91),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_901),
.A2(n_865),
.B(n_503),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_984),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_894),
.Y(n_1117)
);

O2A1O1Ixp5_ASAP7_75t_L g1118 ( 
.A1(n_1061),
.A2(n_865),
.B(n_141),
.C(n_190),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_966),
.A2(n_366),
.B(n_15),
.C(n_16),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_998),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_981),
.B(n_366),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_912),
.B(n_14),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_886),
.B(n_14),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1039),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_SL g1125 ( 
.A1(n_968),
.A2(n_186),
.B(n_184),
.C(n_159),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_901),
.A2(n_158),
.B(n_155),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_950),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_949),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_921),
.A2(n_19),
.B1(n_22),
.B2(n_26),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_995),
.B(n_149),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_910),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_SL g1132 ( 
.A1(n_1032),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_1050),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1056),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_1050),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_967),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_995),
.B(n_98),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_980),
.A2(n_95),
.B(n_147),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1005),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_911),
.B(n_48),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_905),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_980),
.A2(n_108),
.B(n_145),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_960),
.B(n_105),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_885),
.A2(n_50),
.B(n_53),
.C(n_54),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_976),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1009),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_926),
.A2(n_111),
.B(n_144),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_891),
.B(n_80),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_953),
.Y(n_1149)
);

OAI21xp33_ASAP7_75t_L g1150 ( 
.A1(n_961),
.A2(n_54),
.B(n_56),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1035),
.Y(n_1151)
);

INVx3_ASAP7_75t_SL g1152 ( 
.A(n_1017),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1018),
.B(n_58),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_934),
.A2(n_117),
.B(n_131),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_891),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_1155)
);

HB1xp67_ASAP7_75t_L g1156 ( 
.A(n_1036),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_895),
.B(n_119),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1041),
.B(n_60),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_919),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_935),
.A2(n_114),
.B(n_120),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_895),
.B(n_126),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_936),
.A2(n_127),
.B(n_148),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1038),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_919),
.A2(n_65),
.B1(n_68),
.B2(n_897),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_984),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1043),
.A2(n_1008),
.B1(n_1020),
.B2(n_969),
.Y(n_1166)
);

OAI22x1_ASAP7_75t_L g1167 ( 
.A1(n_1042),
.A2(n_994),
.B1(n_987),
.B2(n_1001),
.Y(n_1167)
);

BUFx8_ASAP7_75t_L g1168 ( 
.A(n_895),
.Y(n_1168)
);

BUFx8_ASAP7_75t_L g1169 ( 
.A(n_898),
.Y(n_1169)
);

INVx4_ASAP7_75t_L g1170 ( 
.A(n_898),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_SL g1171 ( 
.A(n_1006),
.B(n_1024),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_989),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_887),
.A2(n_959),
.B(n_906),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_991),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_906),
.A2(n_908),
.B(n_983),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_1034),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_908),
.A2(n_896),
.B(n_922),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1023),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1034),
.B(n_898),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_900),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_896),
.A2(n_957),
.B(n_1054),
.Y(n_1181)
);

AOI21x1_ASAP7_75t_L g1182 ( 
.A1(n_985),
.A2(n_997),
.B(n_982),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_982),
.A2(n_902),
.B(n_985),
.Y(n_1183)
);

AO21x1_ASAP7_75t_L g1184 ( 
.A1(n_925),
.A2(n_1066),
.B(n_1062),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_944),
.A2(n_1055),
.B(n_888),
.C(n_1007),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1002),
.A2(n_1011),
.B(n_1013),
.C(n_1016),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_997),
.A2(n_940),
.B(n_937),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1030),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1033),
.A2(n_965),
.B(n_951),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_971),
.B(n_1045),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_903),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_978),
.B(n_1053),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_903),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1053),
.B(n_958),
.Y(n_1194)
);

O2A1O1Ixp5_ASAP7_75t_L g1195 ( 
.A1(n_970),
.A2(n_975),
.B(n_963),
.C(n_955),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_964),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_974),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_986),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_988),
.B(n_993),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_947),
.A2(n_948),
.B(n_1000),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_979),
.B(n_918),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_924),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_947),
.A2(n_948),
.B(n_1000),
.Y(n_1203)
);

BUFx8_ASAP7_75t_SL g1204 ( 
.A(n_1019),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_930),
.B(n_952),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1029),
.B(n_1021),
.Y(n_1206)
);

NAND3xp33_ASAP7_75t_SL g1207 ( 
.A(n_1057),
.B(n_1046),
.C(n_1047),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1065),
.Y(n_1208)
);

INVx6_ASAP7_75t_L g1209 ( 
.A(n_924),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1031),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_907),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1040),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1048),
.B(n_1051),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_952),
.B(n_999),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1051),
.B(n_1052),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_917),
.A2(n_999),
.B(n_1003),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_954),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1046),
.B(n_1047),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1003),
.A2(n_1025),
.B(n_1012),
.Y(n_1219)
);

AOI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1012),
.A2(n_1025),
.B(n_1014),
.Y(n_1220)
);

INVx8_ASAP7_75t_L g1221 ( 
.A(n_972),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1014),
.B(n_1015),
.Y(n_1222)
);

INVxp67_ASAP7_75t_L g1223 ( 
.A(n_1052),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1095),
.Y(n_1224)
);

INVx2_ASAP7_75t_SL g1225 ( 
.A(n_1145),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1189),
.A2(n_1175),
.B(n_1173),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1106),
.A2(n_1066),
.B(n_1022),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1070),
.A2(n_1089),
.B(n_1158),
.C(n_1153),
.Y(n_1228)
);

NAND3xp33_ASAP7_75t_L g1229 ( 
.A(n_1121),
.B(n_1044),
.C(n_1060),
.Y(n_1229)
);

INVx4_ASAP7_75t_L g1230 ( 
.A(n_1072),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1070),
.A2(n_1015),
.B(n_1022),
.C(n_1026),
.Y(n_1231)
);

O2A1O1Ixp5_ASAP7_75t_SL g1232 ( 
.A1(n_1131),
.A2(n_1026),
.B(n_1027),
.C(n_1037),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1108),
.A2(n_1027),
.B(n_1037),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1094),
.B(n_1064),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1076),
.B(n_1064),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1103),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_SL g1237 ( 
.A(n_1093),
.B(n_1109),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1115),
.A2(n_1182),
.B(n_1220),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1219),
.A2(n_1203),
.B(n_1200),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_SL g1240 ( 
.A(n_1093),
.B(n_1109),
.Y(n_1240)
);

NOR4xp25_ASAP7_75t_L g1241 ( 
.A(n_1150),
.B(n_1131),
.C(n_1124),
.D(n_1129),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1184),
.A2(n_1105),
.A3(n_1183),
.B(n_1222),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1187),
.A2(n_1075),
.B(n_1177),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1119),
.A2(n_1129),
.B(n_1124),
.C(n_1144),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1091),
.A2(n_1080),
.B(n_1186),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1195),
.A2(n_1185),
.B(n_1075),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1068),
.B(n_1135),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1073),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1079),
.B(n_1087),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1074),
.Y(n_1250)
);

O2A1O1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1164),
.A2(n_1141),
.B(n_1190),
.C(n_1134),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1081),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1080),
.A2(n_1100),
.B(n_1181),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1071),
.A2(n_1166),
.B(n_1223),
.Y(n_1254)
);

OA21x2_ASAP7_75t_L g1255 ( 
.A1(n_1216),
.A2(n_1222),
.B(n_1214),
.Y(n_1255)
);

O2A1O1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1164),
.A2(n_1141),
.B(n_1134),
.C(n_1123),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1214),
.A2(n_1205),
.B(n_1218),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1210),
.B(n_1212),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1097),
.B(n_1086),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1105),
.A2(n_1205),
.A3(n_1218),
.B(n_1085),
.Y(n_1260)
);

AO31x2_ASAP7_75t_L g1261 ( 
.A1(n_1085),
.A2(n_1194),
.A3(n_1211),
.B(n_1071),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1082),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1078),
.A2(n_1199),
.B(n_1213),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1199),
.A2(n_1099),
.B(n_1216),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1128),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1069),
.B(n_1112),
.Y(n_1266)
);

AO21x2_ASAP7_75t_L g1267 ( 
.A1(n_1207),
.A2(n_1096),
.B(n_1194),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1084),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1168),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1140),
.A2(n_1122),
.B(n_1159),
.C(n_1155),
.Y(n_1270)
);

NAND3xp33_ASAP7_75t_SL g1271 ( 
.A(n_1104),
.B(n_1206),
.C(n_1136),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1196),
.B(n_1198),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1132),
.A2(n_1221),
.B1(n_1201),
.B2(n_1167),
.Y(n_1273)
);

BUFx4f_ASAP7_75t_L g1274 ( 
.A(n_1098),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1197),
.B(n_1221),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1117),
.Y(n_1276)
);

AOI221x1_ASAP7_75t_L g1277 ( 
.A1(n_1138),
.A2(n_1142),
.B1(n_1126),
.B2(n_1154),
.C(n_1147),
.Y(n_1277)
);

OAI21xp33_ASAP7_75t_L g1278 ( 
.A1(n_1171),
.A2(n_1155),
.B(n_1159),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1120),
.Y(n_1279)
);

CKINVDCx8_ASAP7_75t_R g1280 ( 
.A(n_1127),
.Y(n_1280)
);

O2A1O1Ixp33_ASAP7_75t_SL g1281 ( 
.A1(n_1130),
.A2(n_1137),
.B(n_1148),
.C(n_1125),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1093),
.A2(n_1109),
.B(n_1067),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1093),
.A2(n_1109),
.B(n_1192),
.Y(n_1283)
);

AOI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1215),
.A2(n_1217),
.B(n_1148),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1130),
.A2(n_1137),
.B(n_1162),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1101),
.A2(n_1110),
.B(n_1221),
.C(n_1118),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_1090),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1209),
.A2(n_1092),
.B1(n_1116),
.B2(n_1165),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1192),
.A2(n_1160),
.A3(n_1208),
.B(n_1088),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1088),
.A2(n_1151),
.A3(n_1163),
.B(n_1146),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1111),
.B(n_1139),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1116),
.B(n_1165),
.Y(n_1292)
);

INVx4_ASAP7_75t_L g1293 ( 
.A(n_1072),
.Y(n_1293)
);

NOR2xp67_ASAP7_75t_SL g1294 ( 
.A(n_1176),
.B(n_1072),
.Y(n_1294)
);

AOI31xp67_ASAP7_75t_L g1295 ( 
.A1(n_1157),
.A2(n_1161),
.A3(n_1178),
.B(n_1174),
.Y(n_1295)
);

OAI221xp5_ASAP7_75t_L g1296 ( 
.A1(n_1152),
.A2(n_1156),
.B1(n_1143),
.B2(n_1114),
.C(n_1172),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_1193),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1204),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1201),
.A2(n_1149),
.B(n_1188),
.C(n_1180),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1209),
.Y(n_1300)
);

AO32x2_ASAP7_75t_L g1301 ( 
.A1(n_1170),
.A2(n_1112),
.A3(n_1169),
.B1(n_1168),
.B2(n_1209),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1179),
.B(n_1107),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1202),
.A2(n_1170),
.B(n_1169),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1179),
.A2(n_1191),
.B(n_1107),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1191),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1191),
.B(n_1107),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1113),
.A2(n_1133),
.B(n_1102),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_1113),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_SL g1309 ( 
.A1(n_1113),
.A2(n_938),
.B(n_710),
.C(n_1186),
.Y(n_1309)
);

OR2x6_ASAP7_75t_L g1310 ( 
.A(n_1102),
.B(n_996),
.Y(n_1310)
);

NAND3xp33_ASAP7_75t_L g1311 ( 
.A(n_1089),
.B(n_938),
.C(n_711),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1070),
.B(n_715),
.Y(n_1312)
);

INVxp67_ASAP7_75t_L g1313 ( 
.A(n_1077),
.Y(n_1313)
);

NOR4xp25_ASAP7_75t_L g1314 ( 
.A(n_1150),
.B(n_938),
.C(n_1131),
.D(n_1124),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1070),
.A2(n_938),
.B(n_914),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1070),
.A2(n_938),
.B1(n_1089),
.B2(n_942),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1083),
.A2(n_1115),
.B(n_1182),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1189),
.A2(n_990),
.B(n_942),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1089),
.A2(n_899),
.B1(n_938),
.B2(n_612),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1097),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1209),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1083),
.A2(n_1115),
.B(n_1182),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1136),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1070),
.B(n_715),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1095),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1070),
.A2(n_938),
.B1(n_1089),
.B2(n_942),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1145),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1073),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1189),
.A2(n_938),
.B(n_1195),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1094),
.B(n_899),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1136),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1072),
.Y(n_1332)
);

O2A1O1Ixp33_ASAP7_75t_SL g1333 ( 
.A1(n_1186),
.A2(n_938),
.B(n_710),
.C(n_1144),
.Y(n_1333)
);

INVx3_ASAP7_75t_SL g1334 ( 
.A(n_1136),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1094),
.B(n_899),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1189),
.A2(n_990),
.B(n_942),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1189),
.A2(n_990),
.B(n_942),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1070),
.B(n_720),
.Y(n_1338)
);

NOR2x1_ASAP7_75t_SL g1339 ( 
.A(n_1093),
.B(n_1109),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1070),
.B(n_715),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1070),
.B(n_715),
.Y(n_1341)
);

AO32x2_ASAP7_75t_L g1342 ( 
.A1(n_1131),
.A2(n_1164),
.A3(n_1141),
.B1(n_1129),
.B2(n_1124),
.Y(n_1342)
);

AO21x2_ASAP7_75t_L g1343 ( 
.A1(n_1189),
.A2(n_1175),
.B(n_1216),
.Y(n_1343)
);

INVx5_ASAP7_75t_L g1344 ( 
.A(n_1093),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1089),
.A2(n_938),
.B(n_1190),
.C(n_711),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1070),
.B(n_771),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1070),
.A2(n_938),
.B(n_914),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1184),
.A2(n_1189),
.A3(n_1175),
.B(n_1105),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_1136),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1073),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1070),
.B(n_715),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1136),
.Y(n_1352)
);

O2A1O1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1070),
.A2(n_938),
.B(n_771),
.C(n_758),
.Y(n_1353)
);

CKINVDCx14_ASAP7_75t_R g1354 ( 
.A(n_1127),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1189),
.A2(n_990),
.B(n_942),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1073),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1069),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1094),
.B(n_899),
.Y(n_1358)
);

AO21x2_ASAP7_75t_L g1359 ( 
.A1(n_1189),
.A2(n_1175),
.B(n_1216),
.Y(n_1359)
);

AO32x2_ASAP7_75t_L g1360 ( 
.A1(n_1131),
.A2(n_1164),
.A3(n_1141),
.B1(n_1129),
.B2(n_1124),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1089),
.A2(n_899),
.B1(n_938),
.B2(n_612),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1070),
.B(n_715),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1070),
.B(n_715),
.Y(n_1363)
);

INVxp67_ASAP7_75t_SL g1364 ( 
.A(n_1077),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1089),
.A2(n_899),
.B1(n_938),
.B2(n_612),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1070),
.A2(n_938),
.B(n_914),
.Y(n_1366)
);

AO31x2_ASAP7_75t_L g1367 ( 
.A1(n_1184),
.A2(n_1189),
.A3(n_1175),
.B(n_1105),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1070),
.B(n_715),
.Y(n_1368)
);

AOI221x1_ASAP7_75t_L g1369 ( 
.A1(n_1164),
.A2(n_938),
.B1(n_1131),
.B2(n_1144),
.C(n_1150),
.Y(n_1369)
);

AO31x2_ASAP7_75t_L g1370 ( 
.A1(n_1184),
.A2(n_1189),
.A3(n_1175),
.B(n_1105),
.Y(n_1370)
);

AO31x2_ASAP7_75t_L g1371 ( 
.A1(n_1184),
.A2(n_1189),
.A3(n_1175),
.B(n_1105),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1189),
.A2(n_1216),
.B(n_1175),
.Y(n_1372)
);

A2O1A1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1089),
.A2(n_938),
.B(n_1190),
.C(n_711),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1083),
.A2(n_1115),
.B(n_1182),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1097),
.Y(n_1375)
);

AO21x2_ASAP7_75t_L g1376 ( 
.A1(n_1189),
.A2(n_1175),
.B(n_1216),
.Y(n_1376)
);

BUFx2_ASAP7_75t_R g1377 ( 
.A(n_1127),
.Y(n_1377)
);

NAND3xp33_ASAP7_75t_L g1378 ( 
.A(n_1089),
.B(n_938),
.C(n_711),
.Y(n_1378)
);

O2A1O1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1070),
.A2(n_938),
.B(n_771),
.C(n_758),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1073),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1224),
.Y(n_1381)
);

OAI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1319),
.A2(n_1365),
.B1(n_1361),
.B2(n_1311),
.Y(n_1382)
);

INVx6_ASAP7_75t_L g1383 ( 
.A(n_1344),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1311),
.A2(n_1378),
.B1(n_1319),
.B2(n_1361),
.Y(n_1384)
);

OAI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1365),
.A2(n_1378),
.B1(n_1363),
.B2(n_1324),
.Y(n_1385)
);

BUFx4f_ASAP7_75t_SL g1386 ( 
.A(n_1331),
.Y(n_1386)
);

INVx1_ASAP7_75t_SL g1387 ( 
.A(n_1265),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1250),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_SL g1389 ( 
.A1(n_1273),
.A2(n_1259),
.B1(n_1346),
.B2(n_1314),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1320),
.Y(n_1390)
);

INVx4_ASAP7_75t_L g1391 ( 
.A(n_1344),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1236),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_1349),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1278),
.A2(n_1338),
.B1(n_1271),
.B2(n_1249),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1278),
.A2(n_1326),
.B1(n_1316),
.B2(n_1273),
.Y(n_1395)
);

INVx4_ASAP7_75t_L g1396 ( 
.A(n_1332),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1265),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1375),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1345),
.B(n_1373),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1332),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1252),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1254),
.A2(n_1335),
.B1(n_1330),
.B2(n_1358),
.Y(n_1402)
);

CKINVDCx11_ASAP7_75t_R g1403 ( 
.A(n_1280),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1258),
.B(n_1275),
.Y(n_1404)
);

BUFx12f_ASAP7_75t_L g1405 ( 
.A(n_1323),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1327),
.Y(n_1406)
);

BUFx12f_ASAP7_75t_L g1407 ( 
.A(n_1352),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1262),
.Y(n_1408)
);

BUFx12f_ASAP7_75t_L g1409 ( 
.A(n_1310),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1328),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1235),
.A2(n_1366),
.B1(n_1347),
.B2(n_1315),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1350),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1329),
.A2(n_1351),
.B1(n_1340),
.B2(n_1341),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_1354),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1329),
.A2(n_1246),
.B1(n_1362),
.B2(n_1368),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1312),
.A2(n_1267),
.B1(n_1296),
.B2(n_1234),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1357),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1276),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1287),
.A2(n_1314),
.B1(n_1266),
.B2(n_1241),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1291),
.B(n_1325),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1267),
.A2(n_1343),
.B1(n_1359),
.B2(n_1376),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1302),
.B(n_1300),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1356),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1228),
.A2(n_1272),
.B1(n_1379),
.B2(n_1353),
.Y(n_1424)
);

BUFx12f_ASAP7_75t_L g1425 ( 
.A(n_1310),
.Y(n_1425)
);

OAI22x1_ASAP7_75t_L g1426 ( 
.A1(n_1364),
.A2(n_1279),
.B1(n_1268),
.B2(n_1380),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1301),
.Y(n_1427)
);

AOI22xp5_ASAP7_75t_SL g1428 ( 
.A1(n_1298),
.A2(n_1313),
.B1(n_1269),
.B2(n_1297),
.Y(n_1428)
);

INVx2_ASAP7_75t_SL g1429 ( 
.A(n_1225),
.Y(n_1429)
);

BUFx10_ASAP7_75t_L g1430 ( 
.A(n_1310),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1334),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1343),
.A2(n_1376),
.B1(n_1359),
.B2(n_1288),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1246),
.A2(n_1241),
.B1(n_1360),
.B2(n_1342),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_SL g1434 ( 
.A1(n_1342),
.A2(n_1360),
.B1(n_1372),
.B2(n_1240),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_SL g1435 ( 
.A1(n_1244),
.A2(n_1251),
.B(n_1369),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1229),
.A2(n_1372),
.B1(n_1226),
.B2(n_1292),
.Y(n_1436)
);

OAI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1237),
.A2(n_1240),
.B1(n_1257),
.B2(n_1360),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1229),
.A2(n_1255),
.B1(n_1245),
.B2(n_1264),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1290),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_1247),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1305),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1255),
.A2(n_1321),
.B1(n_1263),
.B2(n_1355),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1295),
.Y(n_1443)
);

OAI21xp33_ASAP7_75t_L g1444 ( 
.A1(n_1270),
.A2(n_1256),
.B(n_1299),
.Y(n_1444)
);

BUFx2_ASAP7_75t_SL g1445 ( 
.A(n_1230),
.Y(n_1445)
);

INVx6_ASAP7_75t_L g1446 ( 
.A(n_1230),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_SL g1447 ( 
.A1(n_1342),
.A2(n_1237),
.B1(n_1274),
.B2(n_1318),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1261),
.B(n_1333),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1286),
.A2(n_1337),
.B1(n_1336),
.B2(n_1308),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1377),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1332),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1293),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1277),
.A2(n_1253),
.B1(n_1306),
.B2(n_1293),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1294),
.A2(n_1233),
.B1(n_1227),
.B2(n_1243),
.Y(n_1454)
);

INVx6_ASAP7_75t_L g1455 ( 
.A(n_1303),
.Y(n_1455)
);

OAI22xp33_ASAP7_75t_R g1456 ( 
.A1(n_1301),
.A2(n_1309),
.B1(n_1307),
.B2(n_1261),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1301),
.Y(n_1457)
);

NAND2x1p5_ASAP7_75t_L g1458 ( 
.A(n_1283),
.B(n_1282),
.Y(n_1458)
);

CKINVDCx11_ASAP7_75t_R g1459 ( 
.A(n_1304),
.Y(n_1459)
);

BUFx5_ASAP7_75t_L g1460 ( 
.A(n_1239),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1289),
.B(n_1260),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1260),
.B(n_1289),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1231),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1260),
.Y(n_1464)
);

INVx6_ASAP7_75t_L g1465 ( 
.A(n_1339),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1242),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_SL g1467 ( 
.A1(n_1285),
.A2(n_1348),
.B1(n_1371),
.B2(n_1367),
.Y(n_1467)
);

INVx6_ASAP7_75t_L g1468 ( 
.A(n_1232),
.Y(n_1468)
);

OAI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1284),
.A2(n_1348),
.B1(n_1371),
.B2(n_1370),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1348),
.A2(n_1371),
.B1(n_1370),
.B2(n_1367),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1367),
.A2(n_1370),
.B1(n_1242),
.B2(n_1238),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_1281),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1317),
.B(n_1322),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_SL g1474 ( 
.A1(n_1374),
.A2(n_1132),
.B1(n_899),
.B2(n_1311),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_1265),
.Y(n_1475)
);

INVx4_ASAP7_75t_L g1476 ( 
.A(n_1344),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1261),
.Y(n_1477)
);

BUFx4f_ASAP7_75t_SL g1478 ( 
.A(n_1331),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1311),
.A2(n_938),
.B1(n_1378),
.B2(n_899),
.Y(n_1479)
);

INVx3_ASAP7_75t_SL g1480 ( 
.A(n_1323),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1311),
.A2(n_938),
.B1(n_1089),
.B2(n_1378),
.Y(n_1481)
);

INVx2_ASAP7_75t_SL g1482 ( 
.A(n_1327),
.Y(n_1482)
);

BUFx2_ASAP7_75t_SL g1483 ( 
.A(n_1331),
.Y(n_1483)
);

BUFx8_ASAP7_75t_L g1484 ( 
.A(n_1269),
.Y(n_1484)
);

BUFx12f_ASAP7_75t_L g1485 ( 
.A(n_1323),
.Y(n_1485)
);

BUFx8_ASAP7_75t_SL g1486 ( 
.A(n_1331),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1248),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1319),
.A2(n_1361),
.B1(n_1365),
.B2(n_1311),
.Y(n_1488)
);

OAI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1319),
.A2(n_1361),
.B1(n_1365),
.B2(n_938),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1248),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_SL g1491 ( 
.A1(n_1311),
.A2(n_1132),
.B1(n_899),
.B2(n_1378),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1323),
.Y(n_1492)
);

AOI21xp33_ASAP7_75t_L g1493 ( 
.A1(n_1228),
.A2(n_938),
.B(n_1311),
.Y(n_1493)
);

INVxp67_ASAP7_75t_SL g1494 ( 
.A(n_1257),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1311),
.A2(n_938),
.B1(n_1378),
.B2(n_899),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1248),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1327),
.Y(n_1497)
);

CKINVDCx11_ASAP7_75t_R g1498 ( 
.A(n_1280),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1319),
.A2(n_1361),
.B1(n_1365),
.B2(n_1311),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1265),
.Y(n_1500)
);

BUFx8_ASAP7_75t_SL g1501 ( 
.A(n_1331),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1311),
.A2(n_1132),
.B1(n_899),
.B2(n_1378),
.Y(n_1502)
);

BUFx8_ASAP7_75t_L g1503 ( 
.A(n_1269),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1316),
.B(n_1326),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1323),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1344),
.Y(n_1506)
);

OAI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1319),
.A2(n_1361),
.B1(n_1365),
.B2(n_938),
.Y(n_1507)
);

INVx4_ASAP7_75t_L g1508 ( 
.A(n_1344),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1345),
.A2(n_938),
.B(n_1373),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1327),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_SL g1511 ( 
.A1(n_1311),
.A2(n_1132),
.B1(n_899),
.B2(n_1378),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1344),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1319),
.A2(n_1361),
.B1(n_1365),
.B2(n_1311),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1319),
.A2(n_1361),
.B1(n_1365),
.B2(n_1311),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1332),
.Y(n_1515)
);

BUFx2_ASAP7_75t_SL g1516 ( 
.A(n_1331),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1224),
.Y(n_1517)
);

INVx3_ASAP7_75t_SL g1518 ( 
.A(n_1323),
.Y(n_1518)
);

INVx5_ASAP7_75t_L g1519 ( 
.A(n_1344),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1455),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1439),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1455),
.Y(n_1522)
);

INVx11_ASAP7_75t_L g1523 ( 
.A(n_1484),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1390),
.Y(n_1524)
);

AND2x2_ASAP7_75t_SL g1525 ( 
.A(n_1384),
.B(n_1411),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1458),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1388),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1387),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1401),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1408),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1433),
.B(n_1434),
.Y(n_1531)
);

INVx2_ASAP7_75t_SL g1532 ( 
.A(n_1465),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1477),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1473),
.A2(n_1454),
.B(n_1438),
.Y(n_1534)
);

OA21x2_ASAP7_75t_L g1535 ( 
.A1(n_1443),
.A2(n_1462),
.B(n_1448),
.Y(n_1535)
);

AO21x2_ASAP7_75t_L g1536 ( 
.A1(n_1509),
.A2(n_1469),
.B(n_1473),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1427),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1433),
.B(n_1434),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1410),
.Y(n_1539)
);

AOI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1424),
.A2(n_1463),
.B(n_1449),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1426),
.Y(n_1541)
);

NAND2x1_ASAP7_75t_L g1542 ( 
.A(n_1465),
.B(n_1442),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1398),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1412),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1423),
.Y(n_1545)
);

AO21x1_ASAP7_75t_L g1546 ( 
.A1(n_1435),
.A2(n_1507),
.B(n_1489),
.Y(n_1546)
);

OR2x6_ASAP7_75t_L g1547 ( 
.A(n_1488),
.B(n_1499),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1513),
.B(n_1514),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1464),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1462),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1466),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1461),
.B(n_1404),
.Y(n_1552)
);

CKINVDCx20_ASAP7_75t_R g1553 ( 
.A(n_1403),
.Y(n_1553)
);

BUFx12f_ASAP7_75t_L g1554 ( 
.A(n_1498),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1448),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1494),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1487),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1494),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1386),
.B(n_1389),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1490),
.Y(n_1560)
);

OA21x2_ASAP7_75t_L g1561 ( 
.A1(n_1421),
.A2(n_1504),
.B(n_1432),
.Y(n_1561)
);

INVx2_ASAP7_75t_SL g1562 ( 
.A(n_1465),
.Y(n_1562)
);

AO21x2_ASAP7_75t_L g1563 ( 
.A1(n_1469),
.A2(n_1453),
.B(n_1493),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_1519),
.Y(n_1564)
);

BUFx3_ASAP7_75t_L g1565 ( 
.A(n_1459),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1496),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_1383),
.Y(n_1567)
);

AO21x2_ASAP7_75t_L g1568 ( 
.A1(n_1453),
.A2(n_1493),
.B(n_1437),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1457),
.B(n_1419),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1415),
.B(n_1447),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1382),
.B(n_1399),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1415),
.B(n_1447),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1437),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1397),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1468),
.Y(n_1575)
);

BUFx10_ASAP7_75t_L g1576 ( 
.A(n_1446),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1475),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1413),
.B(n_1481),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1456),
.Y(n_1579)
);

OAI21x1_ASAP7_75t_L g1580 ( 
.A1(n_1436),
.A2(n_1416),
.B(n_1444),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1470),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1479),
.A2(n_1495),
.B(n_1502),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1489),
.A2(n_1507),
.B(n_1382),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1470),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1468),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1472),
.Y(n_1586)
);

INVx3_ASAP7_75t_L g1587 ( 
.A(n_1468),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1467),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1467),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1460),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1381),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1500),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1430),
.Y(n_1593)
);

OR2x6_ASAP7_75t_L g1594 ( 
.A(n_1391),
.B(n_1476),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_1519),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1395),
.B(n_1402),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1471),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1471),
.B(n_1394),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1392),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1418),
.Y(n_1600)
);

NAND2x1p5_ASAP7_75t_L g1601 ( 
.A(n_1519),
.B(n_1476),
.Y(n_1601)
);

AO21x2_ASAP7_75t_L g1602 ( 
.A1(n_1385),
.A2(n_1460),
.B(n_1441),
.Y(n_1602)
);

OAI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1491),
.A2(n_1502),
.B(n_1511),
.Y(n_1603)
);

NAND2x1p5_ASAP7_75t_L g1604 ( 
.A(n_1391),
.B(n_1508),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1385),
.B(n_1420),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1517),
.Y(n_1606)
);

OAI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1506),
.A2(n_1512),
.B(n_1452),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1474),
.B(n_1511),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1446),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1474),
.Y(n_1610)
);

BUFx2_ASAP7_75t_L g1611 ( 
.A(n_1417),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1386),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1430),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_1486),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1491),
.B(n_1422),
.Y(n_1615)
);

A2O1A1Ixp33_ASAP7_75t_L g1616 ( 
.A1(n_1583),
.A2(n_1603),
.B(n_1582),
.C(n_1608),
.Y(n_1616)
);

OAI21xp33_ASAP7_75t_SL g1617 ( 
.A1(n_1608),
.A2(n_1440),
.B(n_1396),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1547),
.A2(n_1428),
.B1(n_1409),
.B2(n_1425),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1522),
.B(n_1520),
.Y(n_1619)
);

A2O1A1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1548),
.A2(n_1422),
.B(n_1452),
.C(n_1429),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1552),
.B(n_1516),
.Y(n_1621)
);

OA21x2_ASAP7_75t_L g1622 ( 
.A1(n_1534),
.A2(n_1482),
.B(n_1450),
.Y(n_1622)
);

A2O1A1Ixp33_ASAP7_75t_L g1623 ( 
.A1(n_1548),
.A2(n_1445),
.B(n_1451),
.C(n_1431),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1552),
.B(n_1483),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1547),
.A2(n_1518),
.B1(n_1480),
.B2(n_1414),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1578),
.B(n_1480),
.Y(n_1626)
);

INVxp67_ASAP7_75t_L g1627 ( 
.A(n_1541),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1541),
.B(n_1400),
.Y(n_1628)
);

AO32x2_ASAP7_75t_L g1629 ( 
.A1(n_1537),
.A2(n_1396),
.A3(n_1503),
.B1(n_1484),
.B2(n_1515),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1554),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1537),
.B(n_1518),
.Y(n_1631)
);

AOI221xp5_ASAP7_75t_L g1632 ( 
.A1(n_1546),
.A2(n_1510),
.B1(n_1406),
.B2(n_1497),
.C(n_1505),
.Y(n_1632)
);

OA21x2_ASAP7_75t_L g1633 ( 
.A1(n_1534),
.A2(n_1492),
.B(n_1446),
.Y(n_1633)
);

AOI221xp5_ASAP7_75t_L g1634 ( 
.A1(n_1546),
.A2(n_1393),
.B1(n_1400),
.B2(n_1515),
.C(n_1503),
.Y(n_1634)
);

A2O1A1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1525),
.A2(n_1515),
.B(n_1501),
.C(n_1478),
.Y(n_1635)
);

INVxp33_ASAP7_75t_L g1636 ( 
.A(n_1524),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1560),
.Y(n_1637)
);

INVx4_ASAP7_75t_L g1638 ( 
.A(n_1576),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1522),
.B(n_1405),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1566),
.Y(n_1640)
);

INVxp67_ASAP7_75t_L g1641 ( 
.A(n_1543),
.Y(n_1641)
);

OA21x2_ASAP7_75t_L g1642 ( 
.A1(n_1580),
.A2(n_1407),
.B(n_1485),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1571),
.B(n_1556),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1525),
.A2(n_1547),
.B(n_1580),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1547),
.B(n_1605),
.Y(n_1645)
);

AO32x2_ASAP7_75t_L g1646 ( 
.A1(n_1579),
.A2(n_1532),
.A3(n_1562),
.B1(n_1581),
.B2(n_1584),
.Y(n_1646)
);

OA21x2_ASAP7_75t_L g1647 ( 
.A1(n_1540),
.A2(n_1585),
.B(n_1573),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1525),
.A2(n_1540),
.B(n_1571),
.Y(n_1648)
);

A2O1A1Ixp33_ASAP7_75t_L g1649 ( 
.A1(n_1559),
.A2(n_1570),
.B(n_1572),
.C(n_1596),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1527),
.B(n_1529),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1596),
.B(n_1610),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1533),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1558),
.B(n_1573),
.Y(n_1653)
);

AOI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1610),
.A2(n_1598),
.B1(n_1538),
.B2(n_1531),
.C(n_1568),
.Y(n_1654)
);

BUFx3_ASAP7_75t_L g1655 ( 
.A(n_1554),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1523),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1529),
.B(n_1530),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1558),
.A2(n_1542),
.B(n_1536),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1569),
.B(n_1530),
.Y(n_1659)
);

OAI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1542),
.A2(n_1574),
.B(n_1598),
.Y(n_1660)
);

NOR2x1_ASAP7_75t_SL g1661 ( 
.A(n_1564),
.B(n_1595),
.Y(n_1661)
);

AOI211xp5_ASAP7_75t_L g1662 ( 
.A1(n_1615),
.A2(n_1586),
.B(n_1565),
.C(n_1538),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1539),
.B(n_1544),
.Y(n_1663)
);

A2O1A1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1531),
.A2(n_1565),
.B(n_1581),
.C(n_1584),
.Y(n_1664)
);

A2O1A1Ixp33_ASAP7_75t_L g1665 ( 
.A1(n_1565),
.A2(n_1586),
.B(n_1588),
.C(n_1589),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_1545),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1612),
.A2(n_1553),
.B1(n_1568),
.B2(n_1611),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1550),
.B(n_1557),
.Y(n_1668)
);

A2O1A1Ixp33_ASAP7_75t_L g1669 ( 
.A1(n_1588),
.A2(n_1589),
.B(n_1597),
.C(n_1555),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1568),
.A2(n_1611),
.B1(n_1593),
.B2(n_1577),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1528),
.B(n_1592),
.Y(n_1671)
);

BUFx6f_ASAP7_75t_L g1672 ( 
.A(n_1567),
.Y(n_1672)
);

OAI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1585),
.A2(n_1607),
.B(n_1526),
.Y(n_1673)
);

NOR2x1_ASAP7_75t_L g1674 ( 
.A(n_1593),
.B(n_1567),
.Y(n_1674)
);

AOI21xp33_ASAP7_75t_L g1675 ( 
.A1(n_1563),
.A2(n_1561),
.B(n_1602),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1614),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1627),
.B(n_1536),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1652),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1627),
.B(n_1602),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1659),
.B(n_1536),
.Y(n_1680)
);

INVxp67_ASAP7_75t_SL g1681 ( 
.A(n_1652),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1675),
.B(n_1602),
.Y(n_1682)
);

INVx4_ASAP7_75t_L g1683 ( 
.A(n_1638),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1637),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1626),
.B(n_1593),
.Y(n_1685)
);

INVx3_ASAP7_75t_R g1686 ( 
.A(n_1639),
.Y(n_1686)
);

INVxp33_ASAP7_75t_L g1687 ( 
.A(n_1671),
.Y(n_1687)
);

AOI221xp5_ASAP7_75t_L g1688 ( 
.A1(n_1616),
.A2(n_1597),
.B1(n_1563),
.B2(n_1606),
.C(n_1549),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1640),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1666),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1643),
.B(n_1654),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1675),
.B(n_1563),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1673),
.B(n_1590),
.Y(n_1693)
);

INVx2_ASAP7_75t_SL g1694 ( 
.A(n_1650),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1654),
.B(n_1555),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1666),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1622),
.B(n_1535),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1670),
.B(n_1616),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1622),
.B(n_1535),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1658),
.B(n_1653),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1657),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1663),
.B(n_1535),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1668),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1632),
.A2(n_1561),
.B1(n_1575),
.B2(n_1587),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_1672),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1632),
.A2(n_1561),
.B1(n_1575),
.B2(n_1587),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1668),
.Y(n_1707)
);

OAI222xp33_ASAP7_75t_L g1708 ( 
.A1(n_1667),
.A2(n_1594),
.B1(n_1551),
.B2(n_1591),
.C1(n_1600),
.C2(n_1599),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1647),
.B(n_1551),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1646),
.B(n_1521),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1687),
.B(n_1626),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1698),
.A2(n_1649),
.B1(n_1688),
.B2(n_1691),
.C(n_1644),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1678),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1678),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1691),
.B(n_1641),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1684),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1684),
.Y(n_1717)
);

OAI211xp5_ASAP7_75t_L g1718 ( 
.A1(n_1698),
.A2(n_1664),
.B(n_1662),
.C(n_1634),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1684),
.Y(n_1719)
);

BUFx6f_ASAP7_75t_L g1720 ( 
.A(n_1683),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1689),
.Y(n_1721)
);

BUFx3_ASAP7_75t_L g1722 ( 
.A(n_1705),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1693),
.B(n_1661),
.Y(n_1723)
);

AND4x1_ASAP7_75t_L g1724 ( 
.A(n_1688),
.B(n_1634),
.C(n_1635),
.D(n_1623),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1710),
.Y(n_1725)
);

OAI33xp33_ASAP7_75t_L g1726 ( 
.A1(n_1695),
.A2(n_1641),
.A3(n_1618),
.B1(n_1625),
.B2(n_1631),
.B3(n_1645),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1695),
.A2(n_1664),
.B1(n_1648),
.B2(n_1651),
.C(n_1665),
.Y(n_1727)
);

BUFx3_ASAP7_75t_L g1728 ( 
.A(n_1705),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1689),
.Y(n_1729)
);

INVxp67_ASAP7_75t_SL g1730 ( 
.A(n_1690),
.Y(n_1730)
);

NAND4xp25_ASAP7_75t_L g1731 ( 
.A(n_1704),
.B(n_1706),
.C(n_1651),
.D(n_1665),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1710),
.Y(n_1732)
);

INVx4_ASAP7_75t_L g1733 ( 
.A(n_1683),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1689),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1680),
.B(n_1633),
.Y(n_1735)
);

NAND4xp25_ASAP7_75t_L g1736 ( 
.A(n_1704),
.B(n_1671),
.C(n_1635),
.D(n_1660),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1705),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1700),
.B(n_1633),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1680),
.B(n_1629),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1706),
.A2(n_1642),
.B1(n_1625),
.B2(n_1618),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1703),
.B(n_1636),
.Y(n_1741)
);

NAND3xp33_ASAP7_75t_L g1742 ( 
.A(n_1692),
.B(n_1669),
.C(n_1623),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1680),
.B(n_1702),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1702),
.B(n_1629),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1700),
.B(n_1561),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1710),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1702),
.B(n_1629),
.Y(n_1747)
);

BUFx6f_ASAP7_75t_L g1748 ( 
.A(n_1683),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1681),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1693),
.B(n_1619),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1725),
.B(n_1677),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1725),
.B(n_1677),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1745),
.B(n_1700),
.Y(n_1753)
);

BUFx2_ASAP7_75t_L g1754 ( 
.A(n_1723),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1732),
.B(n_1697),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1715),
.B(n_1703),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1716),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1716),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_SL g1759 ( 
.A(n_1731),
.B(n_1708),
.Y(n_1759)
);

BUFx3_ASAP7_75t_L g1760 ( 
.A(n_1722),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1746),
.B(n_1697),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1746),
.B(n_1699),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1717),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1719),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1713),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1749),
.B(n_1707),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1719),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1749),
.B(n_1707),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1711),
.B(n_1630),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1745),
.B(n_1679),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1738),
.B(n_1679),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1721),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1713),
.B(n_1690),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1714),
.B(n_1730),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1744),
.B(n_1699),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1738),
.B(n_1679),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1721),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1729),
.Y(n_1778)
);

INVx3_ASAP7_75t_L g1779 ( 
.A(n_1723),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1714),
.B(n_1696),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1729),
.Y(n_1781)
);

NOR2x1_ASAP7_75t_L g1782 ( 
.A(n_1742),
.B(n_1674),
.Y(n_1782)
);

NOR2xp67_ASAP7_75t_L g1783 ( 
.A(n_1742),
.B(n_1709),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1743),
.B(n_1694),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1734),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1734),
.Y(n_1786)
);

INVx5_ASAP7_75t_L g1787 ( 
.A(n_1720),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1744),
.B(n_1699),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1783),
.Y(n_1789)
);

INVxp67_ASAP7_75t_L g1790 ( 
.A(n_1782),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1754),
.B(n_1747),
.Y(n_1791)
);

INVxp67_ASAP7_75t_L g1792 ( 
.A(n_1782),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1765),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1763),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1774),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1774),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1753),
.B(n_1743),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1773),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1759),
.A2(n_1712),
.B(n_1718),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1757),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1783),
.B(n_1727),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1757),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1753),
.B(n_1694),
.Y(n_1803)
);

AOI32xp33_ASAP7_75t_L g1804 ( 
.A1(n_1759),
.A2(n_1739),
.A3(n_1747),
.B1(n_1740),
.B2(n_1692),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1756),
.B(n_1739),
.Y(n_1805)
);

OAI21xp33_ASAP7_75t_L g1806 ( 
.A1(n_1756),
.A2(n_1731),
.B(n_1736),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1773),
.Y(n_1807)
);

CKINVDCx16_ASAP7_75t_R g1808 ( 
.A(n_1769),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1760),
.B(n_1655),
.Y(n_1809)
);

NAND2xp33_ASAP7_75t_SL g1810 ( 
.A(n_1754),
.B(n_1686),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1780),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1763),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1771),
.B(n_1694),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1760),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1763),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1764),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1779),
.B(n_1723),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1779),
.B(n_1723),
.Y(n_1818)
);

INVxp67_ASAP7_75t_L g1819 ( 
.A(n_1760),
.Y(n_1819)
);

BUFx2_ASAP7_75t_L g1820 ( 
.A(n_1787),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1787),
.B(n_1733),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1764),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1779),
.B(n_1750),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1771),
.B(n_1701),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1780),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1758),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1779),
.B(n_1750),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1776),
.B(n_1701),
.Y(n_1828)
);

NAND2x2_ASAP7_75t_L g1829 ( 
.A(n_1784),
.B(n_1656),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1766),
.B(n_1741),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1787),
.B(n_1733),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1766),
.B(n_1735),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1820),
.B(n_1787),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1806),
.B(n_1735),
.Y(n_1834)
);

OAI21xp33_ASAP7_75t_L g1835 ( 
.A1(n_1801),
.A2(n_1724),
.B(n_1692),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1789),
.Y(n_1836)
);

AOI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1799),
.A2(n_1726),
.B(n_1787),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1791),
.B(n_1814),
.Y(n_1838)
);

NAND4xp25_ASAP7_75t_L g1839 ( 
.A(n_1804),
.B(n_1790),
.C(n_1792),
.D(n_1809),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1810),
.A2(n_1642),
.B1(n_1685),
.B2(n_1617),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1793),
.B(n_1776),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1819),
.B(n_1775),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1808),
.B(n_1775),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1798),
.B(n_1770),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1791),
.B(n_1787),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1830),
.B(n_1523),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1810),
.A2(n_1787),
.B(n_1768),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1795),
.B(n_1775),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1796),
.B(n_1788),
.Y(n_1849)
);

INVx3_ASAP7_75t_L g1850 ( 
.A(n_1821),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1807),
.B(n_1676),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1800),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1800),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1820),
.Y(n_1854)
);

NAND3xp33_ASAP7_75t_L g1855 ( 
.A(n_1811),
.B(n_1724),
.C(n_1682),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1825),
.B(n_1788),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1802),
.Y(n_1857)
);

AND2x4_ASAP7_75t_L g1858 ( 
.A(n_1821),
.B(n_1751),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1823),
.B(n_1788),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1823),
.B(n_1751),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1802),
.Y(n_1861)
);

INVxp67_ASAP7_75t_L g1862 ( 
.A(n_1821),
.Y(n_1862)
);

A2O1A1Ixp33_ASAP7_75t_L g1863 ( 
.A1(n_1831),
.A2(n_1682),
.B(n_1669),
.C(n_1770),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1827),
.B(n_1751),
.Y(n_1864)
);

HB1xp67_ASAP7_75t_L g1865 ( 
.A(n_1803),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1803),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1827),
.B(n_1752),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1826),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1794),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1836),
.B(n_1805),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1835),
.A2(n_1855),
.B(n_1837),
.Y(n_1871)
);

INVx2_ASAP7_75t_SL g1872 ( 
.A(n_1833),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1839),
.A2(n_1834),
.B1(n_1843),
.B2(n_1829),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1845),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1846),
.B(n_1831),
.Y(n_1875)
);

INVx2_ASAP7_75t_SL g1876 ( 
.A(n_1833),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1852),
.Y(n_1877)
);

OA21x2_ASAP7_75t_L g1878 ( 
.A1(n_1847),
.A2(n_1831),
.B(n_1812),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1852),
.Y(n_1879)
);

OAI32xp33_ASAP7_75t_L g1880 ( 
.A1(n_1838),
.A2(n_1829),
.A3(n_1797),
.B1(n_1832),
.B2(n_1824),
.Y(n_1880)
);

NAND2xp33_ASAP7_75t_SL g1881 ( 
.A(n_1838),
.B(n_1686),
.Y(n_1881)
);

AOI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1863),
.A2(n_1768),
.B(n_1682),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1853),
.Y(n_1883)
);

OAI21xp5_ASAP7_75t_L g1884 ( 
.A1(n_1840),
.A2(n_1862),
.B(n_1845),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1853),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1857),
.Y(n_1886)
);

INVxp67_ASAP7_75t_SL g1887 ( 
.A(n_1850),
.Y(n_1887)
);

OAI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1833),
.A2(n_1818),
.B(n_1817),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1861),
.Y(n_1889)
);

AOI222xp33_ASAP7_75t_L g1890 ( 
.A1(n_1842),
.A2(n_1818),
.B1(n_1817),
.B2(n_1621),
.C1(n_1624),
.C2(n_1708),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1865),
.B(n_1797),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1868),
.Y(n_1892)
);

INVxp67_ASAP7_75t_SL g1893 ( 
.A(n_1850),
.Y(n_1893)
);

O2A1O1Ixp33_ASAP7_75t_L g1894 ( 
.A1(n_1854),
.A2(n_1794),
.B(n_1812),
.C(n_1822),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1866),
.A2(n_1720),
.B1(n_1748),
.B2(n_1750),
.Y(n_1895)
);

OAI221xp5_ASAP7_75t_L g1896 ( 
.A1(n_1871),
.A2(n_1850),
.B1(n_1851),
.B2(n_1854),
.C(n_1841),
.Y(n_1896)
);

BUFx2_ASAP7_75t_SL g1897 ( 
.A(n_1887),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1893),
.B(n_1868),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1875),
.B(n_1841),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1892),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1881),
.A2(n_1858),
.B1(n_1849),
.B2(n_1848),
.Y(n_1901)
);

AOI21xp33_ASAP7_75t_R g1902 ( 
.A1(n_1874),
.A2(n_1869),
.B(n_1856),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1874),
.B(n_1859),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1881),
.A2(n_1858),
.B1(n_1859),
.B2(n_1844),
.Y(n_1904)
);

AOI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1873),
.A2(n_1858),
.B1(n_1867),
.B2(n_1864),
.Y(n_1905)
);

OAI322xp33_ASAP7_75t_L g1906 ( 
.A1(n_1882),
.A2(n_1844),
.A3(n_1869),
.B1(n_1824),
.B2(n_1828),
.C1(n_1813),
.C2(n_1860),
.Y(n_1906)
);

OAI21xp5_ASAP7_75t_SL g1907 ( 
.A1(n_1884),
.A2(n_1890),
.B(n_1895),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1888),
.B(n_1872),
.Y(n_1908)
);

OA21x2_ASAP7_75t_L g1909 ( 
.A1(n_1892),
.A2(n_1816),
.B(n_1815),
.Y(n_1909)
);

AOI211xp5_ASAP7_75t_L g1910 ( 
.A1(n_1880),
.A2(n_1867),
.B(n_1864),
.C(n_1860),
.Y(n_1910)
);

INVxp67_ASAP7_75t_L g1911 ( 
.A(n_1872),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1886),
.B(n_1815),
.Y(n_1912)
);

BUFx2_ASAP7_75t_L g1913 ( 
.A(n_1876),
.Y(n_1913)
);

INVx1_ASAP7_75t_SL g1914 ( 
.A(n_1891),
.Y(n_1914)
);

NAND3xp33_ASAP7_75t_L g1915 ( 
.A(n_1876),
.B(n_1822),
.C(n_1816),
.Y(n_1915)
);

INVx1_ASAP7_75t_SL g1916 ( 
.A(n_1897),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1913),
.B(n_1870),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1898),
.Y(n_1918)
);

NOR4xp25_ASAP7_75t_L g1919 ( 
.A(n_1896),
.B(n_1889),
.C(n_1877),
.D(n_1885),
.Y(n_1919)
);

AOI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1907),
.A2(n_1880),
.B(n_1878),
.Y(n_1920)
);

AOI21xp33_ASAP7_75t_SL g1921 ( 
.A1(n_1899),
.A2(n_1878),
.B(n_1889),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1898),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1900),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1908),
.B(n_1878),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1911),
.B(n_1914),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1904),
.B(n_1894),
.Y(n_1926)
);

AOI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1905),
.A2(n_1883),
.B1(n_1879),
.B2(n_1733),
.Y(n_1927)
);

NOR3xp33_ASAP7_75t_L g1928 ( 
.A(n_1916),
.B(n_1903),
.C(n_1906),
.Y(n_1928)
);

AOI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1926),
.A2(n_1901),
.B1(n_1910),
.B2(n_1915),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1925),
.B(n_1912),
.Y(n_1930)
);

NOR2x1_ASAP7_75t_L g1931 ( 
.A(n_1918),
.B(n_1909),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_L g1932 ( 
.A(n_1917),
.B(n_1912),
.Y(n_1932)
);

NOR2x1_ASAP7_75t_L g1933 ( 
.A(n_1922),
.B(n_1909),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1917),
.B(n_1902),
.Y(n_1934)
);

NAND5xp2_ASAP7_75t_L g1935 ( 
.A(n_1920),
.B(n_1601),
.C(n_1604),
.D(n_1620),
.E(n_1628),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1924),
.B(n_1813),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1923),
.Y(n_1937)
);

NOR3xp33_ASAP7_75t_L g1938 ( 
.A(n_1926),
.B(n_1639),
.C(n_1733),
.Y(n_1938)
);

AOI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1921),
.A2(n_1828),
.B(n_1785),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1932),
.B(n_1927),
.Y(n_1940)
);

INVx1_ASAP7_75t_SL g1941 ( 
.A(n_1934),
.Y(n_1941)
);

A2O1A1Ixp33_ASAP7_75t_L g1942 ( 
.A1(n_1929),
.A2(n_1931),
.B(n_1933),
.C(n_1928),
.Y(n_1942)
);

OAI221xp5_ASAP7_75t_SL g1943 ( 
.A1(n_1938),
.A2(n_1919),
.B1(n_1924),
.B2(n_1728),
.C(n_1722),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1936),
.Y(n_1944)
);

O2A1O1Ixp33_ASAP7_75t_L g1945 ( 
.A1(n_1930),
.A2(n_1737),
.B(n_1620),
.C(n_1728),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1944),
.Y(n_1946)
);

OAI211xp5_ASAP7_75t_SL g1947 ( 
.A1(n_1942),
.A2(n_1937),
.B(n_1939),
.C(n_1935),
.Y(n_1947)
);

AOI211x1_ASAP7_75t_SL g1948 ( 
.A1(n_1943),
.A2(n_1764),
.B(n_1785),
.C(n_1720),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1940),
.A2(n_1941),
.B(n_1945),
.Y(n_1949)
);

AOI32xp33_ASAP7_75t_L g1950 ( 
.A1(n_1941),
.A2(n_1728),
.A3(n_1722),
.B1(n_1761),
.B2(n_1762),
.Y(n_1950)
);

BUFx8_ASAP7_75t_SL g1951 ( 
.A(n_1944),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1941),
.B(n_1720),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1951),
.Y(n_1953)
);

NOR2x1_ASAP7_75t_L g1954 ( 
.A(n_1946),
.B(n_1785),
.Y(n_1954)
);

NOR2xp33_ASAP7_75t_L g1955 ( 
.A(n_1947),
.B(n_1720),
.Y(n_1955)
);

XOR2xp5_ASAP7_75t_L g1956 ( 
.A(n_1949),
.B(n_1613),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1952),
.B(n_1784),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1948),
.B(n_1755),
.Y(n_1958)
);

NOR2x1p5_ASAP7_75t_L g1959 ( 
.A(n_1953),
.B(n_1950),
.Y(n_1959)
);

XOR2xp5_ASAP7_75t_L g1960 ( 
.A(n_1956),
.B(n_1613),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1954),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1959),
.B(n_1955),
.Y(n_1962)
);

AOI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1962),
.A2(n_1960),
.B1(n_1961),
.B2(n_1957),
.Y(n_1963)
);

XOR2xp5_ASAP7_75t_L g1964 ( 
.A(n_1963),
.B(n_1958),
.Y(n_1964)
);

XOR2x2_ASAP7_75t_L g1965 ( 
.A(n_1963),
.B(n_1604),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1964),
.B(n_1613),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1965),
.Y(n_1967)
);

OA22x2_ASAP7_75t_L g1968 ( 
.A1(n_1967),
.A2(n_1737),
.B1(n_1781),
.B2(n_1778),
.Y(n_1968)
);

AOI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1966),
.A2(n_1748),
.B1(n_1720),
.B2(n_1755),
.Y(n_1969)
);

AOI221xp5_ASAP7_75t_L g1970 ( 
.A1(n_1969),
.A2(n_1968),
.B1(n_1748),
.B2(n_1781),
.C(n_1778),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_SL g1971 ( 
.A1(n_1970),
.A2(n_1604),
.B(n_1601),
.Y(n_1971)
);

XNOR2xp5_ASAP7_75t_L g1972 ( 
.A(n_1971),
.B(n_1609),
.Y(n_1972)
);

AOI221xp5_ASAP7_75t_L g1973 ( 
.A1(n_1972),
.A2(n_1786),
.B1(n_1777),
.B2(n_1772),
.C(n_1767),
.Y(n_1973)
);

AOI211xp5_ASAP7_75t_L g1974 ( 
.A1(n_1973),
.A2(n_1613),
.B(n_1609),
.C(n_1748),
.Y(n_1974)
);


endmodule