module fake_jpeg_2271_n_589 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_589);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_589;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_13),
.B(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_11),
.B(n_5),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_60),
.Y(n_164)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_61),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_62),
.B(n_67),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_63),
.Y(n_157)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_65),
.Y(n_159)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_16),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_71),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_80),
.Y(n_124)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_29),
.Y(n_76)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_78),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_28),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_82),
.B(n_100),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_83),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_85),
.Y(n_171)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_86),
.Y(n_163)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_89),
.Y(n_180)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_92),
.Y(n_182)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_21),
.B(n_12),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_95),
.B(n_112),
.Y(n_186)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_20),
.B(n_1),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_101),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_26),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_102),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_27),
.B(n_1),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_2),
.Y(n_148)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_106),
.Y(n_184)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_41),
.Y(n_107)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_109),
.Y(n_173)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_21),
.B(n_2),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_19),
.Y(n_113)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_30),
.Y(n_114)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_24),
.B(n_2),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_115),
.B(n_2),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_27),
.Y(n_117)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_30),
.Y(n_119)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_119),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_30),
.Y(n_120)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_73),
.A2(n_44),
.B1(n_30),
.B2(n_48),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_138),
.A2(n_151),
.B1(n_156),
.B2(n_166),
.Y(n_234)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_142),
.Y(n_199)
);

AOI21xp33_ASAP7_75t_L g254 ( 
.A1(n_148),
.A2(n_187),
.B(n_56),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_82),
.A2(n_38),
.B1(n_48),
.B2(n_47),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_100),
.A2(n_38),
.B1(n_48),
.B2(n_47),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_103),
.A2(n_23),
.B1(n_47),
.B2(n_38),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_167),
.Y(n_227)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_69),
.Y(n_169)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_85),
.Y(n_174)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_174),
.Y(n_228)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_59),
.Y(n_178)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_178),
.Y(n_263)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_60),
.Y(n_181)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_83),
.B(n_32),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_185),
.B(n_192),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_83),
.B(n_32),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_186),
.Y(n_224)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_92),
.Y(n_189)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_114),
.Y(n_190)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_88),
.A2(n_23),
.B1(n_70),
.B2(n_79),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_191),
.A2(n_194),
.B1(n_36),
.B2(n_24),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_63),
.B(n_35),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_72),
.A2(n_47),
.B1(n_38),
.B2(n_48),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_78),
.Y(n_195)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_84),
.Y(n_196)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_133),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_200),
.Y(n_271)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_131),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_202),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_166),
.A2(n_106),
.B1(n_102),
.B2(n_108),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_203),
.A2(n_244),
.B1(n_234),
.B2(n_173),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_124),
.A2(n_23),
.B1(n_22),
.B2(n_37),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_204),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_205),
.Y(n_273)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_206),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_207),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_208),
.Y(n_326)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_160),
.Y(n_209)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_209),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_210),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_187),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_211),
.B(n_216),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_71),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_214),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_146),
.A2(n_37),
.B(n_58),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_215),
.A2(n_226),
.B(n_231),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_152),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

INVx8_ASAP7_75t_L g283 ( 
.A(n_217),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_124),
.B(n_31),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_220),
.B(n_224),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_140),
.B(n_119),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_222),
.B(n_223),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_140),
.B(n_119),
.Y(n_223)
);

O2A1O1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_156),
.A2(n_138),
.B(n_151),
.C(n_134),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_135),
.B(n_49),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_230),
.B(n_255),
.Y(n_320)
);

O2A1O1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_139),
.A2(n_98),
.B(n_96),
.C(n_110),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_130),
.Y(n_232)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_232),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_122),
.B(n_51),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_233),
.B(n_239),
.C(n_8),
.Y(n_306)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_162),
.Y(n_235)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_235),
.Y(n_285)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_158),
.Y(n_236)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_236),
.Y(n_323)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_176),
.Y(n_237)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_237),
.Y(n_327)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_123),
.Y(n_238)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_238),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_146),
.B(n_49),
.C(n_19),
.Y(n_239)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_240),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_128),
.B(n_31),
.Y(n_241)
);

NOR3xp33_ASAP7_75t_L g276 ( 
.A(n_241),
.B(n_242),
.C(n_253),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_148),
.B(n_22),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_147),
.A2(n_51),
.B1(n_58),
.B2(n_56),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_243),
.A2(n_258),
.B1(n_262),
.B2(n_268),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_191),
.A2(n_111),
.B1(n_93),
.B2(n_35),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_163),
.A2(n_53),
.B1(n_50),
.B2(n_46),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_245),
.A2(n_264),
.B1(n_173),
.B2(n_149),
.Y(n_275)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_141),
.Y(n_246)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_246),
.Y(n_288)
);

INVx3_ASAP7_75t_SL g247 ( 
.A(n_183),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_161),
.Y(n_248)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_248),
.Y(n_319)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_127),
.Y(n_249)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_249),
.Y(n_292)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_143),
.Y(n_250)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_250),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_157),
.Y(n_251)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_251),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_136),
.A2(n_46),
.B1(n_36),
.B2(n_53),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_252),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_121),
.A2(n_50),
.B(n_42),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_254),
.B(n_256),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_165),
.B(n_42),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_132),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_150),
.Y(n_257)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_257),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_170),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_259),
.B(n_260),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_153),
.Y(n_260)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_137),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_261),
.Y(n_318)
);

INVx11_ASAP7_75t_L g262 ( 
.A(n_168),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_125),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_129),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_266),
.Y(n_300)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_180),
.Y(n_266)
);

O2A1O1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_145),
.A2(n_77),
.B(n_4),
.C(n_6),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_267),
.A2(n_168),
.B(n_144),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_171),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_182),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_269),
.B(n_12),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_226),
.A2(n_164),
.B1(n_179),
.B2(n_197),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_272),
.A2(n_284),
.B1(n_290),
.B2(n_304),
.Y(n_342)
);

OAI21xp33_ASAP7_75t_SL g330 ( 
.A1(n_275),
.A2(n_302),
.B(n_324),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_215),
.B(n_164),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_277),
.B(n_282),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_214),
.B(n_197),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_214),
.B(n_221),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_287),
.B(n_293),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_239),
.A2(n_179),
.B1(n_193),
.B2(n_172),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_233),
.B(n_172),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_233),
.B(n_126),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_294),
.B(n_296),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_238),
.B(n_155),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_297),
.B(n_301),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_203),
.B(n_175),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_299),
.B(n_309),
.Y(n_341)
);

AO22x2_ASAP7_75t_L g301 ( 
.A1(n_244),
.A2(n_144),
.B1(n_10),
.B2(n_11),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_257),
.A2(n_202),
.B1(n_240),
.B2(n_209),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_199),
.A2(n_8),
.B1(n_12),
.B2(n_250),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_305),
.A2(n_315),
.B1(n_273),
.B2(n_289),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_306),
.B(n_206),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_307),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_228),
.B(n_229),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_201),
.B(n_219),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_225),
.Y(n_332)
);

A2O1A1Ixp33_ASAP7_75t_L g314 ( 
.A1(n_267),
.A2(n_231),
.B(n_222),
.C(n_223),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_314),
.A2(n_285),
.B(n_311),
.C(n_292),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_212),
.B(n_218),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_316),
.B(n_322),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_222),
.A2(n_223),
.B1(n_236),
.B2(n_269),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_266),
.A2(n_246),
.B1(n_248),
.B2(n_259),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_316),
.Y(n_329)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_329),
.Y(n_378)
);

OAI32xp33_ASAP7_75t_L g331 ( 
.A1(n_287),
.A2(n_321),
.A3(n_291),
.B1(n_299),
.B2(n_277),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_331),
.B(n_367),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_332),
.Y(n_392)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_286),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g396 ( 
.A(n_333),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_321),
.A2(n_207),
.B(n_213),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_334),
.A2(n_340),
.B(n_295),
.Y(n_382)
);

AO22x1_ASAP7_75t_SL g335 ( 
.A1(n_284),
.A2(n_229),
.B1(n_218),
.B2(n_212),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_335),
.B(n_357),
.Y(n_405)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_309),
.Y(n_336)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_336),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_200),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_337),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_338),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_310),
.Y(n_339)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_339),
.Y(n_389)
);

HB1xp67_ASAP7_75t_SL g340 ( 
.A(n_281),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_297),
.B(n_251),
.Y(n_344)
);

NOR2x1_ASAP7_75t_L g410 ( 
.A(n_344),
.B(n_371),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_312),
.A2(n_237),
.B1(n_261),
.B2(n_263),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_345),
.A2(n_351),
.B1(n_356),
.B2(n_344),
.Y(n_398)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_286),
.Y(n_346)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_346),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_312),
.A2(n_217),
.B1(n_227),
.B2(n_247),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_347),
.Y(n_407)
);

MAJx2_ASAP7_75t_L g348 ( 
.A(n_303),
.B(n_262),
.C(n_210),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_348),
.B(n_349),
.C(n_350),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_274),
.B(n_306),
.C(n_325),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_281),
.B(n_282),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_308),
.A2(n_272),
.B1(n_314),
.B2(n_301),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_352),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_278),
.B(n_276),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_355),
.B(n_373),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_301),
.A2(n_302),
.B1(n_293),
.B2(n_294),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_270),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_270),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_358),
.B(n_364),
.Y(n_393)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_323),
.Y(n_359)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_359),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_301),
.A2(n_281),
.B1(n_304),
.B2(n_318),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_362),
.A2(n_365),
.B1(n_369),
.B2(n_317),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_279),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_363),
.Y(n_379)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_326),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_298),
.A2(n_296),
.B1(n_300),
.B2(n_289),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_366),
.A2(n_271),
.B(n_327),
.Y(n_390)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_323),
.Y(n_368)
);

INVx13_ASAP7_75t_L g380 ( 
.A(n_368),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_327),
.A2(n_280),
.B1(n_326),
.B2(n_273),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_310),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_370),
.Y(n_384)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_322),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_372),
.B(n_357),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_288),
.B(n_319),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_288),
.B(n_319),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_374),
.B(n_317),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_350),
.B(n_311),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_376),
.B(n_391),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_271),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_381),
.B(n_364),
.C(n_372),
.Y(n_424)
);

OAI21xp33_ASAP7_75t_SL g414 ( 
.A1(n_382),
.A2(n_348),
.B(n_360),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_344),
.A2(n_295),
.B(n_280),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_383),
.A2(n_390),
.B(n_394),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_385),
.B(n_403),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_387),
.A2(n_398),
.B1(n_412),
.B2(n_342),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_353),
.B(n_283),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_344),
.A2(n_283),
.B(n_371),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_363),
.Y(n_399)
);

CKINVDCx14_ASAP7_75t_R g415 ( 
.A(n_399),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_366),
.A2(n_371),
.B(n_334),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_402),
.A2(n_410),
.B(n_394),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_370),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g404 ( 
.A(n_343),
.B(n_341),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_409),
.Y(n_423)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_408),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_329),
.B(n_336),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_410),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_361),
.B(n_343),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_413),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_342),
.A2(n_362),
.B1(n_351),
.B2(n_331),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_361),
.B(n_365),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_414),
.A2(n_447),
.B(n_384),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_416),
.A2(n_426),
.B1(n_390),
.B2(n_405),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_406),
.B(n_349),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_417),
.B(n_427),
.C(n_444),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_398),
.A2(n_356),
.B1(n_335),
.B2(n_330),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_419),
.A2(n_435),
.B1(n_439),
.B2(n_405),
.Y(n_475)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_408),
.Y(n_420)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_420),
.Y(n_460)
);

OA22x2_ASAP7_75t_L g422 ( 
.A1(n_402),
.A2(n_345),
.B1(n_335),
.B2(n_360),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_422),
.B(n_434),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_424),
.B(n_427),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_393),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_425),
.B(n_428),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_412),
.A2(n_338),
.B1(n_354),
.B2(n_369),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_406),
.B(n_354),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_393),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_385),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_430),
.B(n_443),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_358),
.Y(n_431)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_431),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_375),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_432),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_383),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_401),
.A2(n_368),
.B1(n_346),
.B2(n_333),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_395),
.Y(n_436)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_436),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_359),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_437),
.B(n_384),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_378),
.B(n_386),
.Y(n_438)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_438),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_401),
.A2(n_404),
.B1(n_411),
.B2(n_413),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_375),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_440),
.Y(n_458)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_395),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_376),
.B(n_381),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_444),
.B(n_387),
.Y(n_469)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_378),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_445),
.B(n_379),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_386),
.B(n_399),
.Y(n_446)
);

CKINVDCx14_ASAP7_75t_R g454 ( 
.A(n_446),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_417),
.B(n_376),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_449),
.B(n_461),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_450),
.B(n_453),
.C(n_463),
.Y(n_478)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_451),
.Y(n_487)
);

INVx13_ASAP7_75t_L g452 ( 
.A(n_415),
.Y(n_452)
);

CKINVDCx14_ASAP7_75t_R g488 ( 
.A(n_452),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_391),
.C(n_404),
.Y(n_453)
);

CKINVDCx14_ASAP7_75t_R g459 ( 
.A(n_418),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_459),
.B(n_476),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_439),
.B(n_382),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_421),
.B(n_410),
.C(n_397),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_466),
.A2(n_419),
.B1(n_416),
.B2(n_426),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_447),
.A2(n_388),
.B(n_405),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_467),
.A2(n_474),
.B(n_388),
.Y(n_503)
);

MAJx2_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_472),
.C(n_473),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_424),
.B(n_379),
.C(n_403),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_470),
.B(n_433),
.C(n_431),
.Y(n_494)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_471),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_423),
.B(n_377),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_423),
.B(n_377),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_475),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_446),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_429),
.B(n_405),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_477),
.B(n_422),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_392),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_480),
.B(n_465),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_481),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_454),
.A2(n_435),
.B1(n_442),
.B2(n_441),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_482),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_448),
.B(n_429),
.Y(n_484)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_484),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_475),
.A2(n_442),
.B1(n_441),
.B2(n_434),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_489),
.B(n_496),
.Y(n_504)
);

XNOR2x1_ASAP7_75t_L g491 ( 
.A(n_461),
.B(n_418),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_491),
.B(n_477),
.Y(n_520)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_456),
.Y(n_492)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_492),
.Y(n_518)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_471),
.Y(n_493)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_493),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_494),
.B(n_502),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_455),
.B(n_433),
.C(n_438),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_495),
.B(n_498),
.C(n_501),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_472),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_497),
.B(n_463),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_455),
.B(n_445),
.C(n_422),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_467),
.A2(n_388),
.B(n_407),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_499),
.A2(n_503),
.B(n_468),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_473),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_500),
.B(n_469),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_450),
.B(n_422),
.C(n_443),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_453),
.B(n_389),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_489),
.A2(n_468),
.B(n_474),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_506),
.B(n_513),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g507 ( 
.A(n_488),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_SL g534 ( 
.A1(n_507),
.A2(n_457),
.B1(n_509),
.B2(n_440),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_487),
.Y(n_510)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_510),
.Y(n_533)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_511),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_512),
.B(n_517),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_490),
.B(n_460),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_483),
.A2(n_460),
.B(n_465),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_514),
.B(n_521),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_515),
.B(n_520),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_502),
.B(n_449),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_495),
.B(n_501),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_522),
.B(n_478),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_498),
.B(n_462),
.C(n_458),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_524),
.B(n_525),
.C(n_497),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_494),
.B(n_462),
.C(n_458),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_526),
.B(n_517),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_527),
.B(n_528),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_519),
.A2(n_481),
.B1(n_486),
.B2(n_482),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_516),
.B(n_478),
.C(n_479),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_530),
.B(n_532),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_516),
.B(n_479),
.C(n_491),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_534),
.A2(n_464),
.B1(n_507),
.B2(n_505),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_522),
.B(n_485),
.C(n_503),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_536),
.B(n_538),
.C(n_515),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_523),
.A2(n_509),
.B1(n_506),
.B2(n_504),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_537),
.A2(n_541),
.B1(n_507),
.B2(n_520),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_508),
.B(n_485),
.C(n_499),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_525),
.A2(n_457),
.B1(n_464),
.B2(n_452),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_518),
.B(n_389),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_542),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_531),
.A2(n_512),
.B(n_524),
.Y(n_544)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_544),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_529),
.B(n_508),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_545),
.B(n_546),
.Y(n_558)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_539),
.Y(n_547)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_547),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_550),
.B(n_552),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_551),
.B(n_530),
.C(n_532),
.Y(n_559)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_541),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_553),
.B(n_554),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_526),
.B(n_432),
.C(n_396),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_537),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_555),
.Y(n_557)
);

NOR2x1_ASAP7_75t_L g556 ( 
.A(n_529),
.B(n_507),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_556),
.B(n_535),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_559),
.B(n_561),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_545),
.B(n_538),
.C(n_536),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_555),
.A2(n_540),
.B1(n_533),
.B2(n_535),
.Y(n_562)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_562),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_564),
.B(n_566),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_554),
.B(n_375),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_557),
.B(n_549),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_570),
.B(n_571),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_558),
.B(n_550),
.C(n_548),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_565),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g580 ( 
.A1(n_572),
.A2(n_380),
.B(n_396),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_560),
.A2(n_544),
.B(n_556),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_573),
.A2(n_557),
.B(n_543),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_561),
.B(n_551),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_574),
.B(n_558),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_576),
.B(n_578),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_568),
.B(n_567),
.C(n_563),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_579),
.B(n_580),
.C(n_575),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_581),
.A2(n_582),
.B(n_569),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_577),
.B(n_571),
.C(n_572),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_583),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_584),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_586),
.B(n_585),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_587),
.B(n_396),
.C(n_380),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_588),
.A2(n_396),
.B(n_380),
.Y(n_589)
);


endmodule