module fake_jpeg_28796_n_513 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_513);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_513;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_6),
.B(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_9),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_54),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_26),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_59),
.B(n_64),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_63),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_18),
.B(n_9),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_18),
.B(n_9),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_89),
.Y(n_103)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_75),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_23),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_82),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_31),
.B(n_8),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_21),
.B(n_8),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_87),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_8),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_26),
.B(n_10),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_27),
.B(n_10),
.C(n_1),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_95),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_27),
.B(n_10),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_96),
.Y(n_115)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_98),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_100),
.Y(n_140)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_50),
.A2(n_28),
.B1(n_30),
.B2(n_47),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_101),
.A2(n_104),
.B1(n_149),
.B2(n_152),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_56),
.A2(n_98),
.B1(n_97),
.B2(n_96),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_28),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_105),
.B(n_153),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_108),
.B(n_120),
.Y(n_210)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_29),
.B(n_30),
.C(n_47),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_109),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_55),
.A2(n_46),
.B1(n_25),
.B2(n_42),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_112),
.A2(n_114),
.B1(n_138),
.B2(n_159),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_83),
.A2(n_46),
.B1(n_49),
.B2(n_48),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_61),
.B(n_29),
.Y(n_120)
);

AND2x4_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_49),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_132),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_71),
.A2(n_38),
.B1(n_48),
.B2(n_36),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_53),
.B(n_37),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_155),
.C(n_22),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_58),
.A2(n_46),
.B1(n_49),
.B2(n_48),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_66),
.A2(n_38),
.B1(n_36),
.B2(n_45),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_143),
.A2(n_22),
.B1(n_63),
.B2(n_0),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_67),
.A2(n_37),
.B1(n_36),
.B2(n_35),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_69),
.A2(n_37),
.B1(n_35),
.B2(n_34),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_61),
.B(n_46),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_72),
.B(n_22),
.C(n_35),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_73),
.A2(n_46),
.B1(n_49),
.B2(n_45),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_46),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_161),
.B(n_170),
.Y(n_232)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_162),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_129),
.A2(n_24),
.B1(n_34),
.B2(n_43),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_165),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_111),
.Y(n_166)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_166),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_103),
.A2(n_24),
.B(n_45),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_168),
.B(n_0),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_140),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_169),
.B(n_182),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_102),
.B(n_49),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_171),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_115),
.B(n_31),
.Y(n_173)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_173),
.B(n_214),
.CI(n_160),
.CON(n_237),
.SN(n_237)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_174),
.Y(n_228)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_175),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_113),
.A2(n_90),
.B1(n_80),
.B2(n_78),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_179),
.A2(n_212),
.B1(n_116),
.B2(n_148),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_180),
.B(n_205),
.Y(n_268)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_181),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_109),
.B(n_113),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_106),
.A2(n_75),
.B1(n_74),
.B2(n_24),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_183),
.A2(n_207),
.B1(n_208),
.B2(n_5),
.Y(n_267)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_185),
.Y(n_254)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_132),
.A2(n_135),
.B1(n_149),
.B2(n_152),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g221 ( 
.A1(n_190),
.A2(n_112),
.B1(n_114),
.B2(n_159),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_110),
.B(n_43),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_191),
.B(n_198),
.Y(n_245)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_192),
.Y(n_255)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_193),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_111),
.Y(n_194)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_194),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_196),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_126),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_155),
.B(n_43),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_199),
.Y(n_248)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_119),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_201),
.Y(n_239)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_139),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_202),
.Y(n_235)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_203),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_127),
.B(n_34),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_215),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_138),
.A2(n_88),
.B(n_84),
.Y(n_205)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_128),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_206),
.A2(n_122),
.B1(n_141),
.B2(n_123),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_106),
.A2(n_49),
.B1(n_31),
.B2(n_2),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_136),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_211),
.Y(n_241)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_128),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_117),
.A2(n_31),
.B1(n_1),
.B2(n_3),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_124),
.B(n_11),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_218),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_127),
.B(n_0),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_127),
.B(n_124),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_116),
.B(n_11),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_1),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_122),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_217),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_139),
.B(n_11),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_136),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_219),
.B(n_5),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_220),
.A2(n_207),
.B1(n_176),
.B2(n_203),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_221),
.B(n_237),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_L g312 ( 
.A1(n_226),
.A2(n_263),
.B(n_244),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_190),
.A2(n_154),
.B1(n_148),
.B2(n_118),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_227),
.A2(n_238),
.B1(n_251),
.B2(n_267),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_236),
.A2(n_195),
.B1(n_175),
.B2(n_217),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_190),
.A2(n_154),
.B1(n_147),
.B2(n_134),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_250),
.B(n_266),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_177),
.A2(n_141),
.B1(n_147),
.B2(n_134),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_172),
.A2(n_123),
.B1(n_130),
.B2(n_6),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_167),
.B(n_164),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_180),
.B(n_173),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_260),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_173),
.B(n_130),
.Y(n_260)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_190),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_261),
.Y(n_291)
);

O2A1O1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_167),
.A2(n_4),
.B(n_5),
.C(n_12),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_263),
.Y(n_310)
);

BUFx24_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_269),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_167),
.B(n_214),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_270),
.A2(n_226),
.B(n_237),
.Y(n_316)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_234),
.Y(n_271)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_272),
.A2(n_294),
.B(n_300),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_273),
.A2(n_276),
.B1(n_279),
.B2(n_285),
.Y(n_322)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_222),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_275),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_221),
.A2(n_176),
.B1(n_205),
.B2(n_214),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_277),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_239),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_278),
.B(n_295),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_221),
.A2(n_179),
.B1(n_178),
.B2(n_174),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_238),
.A2(n_210),
.B1(n_186),
.B2(n_193),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_282),
.A2(n_292),
.B1(n_296),
.B2(n_303),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_221),
.A2(n_202),
.B1(n_206),
.B2(n_211),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_283),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_192),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_284),
.B(n_288),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_220),
.A2(n_188),
.B1(n_197),
.B2(n_163),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_227),
.A2(n_185),
.B1(n_199),
.B2(n_200),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_286),
.A2(n_231),
.B1(n_262),
.B2(n_235),
.Y(n_319)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_234),
.Y(n_287)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_287),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_224),
.B(n_162),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_246),
.Y(n_289)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_289),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_224),
.B(n_184),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_290),
.B(n_293),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_267),
.A2(n_171),
.B1(n_194),
.B2(n_166),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_12),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_264),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_233),
.B(n_15),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_229),
.A2(n_16),
.B1(n_17),
.B2(n_268),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_16),
.C(n_17),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_247),
.C(n_258),
.Y(n_318)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_228),
.Y(n_298)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_298),
.Y(n_327)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_228),
.Y(n_299)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_299),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_264),
.A2(n_17),
.B1(n_256),
.B2(n_259),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_256),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_301),
.Y(n_314)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_246),
.Y(n_302)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_302),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_229),
.A2(n_17),
.B1(n_232),
.B2(n_252),
.Y(n_303)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_222),
.Y(n_304)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_304),
.Y(n_343)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_255),
.Y(n_305)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_305),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_260),
.A2(n_245),
.B1(n_230),
.B2(n_237),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_306),
.B(n_225),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_241),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_308),
.B(n_309),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_243),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_223),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_311),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_247),
.Y(n_317)
);

A2O1A1O1Ixp25_ASAP7_75t_L g368 ( 
.A1(n_316),
.A2(n_269),
.B(n_305),
.C(n_302),
.D(n_287),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_317),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_348),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_319),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_274),
.A2(n_242),
.B1(n_235),
.B2(n_231),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_274),
.A2(n_257),
.B1(n_255),
.B2(n_262),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_291),
.A2(n_282),
.B1(n_303),
.B2(n_281),
.Y(n_325)
);

AO22x1_ASAP7_75t_SL g329 ( 
.A1(n_291),
.A2(n_281),
.B1(n_276),
.B2(n_273),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_329),
.B(n_349),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_265),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_330),
.B(n_337),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_281),
.B(n_257),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_334),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_280),
.B(n_265),
.C(n_249),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_336),
.B(n_352),
.C(n_311),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_307),
.B(n_249),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_271),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_340),
.B(n_344),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_278),
.B(n_225),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_342),
.B(n_248),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_301),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_345),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_306),
.B(n_248),
.Y(n_348)
);

MAJx2_ASAP7_75t_L g351 ( 
.A(n_280),
.B(n_248),
.C(n_254),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_351),
.B(n_318),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_293),
.B(n_240),
.C(n_254),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_313),
.Y(n_354)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_354),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_341),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_355),
.B(n_357),
.Y(n_411)
);

AND2x6_ASAP7_75t_L g357 ( 
.A(n_329),
.B(n_279),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_360),
.B(n_368),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_284),
.Y(n_361)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_361),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_335),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_362),
.B(n_343),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_322),
.A2(n_270),
.B1(n_292),
.B2(n_296),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_363),
.A2(n_366),
.B1(n_377),
.B2(n_345),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_323),
.A2(n_286),
.B1(n_272),
.B2(n_285),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_364),
.A2(n_365),
.B1(n_382),
.B2(n_343),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_325),
.A2(n_310),
.B1(n_308),
.B2(n_290),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_322),
.A2(n_310),
.B1(n_288),
.B2(n_297),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_367),
.Y(n_389)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_313),
.Y(n_369)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_369),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_328),
.B(n_289),
.Y(n_371)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_371),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_333),
.B(n_269),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_372),
.B(n_373),
.C(n_352),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_269),
.C(n_240),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_350),
.A2(n_275),
.B(n_298),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_374),
.A2(n_384),
.B(n_331),
.Y(n_396)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_327),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_375),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_350),
.A2(n_304),
.B(n_299),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_376),
.A2(n_379),
.B(n_380),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_349),
.A2(n_329),
.B1(n_336),
.B2(n_333),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_344),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_378),
.B(n_347),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_334),
.A2(n_316),
.B(n_351),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_324),
.A2(n_315),
.B1(n_334),
.B2(n_346),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_383),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_346),
.A2(n_331),
.B(n_339),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_385),
.B(n_317),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_378),
.B(n_337),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_388),
.B(n_397),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_380),
.B(n_315),
.Y(n_390)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_390),
.Y(n_415)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_391),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_393),
.A2(n_379),
.B(n_376),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_395),
.B(n_399),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_396),
.A2(n_413),
.B(n_388),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_359),
.A2(n_339),
.B1(n_347),
.B2(n_320),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_371),
.B(n_338),
.Y(n_398)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_398),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_359),
.A2(n_338),
.B1(n_320),
.B2(n_326),
.Y(n_400)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_400),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_361),
.B(n_326),
.Y(n_401)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_401),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_327),
.C(n_332),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_402),
.B(n_404),
.C(n_373),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_355),
.B(n_314),
.Y(n_403)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_403),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_358),
.B(n_332),
.C(n_314),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_405),
.A2(n_414),
.B1(n_368),
.B2(n_354),
.Y(n_425)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_406),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_409),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_353),
.B(n_321),
.Y(n_410)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_410),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_370),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_382),
.A2(n_321),
.B1(n_365),
.B2(n_364),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_416),
.B(n_419),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_417),
.B(n_421),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_402),
.B(n_360),
.C(n_358),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_420),
.C(n_429),
.Y(n_447)
);

OA21x2_ASAP7_75t_L g419 ( 
.A1(n_411),
.A2(n_356),
.B(n_357),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_372),
.C(n_381),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_395),
.B(n_387),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_411),
.A2(n_356),
.B1(n_377),
.B2(n_381),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_422),
.A2(n_424),
.B1(n_425),
.B2(n_414),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_390),
.A2(n_363),
.B1(n_366),
.B2(n_384),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_387),
.B(n_374),
.C(n_369),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_399),
.B(n_375),
.C(n_370),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_435),
.B(n_403),
.C(n_391),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_437),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_396),
.A2(n_393),
.B(n_390),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_413),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_415),
.A2(n_405),
.B1(n_408),
.B2(n_389),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_440),
.A2(n_444),
.B1(n_428),
.B2(n_422),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_433),
.B(n_406),
.Y(n_441)
);

CKINVDCx14_ASAP7_75t_R g462 ( 
.A(n_441),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_442),
.A2(n_430),
.B(n_426),
.Y(n_468)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_433),
.Y(n_443)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_443),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_415),
.A2(n_408),
.B1(n_389),
.B2(n_394),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_446),
.A2(n_434),
.B1(n_432),
.B2(n_427),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_450),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_436),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_452),
.Y(n_459)
);

MAJx2_ASAP7_75t_L g450 ( 
.A(n_420),
.B(n_394),
.C(n_398),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_436),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_423),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_453),
.B(n_457),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_417),
.B(n_418),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_456),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_432),
.A2(n_392),
.B1(n_413),
.B2(n_410),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_455),
.B(n_424),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_435),
.B(n_409),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_431),
.B(n_397),
.C(n_400),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_425),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_458),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_460),
.A2(n_448),
.B1(n_412),
.B2(n_421),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_456),
.B(n_431),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_461),
.B(n_463),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_SL g464 ( 
.A1(n_439),
.A2(n_413),
.B1(n_423),
.B2(n_430),
.Y(n_464)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_464),
.Y(n_477)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_468),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_442),
.B(n_444),
.Y(n_469)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_469),
.Y(n_485)
);

OAI221xp5_ASAP7_75t_L g470 ( 
.A1(n_450),
.A2(n_426),
.B1(n_428),
.B2(n_438),
.C(n_416),
.Y(n_470)
);

AOI31xp33_ASAP7_75t_L g482 ( 
.A1(n_470),
.A2(n_451),
.A3(n_437),
.B(n_468),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_473),
.A2(n_446),
.B1(n_434),
.B2(n_427),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_429),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_474),
.B(n_447),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_466),
.B(n_419),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_479),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_471),
.B(n_454),
.C(n_445),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_478),
.B(n_481),
.Y(n_490)
);

FAx1_ASAP7_75t_SL g479 ( 
.A(n_473),
.B(n_451),
.CI(n_440),
.CON(n_479),
.SN(n_479)
);

NOR3xp33_ASAP7_75t_L g480 ( 
.A(n_462),
.B(n_419),
.C(n_451),
.Y(n_480)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_480),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_482),
.A2(n_472),
.B1(n_467),
.B2(n_465),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_483),
.B(n_486),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_463),
.A2(n_401),
.B1(n_447),
.B2(n_412),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_487),
.B(n_469),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_476),
.B(n_471),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_491),
.B(n_492),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_487),
.B(n_459),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_493),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_494),
.A2(n_496),
.B(n_486),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_466),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_490),
.B(n_478),
.C(n_483),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_498),
.A2(n_501),
.B(n_491),
.Y(n_504)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_489),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_499),
.A2(n_477),
.B1(n_412),
.B2(n_407),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_500),
.B(n_488),
.C(n_474),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_495),
.A2(n_484),
.B(n_485),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_503),
.B(n_504),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_497),
.A2(n_488),
.B(n_496),
.Y(n_505)
);

AOI31xp33_ASAP7_75t_L g508 ( 
.A1(n_505),
.A2(n_506),
.A3(n_502),
.B(n_479),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_507),
.C(n_479),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_509),
.A2(n_386),
.B(n_407),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_510),
.B(n_386),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_511),
.B(n_481),
.C(n_445),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_512),
.B(n_461),
.Y(n_513)
);


endmodule