module fake_jpeg_29492_n_93 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_93);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_93;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_42),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_45),
.B1(n_46),
.B2(n_7),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_44),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_1),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_43),
.B(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_54),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_52),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_32),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_18),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_36),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_37),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_12),
.C(n_16),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_8),
.B1(n_30),
.B2(n_15),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_7),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_69),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_37),
.B1(n_30),
.B2(n_8),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_62),
.B1(n_64),
.B2(n_24),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_37),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_65),
.C(n_68),
.Y(n_74)
);

OAI22x1_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_30),
.B1(n_9),
.B2(n_10),
.Y(n_62)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_25),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_53),
.B(n_22),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_23),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_76),
.B(n_81),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_79),
.B(n_80),
.Y(n_85)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_85),
.A2(n_62),
.B1(n_79),
.B2(n_58),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_87),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_84),
.A2(n_79),
.B1(n_67),
.B2(n_71),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_82),
.C(n_75),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_63),
.B1(n_74),
.B2(n_83),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_49),
.B(n_27),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_28),
.Y(n_93)
);


endmodule