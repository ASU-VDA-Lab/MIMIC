module fake_jpeg_23188_n_134 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_11),
.B(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_4),
.B(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_31),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_28),
.Y(n_31)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_34),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_23),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_34),
.Y(n_57)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_37),
.B1(n_32),
.B2(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_33),
.Y(n_54)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_32),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_31),
.A2(n_23),
.B1(n_14),
.B2(n_17),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_47),
.A2(n_22),
.B1(n_15),
.B2(n_19),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_14),
.B1(n_32),
.B2(n_31),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_53),
.Y(n_83)
);

AO22x2_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_30),
.B1(n_33),
.B2(n_23),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_22),
.B(n_49),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_SL g80 ( 
.A1(n_52),
.A2(n_69),
.B(n_70),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_23),
.B(n_30),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_56),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_55)
);

AO21x1_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_49),
.B(n_27),
.Y(n_75)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_1),
.Y(n_79)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_59),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_29),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_68),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_45),
.B1(n_39),
.B2(n_48),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_67),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_35),
.B(n_27),
.C(n_25),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_63),
.B(n_21),
.Y(n_85)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_46),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_17),
.B1(n_26),
.B2(n_16),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_17),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_19),
.B1(n_26),
.B2(n_16),
.Y(n_69)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_2),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_80),
.B1(n_62),
.B2(n_51),
.Y(n_87)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_67),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_15),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_78),
.B(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_79),
.B(n_86),
.Y(n_93)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_10),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_9),
.B(n_12),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_18),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_97),
.B(n_85),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_51),
.B1(n_55),
.B2(n_57),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_95),
.C(n_99),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_51),
.B1(n_50),
.B2(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_92),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_61),
.B1(n_25),
.B2(n_20),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_79),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_20),
.B1(n_18),
.B2(n_5),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_108),
.B(n_99),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_106),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_72),
.C(n_83),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_107),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_81),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_76),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_84),
.B(n_79),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_98),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_89),
.B1(n_96),
.B2(n_75),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_114),
.B(n_109),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_90),
.C(n_87),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_116),
.B(n_101),
.Y(n_121)
);

XOR2x2_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_105),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_121),
.B(n_101),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_91),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_123),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_113),
.B(n_73),
.C(n_86),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_126),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_77),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_10),
.A3(n_11),
.B1(n_5),
.B2(n_7),
.C1(n_2),
.C2(n_3),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_8),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_3),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_132),
.B1(n_127),
.B2(n_128),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_133),
.B(n_3),
.Y(n_134)
);


endmodule