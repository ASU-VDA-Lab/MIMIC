module fake_aes_745_n_1567 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_236, n_340, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_32, n_235, n_243, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_343, n_127, n_291, n_170, n_281, n_341, n_58, n_122, n_187, n_138, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_350, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1567, n_824);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_236;
input n_340;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_32;
input n_235;
input n_243;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_343;
input n_127;
input n_291;
input n_170;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_350;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1567;
output n_824;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1477;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_641;
wire n_379;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_822;
wire n_706;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_815;
wire n_477;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1533;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_1563;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_1557;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_799;
wire n_423;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_606;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_400;
wire n_1455;
wire n_386;
wire n_432;
wire n_1329;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_584;
wire n_1130;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1489;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_458;
wire n_1084;
wire n_618;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_401;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_1518;
wire n_945;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1491;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_374;
wire n_718;
wire n_1484;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_1531;
wire n_371;
wire n_1548;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_63), .Y(n_355) );
INVx1_ASAP7_75t_SL g356 ( .A(n_302), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_19), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_129), .Y(n_358) );
INVxp67_ASAP7_75t_SL g359 ( .A(n_60), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_60), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_42), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_42), .Y(n_362) );
INVxp33_ASAP7_75t_SL g363 ( .A(n_241), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_80), .Y(n_364) );
INVxp33_ASAP7_75t_L g365 ( .A(n_289), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_23), .Y(n_366) );
BUFx3_ASAP7_75t_L g367 ( .A(n_349), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_48), .Y(n_368) );
CKINVDCx16_ASAP7_75t_R g369 ( .A(n_53), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_222), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_172), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_152), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_335), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_321), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_246), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_270), .Y(n_376) );
INVxp33_ASAP7_75t_L g377 ( .A(n_233), .Y(n_377) );
NOR2xp67_ASAP7_75t_L g378 ( .A(n_187), .B(n_101), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_171), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_44), .Y(n_380) );
INVxp67_ASAP7_75t_SL g381 ( .A(n_165), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_210), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_122), .Y(n_383) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_50), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_97), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_155), .Y(n_386) );
INVxp33_ASAP7_75t_SL g387 ( .A(n_193), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_337), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_177), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_135), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_164), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_309), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_296), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_167), .Y(n_394) );
BUFx3_ASAP7_75t_L g395 ( .A(n_31), .Y(n_395) );
INVx4_ASAP7_75t_R g396 ( .A(n_91), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_71), .Y(n_397) );
CKINVDCx16_ASAP7_75t_R g398 ( .A(n_146), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_313), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_95), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_119), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_64), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_170), .Y(n_403) );
CKINVDCx14_ASAP7_75t_R g404 ( .A(n_297), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_33), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_342), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_332), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_127), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_347), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_245), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_200), .Y(n_411) );
INVxp33_ASAP7_75t_L g412 ( .A(n_224), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_66), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_71), .Y(n_414) );
INVx2_ASAP7_75t_SL g415 ( .A(n_35), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_242), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_350), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_261), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_253), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_315), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_304), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_29), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_267), .Y(n_423) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_318), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_129), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_314), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_65), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_41), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_228), .Y(n_429) );
INVxp33_ASAP7_75t_L g430 ( .A(n_243), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_59), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_21), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_190), .Y(n_433) );
INVxp67_ASAP7_75t_SL g434 ( .A(n_119), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_303), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_26), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_182), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_87), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_301), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_131), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_275), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_48), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_126), .Y(n_443) );
CKINVDCx16_ASAP7_75t_R g444 ( .A(n_338), .Y(n_444) );
BUFx5_ASAP7_75t_L g445 ( .A(n_34), .Y(n_445) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_263), .Y(n_446) );
INVxp67_ASAP7_75t_SL g447 ( .A(n_56), .Y(n_447) );
BUFx5_ASAP7_75t_L g448 ( .A(n_197), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_54), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_147), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_310), .Y(n_451) );
INVxp67_ASAP7_75t_L g452 ( .A(n_185), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_49), .Y(n_453) );
CKINVDCx14_ASAP7_75t_R g454 ( .A(n_28), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_51), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_331), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_126), .Y(n_457) );
INVxp33_ASAP7_75t_L g458 ( .A(n_227), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_6), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_305), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_96), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_238), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_74), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_260), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_176), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_68), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_108), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_62), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_323), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_295), .Y(n_470) );
INVxp67_ASAP7_75t_SL g471 ( .A(n_7), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_95), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_325), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_199), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_205), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_192), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_175), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_76), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_217), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_20), .Y(n_480) );
INVxp67_ASAP7_75t_SL g481 ( .A(n_15), .Y(n_481) );
INVxp67_ASAP7_75t_SL g482 ( .A(n_278), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_239), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_85), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_319), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_265), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_183), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_68), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_271), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_268), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_87), .Y(n_491) );
INVxp67_ASAP7_75t_SL g492 ( .A(n_237), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_47), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_336), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_249), .Y(n_495) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_279), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_78), .Y(n_497) );
NOR2xp67_ASAP7_75t_L g498 ( .A(n_206), .B(n_194), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_346), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_215), .Y(n_500) );
INVxp67_ASAP7_75t_SL g501 ( .A(n_308), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_294), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g503 ( .A(n_67), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_84), .Y(n_504) );
NOR2xp67_ASAP7_75t_L g505 ( .A(n_39), .B(n_353), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_254), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_339), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_124), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_135), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_320), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g511 ( .A(n_50), .Y(n_511) );
CKINVDCx16_ASAP7_75t_R g512 ( .A(n_157), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_311), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_120), .Y(n_514) );
BUFx2_ASAP7_75t_L g515 ( .A(n_284), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_272), .Y(n_516) );
INVxp67_ASAP7_75t_L g517 ( .A(n_103), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_280), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_30), .B(n_154), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_273), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_144), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_257), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_139), .Y(n_523) );
INVxp67_ASAP7_75t_SL g524 ( .A(n_12), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_39), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_15), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_44), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_142), .Y(n_528) );
NOR2xp67_ASAP7_75t_L g529 ( .A(n_94), .B(n_45), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_448), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_454), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_398), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_445), .Y(n_533) );
INVx3_ASAP7_75t_L g534 ( .A(n_448), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_515), .B(n_0), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_445), .Y(n_536) );
NAND2xp33_ASAP7_75t_SL g537 ( .A(n_365), .B(n_0), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_448), .Y(n_538) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_371), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_515), .B(n_1), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_367), .Y(n_541) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_371), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_445), .Y(n_543) );
INVx3_ASAP7_75t_L g544 ( .A(n_448), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_448), .Y(n_545) );
AND2x6_ASAP7_75t_L g546 ( .A(n_384), .B(n_143), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_448), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_445), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_362), .B(n_1), .Y(n_549) );
BUFx3_ASAP7_75t_L g550 ( .A(n_367), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_445), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_395), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_445), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_445), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_448), .Y(n_555) );
BUFx2_ASAP7_75t_L g556 ( .A(n_395), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_415), .B(n_2), .Y(n_557) );
INVx5_ASAP7_75t_L g558 ( .A(n_386), .Y(n_558) );
BUFx2_ASAP7_75t_L g559 ( .A(n_404), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_377), .B(n_2), .Y(n_560) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_386), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_415), .B(n_3), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_392), .B(n_3), .Y(n_563) );
AND2x4_ASAP7_75t_L g564 ( .A(n_392), .B(n_4), .Y(n_564) );
INVx2_ASAP7_75t_SL g565 ( .A(n_374), .Y(n_565) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_355), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_445), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_412), .B(n_4), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_382), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_530), .Y(n_570) );
INVx3_ASAP7_75t_L g571 ( .A(n_563), .Y(n_571) );
INVxp67_ASAP7_75t_SL g572 ( .A(n_552), .Y(n_572) );
AO22x2_ASAP7_75t_L g573 ( .A1(n_563), .A2(n_388), .B1(n_389), .B2(n_382), .Y(n_573) );
INVx4_ASAP7_75t_L g574 ( .A(n_530), .Y(n_574) );
AO22x2_ASAP7_75t_L g575 ( .A1(n_563), .A2(n_389), .B1(n_393), .B2(n_388), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_559), .B(n_444), .Y(n_576) );
INVx2_ASAP7_75t_SL g577 ( .A(n_559), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_559), .B(n_496), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_559), .B(n_512), .Y(n_579) );
INVx5_ASAP7_75t_L g580 ( .A(n_546), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_569), .B(n_394), .C(n_393), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_532), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_566), .A2(n_503), .B1(n_511), .B2(n_369), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_530), .Y(n_584) );
AND2x4_ASAP7_75t_L g585 ( .A(n_556), .B(n_390), .Y(n_585) );
AO22x2_ASAP7_75t_L g586 ( .A1(n_563), .A2(n_399), .B1(n_403), .B2(n_394), .Y(n_586) );
AND2x6_ASAP7_75t_L g587 ( .A(n_535), .B(n_399), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_532), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_531), .B(n_500), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_556), .B(n_390), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_556), .B(n_469), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_539), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_531), .B(n_500), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_552), .B(n_430), .Y(n_594) );
AND2x4_ASAP7_75t_SL g595 ( .A(n_535), .B(n_560), .Y(n_595) );
AO22x2_ASAP7_75t_L g596 ( .A1(n_563), .A2(n_406), .B1(n_407), .B2(n_403), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_530), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_539), .Y(n_598) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_539), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_530), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_566), .B(n_458), .Y(n_601) );
CKINVDCx8_ASAP7_75t_R g602 ( .A(n_563), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_560), .B(n_355), .Y(n_603) );
BUFx3_ASAP7_75t_L g604 ( .A(n_550), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_539), .Y(n_605) );
BUFx3_ASAP7_75t_L g606 ( .A(n_550), .Y(n_606) );
NAND2x1p5_ASAP7_75t_L g607 ( .A(n_563), .B(n_406), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_530), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_530), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_534), .Y(n_610) );
INVx3_ASAP7_75t_L g611 ( .A(n_564), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_534), .Y(n_612) );
AND2x4_ASAP7_75t_L g613 ( .A(n_535), .B(n_414), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_534), .Y(n_614) );
AND2x4_ASAP7_75t_L g615 ( .A(n_535), .B(n_414), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_534), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_571), .Y(n_617) );
AND2x6_ASAP7_75t_L g618 ( .A(n_571), .B(n_564), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_594), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_601), .B(n_549), .Y(n_620) );
INVx3_ASAP7_75t_L g621 ( .A(n_571), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_571), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_583), .B(n_549), .Y(n_623) );
AND2x4_ASAP7_75t_L g624 ( .A(n_595), .B(n_549), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_595), .Y(n_625) );
INVx3_ASAP7_75t_L g626 ( .A(n_611), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_595), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_594), .B(n_560), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_613), .B(n_560), .Y(n_629) );
INVx1_ASAP7_75t_SL g630 ( .A(n_576), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_611), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_607), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_607), .Y(n_633) );
BUFx4f_ASAP7_75t_L g634 ( .A(n_587), .Y(n_634) );
INVx2_ASAP7_75t_SL g635 ( .A(n_607), .Y(n_635) );
AOI22xp33_ASAP7_75t_SL g636 ( .A1(n_587), .A2(n_408), .B1(n_431), .B2(n_383), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_611), .Y(n_637) );
AOI22xp5_ASAP7_75t_SL g638 ( .A1(n_582), .A2(n_408), .B1(n_431), .B2(n_383), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_602), .B(n_564), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_611), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_587), .A2(n_568), .B1(n_549), .B2(n_537), .Y(n_641) );
INVx6_ASAP7_75t_L g642 ( .A(n_585), .Y(n_642) );
NAND2x1p5_ASAP7_75t_L g643 ( .A(n_580), .B(n_564), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_585), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_613), .B(n_568), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_585), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_585), .Y(n_647) );
INVx6_ASAP7_75t_L g648 ( .A(n_590), .Y(n_648) );
AND2x4_ASAP7_75t_L g649 ( .A(n_613), .B(n_568), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_604), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_613), .B(n_568), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_604), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_577), .Y(n_653) );
OAI21xp5_ASAP7_75t_L g654 ( .A1(n_570), .A2(n_536), .B(n_533), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_615), .B(n_569), .Y(n_655) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_604), .Y(n_656) );
INVx5_ASAP7_75t_L g657 ( .A(n_574), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_590), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_615), .B(n_569), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_590), .Y(n_660) );
INVx5_ASAP7_75t_L g661 ( .A(n_574), .Y(n_661) );
BUFx12f_ASAP7_75t_L g662 ( .A(n_588), .Y(n_662) );
AND2x4_ASAP7_75t_L g663 ( .A(n_615), .B(n_540), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_615), .B(n_564), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_587), .A2(n_564), .B1(n_537), .B2(n_540), .Y(n_665) );
BUFx2_ASAP7_75t_L g666 ( .A(n_587), .Y(n_666) );
BUFx3_ASAP7_75t_L g667 ( .A(n_606), .Y(n_667) );
BUFx6f_ASAP7_75t_L g668 ( .A(n_606), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_606), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_590), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_592), .Y(n_671) );
INVx2_ASAP7_75t_SL g672 ( .A(n_577), .Y(n_672) );
OR2x6_ASAP7_75t_L g673 ( .A(n_575), .B(n_557), .Y(n_673) );
INVxp67_ASAP7_75t_SL g674 ( .A(n_574), .Y(n_674) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_599), .Y(n_675) );
AND2x4_ASAP7_75t_L g676 ( .A(n_587), .B(n_564), .Y(n_676) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_599), .Y(n_677) );
OR2x2_ASAP7_75t_L g678 ( .A(n_603), .B(n_572), .Y(n_678) );
INVx3_ASAP7_75t_L g679 ( .A(n_602), .Y(n_679) );
BUFx12f_ASAP7_75t_L g680 ( .A(n_587), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g681 ( .A(n_578), .B(n_562), .C(n_557), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_575), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_592), .Y(n_683) );
AND2x4_ASAP7_75t_L g684 ( .A(n_579), .B(n_557), .Y(n_684) );
BUFx3_ASAP7_75t_L g685 ( .A(n_574), .Y(n_685) );
INVxp33_ASAP7_75t_SL g686 ( .A(n_591), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_573), .B(n_562), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_573), .B(n_562), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_575), .Y(n_689) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_575), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_573), .B(n_550), .Y(n_691) );
NAND2x1p5_ASAP7_75t_L g692 ( .A(n_580), .B(n_534), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_589), .B(n_363), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_575), .Y(n_694) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_573), .Y(n_695) );
INVx2_ASAP7_75t_SL g696 ( .A(n_586), .Y(n_696) );
OR2x4_ASAP7_75t_L g697 ( .A(n_593), .B(n_364), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_592), .Y(n_698) );
BUFx8_ASAP7_75t_L g699 ( .A(n_586), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_570), .B(n_533), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_598), .Y(n_701) );
INVx2_ASAP7_75t_SL g702 ( .A(n_586), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_586), .B(n_550), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_584), .B(n_533), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_596), .B(n_358), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_598), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_596), .Y(n_707) );
NOR2xp67_ASAP7_75t_L g708 ( .A(n_581), .B(n_534), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_673), .A2(n_596), .B1(n_581), .B2(n_451), .Y(n_709) );
BUFx3_ASAP7_75t_L g710 ( .A(n_662), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_673), .A2(n_596), .B1(n_451), .B2(n_474), .Y(n_711) );
INVx3_ASAP7_75t_L g712 ( .A(n_680), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_621), .Y(n_713) );
INVx5_ASAP7_75t_L g714 ( .A(n_680), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_621), .Y(n_715) );
INVx5_ASAP7_75t_L g716 ( .A(n_673), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_621), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_619), .B(n_449), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_673), .A2(n_473), .B1(n_486), .B2(n_474), .Y(n_719) );
BUFx10_ASAP7_75t_L g720 ( .A(n_697), .Y(n_720) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_662), .Y(n_721) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_635), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_620), .B(n_449), .Y(n_723) );
OR2x6_ASAP7_75t_L g724 ( .A(n_635), .B(n_529), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_638), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_642), .Y(n_726) );
INVx4_ASAP7_75t_L g727 ( .A(n_634), .Y(n_727) );
AND2x4_ASAP7_75t_L g728 ( .A(n_624), .B(n_359), .Y(n_728) );
BUFx3_ASAP7_75t_L g729 ( .A(n_699), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_682), .A2(n_538), .B1(n_547), .B2(n_545), .Y(n_730) );
INVxp67_ASAP7_75t_L g731 ( .A(n_653), .Y(n_731) );
NAND2xp33_ASAP7_75t_L g732 ( .A(n_696), .B(n_546), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_626), .Y(n_733) );
NOR2xp33_ASAP7_75t_R g734 ( .A(n_699), .B(n_473), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_642), .Y(n_735) );
BUFx6f_ASAP7_75t_L g736 ( .A(n_634), .Y(n_736) );
INVx2_ASAP7_75t_SL g737 ( .A(n_697), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_626), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_642), .Y(n_739) );
AND2x4_ASAP7_75t_L g740 ( .A(n_624), .B(n_434), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_689), .A2(n_538), .B1(n_547), .B2(n_545), .Y(n_741) );
BUFx10_ASAP7_75t_L g742 ( .A(n_684), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_626), .Y(n_743) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_699), .Y(n_744) );
INVx3_ASAP7_75t_L g745 ( .A(n_657), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_642), .Y(n_746) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_636), .A2(n_686), .B1(n_623), .B2(n_630), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_686), .A2(n_490), .B1(n_486), .B2(n_360), .Y(n_748) );
BUFx2_ASAP7_75t_L g749 ( .A(n_624), .Y(n_749) );
AOI22x1_ASAP7_75t_L g750 ( .A1(n_617), .A2(n_541), .B1(n_565), .B2(n_598), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_648), .Y(n_751) );
OR2x2_ASAP7_75t_L g752 ( .A(n_620), .B(n_358), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_648), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_694), .A2(n_538), .B1(n_547), .B2(n_545), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_705), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_649), .B(n_584), .Y(n_756) );
BUFx2_ASAP7_75t_L g757 ( .A(n_690), .Y(n_757) );
OR2x2_ASAP7_75t_L g758 ( .A(n_623), .B(n_360), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_649), .B(n_597), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_617), .Y(n_760) );
INVx3_ASAP7_75t_L g761 ( .A(n_657), .Y(n_761) );
AOI21xp5_ASAP7_75t_SL g762 ( .A1(n_696), .A2(n_550), .B(n_424), .Y(n_762) );
BUFx6f_ASAP7_75t_L g763 ( .A(n_634), .Y(n_763) );
BUFx6f_ASAP7_75t_L g764 ( .A(n_632), .Y(n_764) );
INVxp67_ASAP7_75t_SL g765 ( .A(n_695), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_622), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_649), .B(n_597), .Y(n_767) );
AOI21xp5_ASAP7_75t_L g768 ( .A1(n_700), .A2(n_608), .B(n_600), .Y(n_768) );
BUFx2_ASAP7_75t_L g769 ( .A(n_633), .Y(n_769) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_702), .Y(n_770) );
CKINVDCx5p33_ASAP7_75t_R g771 ( .A(n_705), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_648), .Y(n_772) );
BUFx6f_ASAP7_75t_L g773 ( .A(n_657), .Y(n_773) );
INVx2_ASAP7_75t_SL g774 ( .A(n_678), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_702), .A2(n_490), .B1(n_443), .B2(n_463), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_641), .A2(n_443), .B1(n_463), .B2(n_427), .Y(n_776) );
AND2x4_ASAP7_75t_L g777 ( .A(n_625), .B(n_447), .Y(n_777) );
BUFx6f_ASAP7_75t_L g778 ( .A(n_657), .Y(n_778) );
BUFx6f_ASAP7_75t_L g779 ( .A(n_657), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_684), .B(n_600), .Y(n_780) );
AND2x4_ASAP7_75t_L g781 ( .A(n_627), .B(n_471), .Y(n_781) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_676), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_707), .A2(n_538), .B1(n_547), .B2(n_545), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_648), .Y(n_784) );
BUFx6f_ASAP7_75t_L g785 ( .A(n_661), .Y(n_785) );
INVx6_ASAP7_75t_L g786 ( .A(n_656), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_622), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_687), .A2(n_357), .B1(n_380), .B2(n_361), .Y(n_788) );
AND2x4_ASAP7_75t_L g789 ( .A(n_684), .B(n_481), .Y(n_789) );
O2A1O1Ixp33_ASAP7_75t_L g790 ( .A1(n_628), .A2(n_357), .B(n_380), .C(n_361), .Y(n_790) );
NAND2xp5_ASAP7_75t_SL g791 ( .A(n_661), .B(n_608), .Y(n_791) );
AND2x4_ASAP7_75t_L g792 ( .A(n_663), .B(n_524), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_688), .A2(n_397), .B1(n_400), .B2(n_385), .Y(n_793) );
INVxp67_ASAP7_75t_SL g794 ( .A(n_666), .Y(n_794) );
INVx3_ASAP7_75t_L g795 ( .A(n_661), .Y(n_795) );
BUFx6f_ASAP7_75t_L g796 ( .A(n_661), .Y(n_796) );
INVx2_ASAP7_75t_SL g797 ( .A(n_678), .Y(n_797) );
BUFx2_ASAP7_75t_SL g798 ( .A(n_676), .Y(n_798) );
AND2x2_ASAP7_75t_L g799 ( .A(n_629), .B(n_427), .Y(n_799) );
INVx5_ASAP7_75t_L g800 ( .A(n_666), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_681), .B(n_363), .Y(n_801) );
BUFx2_ASAP7_75t_L g802 ( .A(n_676), .Y(n_802) );
INVx8_ASAP7_75t_L g803 ( .A(n_618), .Y(n_803) );
AND2x4_ASAP7_75t_L g804 ( .A(n_663), .B(n_366), .Y(n_804) );
CKINVDCx8_ASAP7_75t_R g805 ( .A(n_663), .Y(n_805) );
NOR3xp33_ASAP7_75t_L g806 ( .A(n_693), .B(n_517), .C(n_422), .Y(n_806) );
NOR2xp67_ASAP7_75t_SL g807 ( .A(n_661), .B(n_580), .Y(n_807) );
OR2x6_ASAP7_75t_L g808 ( .A(n_672), .B(n_385), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_644), .Y(n_809) );
INVx2_ASAP7_75t_SL g810 ( .A(n_672), .Y(n_810) );
INVx2_ASAP7_75t_SL g811 ( .A(n_655), .Y(n_811) );
NAND3xp33_ASAP7_75t_L g812 ( .A(n_665), .B(n_484), .C(n_466), .Y(n_812) );
INVx3_ASAP7_75t_L g813 ( .A(n_685), .Y(n_813) );
HAxp5_ASAP7_75t_L g814 ( .A(n_645), .B(n_466), .CON(n_814), .SN(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_631), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_646), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_651), .B(n_647), .Y(n_817) );
BUFx3_ASAP7_75t_L g818 ( .A(n_658), .Y(n_818) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_679), .Y(n_819) );
INVx3_ASAP7_75t_L g820 ( .A(n_685), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_631), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_660), .Y(n_822) );
AND2x4_ASAP7_75t_L g823 ( .A(n_670), .B(n_368), .Y(n_823) );
UNKNOWN g824 ( );
INVx1_ASAP7_75t_L g825 ( .A(n_664), .Y(n_825) );
INVx3_ASAP7_75t_L g826 ( .A(n_667), .Y(n_826) );
NAND2xp5_ASAP7_75t_SL g827 ( .A(n_679), .B(n_609), .Y(n_827) );
INVx1_ASAP7_75t_SL g828 ( .A(n_618), .Y(n_828) );
AND2x4_ASAP7_75t_L g829 ( .A(n_679), .B(n_425), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_639), .A2(n_497), .B1(n_523), .B2(n_484), .Y(n_830) );
INVx1_ASAP7_75t_SL g831 ( .A(n_618), .Y(n_831) );
BUFx10_ASAP7_75t_L g832 ( .A(n_618), .Y(n_832) );
INVx5_ASAP7_75t_L g833 ( .A(n_618), .Y(n_833) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_674), .Y(n_834) );
OAI21xp33_ASAP7_75t_L g835 ( .A1(n_639), .A2(n_616), .B(n_610), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_691), .A2(n_397), .B1(n_401), .B2(n_400), .Y(n_836) );
INVx2_ASAP7_75t_SL g837 ( .A(n_618), .Y(n_837) );
OR2x2_ASAP7_75t_L g838 ( .A(n_703), .B(n_497), .Y(n_838) );
OR2x6_ASAP7_75t_L g839 ( .A(n_643), .B(n_401), .Y(n_839) );
INVx3_ASAP7_75t_L g840 ( .A(n_667), .Y(n_840) );
INVx2_ASAP7_75t_SL g841 ( .A(n_643), .Y(n_841) );
INVx2_ASAP7_75t_SL g842 ( .A(n_643), .Y(n_842) );
INVx3_ASAP7_75t_L g843 ( .A(n_656), .Y(n_843) );
AND2x4_ASAP7_75t_L g844 ( .A(n_637), .B(n_428), .Y(n_844) );
INVx4_ASAP7_75t_L g845 ( .A(n_656), .Y(n_845) );
BUFx6f_ASAP7_75t_L g846 ( .A(n_656), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_656), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g848 ( .A1(n_640), .A2(n_527), .B1(n_523), .B2(n_387), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_774), .B(n_527), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_797), .B(n_654), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_773), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_808), .A2(n_387), .B1(n_668), .B2(n_652), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_747), .A2(n_384), .B1(n_436), .B2(n_432), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_709), .A2(n_384), .B1(n_440), .B2(n_438), .Y(n_854) );
OAI21xp5_ASAP7_75t_L g855 ( .A1(n_768), .A2(n_704), .B(n_700), .Y(n_855) );
AND2x4_ASAP7_75t_L g856 ( .A(n_731), .B(n_668), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_773), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_709), .A2(n_384), .B1(n_453), .B2(n_442), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_804), .A2(n_384), .B1(n_457), .B2(n_455), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g860 ( .A1(n_711), .A2(n_708), .B1(n_704), .B2(n_650), .Y(n_860) );
OR2x6_ASAP7_75t_L g861 ( .A(n_803), .B(n_692), .Y(n_861) );
BUFx3_ASAP7_75t_L g862 ( .A(n_710), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_844), .Y(n_863) );
BUFx4f_ASAP7_75t_L g864 ( .A(n_839), .Y(n_864) );
NOR2xp33_ASAP7_75t_L g865 ( .A(n_805), .B(n_650), .Y(n_865) );
AND2x4_ASAP7_75t_L g866 ( .A(n_731), .B(n_668), .Y(n_866) );
AOI21xp5_ASAP7_75t_L g867 ( .A1(n_768), .A2(n_669), .B(n_652), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_723), .B(n_402), .Y(n_868) );
AOI21xp33_ASAP7_75t_L g869 ( .A1(n_801), .A2(n_669), .B(n_668), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_773), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_844), .Y(n_871) );
INVx2_ASAP7_75t_SL g872 ( .A(n_734), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_808), .A2(n_668), .B1(n_565), .B2(n_541), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_823), .Y(n_874) );
CKINVDCx14_ASAP7_75t_R g875 ( .A(n_734), .Y(n_875) );
INVx6_ASAP7_75t_L g876 ( .A(n_714), .Y(n_876) );
INVx2_ASAP7_75t_L g877 ( .A(n_773), .Y(n_877) );
BUFx3_ASAP7_75t_L g878 ( .A(n_721), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_811), .B(n_459), .Y(n_879) );
OR2x6_ASAP7_75t_L g880 ( .A(n_803), .B(n_692), .Y(n_880) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_808), .A2(n_565), .B1(n_541), .B2(n_521), .Y(n_881) );
CKINVDCx20_ASAP7_75t_R g882 ( .A(n_725), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_804), .A2(n_467), .B1(n_468), .B2(n_461), .Y(n_883) );
OAI22xp33_ASAP7_75t_L g884 ( .A1(n_711), .A2(n_405), .B1(n_413), .B2(n_402), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_839), .A2(n_565), .B1(n_541), .B2(n_521), .Y(n_885) );
OR2x2_ASAP7_75t_L g886 ( .A(n_748), .B(n_405), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_823), .Y(n_887) );
OAI22xp33_ASAP7_75t_L g888 ( .A1(n_719), .A2(n_514), .B1(n_526), .B2(n_413), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_799), .B(n_472), .Y(n_889) );
BUFx4f_ASAP7_75t_SL g890 ( .A(n_729), .Y(n_890) );
NOR2xp67_ASAP7_75t_L g891 ( .A(n_719), .B(n_5), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_814), .B(n_514), .Y(n_892) );
BUFx12f_ASAP7_75t_L g893 ( .A(n_720), .Y(n_893) );
AOI21xp5_ASAP7_75t_L g894 ( .A1(n_827), .A2(n_683), .B(n_671), .Y(n_894) );
INVx3_ASAP7_75t_L g895 ( .A(n_778), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_829), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_825), .A2(n_488), .B1(n_491), .B2(n_478), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_829), .Y(n_898) );
NAND2x1p5_ASAP7_75t_L g899 ( .A(n_714), .B(n_580), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g900 ( .A1(n_839), .A2(n_534), .B1(n_544), .B2(n_452), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_769), .B(n_493), .Y(n_901) );
OR2x2_ASAP7_75t_L g902 ( .A(n_752), .B(n_526), .Y(n_902) );
NOR2x1_ASAP7_75t_SL g903 ( .A(n_833), .B(n_580), .Y(n_903) );
BUFx3_ASAP7_75t_L g904 ( .A(n_764), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_817), .B(n_508), .Y(n_905) );
AOI22xp33_ASAP7_75t_SL g906 ( .A1(n_755), .A2(n_480), .B1(n_509), .B2(n_504), .Y(n_906) );
INVx3_ASAP7_75t_L g907 ( .A(n_778), .Y(n_907) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_765), .A2(n_544), .B1(n_381), .B2(n_482), .Y(n_908) );
BUFx6f_ASAP7_75t_L g909 ( .A(n_778), .Y(n_909) );
OR2x2_ASAP7_75t_L g910 ( .A(n_758), .B(n_480), .Y(n_910) );
OAI21x1_ASAP7_75t_L g911 ( .A1(n_750), .A2(n_683), .B(n_671), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_817), .B(n_609), .Y(n_912) );
OAI22xp33_ASAP7_75t_L g913 ( .A1(n_716), .A2(n_509), .B1(n_525), .B2(n_504), .Y(n_913) );
BUFx6f_ASAP7_75t_L g914 ( .A(n_778), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_779), .Y(n_915) );
OAI22xp33_ASAP7_75t_L g916 ( .A1(n_716), .A2(n_771), .B1(n_744), .B2(n_765), .Y(n_916) );
AOI221xp5_ASAP7_75t_L g917 ( .A1(n_806), .A2(n_525), .B1(n_536), .B2(n_548), .C(n_543), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_789), .B(n_610), .Y(n_918) );
HB1xp67_ASAP7_75t_L g919 ( .A(n_834), .Y(n_919) );
AOI21xp5_ASAP7_75t_L g920 ( .A1(n_827), .A2(n_701), .B(n_698), .Y(n_920) );
INVx3_ASAP7_75t_L g921 ( .A(n_779), .Y(n_921) );
AOI21xp5_ASAP7_75t_L g922 ( .A1(n_791), .A2(n_701), .B(n_698), .Y(n_922) );
AOI221xp5_ASAP7_75t_L g923 ( .A1(n_806), .A2(n_548), .B1(n_551), .B2(n_543), .C(n_536), .Y(n_923) );
AND2x2_ASAP7_75t_L g924 ( .A(n_814), .B(n_718), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_789), .B(n_612), .Y(n_925) );
OAI22xp5_ASAP7_75t_SL g926 ( .A1(n_744), .A2(n_492), .B1(n_501), .B2(n_446), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_792), .B(n_612), .Y(n_927) );
AOI22xp5_ASAP7_75t_L g928 ( .A1(n_775), .A2(n_816), .B1(n_728), .B2(n_740), .Y(n_928) );
INVx2_ASAP7_75t_SL g929 ( .A(n_714), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_728), .B(n_544), .Y(n_930) );
AND2x4_ASAP7_75t_L g931 ( .A(n_714), .B(n_378), .Y(n_931) );
INVx1_ASAP7_75t_SL g932 ( .A(n_764), .Y(n_932) );
OAI21xp5_ASAP7_75t_L g933 ( .A1(n_730), .A2(n_616), .B(n_614), .Y(n_933) );
AOI222xp33_ASAP7_75t_L g934 ( .A1(n_824), .A2(n_505), .B1(n_411), .B2(n_410), .C1(n_409), .C2(n_407), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_809), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_792), .B(n_614), .Y(n_936) );
AOI221xp5_ASAP7_75t_L g937 ( .A1(n_790), .A2(n_543), .B1(n_553), .B2(n_551), .C(n_548), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_716), .A2(n_544), .B1(n_539), .B2(n_542), .Y(n_938) );
OAI211xp5_ASAP7_75t_SL g939 ( .A1(n_790), .A2(n_776), .B(n_848), .C(n_830), .Y(n_939) );
AND2x4_ASAP7_75t_L g940 ( .A(n_833), .B(n_409), .Y(n_940) );
INVx2_ASAP7_75t_L g941 ( .A(n_779), .Y(n_941) );
AND2x2_ASAP7_75t_L g942 ( .A(n_740), .B(n_544), .Y(n_942) );
CKINVDCx5p33_ASAP7_75t_R g943 ( .A(n_720), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_822), .Y(n_944) );
O2A1O1Ixp5_ASAP7_75t_L g945 ( .A1(n_788), .A2(n_450), .B(n_502), .C(n_429), .Y(n_945) );
CKINVDCx14_ASAP7_75t_R g946 ( .A(n_724), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_777), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_777), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_716), .A2(n_544), .B1(n_539), .B2(n_542), .Y(n_949) );
AO31x2_ASAP7_75t_L g950 ( .A1(n_788), .A2(n_793), .A3(n_836), .B(n_545), .Y(n_950) );
AO21x2_ASAP7_75t_L g951 ( .A1(n_793), .A2(n_498), .B(n_411), .Y(n_951) );
AOI22xp33_ASAP7_75t_SL g952 ( .A1(n_803), .A2(n_448), .B1(n_391), .B2(n_374), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_749), .A2(n_544), .B1(n_539), .B2(n_542), .Y(n_953) );
BUFx2_ASAP7_75t_L g954 ( .A(n_764), .Y(n_954) );
OR2x6_ASAP7_75t_L g955 ( .A(n_798), .B(n_692), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_781), .Y(n_956) );
AOI221xp5_ASAP7_75t_L g957 ( .A1(n_836), .A2(n_554), .B1(n_567), .B2(n_553), .C(n_551), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_801), .A2(n_539), .B1(n_561), .B2(n_542), .Y(n_958) );
OAI22xp5_ASAP7_75t_L g959 ( .A1(n_794), .A2(n_558), .B1(n_410), .B2(n_513), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_742), .B(n_538), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_812), .A2(n_542), .B1(n_561), .B2(n_539), .Y(n_961) );
OAI22xp5_ASAP7_75t_SL g962 ( .A1(n_737), .A2(n_423), .B1(n_356), .B2(n_519), .Y(n_962) );
AOI21xp5_ASAP7_75t_L g963 ( .A1(n_791), .A2(n_706), .B(n_677), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_838), .A2(n_542), .B1(n_561), .B2(n_539), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_781), .Y(n_965) );
INVx6_ASAP7_75t_L g966 ( .A(n_764), .Y(n_966) );
OAI222xp33_ASAP7_75t_L g967 ( .A1(n_724), .A2(n_528), .B1(n_522), .B2(n_520), .C1(n_516), .C2(n_513), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_818), .Y(n_968) );
OAI22xp33_ASAP7_75t_L g969 ( .A1(n_757), .A2(n_558), .B1(n_555), .B2(n_547), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_802), .A2(n_782), .B1(n_834), .B2(n_742), .Y(n_970) );
OR2x6_ASAP7_75t_L g971 ( .A(n_722), .B(n_510), .Y(n_971) );
INVx2_ASAP7_75t_L g972 ( .A(n_779), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_726), .Y(n_973) );
BUFx2_ASAP7_75t_L g974 ( .A(n_722), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_735), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_739), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_782), .B(n_555), .Y(n_977) );
OAI21x1_ASAP7_75t_L g978 ( .A1(n_843), .A2(n_706), .B(n_605), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_756), .A2(n_561), .B1(n_542), .B2(n_546), .Y(n_979) );
OAI22xp33_ASAP7_75t_L g980 ( .A1(n_794), .A2(n_558), .B1(n_555), .B2(n_510), .Y(n_980) );
INVx5_ASAP7_75t_L g981 ( .A(n_785), .Y(n_981) );
AOI22xp5_ASAP7_75t_L g982 ( .A1(n_819), .A2(n_372), .B1(n_373), .B2(n_370), .Y(n_982) );
AOI21xp5_ASAP7_75t_L g983 ( .A1(n_780), .A2(n_677), .B(n_675), .Y(n_983) );
AND2x4_ASAP7_75t_L g984 ( .A(n_833), .B(n_516), .Y(n_984) );
BUFx2_ASAP7_75t_L g985 ( .A(n_785), .Y(n_985) );
INVx2_ASAP7_75t_L g986 ( .A(n_785), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_780), .B(n_756), .Y(n_987) );
AND2x2_ASAP7_75t_L g988 ( .A(n_746), .B(n_555), .Y(n_988) );
BUFx3_ASAP7_75t_L g989 ( .A(n_785), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_759), .A2(n_561), .B1(n_542), .B2(n_546), .Y(n_990) );
AOI22xp33_ASAP7_75t_SL g991 ( .A1(n_724), .A2(n_391), .B1(n_522), .B2(n_520), .Y(n_991) );
O2A1O1Ixp33_ASAP7_75t_SL g992 ( .A1(n_770), .A2(n_555), .B(n_554), .C(n_553), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_796), .Y(n_993) );
INVx6_ASAP7_75t_L g994 ( .A(n_796), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_751), .Y(n_995) );
AND2x4_ASAP7_75t_L g996 ( .A(n_833), .B(n_528), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_759), .A2(n_561), .B1(n_542), .B2(n_546), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_767), .A2(n_561), .B1(n_542), .B2(n_546), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_753), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_767), .A2(n_561), .B1(n_546), .B2(n_554), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_772), .Y(n_1001) );
INVx2_ASAP7_75t_L g1002 ( .A(n_796), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_784), .B(n_558), .Y(n_1003) );
BUFx10_ASAP7_75t_L g1004 ( .A(n_796), .Y(n_1004) );
INVx1_ASAP7_75t_SL g1005 ( .A(n_841), .Y(n_1005) );
BUFx8_ASAP7_75t_SL g1006 ( .A(n_712), .Y(n_1006) );
INVx1_ASAP7_75t_SL g1007 ( .A(n_842), .Y(n_1007) );
INVx1_ASAP7_75t_SL g1008 ( .A(n_745), .Y(n_1008) );
AND2x4_ASAP7_75t_L g1009 ( .A(n_712), .B(n_580), .Y(n_1009) );
OAI22xp33_ASAP7_75t_L g1010 ( .A1(n_864), .A2(n_810), .B1(n_831), .B2(n_828), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_924), .B(n_819), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_864), .A2(n_837), .B1(n_835), .B2(n_732), .Y(n_1012) );
CKINVDCx5p33_ASAP7_75t_R g1013 ( .A(n_875), .Y(n_1013) );
AOI221xp5_ASAP7_75t_SL g1014 ( .A1(n_884), .A2(n_783), .B1(n_754), .B2(n_741), .C(n_730), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g1015 ( .A1(n_971), .A2(n_770), .B1(n_741), .B2(n_754), .Y(n_1015) );
AOI222xp33_ASAP7_75t_L g1016 ( .A1(n_888), .A2(n_546), .B1(n_375), .B2(n_506), .C1(n_376), .C2(n_421), .Y(n_1016) );
CKINVDCx8_ASAP7_75t_R g1017 ( .A(n_981), .Y(n_1017) );
INVx2_ASAP7_75t_L g1018 ( .A(n_978), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_891), .A2(n_713), .B1(n_717), .B2(n_715), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g1020 ( .A1(n_946), .A2(n_971), .B1(n_872), .B2(n_974), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_919), .Y(n_1021) );
CKINVDCx5p33_ASAP7_75t_R g1022 ( .A(n_890), .Y(n_1022) );
OAI22xp5_ASAP7_75t_SL g1023 ( .A1(n_882), .A2(n_800), .B1(n_727), .B2(n_761), .Y(n_1023) );
NOR2xp33_ASAP7_75t_L g1024 ( .A(n_928), .B(n_745), .Y(n_1024) );
INVx6_ASAP7_75t_L g1025 ( .A(n_1004), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_884), .A2(n_738), .B1(n_743), .B2(n_733), .Y(n_1026) );
OR2x2_ASAP7_75t_L g1027 ( .A(n_919), .B(n_845), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_939), .A2(n_800), .B1(n_832), .B2(n_820), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_939), .A2(n_800), .B1(n_832), .B2(n_820), .Y(n_1029) );
AOI21x1_ASAP7_75t_L g1030 ( .A1(n_983), .A2(n_847), .B(n_605), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_935), .Y(n_1031) );
A2O1A1Ixp33_ASAP7_75t_L g1032 ( .A1(n_854), .A2(n_760), .B(n_787), .C(n_766), .Y(n_1032) );
AOI22xp33_ASAP7_75t_SL g1033 ( .A1(n_971), .A2(n_800), .B1(n_795), .B2(n_761), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_906), .A2(n_853), .B1(n_892), .B2(n_888), .Y(n_1034) );
INVx2_ASAP7_75t_L g1035 ( .A(n_909), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_906), .A2(n_813), .B1(n_795), .B2(n_826), .Y(n_1036) );
AOI211xp5_ASAP7_75t_L g1037 ( .A1(n_962), .A2(n_416), .B(n_417), .C(n_379), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_853), .A2(n_813), .B1(n_840), .B2(n_826), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_854), .A2(n_783), .B1(n_840), .B2(n_821), .Y(n_1039) );
AOI22xp5_ASAP7_75t_SL g1040 ( .A1(n_943), .A2(n_546), .B1(n_727), .B2(n_418), .Y(n_1040) );
OAI221xp5_ASAP7_75t_L g1041 ( .A1(n_883), .A2(n_762), .B1(n_815), .B2(n_420), .C(n_433), .Y(n_1041) );
AOI21xp5_ASAP7_75t_L g1042 ( .A1(n_963), .A2(n_846), .B(n_843), .Y(n_1042) );
AOI221xp5_ASAP7_75t_L g1043 ( .A1(n_868), .A2(n_567), .B1(n_561), .B2(n_426), .C(n_437), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_858), .A2(n_845), .B1(n_736), .B2(n_763), .Y(n_1044) );
OA21x2_ASAP7_75t_L g1045 ( .A1(n_945), .A2(n_605), .B(n_450), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_858), .A2(n_736), .B1(n_763), .B2(n_786), .Y(n_1046) );
OAI21xp33_ASAP7_75t_L g1047 ( .A1(n_991), .A2(n_567), .B(n_502), .Y(n_1047) );
INVx2_ASAP7_75t_L g1048 ( .A(n_909), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_987), .A2(n_786), .B1(n_846), .B2(n_736), .Y(n_1049) );
CKINVDCx20_ASAP7_75t_R g1050 ( .A(n_890), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_897), .B(n_786), .Y(n_1051) );
AOI22xp33_ASAP7_75t_SL g1052 ( .A1(n_881), .A2(n_736), .B1(n_763), .B2(n_846), .Y(n_1052) );
AOI21xp33_ASAP7_75t_L g1053 ( .A1(n_916), .A2(n_846), .B(n_763), .Y(n_1053) );
AOI22xp33_ASAP7_75t_SL g1054 ( .A1(n_852), .A2(n_546), .B1(n_558), .B2(n_419), .Y(n_1054) );
OAI22xp5_ASAP7_75t_L g1055 ( .A1(n_850), .A2(n_558), .B1(n_439), .B2(n_441), .Y(n_1055) );
AOI222xp33_ASAP7_75t_L g1056 ( .A1(n_889), .A2(n_546), .B1(n_483), .B2(n_435), .C1(n_479), .C2(n_456), .Y(n_1056) );
INVxp67_ASAP7_75t_L g1057 ( .A(n_849), .Y(n_1057) );
INVx1_ASAP7_75t_SL g1058 ( .A(n_862), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_950), .B(n_558), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_991), .A2(n_546), .B1(n_462), .B2(n_464), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_944), .Y(n_1061) );
OAI211xp5_ASAP7_75t_L g1062 ( .A1(n_934), .A2(n_465), .B(n_470), .C(n_460), .Y(n_1062) );
NOR2xp33_ASAP7_75t_L g1063 ( .A(n_886), .B(n_475), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_947), .Y(n_1064) );
OAI21xp5_ASAP7_75t_L g1065 ( .A1(n_945), .A2(n_807), .B(n_477), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_917), .A2(n_546), .B1(n_485), .B2(n_487), .Y(n_1066) );
OAI222xp33_ASAP7_75t_L g1067 ( .A1(n_916), .A2(n_495), .B1(n_507), .B2(n_476), .C1(n_489), .C2(n_494), .Y(n_1067) );
OAI22xp5_ASAP7_75t_L g1068 ( .A1(n_913), .A2(n_558), .B1(n_499), .B2(n_518), .Y(n_1068) );
OAI21xp5_ASAP7_75t_L g1069 ( .A1(n_923), .A2(n_518), .B(n_429), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_950), .B(n_558), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_926), .A2(n_546), .B1(n_561), .B2(n_558), .Y(n_1071) );
NOR2x1_ASAP7_75t_SL g1072 ( .A(n_955), .B(n_558), .Y(n_1072) );
NOR2xp67_ASAP7_75t_L g1073 ( .A(n_893), .B(n_5), .Y(n_1073) );
OAI22xp5_ASAP7_75t_L g1074 ( .A1(n_913), .A2(n_396), .B1(n_677), .B2(n_675), .Y(n_1074) );
INVx2_ASAP7_75t_L g1075 ( .A(n_909), .Y(n_1075) );
BUFx2_ASAP7_75t_L g1076 ( .A(n_955), .Y(n_1076) );
INVx2_ASAP7_75t_L g1077 ( .A(n_909), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_863), .A2(n_599), .B1(n_677), .B2(n_675), .Y(n_1078) );
OAI221xp5_ASAP7_75t_L g1079 ( .A1(n_883), .A2(n_599), .B1(n_677), .B2(n_675), .C(n_9), .Y(n_1079) );
AOI21xp5_ASAP7_75t_L g1080 ( .A1(n_867), .A2(n_675), .B(n_599), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_871), .A2(n_874), .B1(n_887), .B2(n_896), .Y(n_1081) );
OAI21xp5_ASAP7_75t_SL g1082 ( .A1(n_967), .A2(n_6), .B(n_7), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_948), .Y(n_1083) );
AOI221xp5_ASAP7_75t_L g1084 ( .A1(n_897), .A2(n_599), .B1(n_9), .B2(n_10), .C(n_11), .Y(n_1084) );
OAI211xp5_ASAP7_75t_L g1085 ( .A1(n_859), .A2(n_11), .B(n_8), .C(n_10), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_950), .B(n_8), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_956), .Y(n_1087) );
HB1xp67_ASAP7_75t_L g1088 ( .A(n_1005), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_898), .A2(n_14), .B1(n_12), .B2(n_13), .Y(n_1089) );
OR2x2_ASAP7_75t_L g1090 ( .A(n_950), .B(n_13), .Y(n_1090) );
AOI22xp33_ASAP7_75t_SL g1091 ( .A1(n_885), .A2(n_17), .B1(n_14), .B2(n_16), .Y(n_1091) );
A2O1A1Ixp33_ASAP7_75t_SL g1092 ( .A1(n_964), .A2(n_18), .B(n_16), .C(n_17), .Y(n_1092) );
INVx2_ASAP7_75t_L g1093 ( .A(n_914), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_902), .A2(n_20), .B1(n_18), .B2(n_19), .Y(n_1094) );
CKINVDCx5p33_ASAP7_75t_R g1095 ( .A(n_1006), .Y(n_1095) );
AND2x4_ASAP7_75t_L g1096 ( .A(n_861), .B(n_21), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1097 ( .A(n_965), .B(n_22), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_910), .A2(n_24), .B1(n_22), .B2(n_23), .Y(n_1098) );
AO21x2_ASAP7_75t_L g1099 ( .A1(n_951), .A2(n_24), .B(n_25), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_970), .A2(n_27), .B1(n_25), .B2(n_26), .Y(n_1100) );
INVxp33_ASAP7_75t_L g1101 ( .A(n_985), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_977), .B(n_27), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_930), .B(n_28), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_970), .A2(n_31), .B1(n_29), .B2(n_30), .Y(n_1104) );
HB1xp67_ASAP7_75t_L g1105 ( .A(n_1007), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_879), .Y(n_1106) );
AO21x2_ASAP7_75t_L g1107 ( .A1(n_951), .A2(n_32), .B(n_33), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_859), .A2(n_35), .B1(n_32), .B2(n_34), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_973), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_940), .A2(n_996), .B1(n_984), .B2(n_866), .Y(n_1110) );
INVx3_ASAP7_75t_L g1111 ( .A(n_981), .Y(n_1111) );
OAI221xp5_ASAP7_75t_L g1112 ( .A1(n_905), .A2(n_36), .B1(n_37), .B2(n_38), .C(n_40), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_942), .B(n_36), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_940), .A2(n_40), .B1(n_37), .B2(n_38), .Y(n_1114) );
HB1xp67_ASAP7_75t_L g1115 ( .A(n_981), .Y(n_1115) );
AOI22xp33_ASAP7_75t_SL g1116 ( .A1(n_876), .A2(n_931), .B1(n_900), .B2(n_984), .Y(n_1116) );
BUFx3_ASAP7_75t_L g1117 ( .A(n_981), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_996), .A2(n_45), .B1(n_41), .B2(n_43), .Y(n_1118) );
AOI221xp5_ASAP7_75t_L g1119 ( .A1(n_967), .A2(n_43), .B1(n_46), .B2(n_47), .C(n_49), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_960), .B(n_46), .Y(n_1120) );
OAI22xp33_ASAP7_75t_L g1121 ( .A1(n_955), .A2(n_53), .B1(n_51), .B2(n_52), .Y(n_1121) );
AOI22xp33_ASAP7_75t_SL g1122 ( .A1(n_876), .A2(n_52), .B1(n_54), .B2(n_55), .Y(n_1122) );
INVx2_ASAP7_75t_L g1123 ( .A(n_914), .Y(n_1123) );
OAI221xp5_ASAP7_75t_L g1124 ( .A1(n_901), .A2(n_55), .B1(n_56), .B2(n_57), .C(n_58), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_912), .B(n_57), .Y(n_1125) );
INVx2_ASAP7_75t_L g1126 ( .A(n_914), .Y(n_1126) );
OAI332xp33_ASAP7_75t_L g1127 ( .A1(n_968), .A2(n_58), .A3(n_59), .B1(n_61), .B2(n_62), .B3(n_63), .C1(n_64), .C2(n_65), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_982), .B(n_61), .Y(n_1128) );
INVx2_ASAP7_75t_L g1129 ( .A(n_914), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_861), .B(n_66), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g1131 ( .A1(n_856), .A2(n_67), .B1(n_69), .B2(n_70), .Y(n_1131) );
INVxp67_ASAP7_75t_SL g1132 ( .A(n_980), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_861), .B(n_69), .Y(n_1133) );
OAI22xp5_ASAP7_75t_L g1134 ( .A1(n_980), .A2(n_70), .B1(n_72), .B2(n_73), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1135 ( .A1(n_880), .A2(n_72), .B1(n_73), .B2(n_74), .Y(n_1135) );
AOI221xp5_ASAP7_75t_L g1136 ( .A1(n_937), .A2(n_75), .B1(n_76), .B2(n_77), .C(n_78), .Y(n_1136) );
INVx8_ASAP7_75t_L g1137 ( .A(n_880), .Y(n_1137) );
AND2x4_ASAP7_75t_L g1138 ( .A(n_880), .B(n_75), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_975), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_856), .A2(n_77), .B1(n_79), .B2(n_80), .Y(n_1140) );
HB1xp67_ASAP7_75t_L g1141 ( .A(n_866), .Y(n_1141) );
OAI22xp5_ASAP7_75t_SL g1142 ( .A1(n_878), .A2(n_79), .B1(n_81), .B2(n_82), .Y(n_1142) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_865), .A2(n_931), .B1(n_908), .B2(n_976), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_995), .Y(n_1144) );
AOI22xp5_ASAP7_75t_SL g1145 ( .A1(n_929), .A2(n_81), .B1(n_82), .B2(n_83), .Y(n_1145) );
A2O1A1Ixp33_ASAP7_75t_L g1146 ( .A1(n_957), .A2(n_83), .B(n_84), .C(n_85), .Y(n_1146) );
AOI21xp5_ASAP7_75t_L g1147 ( .A1(n_922), .A2(n_148), .B(n_145), .Y(n_1147) );
NAND3xp33_ASAP7_75t_L g1148 ( .A(n_952), .B(n_86), .C(n_88), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g1149 ( .A1(n_865), .A2(n_86), .B1(n_88), .B2(n_89), .Y(n_1149) );
AO21x2_ASAP7_75t_L g1150 ( .A1(n_869), .A2(n_89), .B(n_90), .Y(n_1150) );
OR2x2_ASAP7_75t_L g1151 ( .A(n_954), .B(n_90), .Y(n_1151) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_999), .A2(n_91), .B1(n_92), .B2(n_93), .Y(n_1152) );
OR2x2_ASAP7_75t_L g1153 ( .A(n_1008), .B(n_92), .Y(n_1153) );
OR2x6_ASAP7_75t_L g1154 ( .A(n_876), .B(n_93), .Y(n_1154) );
INVx2_ASAP7_75t_L g1155 ( .A(n_988), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1001), .Y(n_1156) );
AOI221xp5_ASAP7_75t_L g1157 ( .A1(n_927), .A2(n_94), .B1(n_96), .B2(n_97), .C(n_98), .Y(n_1157) );
INVxp67_ASAP7_75t_L g1158 ( .A(n_1004), .Y(n_1158) );
HB1xp67_ASAP7_75t_L g1159 ( .A(n_989), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_918), .B(n_98), .Y(n_1160) );
NAND3xp33_ASAP7_75t_L g1161 ( .A(n_1037), .B(n_952), .C(n_958), .Y(n_1161) );
NAND3xp33_ASAP7_75t_SL g1162 ( .A(n_1082), .B(n_958), .C(n_979), .Y(n_1162) );
AO21x2_ASAP7_75t_L g1163 ( .A1(n_1018), .A2(n_873), .B(n_860), .Y(n_1163) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1031), .Y(n_1164) );
OAI211xp5_ASAP7_75t_L g1165 ( .A1(n_1034), .A2(n_998), .B(n_997), .C(n_990), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1061), .Y(n_1166) );
AOI22xp33_ASAP7_75t_SL g1167 ( .A1(n_1137), .A2(n_994), .B1(n_966), .B2(n_904), .Y(n_1167) );
OR2x6_ASAP7_75t_L g1168 ( .A(n_1137), .B(n_966), .Y(n_1168) );
AO21x2_ASAP7_75t_L g1169 ( .A1(n_1018), .A2(n_969), .B(n_992), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_1086), .A2(n_964), .B1(n_959), .B2(n_1003), .Y(n_1170) );
AOI221xp5_ASAP7_75t_L g1171 ( .A1(n_1063), .A2(n_936), .B1(n_925), .B2(n_990), .C(n_998), .Y(n_1171) );
OAI22xp33_ASAP7_75t_L g1172 ( .A1(n_1154), .A2(n_969), .B1(n_932), .B2(n_907), .Y(n_1172) );
NAND4xp25_ASAP7_75t_L g1173 ( .A(n_1016), .B(n_997), .C(n_979), .D(n_1000), .Y(n_1173) );
AOI221xp5_ASAP7_75t_L g1174 ( .A1(n_1106), .A2(n_1000), .B1(n_961), .B2(n_953), .C(n_855), .Y(n_1174) );
OAI33xp33_ASAP7_75t_L g1175 ( .A1(n_1142), .A2(n_99), .A3(n_100), .B1(n_101), .B2(n_102), .B3(n_103), .Y(n_1175) );
OAI211xp5_ASAP7_75t_L g1176 ( .A1(n_1020), .A2(n_961), .B(n_949), .C(n_938), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1177 ( .A(n_1088), .B(n_895), .Y(n_1177) );
AOI221xp5_ASAP7_75t_L g1178 ( .A1(n_1127), .A2(n_953), .B1(n_938), .B2(n_949), .C(n_933), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1021), .Y(n_1179) );
OAI33xp33_ASAP7_75t_L g1180 ( .A1(n_1121), .A2(n_1135), .A3(n_1100), .B1(n_1134), .B2(n_1057), .B3(n_1153), .Y(n_1180) );
INVx2_ASAP7_75t_L g1181 ( .A(n_1030), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1109), .Y(n_1182) );
BUFx3_ASAP7_75t_L g1183 ( .A(n_1017), .Y(n_1183) );
NAND3xp33_ASAP7_75t_L g1184 ( .A(n_1157), .B(n_857), .C(n_851), .Y(n_1184) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_1086), .A2(n_994), .B1(n_895), .B2(n_907), .Y(n_1185) );
AOI221xp5_ASAP7_75t_L g1186 ( .A1(n_1062), .A2(n_1009), .B1(n_894), .B2(n_920), .C(n_921), .Y(n_1186) );
NAND3xp33_ASAP7_75t_L g1187 ( .A(n_1056), .B(n_877), .C(n_870), .Y(n_1187) );
OAI22xp33_ASAP7_75t_L g1188 ( .A1(n_1154), .A2(n_921), .B1(n_994), .B2(n_966), .Y(n_1188) );
AOI22xp5_ASAP7_75t_L g1189 ( .A1(n_1024), .A2(n_1009), .B1(n_1002), .B2(n_993), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_1132), .A2(n_986), .B1(n_972), .B2(n_941), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1139), .Y(n_1191) );
OAI211xp5_ASAP7_75t_L g1192 ( .A1(n_1094), .A2(n_915), .B(n_911), .C(n_102), .Y(n_1192) );
AOI222xp33_ASAP7_75t_L g1193 ( .A1(n_1119), .A2(n_903), .B1(n_100), .B2(n_104), .C1(n_105), .C2(n_106), .Y(n_1193) );
OA21x2_ASAP7_75t_L g1194 ( .A1(n_1080), .A2(n_150), .B(n_149), .Y(n_1194) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1144), .Y(n_1195) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1030), .Y(n_1196) );
OR2x2_ASAP7_75t_L g1197 ( .A(n_1105), .B(n_99), .Y(n_1197) );
NAND3xp33_ASAP7_75t_L g1198 ( .A(n_1122), .B(n_104), .C(n_105), .Y(n_1198) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_1096), .A2(n_899), .B1(n_107), .B2(n_108), .Y(n_1199) );
INVx2_ASAP7_75t_L g1200 ( .A(n_1035), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1130), .B(n_106), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_1011), .B(n_107), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_1096), .A2(n_899), .B1(n_110), .B2(n_111), .Y(n_1203) );
OAI221xp5_ASAP7_75t_L g1204 ( .A1(n_1143), .A2(n_109), .B1(n_110), .B2(n_111), .C(n_112), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1130), .B(n_1133), .Y(n_1205) );
AOI21xp33_ASAP7_75t_L g1206 ( .A1(n_1019), .A2(n_109), .B(n_112), .Y(n_1206) );
INVx3_ASAP7_75t_L g1207 ( .A(n_1017), .Y(n_1207) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_1096), .A2(n_113), .B1(n_114), .B2(n_115), .Y(n_1208) );
AOI33xp33_ASAP7_75t_L g1209 ( .A1(n_1098), .A2(n_113), .A3(n_114), .B1(n_115), .B2(n_116), .B3(n_117), .Y(n_1209) );
AOI22xp33_ASAP7_75t_L g1210 ( .A1(n_1138), .A2(n_116), .B1(n_117), .B2(n_118), .Y(n_1210) );
OAI21xp5_ASAP7_75t_L g1211 ( .A1(n_1079), .A2(n_1065), .B(n_1067), .Y(n_1211) );
INVx2_ASAP7_75t_L g1212 ( .A(n_1035), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1156), .Y(n_1213) );
AOI22xp33_ASAP7_75t_L g1214 ( .A1(n_1138), .A2(n_118), .B1(n_120), .B2(n_121), .Y(n_1214) );
AO21x2_ASAP7_75t_L g1215 ( .A1(n_1092), .A2(n_121), .B(n_122), .Y(n_1215) );
AO21x2_ASAP7_75t_L g1216 ( .A1(n_1092), .A2(n_123), .B(n_124), .Y(n_1216) );
NAND3xp33_ASAP7_75t_L g1217 ( .A(n_1112), .B(n_123), .C(n_125), .Y(n_1217) );
AOI22xp5_ASAP7_75t_L g1218 ( .A1(n_1138), .A2(n_125), .B1(n_127), .B2(n_128), .Y(n_1218) );
AOI221xp5_ASAP7_75t_L g1219 ( .A1(n_1124), .A2(n_128), .B1(n_130), .B2(n_131), .C(n_132), .Y(n_1219) );
AOI221xp5_ASAP7_75t_L g1220 ( .A1(n_1146), .A2(n_130), .B1(n_132), .B2(n_133), .C(n_134), .Y(n_1220) );
OAI22xp5_ASAP7_75t_L g1221 ( .A1(n_1154), .A2(n_133), .B1(n_134), .B2(n_136), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1153), .Y(n_1222) );
OAI21xp5_ASAP7_75t_L g1223 ( .A1(n_1074), .A2(n_136), .B(n_137), .Y(n_1223) );
OAI22xp5_ASAP7_75t_L g1224 ( .A1(n_1154), .A2(n_137), .B1(n_138), .B2(n_139), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1064), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1083), .Y(n_1226) );
OAI21xp5_ASAP7_75t_L g1227 ( .A1(n_1032), .A2(n_138), .B(n_140), .Y(n_1227) );
AO21x2_ASAP7_75t_L g1228 ( .A1(n_1090), .A2(n_140), .B(n_141), .Y(n_1228) );
AOI33xp33_ASAP7_75t_L g1229 ( .A1(n_1091), .A2(n_141), .A3(n_151), .B1(n_153), .B2(n_156), .B3(n_158), .Y(n_1229) );
NOR2xp33_ASAP7_75t_L g1230 ( .A(n_1128), .B(n_159), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_1125), .A2(n_160), .B1(n_161), .B2(n_162), .Y(n_1231) );
OA21x2_ASAP7_75t_L g1232 ( .A1(n_1090), .A2(n_163), .B(n_166), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1160), .B(n_354), .Y(n_1233) );
AOI22xp33_ASAP7_75t_SL g1234 ( .A1(n_1137), .A2(n_168), .B1(n_169), .B2(n_173), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1133), .B(n_352), .Y(n_1235) );
OAI321xp33_ASAP7_75t_L g1236 ( .A1(n_1148), .A2(n_174), .A3(n_178), .B1(n_179), .B2(n_180), .C(n_181), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1103), .B(n_184), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g1238 ( .A1(n_1125), .A2(n_186), .B1(n_188), .B2(n_189), .Y(n_1238) );
OR2x2_ASAP7_75t_L g1239 ( .A(n_1027), .B(n_351), .Y(n_1239) );
OAI221xp5_ASAP7_75t_L g1240 ( .A1(n_1116), .A2(n_191), .B1(n_195), .B2(n_196), .C(n_198), .Y(n_1240) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_1160), .A2(n_201), .B1(n_202), .B2(n_203), .Y(n_1241) );
INVx2_ASAP7_75t_L g1242 ( .A(n_1155), .Y(n_1242) );
INVx3_ASAP7_75t_L g1243 ( .A(n_1137), .Y(n_1243) );
AOI21xp5_ASAP7_75t_L g1244 ( .A1(n_1042), .A2(n_204), .B(n_207), .Y(n_1244) );
INVx2_ASAP7_75t_SL g1245 ( .A(n_1022), .Y(n_1245) );
AOI22xp33_ASAP7_75t_L g1246 ( .A1(n_1103), .A2(n_208), .B1(n_209), .B2(n_211), .Y(n_1246) );
AOI22xp5_ASAP7_75t_L g1247 ( .A1(n_1015), .A2(n_212), .B1(n_213), .B2(n_214), .Y(n_1247) );
OAI22xp5_ASAP7_75t_L g1248 ( .A1(n_1036), .A2(n_216), .B1(n_218), .B2(n_219), .Y(n_1248) );
AOI221xp5_ASAP7_75t_L g1249 ( .A1(n_1146), .A2(n_1136), .B1(n_1084), .B2(n_1087), .C(n_1043), .Y(n_1249) );
HB1xp67_ASAP7_75t_L g1250 ( .A(n_1027), .Y(n_1250) );
BUFx2_ASAP7_75t_L g1251 ( .A(n_1117), .Y(n_1251) );
AOI221xp5_ASAP7_75t_L g1252 ( .A1(n_1081), .A2(n_1104), .B1(n_1108), .B2(n_1149), .C(n_1068), .Y(n_1252) );
NOR2xp33_ASAP7_75t_L g1253 ( .A(n_1051), .B(n_220), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1102), .B(n_348), .Y(n_1254) );
AOI221xp5_ASAP7_75t_L g1255 ( .A1(n_1071), .A2(n_221), .B1(n_223), .B2(n_225), .C(n_226), .Y(n_1255) );
AOI22xp33_ASAP7_75t_L g1256 ( .A1(n_1113), .A2(n_1102), .B1(n_1120), .B2(n_1107), .Y(n_1256) );
OAI22xp33_ASAP7_75t_L g1257 ( .A1(n_1076), .A2(n_229), .B1(n_230), .B2(n_231), .Y(n_1257) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1151), .B(n_345), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1113), .B(n_232), .Y(n_1259) );
AOI22xp33_ASAP7_75t_L g1260 ( .A1(n_1120), .A2(n_234), .B1(n_235), .B2(n_236), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1145), .B(n_240), .Y(n_1261) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1151), .Y(n_1262) );
OAI22xp33_ASAP7_75t_L g1263 ( .A1(n_1076), .A2(n_244), .B1(n_247), .B2(n_248), .Y(n_1263) );
OAI22xp5_ASAP7_75t_L g1264 ( .A1(n_1033), .A2(n_250), .B1(n_251), .B2(n_252), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1097), .Y(n_1265) );
INVx2_ASAP7_75t_L g1266 ( .A(n_1048), .Y(n_1266) );
OR2x2_ASAP7_75t_L g1267 ( .A(n_1058), .B(n_344), .Y(n_1267) );
NOR2x1_ASAP7_75t_SL g1268 ( .A(n_1117), .B(n_255), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1158), .B(n_256), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1101), .B(n_258), .Y(n_1270) );
CKINVDCx5p33_ASAP7_75t_R g1271 ( .A(n_1050), .Y(n_1271) );
OAI332xp33_ASAP7_75t_L g1272 ( .A1(n_1023), .A2(n_259), .A3(n_262), .B1(n_264), .B2(n_266), .B3(n_269), .C1(n_274), .C2(n_276), .Y(n_1272) );
AOI22xp33_ASAP7_75t_L g1273 ( .A1(n_1099), .A2(n_277), .B1(n_281), .B2(n_282), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1101), .B(n_283), .Y(n_1274) );
OAI22xp5_ASAP7_75t_L g1275 ( .A1(n_1110), .A2(n_285), .B1(n_286), .B2(n_287), .Y(n_1275) );
INVx2_ASAP7_75t_L g1276 ( .A(n_1048), .Y(n_1276) );
INVx2_ASAP7_75t_L g1277 ( .A(n_1075), .Y(n_1277) );
INVx2_ASAP7_75t_SL g1278 ( .A(n_1022), .Y(n_1278) );
OA222x2_ASAP7_75t_L g1279 ( .A1(n_1111), .A2(n_288), .B1(n_290), .B2(n_291), .C1(n_292), .C2(n_293), .Y(n_1279) );
OAI33xp33_ASAP7_75t_L g1280 ( .A1(n_1055), .A2(n_298), .A3(n_299), .B1(n_300), .B2(n_306), .B3(n_307), .Y(n_1280) );
OAI221xp5_ASAP7_75t_L g1281 ( .A1(n_1060), .A2(n_312), .B1(n_316), .B2(n_317), .C(n_322), .Y(n_1281) );
NOR2xp33_ASAP7_75t_L g1282 ( .A(n_1041), .B(n_324), .Y(n_1282) );
OAI31xp33_ASAP7_75t_L g1283 ( .A1(n_1261), .A2(n_1085), .A3(n_1047), .B(n_1010), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1164), .Y(n_1284) );
OAI221xp5_ASAP7_75t_L g1285 ( .A1(n_1199), .A2(n_1073), .B1(n_1114), .B2(n_1118), .C(n_1140), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1205), .B(n_1059), .Y(n_1286) );
OAI22xp5_ASAP7_75t_SL g1287 ( .A1(n_1271), .A2(n_1050), .B1(n_1095), .B2(n_1013), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1262), .B(n_1155), .Y(n_1288) );
INVx2_ASAP7_75t_L g1289 ( .A(n_1181), .Y(n_1289) );
NAND3xp33_ASAP7_75t_L g1290 ( .A(n_1208), .B(n_1152), .C(n_1089), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1166), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1182), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1242), .B(n_1059), .Y(n_1293) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1191), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1250), .B(n_1070), .Y(n_1295) );
INVxp67_ASAP7_75t_L g1296 ( .A(n_1251), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1195), .B(n_1070), .Y(n_1297) );
AOI33xp33_ASAP7_75t_L g1298 ( .A1(n_1208), .A2(n_1131), .A3(n_1054), .B1(n_1066), .B2(n_1026), .B3(n_1038), .Y(n_1298) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1213), .Y(n_1299) );
NAND3xp33_ASAP7_75t_L g1300 ( .A(n_1210), .B(n_1069), .C(n_1040), .Y(n_1300) );
BUFx3_ASAP7_75t_L g1301 ( .A(n_1183), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1222), .B(n_1099), .Y(n_1302) );
OAI33xp33_ASAP7_75t_L g1303 ( .A1(n_1221), .A2(n_1013), .A3(n_1039), .B1(n_1095), .B2(n_1049), .B3(n_1099), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1200), .B(n_1107), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1200), .B(n_1107), .Y(n_1305) );
OAI22xp5_ASAP7_75t_L g1306 ( .A1(n_1199), .A2(n_1029), .B1(n_1028), .B2(n_1052), .Y(n_1306) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_1179), .B(n_1141), .Y(n_1307) );
AOI222xp33_ASAP7_75t_L g1308 ( .A1(n_1178), .A2(n_1072), .B1(n_1115), .B2(n_1012), .C1(n_1111), .C2(n_1159), .Y(n_1308) );
AOI22xp5_ASAP7_75t_L g1309 ( .A1(n_1161), .A2(n_1014), .B1(n_1025), .B2(n_1046), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1212), .B(n_1129), .Y(n_1310) );
INVxp67_ASAP7_75t_SL g1311 ( .A(n_1172), .Y(n_1311) );
INVx2_ASAP7_75t_L g1312 ( .A(n_1196), .Y(n_1312) );
INVx8_ASAP7_75t_L g1313 ( .A(n_1168), .Y(n_1313) );
OAI33xp33_ASAP7_75t_L g1314 ( .A1(n_1224), .A2(n_1150), .A3(n_1129), .B1(n_1126), .B2(n_1123), .B3(n_1075), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1225), .Y(n_1315) );
OAI221xp5_ASAP7_75t_L g1316 ( .A1(n_1203), .A2(n_1044), .B1(n_1111), .B2(n_1053), .C(n_1025), .Y(n_1316) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1226), .Y(n_1317) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1177), .Y(n_1318) );
INVxp67_ASAP7_75t_SL g1319 ( .A(n_1172), .Y(n_1319) );
INVx2_ASAP7_75t_SL g1320 ( .A(n_1183), .Y(n_1320) );
NAND2x1p5_ASAP7_75t_SL g1321 ( .A(n_1237), .B(n_1126), .Y(n_1321) );
NAND3xp33_ASAP7_75t_L g1322 ( .A(n_1210), .B(n_1147), .C(n_1032), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1201), .B(n_1072), .Y(n_1323) );
INVx2_ASAP7_75t_L g1324 ( .A(n_1196), .Y(n_1324) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1228), .Y(n_1325) );
AOI33xp33_ASAP7_75t_L g1326 ( .A1(n_1214), .A2(n_1078), .A3(n_1123), .B1(n_1093), .B2(n_1077), .B3(n_1150), .Y(n_1326) );
NOR3xp33_ASAP7_75t_SL g1327 ( .A(n_1175), .B(n_1025), .C(n_1150), .Y(n_1327) );
AND2x4_ASAP7_75t_L g1328 ( .A(n_1212), .B(n_1093), .Y(n_1328) );
AND2x4_ASAP7_75t_SL g1329 ( .A(n_1243), .B(n_1077), .Y(n_1329) );
OAI221xp5_ASAP7_75t_L g1330 ( .A1(n_1203), .A2(n_1025), .B1(n_1045), .B2(n_328), .C(n_329), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1266), .B(n_1045), .Y(n_1331) );
NAND2xp5_ASAP7_75t_L g1332 ( .A(n_1265), .B(n_1045), .Y(n_1332) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1228), .Y(n_1333) );
OAI31xp33_ASAP7_75t_L g1334 ( .A1(n_1204), .A2(n_326), .A3(n_327), .B(n_330), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1197), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1202), .B(n_343), .Y(n_1336) );
INVx2_ASAP7_75t_L g1337 ( .A(n_1266), .Y(n_1337) );
OAI33xp33_ASAP7_75t_L g1338 ( .A1(n_1257), .A2(n_333), .A3(n_334), .B1(n_340), .B2(n_341), .B3(n_1263), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1235), .B(n_1209), .Y(n_1339) );
INVxp33_ASAP7_75t_L g1340 ( .A(n_1259), .Y(n_1340) );
OR2x6_ASAP7_75t_L g1341 ( .A(n_1168), .B(n_1227), .Y(n_1341) );
NAND2xp5_ASAP7_75t_L g1342 ( .A(n_1209), .B(n_1256), .Y(n_1342) );
AOI22xp5_ASAP7_75t_L g1343 ( .A1(n_1180), .A2(n_1193), .B1(n_1282), .B2(n_1252), .Y(n_1343) );
OAI22xp5_ASAP7_75t_L g1344 ( .A1(n_1214), .A2(n_1218), .B1(n_1258), .B2(n_1260), .Y(n_1344) );
NAND3xp33_ASAP7_75t_L g1345 ( .A(n_1256), .B(n_1219), .C(n_1220), .Y(n_1345) );
NAND4xp25_ASAP7_75t_L g1346 ( .A(n_1217), .B(n_1198), .C(n_1249), .D(n_1273), .Y(n_1346) );
AOI21xp5_ASAP7_75t_L g1347 ( .A1(n_1188), .A2(n_1263), .B(n_1257), .Y(n_1347) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1276), .B(n_1277), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1276), .B(n_1277), .Y(n_1349) );
AND4x1_ASAP7_75t_L g1350 ( .A(n_1229), .B(n_1211), .C(n_1246), .D(n_1260), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_1185), .B(n_1190), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1243), .B(n_1189), .Y(n_1352) );
BUFx3_ASAP7_75t_L g1353 ( .A(n_1207), .Y(n_1353) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1239), .Y(n_1354) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1185), .B(n_1190), .Y(n_1355) );
INVx2_ASAP7_75t_L g1356 ( .A(n_1232), .Y(n_1356) );
INVxp67_ASAP7_75t_L g1357 ( .A(n_1267), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1232), .B(n_1279), .Y(n_1358) );
NAND4xp25_ASAP7_75t_L g1359 ( .A(n_1273), .B(n_1229), .C(n_1173), .D(n_1171), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1163), .B(n_1169), .Y(n_1360) );
OR2x2_ASAP7_75t_L g1361 ( .A(n_1207), .B(n_1168), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1269), .B(n_1270), .Y(n_1362) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1274), .Y(n_1363) );
AOI33xp33_ASAP7_75t_L g1364 ( .A1(n_1245), .A2(n_1278), .A3(n_1238), .B1(n_1231), .B2(n_1170), .B3(n_1241), .Y(n_1364) );
AOI22xp33_ASAP7_75t_L g1365 ( .A1(n_1162), .A2(n_1282), .B1(n_1223), .B2(n_1170), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1163), .B(n_1169), .Y(n_1366) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1187), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1230), .B(n_1233), .Y(n_1368) );
OAI321xp33_ASAP7_75t_L g1369 ( .A1(n_1188), .A2(n_1240), .A3(n_1238), .B1(n_1231), .B2(n_1241), .C(n_1246), .Y(n_1369) );
AOI211xp5_ASAP7_75t_SL g1370 ( .A1(n_1272), .A2(n_1165), .B(n_1176), .C(n_1236), .Y(n_1370) );
AOI22xp5_ASAP7_75t_L g1371 ( .A1(n_1230), .A2(n_1253), .B1(n_1192), .B2(n_1174), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1253), .B(n_1215), .Y(n_1372) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1184), .Y(n_1373) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1215), .Y(n_1374) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1318), .B(n_1254), .Y(n_1375) );
OR2x2_ASAP7_75t_L g1376 ( .A(n_1295), .B(n_1216), .Y(n_1376) );
NAND2xp5_ASAP7_75t_L g1377 ( .A(n_1335), .B(n_1216), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1304), .B(n_1194), .Y(n_1378) );
INVx1_ASAP7_75t_SL g1379 ( .A(n_1287), .Y(n_1379) );
NAND2xp5_ASAP7_75t_L g1380 ( .A(n_1284), .B(n_1206), .Y(n_1380) );
OR2x2_ASAP7_75t_L g1381 ( .A(n_1295), .B(n_1167), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1304), .B(n_1194), .Y(n_1382) );
NAND2xp5_ASAP7_75t_L g1383 ( .A(n_1291), .B(n_1186), .Y(n_1383) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1292), .Y(n_1384) );
INVx2_ASAP7_75t_L g1385 ( .A(n_1289), .Y(n_1385) );
NAND2xp5_ASAP7_75t_L g1386 ( .A(n_1294), .B(n_1247), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1305), .B(n_1194), .Y(n_1387) );
HB1xp67_ASAP7_75t_L g1388 ( .A(n_1337), .Y(n_1388) );
OR2x2_ASAP7_75t_L g1389 ( .A(n_1286), .B(n_1297), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1305), .B(n_1268), .Y(n_1390) );
AND2x2_ASAP7_75t_L g1391 ( .A(n_1286), .B(n_1234), .Y(n_1391) );
HB1xp67_ASAP7_75t_L g1392 ( .A(n_1337), .Y(n_1392) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1299), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1394 ( .A(n_1315), .B(n_1317), .Y(n_1394) );
OR2x6_ASAP7_75t_L g1395 ( .A(n_1341), .B(n_1244), .Y(n_1395) );
OR2x2_ASAP7_75t_L g1396 ( .A(n_1297), .B(n_1264), .Y(n_1396) );
INVx1_ASAP7_75t_SL g1397 ( .A(n_1329), .Y(n_1397) );
INVx1_ASAP7_75t_SL g1398 ( .A(n_1329), .Y(n_1398) );
OR2x2_ASAP7_75t_L g1399 ( .A(n_1296), .B(n_1275), .Y(n_1399) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1307), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1348), .B(n_1255), .Y(n_1401) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1288), .Y(n_1402) );
NAND2xp5_ASAP7_75t_L g1403 ( .A(n_1354), .B(n_1248), .Y(n_1403) );
AOI21xp5_ASAP7_75t_L g1404 ( .A1(n_1347), .A2(n_1280), .B(n_1281), .Y(n_1404) );
INVxp67_ASAP7_75t_L g1405 ( .A(n_1323), .Y(n_1405) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1293), .B(n_1342), .Y(n_1406) );
INVx5_ASAP7_75t_L g1407 ( .A(n_1313), .Y(n_1407) );
INVx2_ASAP7_75t_SL g1408 ( .A(n_1301), .Y(n_1408) );
AND2x4_ASAP7_75t_L g1409 ( .A(n_1348), .B(n_1349), .Y(n_1409) );
INVxp67_ASAP7_75t_L g1410 ( .A(n_1352), .Y(n_1410) );
OR2x2_ASAP7_75t_L g1411 ( .A(n_1302), .B(n_1340), .Y(n_1411) );
OAI21xp33_ASAP7_75t_L g1412 ( .A1(n_1358), .A2(n_1367), .B(n_1364), .Y(n_1412) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1332), .Y(n_1413) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_1363), .B(n_1357), .Y(n_1414) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1325), .Y(n_1415) );
INVx2_ASAP7_75t_SL g1416 ( .A(n_1301), .Y(n_1416) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1333), .Y(n_1417) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1310), .Y(n_1418) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1310), .Y(n_1419) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_1339), .B(n_1343), .Y(n_1420) );
NAND2xp5_ASAP7_75t_L g1421 ( .A(n_1340), .B(n_1365), .Y(n_1421) );
AOI211x1_ASAP7_75t_L g1422 ( .A1(n_1350), .A2(n_1359), .B(n_1285), .C(n_1358), .Y(n_1422) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1320), .Y(n_1423) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1320), .Y(n_1424) );
OR2x2_ASAP7_75t_L g1425 ( .A(n_1351), .B(n_1355), .Y(n_1425) );
AND2x4_ASAP7_75t_L g1426 ( .A(n_1341), .B(n_1328), .Y(n_1426) );
NAND2xp5_ASAP7_75t_SL g1427 ( .A(n_1326), .B(n_1364), .Y(n_1427) );
NAND2xp5_ASAP7_75t_L g1428 ( .A(n_1365), .B(n_1362), .Y(n_1428) );
AND2x4_ASAP7_75t_L g1429 ( .A(n_1341), .B(n_1328), .Y(n_1429) );
OR2x2_ASAP7_75t_L g1430 ( .A(n_1351), .B(n_1355), .Y(n_1430) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_1312), .B(n_1324), .Y(n_1431) );
OR2x2_ASAP7_75t_L g1432 ( .A(n_1321), .B(n_1319), .Y(n_1432) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_1312), .B(n_1324), .Y(n_1433) );
AOI22xp33_ASAP7_75t_SL g1434 ( .A1(n_1313), .A2(n_1341), .B1(n_1311), .B2(n_1344), .Y(n_1434) );
NAND2xp5_ASAP7_75t_L g1435 ( .A(n_1373), .B(n_1368), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1360), .B(n_1366), .Y(n_1436) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_1308), .B(n_1371), .Y(n_1437) );
NOR2xp33_ASAP7_75t_L g1438 ( .A(n_1346), .B(n_1300), .Y(n_1438) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1353), .Y(n_1439) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1353), .Y(n_1440) );
NAND2xp5_ASAP7_75t_L g1441 ( .A(n_1425), .B(n_1372), .Y(n_1441) );
AND2x2_ASAP7_75t_L g1442 ( .A(n_1436), .B(n_1366), .Y(n_1442) );
NAND2xp5_ASAP7_75t_L g1443 ( .A(n_1430), .B(n_1372), .Y(n_1443) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1415), .Y(n_1444) );
OR2x2_ASAP7_75t_L g1445 ( .A(n_1411), .B(n_1374), .Y(n_1445) );
OR2x2_ASAP7_75t_L g1446 ( .A(n_1436), .B(n_1321), .Y(n_1446) );
OR2x2_ASAP7_75t_L g1447 ( .A(n_1409), .B(n_1360), .Y(n_1447) );
INVx2_ASAP7_75t_L g1448 ( .A(n_1385), .Y(n_1448) );
HB1xp67_ASAP7_75t_L g1449 ( .A(n_1388), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_1409), .B(n_1356), .Y(n_1450) );
INVx2_ASAP7_75t_L g1451 ( .A(n_1385), .Y(n_1451) );
NAND2xp5_ASAP7_75t_L g1452 ( .A(n_1400), .B(n_1345), .Y(n_1452) );
NAND2xp5_ASAP7_75t_L g1453 ( .A(n_1406), .B(n_1309), .Y(n_1453) );
AND2x2_ASAP7_75t_L g1454 ( .A(n_1409), .B(n_1356), .Y(n_1454) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1417), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_1435), .B(n_1370), .Y(n_1456) );
NAND2xp5_ASAP7_75t_L g1457 ( .A(n_1410), .B(n_1326), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1418), .B(n_1419), .Y(n_1458) );
NOR2x1_ASAP7_75t_L g1459 ( .A(n_1379), .B(n_1397), .Y(n_1459) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1384), .Y(n_1460) );
OAI21xp5_ASAP7_75t_L g1461 ( .A1(n_1438), .A2(n_1327), .B(n_1369), .Y(n_1461) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1393), .Y(n_1462) );
NAND2xp5_ASAP7_75t_L g1463 ( .A(n_1402), .B(n_1306), .Y(n_1463) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1394), .Y(n_1464) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1388), .Y(n_1465) );
NAND2xp5_ASAP7_75t_SL g1466 ( .A(n_1422), .B(n_1283), .Y(n_1466) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1392), .Y(n_1467) );
AND2x4_ASAP7_75t_L g1468 ( .A(n_1426), .B(n_1331), .Y(n_1468) );
NAND2x1_ASAP7_75t_L g1469 ( .A(n_1426), .B(n_1361), .Y(n_1469) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1414), .Y(n_1470) );
OAI21xp33_ASAP7_75t_SL g1471 ( .A1(n_1427), .A2(n_1334), .B(n_1316), .Y(n_1471) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1392), .Y(n_1472) );
INVx1_ASAP7_75t_SL g1473 ( .A(n_1398), .Y(n_1473) );
AOI211x1_ASAP7_75t_SL g1474 ( .A1(n_1427), .A2(n_1290), .B(n_1336), .C(n_1322), .Y(n_1474) );
NAND2xp5_ASAP7_75t_L g1475 ( .A(n_1428), .B(n_1298), .Y(n_1475) );
OR2x2_ASAP7_75t_L g1476 ( .A(n_1389), .B(n_1313), .Y(n_1476) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1423), .Y(n_1477) );
OR2x2_ASAP7_75t_L g1478 ( .A(n_1376), .B(n_1330), .Y(n_1478) );
NOR2xp33_ASAP7_75t_L g1479 ( .A(n_1420), .B(n_1303), .Y(n_1479) );
NAND2xp5_ASAP7_75t_L g1480 ( .A(n_1421), .B(n_1405), .Y(n_1480) );
NOR2x1_ASAP7_75t_L g1481 ( .A(n_1424), .B(n_1338), .Y(n_1481) );
INVxp67_ASAP7_75t_L g1482 ( .A(n_1408), .Y(n_1482) );
INVx3_ASAP7_75t_L g1483 ( .A(n_1426), .Y(n_1483) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1465), .Y(n_1484) );
OR2x2_ASAP7_75t_L g1485 ( .A(n_1441), .B(n_1432), .Y(n_1485) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1465), .Y(n_1486) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1467), .Y(n_1487) );
NAND2xp5_ASAP7_75t_L g1488 ( .A(n_1443), .B(n_1412), .Y(n_1488) );
INVx2_ASAP7_75t_L g1489 ( .A(n_1448), .Y(n_1489) );
AND2x2_ASAP7_75t_L g1490 ( .A(n_1442), .B(n_1429), .Y(n_1490) );
NAND2xp5_ASAP7_75t_L g1491 ( .A(n_1479), .B(n_1377), .Y(n_1491) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1467), .Y(n_1492) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1472), .Y(n_1493) );
NAND2xp5_ASAP7_75t_SL g1494 ( .A(n_1459), .B(n_1434), .Y(n_1494) );
NAND2xp5_ASAP7_75t_L g1495 ( .A(n_1470), .B(n_1383), .Y(n_1495) );
NAND2xp5_ASAP7_75t_SL g1496 ( .A(n_1473), .B(n_1407), .Y(n_1496) );
INVx1_ASAP7_75t_SL g1497 ( .A(n_1449), .Y(n_1497) );
OR2x2_ASAP7_75t_L g1498 ( .A(n_1445), .B(n_1413), .Y(n_1498) );
AOI221xp5_ASAP7_75t_L g1499 ( .A1(n_1466), .A2(n_1437), .B1(n_1375), .B2(n_1380), .C(n_1391), .Y(n_1499) );
INVxp67_ASAP7_75t_L g1500 ( .A(n_1452), .Y(n_1500) );
INVx1_ASAP7_75t_L g1501 ( .A(n_1472), .Y(n_1501) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1444), .Y(n_1502) );
INVx2_ASAP7_75t_L g1503 ( .A(n_1448), .Y(n_1503) );
OAI32xp33_ASAP7_75t_L g1504 ( .A1(n_1476), .A2(n_1381), .A3(n_1416), .B1(n_1399), .B2(n_1391), .Y(n_1504) );
NAND2xp5_ASAP7_75t_L g1505 ( .A(n_1457), .B(n_1416), .Y(n_1505) );
INVx2_ASAP7_75t_L g1506 ( .A(n_1451), .Y(n_1506) );
NAND2xp5_ASAP7_75t_L g1507 ( .A(n_1480), .B(n_1440), .Y(n_1507) );
NAND2xp5_ASAP7_75t_L g1508 ( .A(n_1464), .B(n_1439), .Y(n_1508) );
NAND2xp5_ASAP7_75t_L g1509 ( .A(n_1453), .B(n_1433), .Y(n_1509) );
NAND2xp5_ASAP7_75t_L g1510 ( .A(n_1458), .B(n_1433), .Y(n_1510) );
OAI22xp5_ASAP7_75t_L g1511 ( .A1(n_1476), .A2(n_1407), .B1(n_1429), .B2(n_1395), .Y(n_1511) );
NAND2xp5_ASAP7_75t_L g1512 ( .A(n_1458), .B(n_1431), .Y(n_1512) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1444), .Y(n_1513) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1455), .Y(n_1514) );
XNOR2xp5_ASAP7_75t_L g1515 ( .A(n_1456), .B(n_1429), .Y(n_1515) );
OAI21xp33_ASAP7_75t_L g1516 ( .A1(n_1461), .A2(n_1395), .B(n_1404), .Y(n_1516) );
XNOR2xp5_ASAP7_75t_L g1517 ( .A(n_1474), .B(n_1396), .Y(n_1517) );
XNOR2x1_ASAP7_75t_L g1518 ( .A(n_1475), .B(n_1401), .Y(n_1518) );
NAND2xp5_ASAP7_75t_L g1519 ( .A(n_1463), .B(n_1387), .Y(n_1519) );
O2A1O1Ixp5_ASAP7_75t_L g1520 ( .A1(n_1469), .A2(n_1403), .B(n_1386), .C(n_1314), .Y(n_1520) );
NAND2xp5_ASAP7_75t_SL g1521 ( .A(n_1482), .B(n_1407), .Y(n_1521) );
XNOR2xp5_ASAP7_75t_L g1522 ( .A(n_1447), .B(n_1390), .Y(n_1522) );
NAND2xp5_ASAP7_75t_L g1523 ( .A(n_1477), .B(n_1378), .Y(n_1523) );
XNOR2xp5_ASAP7_75t_L g1524 ( .A(n_1447), .B(n_1390), .Y(n_1524) );
AND2x2_ASAP7_75t_L g1525 ( .A(n_1450), .B(n_1378), .Y(n_1525) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1462), .Y(n_1526) );
INVx2_ASAP7_75t_L g1527 ( .A(n_1451), .Y(n_1527) );
NAND2xp5_ASAP7_75t_SL g1528 ( .A(n_1481), .B(n_1407), .Y(n_1528) );
XNOR2x1_ASAP7_75t_L g1529 ( .A(n_1446), .B(n_1401), .Y(n_1529) );
AOI21xp33_ASAP7_75t_L g1530 ( .A1(n_1471), .A2(n_1395), .B(n_1382), .Y(n_1530) );
INVx1_ASAP7_75t_L g1531 ( .A(n_1462), .Y(n_1531) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1460), .Y(n_1532) );
XNOR2xp5_ASAP7_75t_L g1533 ( .A(n_1468), .B(n_1395), .Y(n_1533) );
OAI211xp5_ASAP7_75t_SL g1534 ( .A1(n_1478), .A2(n_1446), .B(n_1445), .C(n_1483), .Y(n_1534) );
AOI22xp5_ASAP7_75t_L g1535 ( .A1(n_1494), .A2(n_1516), .B1(n_1517), .B2(n_1529), .Y(n_1535) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1485), .Y(n_1536) );
AOI21xp5_ASAP7_75t_L g1537 ( .A1(n_1528), .A2(n_1504), .B(n_1521), .Y(n_1537) );
NAND2xp5_ASAP7_75t_SL g1538 ( .A(n_1528), .B(n_1521), .Y(n_1538) );
AND2x4_ASAP7_75t_L g1539 ( .A(n_1490), .B(n_1483), .Y(n_1539) );
CKINVDCx20_ASAP7_75t_R g1540 ( .A(n_1500), .Y(n_1540) );
NAND3xp33_ASAP7_75t_SL g1541 ( .A(n_1499), .B(n_1497), .C(n_1496), .Y(n_1541) );
OAI31xp33_ASAP7_75t_L g1542 ( .A1(n_1534), .A2(n_1529), .A3(n_1518), .B(n_1530), .Y(n_1542) );
OAI221xp5_ASAP7_75t_SL g1543 ( .A1(n_1491), .A2(n_1515), .B1(n_1533), .B2(n_1488), .C(n_1522), .Y(n_1543) );
AOI22xp5_ASAP7_75t_L g1544 ( .A1(n_1505), .A2(n_1519), .B1(n_1511), .B2(n_1495), .Y(n_1544) );
A2O1A1Ixp33_ASAP7_75t_L g1545 ( .A1(n_1504), .A2(n_1520), .B(n_1483), .C(n_1498), .Y(n_1545) );
OAI221xp5_ASAP7_75t_L g1546 ( .A1(n_1542), .A2(n_1507), .B1(n_1524), .B2(n_1508), .C(n_1498), .Y(n_1546) );
OAI211xp5_ASAP7_75t_L g1547 ( .A1(n_1535), .A2(n_1478), .B(n_1509), .C(n_1532), .Y(n_1547) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1536), .Y(n_1548) );
AOI22xp5_ASAP7_75t_L g1549 ( .A1(n_1541), .A2(n_1523), .B1(n_1531), .B2(n_1526), .Y(n_1549) );
OAI22xp5_ASAP7_75t_L g1550 ( .A1(n_1543), .A2(n_1512), .B1(n_1510), .B2(n_1525), .Y(n_1550) );
OA22x2_ASAP7_75t_L g1551 ( .A1(n_1544), .A2(n_1484), .B1(n_1492), .B2(n_1501), .Y(n_1551) );
NAND4xp25_ASAP7_75t_SL g1552 ( .A(n_1537), .B(n_1450), .C(n_1454), .D(n_1514), .Y(n_1552) );
AOI311xp33_ASAP7_75t_L g1553 ( .A1(n_1546), .A2(n_1545), .A3(n_1540), .B(n_1493), .C(n_1487), .Y(n_1553) );
NAND3xp33_ASAP7_75t_SL g1554 ( .A(n_1547), .B(n_1540), .C(n_1538), .Y(n_1554) );
OAI22xp5_ASAP7_75t_SL g1555 ( .A1(n_1549), .A2(n_1539), .B1(n_1468), .B2(n_1502), .Y(n_1555) );
INVx1_ASAP7_75t_L g1556 ( .A(n_1548), .Y(n_1556) );
OA22x2_ASAP7_75t_L g1557 ( .A1(n_1555), .A2(n_1550), .B1(n_1551), .B2(n_1552), .Y(n_1557) );
OA22x2_ASAP7_75t_L g1558 ( .A1(n_1553), .A2(n_1539), .B1(n_1486), .B2(n_1502), .Y(n_1558) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1556), .Y(n_1559) );
NOR3xp33_ASAP7_75t_L g1560 ( .A(n_1554), .B(n_1513), .C(n_1527), .Y(n_1560) );
INVxp33_ASAP7_75t_SL g1561 ( .A(n_1560), .Y(n_1561) );
OR4x1_ASAP7_75t_L g1562 ( .A(n_1559), .B(n_1489), .C(n_1503), .D(n_1506), .Y(n_1562) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1562), .Y(n_1563) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1561), .Y(n_1564) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1563), .Y(n_1565) );
OAI22xp33_ASAP7_75t_L g1566 ( .A1(n_1565), .A2(n_1557), .B1(n_1558), .B2(n_1564), .Y(n_1566) );
AOI21xp5_ASAP7_75t_L g1567 ( .A1(n_1566), .A2(n_1489), .B(n_1506), .Y(n_1567) );
endmodule