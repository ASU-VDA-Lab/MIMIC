module fake_jpeg_7818_n_80 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_80);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_80;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_8),
.B(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_21),
.Y(n_25)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_14),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_22),
.Y(n_27)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

AND2x6_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_3),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_34),
.B1(n_10),
.B2(n_15),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_22),
.B(n_27),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_10),
.B(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_23),
.A2(n_19),
.B1(n_16),
.B2(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_24),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_41),
.B1(n_10),
.B2(n_15),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_48),
.Y(n_53)
);

NOR4xp25_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_17),
.C(n_8),
.D(n_12),
.Y(n_47)
);

A2O1A1O1Ixp25_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_11),
.B(n_26),
.C(n_13),
.D(n_9),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_31),
.C(n_28),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_9),
.Y(n_57)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_44),
.C(n_4),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_57),
.B(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_31),
.B1(n_26),
.B2(n_11),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_58),
.Y(n_63)
);

A2O1A1O1Ixp25_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_26),
.B(n_11),
.C(n_5),
.D(n_6),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_SL g61 ( 
.A(n_59),
.B(n_51),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_55),
.B(n_4),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_62),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_59),
.B1(n_53),
.B2(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_69),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_3),
.B(n_4),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_62),
.Y(n_70)
);

OAI21x1_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_3),
.B(n_5),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_72),
.B(n_64),
.Y(n_73)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_74),
.B(n_75),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_61),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_71),
.C(n_5),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_7),
.C(n_77),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_7),
.Y(n_80)
);


endmodule