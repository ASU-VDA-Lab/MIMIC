module fake_netlist_6_3786_n_1816 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1816);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1816;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1605;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_5),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_170),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_10),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_7),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_56),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_141),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_149),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_119),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_98),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_13),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_97),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_100),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_22),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_49),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_151),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_19),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_127),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_52),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_52),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_140),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_1),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_53),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_115),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_91),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_46),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_99),
.Y(n_199)
);

INVxp33_ASAP7_75t_SL g200 ( 
.A(n_122),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_8),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_102),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_35),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_7),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_106),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_92),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_66),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_23),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_138),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_128),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_31),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_120),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_28),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_153),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_14),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_161),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_143),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_152),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_94),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_164),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_77),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_57),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_123),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_55),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_18),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_18),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_150),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_57),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_165),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_126),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_33),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_43),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_118),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_55),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_47),
.Y(n_237)
);

INVxp33_ASAP7_75t_SL g238 ( 
.A(n_5),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_111),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_41),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_56),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_41),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_95),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_12),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_42),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g246 ( 
.A(n_136),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_112),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_26),
.Y(n_248)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_40),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_1),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_8),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_74),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_61),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_110),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_43),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_6),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_158),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_33),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_86),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_145),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_129),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_134),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_70),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_75),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_109),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_54),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_107),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_34),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_60),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_46),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_23),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_51),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_53),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_137),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_79),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_89),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_84),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_47),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_116),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_16),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_121),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_117),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_113),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_80),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_64),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_4),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_76),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_103),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_142),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_162),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_159),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_0),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_65),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_108),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_22),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_124),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_90),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_35),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_26),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_169),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_15),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_48),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_32),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_20),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_30),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_44),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_156),
.Y(n_307)
);

CKINVDCx11_ASAP7_75t_R g308 ( 
.A(n_16),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_69),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_17),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_32),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_62),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_29),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_54),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_50),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_96),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_73),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_38),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_36),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_25),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_24),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_63),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_105),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_20),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_81),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_68),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_14),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_146),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_0),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_38),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_4),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_40),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_101),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_11),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_67),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_49),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_83),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_45),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_135),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_88),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_133),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_9),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_177),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_177),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_300),
.B(n_2),
.Y(n_345)
);

NOR2xp67_ASAP7_75t_L g346 ( 
.A(n_237),
.B(n_2),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_318),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_233),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_215),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_177),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_267),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_283),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_287),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_176),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_308),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_177),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_222),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_227),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_177),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_177),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_177),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_177),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_323),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_249),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_283),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_305),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_212),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_249),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_174),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_216),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_249),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_249),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_186),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_224),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_213),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_R g376 ( 
.A(n_217),
.B(n_167),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_249),
.B(n_3),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_200),
.B(n_3),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_223),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_230),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_236),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_242),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_220),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_225),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_176),
.B(n_6),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_244),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_249),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_231),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_249),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_249),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_255),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_335),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_342),
.Y(n_393)
);

BUFx6f_ASAP7_75t_SL g394 ( 
.A(n_220),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_235),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_173),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_256),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_239),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_192),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_192),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_243),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_258),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_173),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_299),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_299),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_342),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_272),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_273),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_191),
.B(n_9),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_175),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_280),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_195),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_200),
.B(n_10),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_220),
.Y(n_414)
);

INVxp33_ASAP7_75t_SL g415 ( 
.A(n_183),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_204),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_183),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_292),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_282),
.B(n_11),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_282),
.B(n_12),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_205),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_187),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_214),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_226),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_175),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_329),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_247),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_240),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_403),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_375),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_403),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_379),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_360),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_410),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_343),
.Y(n_435)
);

NAND2xp33_ASAP7_75t_R g436 ( 
.A(n_367),
.B(n_238),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_410),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_358),
.B(n_257),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_384),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_360),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_361),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_388),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_361),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_395),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_344),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_362),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_362),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_364),
.Y(n_448)
);

OA21x2_ASAP7_75t_L g449 ( 
.A1(n_377),
.A2(n_329),
.B(n_245),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_350),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_356),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_364),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_398),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_401),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_368),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_359),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_R g457 ( 
.A(n_369),
.B(n_259),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_352),
.B(n_178),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_371),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_366),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_368),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_372),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_387),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_358),
.B(n_260),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_389),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_390),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_427),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_367),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_370),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_370),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_374),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_385),
.B(n_181),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_396),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_374),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_425),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_385),
.B(n_335),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_348),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_383),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_425),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_392),
.B(n_178),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_426),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_426),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_412),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_416),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_421),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_349),
.Y(n_487)
);

NAND2xp33_ASAP7_75t_SL g488 ( 
.A(n_420),
.B(n_194),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_419),
.B(n_179),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_423),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_424),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_428),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_422),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_366),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_422),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_365),
.B(n_179),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_365),
.B(n_341),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_393),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_380),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_417),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_399),
.B(n_180),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_400),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_409),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_404),
.B(n_341),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_380),
.Y(n_505)
);

AND2x2_ASAP7_75t_SL g506 ( 
.A(n_449),
.B(n_378),
.Y(n_506)
);

OR2x6_ASAP7_75t_L g507 ( 
.A(n_503),
.B(n_346),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_438),
.B(n_415),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_477),
.B(n_440),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_435),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_477),
.B(n_381),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_477),
.B(n_381),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_440),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_445),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_487),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_464),
.B(n_414),
.Y(n_516)
);

CKINVDCx11_ASAP7_75t_R g517 ( 
.A(n_479),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_503),
.A2(n_345),
.B1(n_413),
.B2(n_347),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g519 ( 
.A(n_460),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_441),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_445),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_491),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_441),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_445),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_503),
.B(n_382),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_436),
.A2(n_363),
.B1(n_357),
.B2(n_408),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_503),
.A2(n_194),
.B1(n_234),
.B2(n_310),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_491),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_445),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_445),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_443),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_497),
.B(n_405),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_443),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_489),
.B(n_382),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_497),
.Y(n_535)
);

INVxp33_ASAP7_75t_L g536 ( 
.A(n_478),
.Y(n_536)
);

INVxp33_ASAP7_75t_L g537 ( 
.A(n_478),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_477),
.B(n_386),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_447),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_479),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_445),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_489),
.B(n_386),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_447),
.B(n_391),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_448),
.B(n_391),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_497),
.B(n_406),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_450),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_451),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_504),
.B(n_354),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_458),
.B(n_397),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_448),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_496),
.B(n_354),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_449),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_455),
.B(n_397),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_455),
.B(n_402),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_504),
.B(n_373),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_450),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_461),
.B(n_458),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_491),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_481),
.B(n_402),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_481),
.A2(n_418),
.B1(n_411),
.B2(n_408),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_491),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_504),
.B(n_407),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_461),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_450),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_498),
.B(n_172),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_462),
.B(n_407),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_462),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_449),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_498),
.B(n_411),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_496),
.B(n_418),
.Y(n_570)
);

AND2x6_ASAP7_75t_L g571 ( 
.A(n_433),
.B(n_219),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_463),
.B(n_262),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_459),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_502),
.B(n_409),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_463),
.B(n_466),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_466),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_501),
.B(n_394),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_459),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_433),
.B(n_263),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_502),
.B(n_182),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_451),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_449),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_433),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_SL g584 ( 
.A1(n_493),
.A2(n_394),
.B1(n_306),
.B2(n_248),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_488),
.A2(n_394),
.B1(n_238),
.B2(n_351),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_501),
.B(n_234),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_459),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_469),
.B(n_355),
.Y(n_588)
);

BUFx8_ASAP7_75t_SL g589 ( 
.A(n_460),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_446),
.B(n_265),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_446),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_451),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_465),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_451),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_446),
.B(n_274),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_491),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_500),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_446),
.B(n_275),
.Y(n_598)
);

BUFx4f_ASAP7_75t_L g599 ( 
.A(n_449),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_465),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_500),
.A2(n_353),
.B1(n_193),
.B2(n_184),
.Y(n_601)
);

NAND2xp33_ASAP7_75t_L g602 ( 
.A(n_473),
.B(n_181),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_470),
.B(n_355),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_465),
.Y(n_604)
);

NAND2x1p5_ASAP7_75t_L g605 ( 
.A(n_452),
.B(n_185),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_483),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_452),
.B(n_276),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_452),
.B(n_277),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_473),
.A2(n_310),
.B1(n_320),
.B2(n_338),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_484),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_457),
.B(n_376),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_484),
.Y(n_612)
);

BUFx4f_ASAP7_75t_L g613 ( 
.A(n_451),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_452),
.B(n_279),
.Y(n_614)
);

INVx4_ASAP7_75t_SL g615 ( 
.A(n_473),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_483),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_451),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_491),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_456),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_456),
.Y(n_620)
);

INVxp67_ASAP7_75t_SL g621 ( 
.A(n_456),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_456),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_456),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_473),
.B(n_285),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_456),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_L g626 ( 
.A(n_473),
.B(n_181),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_473),
.B(n_288),
.Y(n_627)
);

AND2x2_ASAP7_75t_SL g628 ( 
.A(n_494),
.B(n_219),
.Y(n_628)
);

AND2x6_ASAP7_75t_L g629 ( 
.A(n_486),
.B(n_181),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_483),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_430),
.B(n_189),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_432),
.B(n_311),
.Y(n_632)
);

AND2x6_ASAP7_75t_L g633 ( 
.A(n_486),
.B(n_181),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_473),
.B(n_476),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_490),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_471),
.B(n_281),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_473),
.B(n_289),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_483),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_483),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_472),
.B(n_180),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_476),
.B(n_290),
.Y(n_641)
);

AND3x2_ASAP7_75t_L g642 ( 
.A(n_494),
.B(n_246),
.C(n_199),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_483),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_476),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_439),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_467),
.B(n_320),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_467),
.B(n_241),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_442),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_492),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_476),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_485),
.B(n_291),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_475),
.B(n_184),
.Y(n_652)
);

AND2x2_ASAP7_75t_SL g653 ( 
.A(n_493),
.B(n_296),
.Y(n_653)
);

AND2x4_ASAP7_75t_SL g654 ( 
.A(n_495),
.B(n_281),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_557),
.B(n_202),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_535),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_535),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_534),
.B(n_203),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_542),
.B(n_206),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_551),
.B(n_495),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_510),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_508),
.B(n_551),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_597),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_509),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_653),
.B(n_499),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_610),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_653),
.B(n_628),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_543),
.B(n_544),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_548),
.B(n_505),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_553),
.B(n_198),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_506),
.B(n_296),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_570),
.B(n_211),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_506),
.B(n_296),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_531),
.B(n_218),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_599),
.B(n_296),
.Y(n_675)
);

INVxp67_ASAP7_75t_L g676 ( 
.A(n_597),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_552),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_531),
.B(n_221),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_650),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_612),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_533),
.B(n_539),
.Y(n_681)
);

OAI22xp33_ASAP7_75t_L g682 ( 
.A1(n_586),
.A2(n_301),
.B1(n_209),
.B2(n_228),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_533),
.B(n_229),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_554),
.B(n_492),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_539),
.B(n_232),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_513),
.B(n_253),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_548),
.B(n_444),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_532),
.B(n_485),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_635),
.Y(n_689)
);

AOI221xp5_ASAP7_75t_L g690 ( 
.A1(n_518),
.A2(n_250),
.B1(n_201),
.B2(n_187),
.C(n_295),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_628),
.A2(n_293),
.B1(n_340),
.B2(n_297),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_525),
.B(n_453),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_599),
.B(n_650),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_599),
.B(n_296),
.Y(n_694)
);

NOR3xp33_ASAP7_75t_L g695 ( 
.A(n_516),
.B(n_454),
.C(n_468),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_520),
.B(n_254),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_650),
.B(n_261),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_546),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_511),
.A2(n_512),
.B1(n_538),
.B2(n_507),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_560),
.B(n_210),
.C(n_340),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_566),
.B(n_188),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_523),
.B(n_264),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_549),
.B(n_188),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_649),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_634),
.B(n_269),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_552),
.B(n_284),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_532),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_519),
.B(n_201),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_SL g709 ( 
.A(n_648),
.B(n_281),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_568),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_546),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_556),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_550),
.B(n_317),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_559),
.A2(n_207),
.B1(n_190),
.B2(n_337),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_563),
.B(n_325),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_644),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_545),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_545),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_507),
.A2(n_586),
.B1(n_568),
.B2(n_582),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_567),
.B(n_333),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_576),
.B(n_575),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_582),
.B(n_339),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_569),
.B(n_190),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_583),
.B(n_591),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_583),
.B(n_485),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_621),
.A2(n_482),
.B(n_480),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_640),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_L g728 ( 
.A(n_584),
.B(n_286),
.C(n_251),
.Y(n_728)
);

OAI221xp5_ASAP7_75t_L g729 ( 
.A1(n_527),
.A2(n_268),
.B1(n_302),
.B2(n_298),
.C(n_278),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_591),
.B(n_480),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_L g731 ( 
.A(n_571),
.B(n_193),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_556),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_572),
.B(n_480),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_555),
.B(n_474),
.Y(n_734)
);

BUFx8_ASAP7_75t_L g735 ( 
.A(n_562),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_507),
.A2(n_586),
.B1(n_562),
.B2(n_609),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_641),
.B(n_482),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_507),
.A2(n_196),
.B1(n_312),
.B2(n_316),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_577),
.B(n_482),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_586),
.A2(n_196),
.B1(n_197),
.B2(n_207),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_579),
.B(n_429),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_555),
.B(n_474),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_647),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_571),
.A2(n_319),
.B1(n_321),
.B2(n_266),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_SL g745 ( 
.A(n_645),
.B(n_588),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_569),
.A2(n_197),
.B1(n_208),
.B2(n_210),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_590),
.B(n_431),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_595),
.A2(n_607),
.B(n_598),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_652),
.B(n_208),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_608),
.A2(n_252),
.B1(n_297),
.B2(n_307),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_647),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_565),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_565),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_571),
.A2(n_330),
.B1(n_270),
.B2(n_271),
.Y(n_754)
);

OR2x6_ASAP7_75t_L g755 ( 
.A(n_574),
.B(n_636),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_571),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_614),
.B(n_431),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_571),
.A2(n_303),
.B1(n_336),
.B2(n_295),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_651),
.B(n_434),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_622),
.B(n_434),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_565),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_615),
.B(n_252),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_580),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_645),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_536),
.B(n_250),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_611),
.B(n_307),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_564),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_615),
.B(n_322),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_622),
.B(n_437),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_654),
.B(n_322),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_571),
.A2(n_324),
.B1(n_304),
.B2(n_334),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_521),
.B(n_437),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_580),
.A2(n_337),
.B(n_309),
.C(n_312),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_615),
.B(n_605),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_564),
.Y(n_775)
);

NAND3xp33_ASAP7_75t_L g776 ( 
.A(n_601),
.B(n_316),
.C(n_309),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_521),
.B(n_326),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_L g778 ( 
.A(n_605),
.B(n_326),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_654),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_521),
.B(n_328),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_541),
.B(n_328),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_615),
.B(n_294),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_646),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_573),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_536),
.B(n_334),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_541),
.B(n_294),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_646),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_605),
.B(n_294),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_573),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_618),
.B(n_332),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_541),
.B(n_332),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_618),
.B(n_606),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_642),
.B(n_78),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_578),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_578),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_581),
.B(n_331),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_537),
.B(n_331),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_602),
.A2(n_327),
.B1(n_324),
.B2(n_315),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_SL g799 ( 
.A(n_603),
.B(n_327),
.Y(n_799)
);

A2O1A1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_587),
.A2(n_315),
.B(n_314),
.C(n_313),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_537),
.B(n_314),
.Y(n_801)
);

NOR2xp67_ASAP7_75t_SL g802 ( 
.A(n_522),
.B(n_313),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_585),
.B(n_304),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_587),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_606),
.B(n_58),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_593),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_593),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_581),
.B(n_166),
.Y(n_808)
);

NAND3xp33_ASAP7_75t_L g809 ( 
.A(n_526),
.B(n_624),
.C(n_637),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_581),
.B(n_163),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_631),
.B(n_13),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_600),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_631),
.B(n_15),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_594),
.B(n_17),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_600),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_594),
.B(n_19),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_667),
.A2(n_602),
.B(n_626),
.C(n_627),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_727),
.B(n_632),
.Y(n_818)
);

CKINVDCx8_ASAP7_75t_R g819 ( 
.A(n_764),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_716),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_SL g821 ( 
.A(n_662),
.B(n_540),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_668),
.B(n_594),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_688),
.Y(n_823)
);

OAI21xp33_ASAP7_75t_L g824 ( 
.A1(n_662),
.A2(n_632),
.B(n_540),
.Y(n_824)
);

AOI21x1_ASAP7_75t_L g825 ( 
.A1(n_675),
.A2(n_694),
.B(n_673),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_733),
.A2(n_613),
.B(n_514),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_668),
.B(n_623),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_735),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_688),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_737),
.A2(n_613),
.B(n_675),
.Y(n_830)
);

A2O1A1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_670),
.A2(n_626),
.B(n_604),
.C(n_623),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_735),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_SL g833 ( 
.A1(n_671),
.A2(n_643),
.B(n_616),
.C(n_630),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_694),
.A2(n_613),
.B(n_530),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_677),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_671),
.A2(n_604),
.B(n_630),
.C(n_643),
.Y(n_836)
);

AOI21x1_ASAP7_75t_L g837 ( 
.A1(n_673),
.A2(n_616),
.B(n_617),
.Y(n_837)
);

AO21x1_ASAP7_75t_L g838 ( 
.A1(n_719),
.A2(n_514),
.B(n_524),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_664),
.B(n_623),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_684),
.B(n_721),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_748),
.A2(n_693),
.B(n_741),
.Y(n_841)
);

INVx11_ASAP7_75t_L g842 ( 
.A(n_663),
.Y(n_842)
);

BUFx4f_ASAP7_75t_L g843 ( 
.A(n_755),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_684),
.B(n_617),
.Y(n_844)
);

OR2x6_ASAP7_75t_SL g845 ( 
.A(n_811),
.B(n_517),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_665),
.B(n_515),
.Y(n_846)
);

AO22x1_ASAP7_75t_L g847 ( 
.A1(n_803),
.A2(n_633),
.B1(n_629),
.B2(n_589),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_679),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_658),
.A2(n_515),
.B1(n_625),
.B2(n_620),
.Y(n_849)
);

AND2x2_ASAP7_75t_SL g850 ( 
.A(n_813),
.B(n_589),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_679),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_659),
.A2(n_638),
.B(n_620),
.C(n_625),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_693),
.A2(n_514),
.B(n_524),
.Y(n_853)
);

A2O1A1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_670),
.A2(n_619),
.B(n_638),
.C(n_528),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_672),
.B(n_619),
.Y(n_855)
);

AOI21x1_ASAP7_75t_L g856 ( 
.A1(n_792),
.A2(n_524),
.B(n_529),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_749),
.B(n_638),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_656),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_809),
.A2(n_558),
.B1(n_528),
.B2(n_522),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_716),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_676),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_747),
.A2(n_529),
.B(n_530),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_699),
.A2(n_547),
.B1(n_592),
.B2(n_639),
.Y(n_863)
);

O2A1O1Ixp5_ASAP7_75t_L g864 ( 
.A1(n_739),
.A2(n_722),
.B(n_706),
.C(n_705),
.Y(n_864)
);

NOR3xp33_ASAP7_75t_L g865 ( 
.A(n_665),
.B(n_517),
.C(n_592),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_677),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_706),
.A2(n_547),
.B(n_592),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_757),
.A2(n_547),
.B(n_639),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_677),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_661),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_749),
.B(n_561),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_701),
.B(n_681),
.Y(n_872)
);

OR2x6_ASAP7_75t_L g873 ( 
.A(n_779),
.B(n_596),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_758),
.A2(n_596),
.B1(n_561),
.B2(n_558),
.Y(n_874)
);

AND2x6_ASAP7_75t_L g875 ( 
.A(n_677),
.B(n_522),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_701),
.B(n_561),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_774),
.A2(n_639),
.B(n_561),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_669),
.B(n_522),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_734),
.B(n_596),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_742),
.B(n_596),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_774),
.A2(n_558),
.B(n_528),
.Y(n_881)
);

INVx11_ASAP7_75t_L g882 ( 
.A(n_745),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_710),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_657),
.Y(n_884)
);

OAI21x1_ASAP7_75t_L g885 ( 
.A1(n_724),
.A2(n_558),
.B(n_528),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_710),
.Y(n_886)
);

AOI21x1_ASAP7_75t_L g887 ( 
.A1(n_792),
.A2(n_558),
.B(n_528),
.Y(n_887)
);

AOI21x1_ASAP7_75t_L g888 ( 
.A1(n_722),
.A2(n_522),
.B(n_633),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_759),
.A2(n_633),
.B(n_629),
.Y(n_889)
);

NOR2x1_ASAP7_75t_L g890 ( 
.A(n_692),
.B(n_633),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_710),
.B(n_633),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_772),
.A2(n_633),
.B(n_629),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_666),
.Y(n_893)
);

NOR2xp67_ASAP7_75t_L g894 ( 
.A(n_766),
.B(n_71),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_680),
.Y(n_895)
);

NAND3xp33_ASAP7_75t_L g896 ( 
.A(n_703),
.B(n_21),
.C(n_24),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_799),
.B(n_21),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_703),
.A2(n_629),
.B(n_27),
.C(n_28),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_743),
.B(n_629),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_725),
.A2(n_629),
.B(n_82),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_660),
.B(n_25),
.Y(n_901)
);

AO22x1_ASAP7_75t_L g902 ( 
.A1(n_803),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_902)
);

AO32x1_ASAP7_75t_L g903 ( 
.A1(n_736),
.A2(n_31),
.A3(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_777),
.A2(n_93),
.B(n_157),
.Y(n_904)
);

CKINVDCx6p67_ASAP7_75t_R g905 ( 
.A(n_687),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_780),
.A2(n_781),
.B(n_778),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_655),
.B(n_37),
.Y(n_907)
);

AOI22x1_ASAP7_75t_L g908 ( 
.A1(n_689),
.A2(n_104),
.B1(n_155),
.B2(n_154),
.Y(n_908)
);

OA21x2_ASAP7_75t_L g909 ( 
.A1(n_730),
.A2(n_85),
.B(n_148),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_698),
.Y(n_910)
);

AOI22x1_ASAP7_75t_L g911 ( 
.A1(n_704),
.A2(n_72),
.B1(n_147),
.B2(n_139),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_751),
.B(n_39),
.Y(n_912)
);

INVxp67_ASAP7_75t_SL g913 ( 
.A(n_756),
.Y(n_913)
);

OAI21x1_ASAP7_75t_L g914 ( 
.A1(n_808),
.A2(n_59),
.B(n_132),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_760),
.A2(n_160),
.B(n_130),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_769),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_723),
.B(n_783),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_723),
.B(n_39),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_705),
.A2(n_125),
.B(n_114),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_787),
.B(n_42),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_785),
.B(n_44),
.Y(n_921)
);

NAND2xp33_ASAP7_75t_L g922 ( 
.A(n_756),
.B(n_87),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_752),
.B(n_45),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_766),
.B(n_48),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_753),
.A2(n_50),
.B(n_51),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_789),
.Y(n_926)
);

INVx4_ASAP7_75t_L g927 ( 
.A(n_755),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_726),
.A2(n_707),
.B(n_717),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_761),
.B(n_763),
.Y(n_929)
);

INVx11_ASAP7_75t_L g930 ( 
.A(n_695),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_762),
.A2(n_768),
.B(n_796),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_708),
.B(n_770),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_718),
.B(n_674),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_785),
.Y(n_934)
);

INVx1_ASAP7_75t_SL g935 ( 
.A(n_765),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_793),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_791),
.A2(n_810),
.B(n_697),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_678),
.B(n_683),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_758),
.A2(n_771),
.B1(n_691),
.B2(n_754),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_697),
.A2(n_731),
.B(n_782),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_685),
.B(n_720),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_814),
.A2(n_816),
.B(n_812),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_686),
.B(n_715),
.Y(n_943)
);

AOI21xp33_ASAP7_75t_L g944 ( 
.A1(n_771),
.A2(n_816),
.B(n_814),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_806),
.Y(n_945)
);

BUFx12f_ASAP7_75t_L g946 ( 
.A(n_793),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_696),
.B(n_702),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_755),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_797),
.B(n_801),
.Y(n_949)
);

AO21x1_ASAP7_75t_L g950 ( 
.A1(n_788),
.A2(n_805),
.B(n_790),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_713),
.B(n_807),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_711),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_790),
.A2(n_773),
.B(n_815),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_770),
.B(n_700),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_712),
.A2(n_775),
.B(n_804),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_782),
.A2(n_786),
.B(n_795),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_797),
.B(n_801),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_732),
.B(n_767),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_784),
.B(n_794),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_788),
.A2(n_738),
.B1(n_750),
.B2(n_776),
.Y(n_960)
);

AOI21x1_ASAP7_75t_L g961 ( 
.A1(n_805),
.A2(n_802),
.B(n_740),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_744),
.A2(n_754),
.B(n_800),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_746),
.B(n_714),
.Y(n_963)
);

AO21x1_ASAP7_75t_L g964 ( 
.A1(n_728),
.A2(n_682),
.B(n_709),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_744),
.B(n_690),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_798),
.B(n_729),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_798),
.B(n_668),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_667),
.A2(n_673),
.B(n_671),
.C(n_658),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_733),
.A2(n_613),
.B(n_737),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_733),
.A2(n_613),
.B(n_737),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_669),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_716),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_688),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_671),
.A2(n_599),
.B(n_673),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_727),
.B(n_662),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_724),
.A2(n_748),
.B(n_792),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_733),
.A2(n_613),
.B(n_737),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_688),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_679),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_727),
.B(n_662),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_688),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_727),
.B(n_662),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_733),
.A2(n_613),
.B(n_737),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_677),
.Y(n_984)
);

NOR2xp67_ASAP7_75t_L g985 ( 
.A(n_764),
.B(n_727),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_727),
.B(n_662),
.Y(n_986)
);

AND2x6_ASAP7_75t_L g987 ( 
.A(n_677),
.B(n_710),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_733),
.A2(n_613),
.B(n_737),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_733),
.A2(n_613),
.B(n_737),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_663),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_677),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_688),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_671),
.A2(n_599),
.B(n_673),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_733),
.A2(n_613),
.B(n_737),
.Y(n_994)
);

AOI21x1_ASAP7_75t_L g995 ( 
.A1(n_675),
.A2(n_694),
.B(n_673),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_664),
.B(n_668),
.Y(n_996)
);

OAI21x1_ASAP7_75t_L g997 ( 
.A1(n_885),
.A2(n_887),
.B(n_856),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_841),
.A2(n_830),
.B(n_996),
.Y(n_998)
);

CKINVDCx6p67_ASAP7_75t_R g999 ( 
.A(n_946),
.Y(n_999)
);

OAI21x1_ASAP7_75t_L g1000 ( 
.A1(n_976),
.A2(n_853),
.B(n_837),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_957),
.A2(n_918),
.B(n_963),
.C(n_840),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_881),
.A2(n_877),
.B(n_836),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_834),
.A2(n_956),
.B(n_888),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_996),
.A2(n_968),
.B(n_876),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_871),
.A2(n_970),
.B(n_969),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_936),
.B(n_878),
.Y(n_1006)
);

INVx6_ASAP7_75t_L g1007 ( 
.A(n_936),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_840),
.B(n_872),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_937),
.A2(n_955),
.B(n_826),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_949),
.B(n_934),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_974),
.A2(n_993),
.B(n_944),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_977),
.A2(n_988),
.B(n_983),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_893),
.Y(n_1013)
);

OR2x6_ASAP7_75t_L g1014 ( 
.A(n_936),
.B(n_927),
.Y(n_1014)
);

OA21x2_ASAP7_75t_L g1015 ( 
.A1(n_974),
.A2(n_993),
.B(n_942),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_967),
.A2(n_954),
.B(n_944),
.C(n_939),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_975),
.A2(n_982),
.B1(n_980),
.B2(n_986),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_916),
.B(n_917),
.Y(n_1018)
);

AOI211x1_ASAP7_75t_L g1019 ( 
.A1(n_902),
.A2(n_939),
.B(n_965),
.C(n_924),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_SL g1020 ( 
.A1(n_818),
.A2(n_828),
.B1(n_832),
.B2(n_897),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_965),
.A2(n_966),
.B1(n_960),
.B2(n_894),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_835),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_SL g1023 ( 
.A1(n_874),
.A2(n_984),
.B(n_866),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_955),
.A2(n_867),
.B(n_931),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_823),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_940),
.A2(n_906),
.B(n_989),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_819),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_895),
.Y(n_1028)
);

NAND2x1_ASAP7_75t_L g1029 ( 
.A(n_987),
.B(n_875),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_929),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_966),
.A2(n_932),
.B(n_921),
.C(n_864),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_994),
.A2(n_938),
.B(n_822),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_971),
.A2(n_821),
.B1(n_846),
.B2(n_824),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_829),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_835),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_827),
.B(n_941),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_849),
.A2(n_901),
.B(n_907),
.C(n_920),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_825),
.A2(n_995),
.B(n_962),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_928),
.A2(n_862),
.B(n_868),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_953),
.A2(n_933),
.B(n_947),
.C(n_943),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_874),
.A2(n_859),
.B(n_839),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_857),
.A2(n_855),
.B(n_879),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_953),
.A2(n_817),
.B(n_923),
.C(n_992),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_973),
.A2(n_978),
.B(n_981),
.C(n_843),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_926),
.Y(n_1045)
);

O2A1O1Ixp5_ASAP7_75t_L g1046 ( 
.A1(n_950),
.A2(n_942),
.B(n_838),
.C(n_961),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_945),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_844),
.B(n_880),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_843),
.A2(n_912),
.B1(n_896),
.B2(n_882),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_831),
.A2(n_854),
.B(n_852),
.Y(n_1050)
);

AO21x2_ASAP7_75t_L g1051 ( 
.A1(n_863),
.A2(n_833),
.B(n_951),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_848),
.B(n_851),
.Y(n_1052)
);

INVx3_ASAP7_75t_SL g1053 ( 
.A(n_905),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_958),
.A2(n_959),
.B(n_914),
.Y(n_1054)
);

OA22x2_ASAP7_75t_L g1055 ( 
.A1(n_935),
.A2(n_948),
.B1(n_990),
.B2(n_861),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_979),
.B(n_987),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_858),
.Y(n_1057)
);

INVxp67_ASAP7_75t_SL g1058 ( 
.A(n_835),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_935),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_948),
.A2(n_884),
.B1(n_979),
.B2(n_869),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_899),
.A2(n_889),
.B(n_892),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_913),
.A2(n_891),
.B(n_899),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_927),
.B(n_984),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_SL g1064 ( 
.A1(n_925),
.A2(n_904),
.B(n_919),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_820),
.A2(n_972),
.B(n_860),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_952),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_870),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_987),
.B(n_886),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_849),
.A2(n_910),
.B(n_898),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_964),
.A2(n_865),
.B1(n_821),
.B2(n_890),
.Y(n_1070)
);

AO31x2_ASAP7_75t_L g1071 ( 
.A1(n_900),
.A2(n_915),
.A3(n_903),
.B(n_909),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_845),
.Y(n_1072)
);

OA21x2_ASAP7_75t_L g1073 ( 
.A1(n_908),
.A2(n_911),
.B(n_903),
.Y(n_1073)
);

NOR2x1_ASAP7_75t_SL g1074 ( 
.A(n_866),
.B(n_883),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_909),
.A2(n_875),
.B(n_873),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_875),
.A2(n_873),
.B(n_922),
.Y(n_1076)
);

OAI21xp33_ASAP7_75t_L g1077 ( 
.A1(n_985),
.A2(n_850),
.B(n_873),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_866),
.B(n_883),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_869),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_842),
.B(n_930),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_869),
.B(n_883),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_991),
.B(n_875),
.Y(n_1082)
);

AO31x2_ASAP7_75t_L g1083 ( 
.A1(n_903),
.A2(n_838),
.A3(n_950),
.B(n_854),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_991),
.B(n_847),
.Y(n_1084)
);

AO31x2_ASAP7_75t_L g1085 ( 
.A1(n_991),
.A2(n_838),
.A3(n_950),
.B(n_854),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_861),
.Y(n_1086)
);

NAND2x1p5_ASAP7_75t_L g1087 ( 
.A(n_984),
.B(n_835),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_840),
.B(n_996),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_835),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_835),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_885),
.A2(n_887),
.B(n_856),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_974),
.A2(n_993),
.B(n_944),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_893),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_885),
.A2(n_887),
.B(n_856),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_987),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_987),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_885),
.A2(n_887),
.B(n_856),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_840),
.A2(n_996),
.B1(n_967),
.B2(n_939),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_893),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_975),
.B(n_980),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_885),
.A2(n_887),
.B(n_856),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_819),
.Y(n_1102)
);

AO21x1_ASAP7_75t_L g1103 ( 
.A1(n_944),
.A2(n_918),
.B(n_967),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_835),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_885),
.A2(n_887),
.B(n_856),
.Y(n_1105)
);

NAND2x1_ASAP7_75t_L g1106 ( 
.A(n_987),
.B(n_875),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_840),
.B(n_996),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_974),
.A2(n_993),
.B(n_944),
.Y(n_1108)
);

HB1xp67_ASAP7_75t_L g1109 ( 
.A(n_861),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_840),
.B(n_996),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_840),
.A2(n_996),
.B1(n_967),
.B2(n_939),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_838),
.A2(n_950),
.A3(n_854),
.B(n_831),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_840),
.B(n_996),
.Y(n_1113)
);

NAND2x2_ASAP7_75t_L g1114 ( 
.A(n_920),
.B(n_779),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_885),
.A2(n_887),
.B(n_856),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_967),
.A2(n_918),
.B(n_957),
.C(n_924),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_835),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_823),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_975),
.B(n_980),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_885),
.A2(n_887),
.B(n_856),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_835),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_835),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_840),
.B(n_996),
.Y(n_1123)
);

AO31x2_ASAP7_75t_L g1124 ( 
.A1(n_838),
.A2(n_950),
.A3(n_854),
.B(n_831),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_885),
.A2(n_887),
.B(n_856),
.Y(n_1125)
);

AO21x1_ASAP7_75t_L g1126 ( 
.A1(n_944),
.A2(n_918),
.B(n_967),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_885),
.A2(n_887),
.B(n_856),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_935),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_957),
.B(n_996),
.Y(n_1129)
);

AND2x2_ASAP7_75t_SL g1130 ( 
.A(n_821),
.B(n_628),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_975),
.B(n_980),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_885),
.A2(n_887),
.B(n_856),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_957),
.B(n_996),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_885),
.A2(n_887),
.B(n_856),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_974),
.A2(n_993),
.B(n_944),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_823),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_840),
.B(n_996),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_957),
.A2(n_918),
.B(n_963),
.C(n_668),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_840),
.B(n_996),
.Y(n_1139)
);

BUFx4_ASAP7_75t_SL g1140 ( 
.A(n_1027),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_1059),
.Y(n_1141)
);

OR2x6_ASAP7_75t_L g1142 ( 
.A(n_1014),
.B(n_1095),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1100),
.B(n_1131),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1028),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_1014),
.B(n_1063),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_1128),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1008),
.B(n_1088),
.Y(n_1147)
);

BUFx5_ASAP7_75t_L g1148 ( 
.A(n_1078),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1093),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1099),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_1022),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1008),
.B(n_1088),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1032),
.A2(n_998),
.B(n_1040),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1138),
.A2(n_1001),
.B1(n_1113),
.B2(n_1123),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_SL g1155 ( 
.A1(n_1020),
.A2(n_1119),
.B1(n_1130),
.B2(n_1017),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1107),
.A2(n_1139),
.B1(n_1123),
.B2(n_1113),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1107),
.B(n_1110),
.Y(n_1157)
);

AND2x6_ASAP7_75t_L g1158 ( 
.A(n_1078),
.B(n_1081),
.Y(n_1158)
);

BUFx12f_ASAP7_75t_L g1159 ( 
.A(n_1102),
.Y(n_1159)
);

OAI22xp33_ASAP7_75t_SL g1160 ( 
.A1(n_1129),
.A2(n_1133),
.B1(n_1137),
.B2(n_1110),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1128),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1109),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1137),
.A2(n_1139),
.B1(n_1018),
.B2(n_1016),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_1086),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1018),
.B(n_1036),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1055),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1032),
.A2(n_998),
.B(n_1004),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_1055),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_1079),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1036),
.B(n_1098),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_1010),
.B(n_1033),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1098),
.B(n_1111),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1030),
.B(n_1049),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_1060),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_1014),
.B(n_1095),
.Y(n_1175)
);

OR2x6_ASAP7_75t_L g1176 ( 
.A(n_1096),
.B(n_1023),
.Y(n_1176)
);

NOR2x1_ASAP7_75t_R g1177 ( 
.A(n_1072),
.B(n_1007),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1063),
.B(n_1006),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1045),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1111),
.B(n_1019),
.Y(n_1180)
);

INVxp67_ASAP7_75t_SL g1181 ( 
.A(n_1074),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1006),
.B(n_1025),
.Y(n_1182)
);

NOR2xp67_ASAP7_75t_L g1183 ( 
.A(n_1080),
.B(n_1049),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1118),
.B(n_1136),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1057),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1021),
.A2(n_1116),
.B1(n_1031),
.B2(n_1047),
.Y(n_1186)
);

NOR2xp67_ASAP7_75t_L g1187 ( 
.A(n_1067),
.B(n_1066),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1081),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1034),
.B(n_1044),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1096),
.Y(n_1190)
);

INVx4_ASAP7_75t_L g1191 ( 
.A(n_1022),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1037),
.A2(n_1021),
.B(n_1135),
.C(n_1092),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1048),
.B(n_1103),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1077),
.A2(n_1070),
.B1(n_1126),
.B2(n_1060),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1048),
.B(n_1042),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1065),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1026),
.A2(n_1005),
.B(n_1012),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1022),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1053),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1005),
.A2(n_1012),
.B(n_1043),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1117),
.B(n_1122),
.Y(n_1201)
);

INVx1_ASAP7_75t_SL g1202 ( 
.A(n_1035),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1007),
.B(n_1069),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1007),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1011),
.A2(n_1108),
.B1(n_1015),
.B2(n_1069),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1039),
.A2(n_1050),
.B(n_1024),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1050),
.A2(n_1038),
.B(n_1009),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1015),
.B(n_1052),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_999),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1046),
.A2(n_1041),
.B(n_1062),
.C(n_1038),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1035),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1058),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_1035),
.Y(n_1213)
);

BUFx12f_ASAP7_75t_L g1214 ( 
.A(n_1089),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1114),
.A2(n_1084),
.B1(n_1073),
.B2(n_1122),
.Y(n_1215)
);

NOR2x1_ASAP7_75t_L g1216 ( 
.A(n_1082),
.B(n_1068),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1089),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1089),
.B(n_1090),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1090),
.B(n_1104),
.Y(n_1219)
);

CKINVDCx11_ASAP7_75t_R g1220 ( 
.A(n_1104),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1104),
.B(n_1121),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1121),
.Y(n_1222)
);

INVx1_ASAP7_75t_SL g1223 ( 
.A(n_1121),
.Y(n_1223)
);

CKINVDCx8_ASAP7_75t_R g1224 ( 
.A(n_1087),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1029),
.A2(n_1106),
.B1(n_1082),
.B2(n_1056),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1076),
.B(n_1068),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1087),
.B(n_1085),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1051),
.B(n_1061),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1064),
.A2(n_1061),
.B(n_1003),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1085),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1054),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1085),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1075),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1000),
.A2(n_1002),
.B(n_997),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1091),
.A2(n_1101),
.B(n_1134),
.Y(n_1235)
);

AND2x2_ASAP7_75t_SL g1236 ( 
.A(n_1083),
.B(n_1124),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1112),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1124),
.B(n_1083),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1083),
.B(n_1071),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1071),
.B(n_1094),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1097),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1105),
.B(n_1115),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1120),
.B(n_1125),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1127),
.Y(n_1244)
);

OR2x2_ASAP7_75t_L g1245 ( 
.A(n_1132),
.B(n_660),
.Y(n_1245)
);

OAI21xp33_ASAP7_75t_L g1246 ( 
.A1(n_1138),
.A2(n_957),
.B(n_662),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1100),
.B(n_1131),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1013),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1022),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1138),
.A2(n_1001),
.B1(n_1107),
.B2(n_1088),
.Y(n_1250)
);

NOR2x1_ASAP7_75t_SL g1251 ( 
.A(n_1095),
.B(n_1096),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1138),
.A2(n_1001),
.B1(n_1107),
.B2(n_1088),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1008),
.B(n_1088),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_1014),
.B(n_1063),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1119),
.B(n_975),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1130),
.B(n_821),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1027),
.Y(n_1257)
);

O2A1O1Ixp5_ASAP7_75t_L g1258 ( 
.A1(n_1138),
.A2(n_918),
.B(n_944),
.C(n_957),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1059),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1008),
.B(n_1088),
.Y(n_1260)
);

NOR2xp67_ASAP7_75t_L g1261 ( 
.A(n_1080),
.B(n_764),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1014),
.B(n_1063),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1027),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1013),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1014),
.B(n_1063),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1008),
.B(n_1088),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1138),
.A2(n_1001),
.B1(n_1107),
.B2(n_1088),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1095),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1014),
.B(n_1063),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1053),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1130),
.A2(n_963),
.B1(n_957),
.B2(n_918),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1008),
.B(n_1088),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1059),
.Y(n_1273)
);

NOR2xp67_ASAP7_75t_L g1274 ( 
.A(n_1080),
.B(n_764),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1059),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1013),
.Y(n_1276)
);

INVx5_ASAP7_75t_L g1277 ( 
.A(n_1095),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1100),
.B(n_1131),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1013),
.Y(n_1279)
);

INVx11_ASAP7_75t_L g1280 ( 
.A(n_1214),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1185),
.Y(n_1281)
);

BUFx2_ASAP7_75t_SL g1282 ( 
.A(n_1277),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1155),
.A2(n_1255),
.B1(n_1172),
.B2(n_1173),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1248),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1146),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1276),
.Y(n_1286)
);

AOI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1234),
.A2(n_1206),
.B(n_1235),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1203),
.B(n_1165),
.Y(n_1288)
);

AO21x1_ASAP7_75t_L g1289 ( 
.A1(n_1172),
.A2(n_1186),
.B(n_1154),
.Y(n_1289)
);

CKINVDCx20_ASAP7_75t_R g1290 ( 
.A(n_1209),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1144),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1149),
.Y(n_1292)
);

AOI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1271),
.A2(n_1183),
.B1(n_1246),
.B2(n_1256),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1150),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1217),
.Y(n_1295)
);

AOI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1171),
.A2(n_1261),
.B1(n_1274),
.B2(n_1247),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1220),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1277),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1179),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1264),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1143),
.B(n_1278),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1161),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1279),
.Y(n_1303)
);

AOI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1154),
.A2(n_1252),
.B1(n_1267),
.B2(n_1250),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1166),
.A2(n_1168),
.B1(n_1189),
.B2(n_1267),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1165),
.B(n_1147),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1184),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1277),
.Y(n_1308)
);

OR2x6_ASAP7_75t_L g1309 ( 
.A(n_1176),
.B(n_1207),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1187),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1147),
.B(n_1152),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_1257),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1145),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1275),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_1145),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1176),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1140),
.Y(n_1317)
);

OR2x6_ASAP7_75t_L g1318 ( 
.A(n_1176),
.B(n_1186),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1190),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1152),
.B(n_1253),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1254),
.B(n_1262),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1253),
.B(n_1260),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1260),
.B(n_1266),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1189),
.A2(n_1252),
.B1(n_1250),
.B2(n_1163),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_SL g1325 ( 
.A1(n_1170),
.A2(n_1163),
.B1(n_1180),
.B2(n_1160),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1222),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1229),
.A2(n_1167),
.B(n_1197),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1158),
.Y(n_1328)
);

INVx6_ASAP7_75t_L g1329 ( 
.A(n_1142),
.Y(n_1329)
);

BUFx2_ASAP7_75t_R g1330 ( 
.A(n_1263),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1212),
.Y(n_1331)
);

BUFx12f_ASAP7_75t_L g1332 ( 
.A(n_1159),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1156),
.A2(n_1182),
.B1(n_1178),
.B2(n_1194),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1266),
.A2(n_1272),
.B1(n_1157),
.B2(n_1156),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1245),
.Y(n_1335)
);

AO21x1_ASAP7_75t_L g1336 ( 
.A1(n_1170),
.A2(n_1228),
.B(n_1205),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1254),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1174),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1272),
.B(n_1157),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1208),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1162),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1208),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1216),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1200),
.A2(n_1153),
.B(n_1243),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1258),
.A2(n_1195),
.B(n_1192),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1180),
.B(n_1236),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1193),
.B(n_1239),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1243),
.A2(n_1231),
.B(n_1196),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1227),
.Y(n_1349)
);

AO21x2_ASAP7_75t_L g1350 ( 
.A1(n_1210),
.A2(n_1240),
.B(n_1193),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1215),
.B(n_1232),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1158),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_SL g1353 ( 
.A1(n_1205),
.A2(n_1164),
.B1(n_1273),
.B2(n_1259),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1178),
.B(n_1148),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1141),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1226),
.A2(n_1195),
.B1(n_1269),
.B2(n_1265),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1262),
.B(n_1269),
.Y(n_1357)
);

OAI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1142),
.A2(n_1175),
.B1(n_1199),
.B2(n_1270),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1211),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1218),
.Y(n_1360)
);

OAI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1142),
.A2(n_1175),
.B1(n_1224),
.B2(n_1169),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1265),
.B(n_1188),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1158),
.Y(n_1363)
);

BUFx2_ASAP7_75t_SL g1364 ( 
.A(n_1148),
.Y(n_1364)
);

NAND2x1p5_ASAP7_75t_L g1365 ( 
.A(n_1226),
.B(n_1230),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1230),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1175),
.A2(n_1237),
.B1(n_1158),
.B2(n_1148),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1219),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_SL g1369 ( 
.A1(n_1181),
.A2(n_1251),
.B1(n_1268),
.B2(n_1225),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1268),
.B(n_1221),
.Y(n_1370)
);

BUFx2_ASAP7_75t_SL g1371 ( 
.A(n_1191),
.Y(n_1371)
);

INVx1_ASAP7_75t_SL g1372 ( 
.A(n_1198),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1237),
.A2(n_1148),
.B1(n_1201),
.B2(n_1225),
.Y(n_1373)
);

OA21x2_ASAP7_75t_L g1374 ( 
.A1(n_1240),
.A2(n_1238),
.B(n_1244),
.Y(n_1374)
);

AO21x1_ASAP7_75t_L g1375 ( 
.A1(n_1238),
.A2(n_1242),
.B(n_1201),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1241),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1202),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_SL g1378 ( 
.A1(n_1148),
.A2(n_1204),
.B1(n_1223),
.B2(n_1202),
.Y(n_1378)
);

OR2x6_ASAP7_75t_L g1379 ( 
.A(n_1233),
.B(n_1242),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1151),
.Y(n_1380)
);

NAND2x1p5_ASAP7_75t_L g1381 ( 
.A(n_1233),
.B(n_1213),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1151),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1249),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1213),
.A2(n_1223),
.B1(n_1249),
.B2(n_1177),
.Y(n_1384)
);

AOI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1234),
.A2(n_1206),
.B(n_1235),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1271),
.A2(n_1130),
.B1(n_957),
.B2(n_897),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1172),
.B(n_1180),
.Y(n_1387)
);

CKINVDCx20_ASAP7_75t_R g1388 ( 
.A(n_1209),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1145),
.B(n_1254),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1277),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1203),
.B(n_1165),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1161),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1258),
.A2(n_1138),
.B(n_957),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1140),
.Y(n_1394)
);

NOR2x1_ASAP7_75t_R g1395 ( 
.A(n_1317),
.B(n_1394),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1379),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1316),
.Y(n_1397)
);

OA21x2_ASAP7_75t_L g1398 ( 
.A1(n_1327),
.A2(n_1345),
.B(n_1336),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1393),
.A2(n_1304),
.B(n_1283),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1346),
.B(n_1347),
.Y(n_1400)
);

BUFx2_ASAP7_75t_L g1401 ( 
.A(n_1349),
.Y(n_1401)
);

OR2x6_ASAP7_75t_L g1402 ( 
.A(n_1318),
.B(n_1309),
.Y(n_1402)
);

NOR2x1_ASAP7_75t_R g1403 ( 
.A(n_1317),
.B(n_1394),
.Y(n_1403)
);

NOR2xp67_ASAP7_75t_R g1404 ( 
.A(n_1329),
.B(n_1328),
.Y(n_1404)
);

INVxp67_ASAP7_75t_L g1405 ( 
.A(n_1302),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1379),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1379),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1340),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1316),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1327),
.A2(n_1336),
.B(n_1344),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1312),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1342),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1329),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1302),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1379),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1288),
.B(n_1391),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1329),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1348),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1288),
.B(n_1391),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1374),
.Y(n_1420)
);

INVxp67_ASAP7_75t_SL g1421 ( 
.A(n_1289),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1366),
.Y(n_1422)
);

INVx4_ASAP7_75t_SL g1423 ( 
.A(n_1329),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1365),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1374),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1322),
.B(n_1323),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1374),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1392),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1322),
.B(n_1323),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1339),
.B(n_1335),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1285),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_SL g1432 ( 
.A1(n_1334),
.A2(n_1318),
.B(n_1306),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1350),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1375),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1381),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1375),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1338),
.B(n_1351),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1365),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1365),
.Y(n_1439)
);

INVxp67_ASAP7_75t_L g1440 ( 
.A(n_1314),
.Y(n_1440)
);

OR2x6_ASAP7_75t_L g1441 ( 
.A(n_1318),
.B(n_1309),
.Y(n_1441)
);

AOI21xp33_ASAP7_75t_L g1442 ( 
.A1(n_1386),
.A2(n_1324),
.B(n_1293),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1333),
.A2(n_1296),
.B1(n_1305),
.B2(n_1361),
.Y(n_1443)
);

AOI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1287),
.A2(n_1385),
.B(n_1309),
.Y(n_1444)
);

AOI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1309),
.A2(n_1318),
.B(n_1343),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1339),
.B(n_1351),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1377),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1325),
.B(n_1387),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1291),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1387),
.B(n_1286),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1360),
.Y(n_1451)
);

AO21x2_ASAP7_75t_L g1452 ( 
.A1(n_1376),
.A2(n_1300),
.B(n_1294),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1311),
.B(n_1320),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1353),
.B(n_1356),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1292),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1299),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1373),
.A2(n_1303),
.B(n_1367),
.Y(n_1457)
);

BUFx8_ASAP7_75t_SL g1458 ( 
.A(n_1312),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1331),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1368),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1310),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1359),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1354),
.B(n_1328),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1281),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1284),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1437),
.B(n_1301),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1399),
.A2(n_1358),
.B1(n_1389),
.B2(n_1321),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1398),
.B(n_1326),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1400),
.B(n_1354),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1421),
.B(n_1307),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1438),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1421),
.B(n_1369),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1398),
.B(n_1364),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1398),
.B(n_1364),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1408),
.B(n_1341),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1452),
.Y(n_1476)
);

AO21x2_ASAP7_75t_L g1477 ( 
.A1(n_1444),
.A2(n_1362),
.B(n_1357),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1408),
.B(n_1378),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1435),
.Y(n_1479)
);

BUFx4f_ASAP7_75t_L g1480 ( 
.A(n_1402),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1438),
.B(n_1352),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1398),
.B(n_1370),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1398),
.B(n_1370),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1452),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1412),
.B(n_1355),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1400),
.B(n_1370),
.Y(n_1486)
);

CKINVDCx8_ASAP7_75t_R g1487 ( 
.A(n_1423),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1412),
.B(n_1372),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1439),
.B(n_1424),
.Y(n_1489)
);

OAI322xp33_ASAP7_75t_L g1490 ( 
.A1(n_1443),
.A2(n_1453),
.A3(n_1448),
.B1(n_1432),
.B2(n_1454),
.C1(n_1437),
.C2(n_1440),
.Y(n_1490)
);

AOI221xp5_ASAP7_75t_L g1491 ( 
.A1(n_1399),
.A2(n_1295),
.B1(n_1315),
.B2(n_1297),
.C(n_1389),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1420),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1422),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1434),
.B(n_1295),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1442),
.A2(n_1443),
.B1(n_1454),
.B2(n_1448),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1416),
.B(n_1383),
.Y(n_1496)
);

AOI221xp5_ASAP7_75t_L g1497 ( 
.A1(n_1442),
.A2(n_1315),
.B1(n_1297),
.B2(n_1337),
.C(n_1313),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1424),
.B(n_1352),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1433),
.B(n_1434),
.Y(n_1499)
);

NOR2x1_ASAP7_75t_L g1500 ( 
.A(n_1432),
.B(n_1282),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1424),
.B(n_1363),
.Y(n_1501)
);

AO21x2_ASAP7_75t_L g1502 ( 
.A1(n_1444),
.A2(n_1384),
.B(n_1282),
.Y(n_1502)
);

OAI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1453),
.A2(n_1337),
.B1(n_1313),
.B2(n_1298),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1450),
.B(n_1319),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1396),
.B(n_1415),
.Y(n_1505)
);

OAI21xp33_ASAP7_75t_L g1506 ( 
.A1(n_1495),
.A2(n_1446),
.B(n_1436),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_SL g1507 ( 
.A1(n_1491),
.A2(n_1467),
.B(n_1497),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1467),
.A2(n_1441),
.B1(n_1402),
.B2(n_1405),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_SL g1509 ( 
.A1(n_1491),
.A2(n_1445),
.B(n_1446),
.Y(n_1509)
);

AND4x1_ASAP7_75t_L g1510 ( 
.A(n_1497),
.B(n_1395),
.C(n_1403),
.D(n_1458),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1482),
.B(n_1402),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1482),
.B(n_1402),
.Y(n_1512)
);

NAND3xp33_ASAP7_75t_L g1513 ( 
.A(n_1472),
.B(n_1461),
.C(n_1440),
.Y(n_1513)
);

OAI221xp5_ASAP7_75t_L g1514 ( 
.A1(n_1472),
.A2(n_1431),
.B1(n_1461),
.B2(n_1405),
.C(n_1414),
.Y(n_1514)
);

NAND3xp33_ASAP7_75t_L g1515 ( 
.A(n_1470),
.B(n_1457),
.C(n_1428),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1466),
.B(n_1431),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1469),
.B(n_1414),
.Y(n_1517)
);

OAI21xp33_ASAP7_75t_L g1518 ( 
.A1(n_1494),
.A2(n_1450),
.B(n_1419),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1469),
.B(n_1426),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1504),
.B(n_1426),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1504),
.B(n_1429),
.Y(n_1521)
);

OAI211xp5_ASAP7_75t_L g1522 ( 
.A1(n_1488),
.A2(n_1462),
.B(n_1451),
.C(n_1460),
.Y(n_1522)
);

NAND3xp33_ASAP7_75t_L g1523 ( 
.A(n_1470),
.B(n_1457),
.C(n_1447),
.Y(n_1523)
);

NAND2xp33_ASAP7_75t_SL g1524 ( 
.A(n_1478),
.B(n_1411),
.Y(n_1524)
);

OA21x2_ASAP7_75t_L g1525 ( 
.A1(n_1476),
.A2(n_1425),
.B(n_1427),
.Y(n_1525)
);

NAND4xp25_ASAP7_75t_L g1526 ( 
.A(n_1475),
.B(n_1401),
.C(n_1459),
.D(n_1449),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1482),
.B(n_1402),
.Y(n_1527)
);

OAI21xp5_ASAP7_75t_SL g1528 ( 
.A1(n_1500),
.A2(n_1445),
.B(n_1503),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1487),
.A2(n_1402),
.B1(n_1441),
.B2(n_1413),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1483),
.B(n_1441),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1483),
.B(n_1441),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1487),
.A2(n_1441),
.B1(n_1413),
.B2(n_1417),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1485),
.B(n_1429),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1500),
.B(n_1397),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1503),
.B(n_1397),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1471),
.B(n_1419),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1471),
.B(n_1425),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1466),
.B(n_1430),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1480),
.A2(n_1404),
.B(n_1410),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1505),
.B(n_1396),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1505),
.B(n_1427),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1505),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1488),
.B(n_1459),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1475),
.B(n_1401),
.Y(n_1544)
);

OAI211xp5_ASAP7_75t_L g1545 ( 
.A1(n_1478),
.A2(n_1449),
.B(n_1465),
.C(n_1464),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1487),
.A2(n_1413),
.B1(n_1417),
.B2(n_1337),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1480),
.A2(n_1463),
.B1(n_1498),
.B2(n_1501),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1480),
.A2(n_1417),
.B1(n_1337),
.B2(n_1313),
.Y(n_1548)
);

NAND3xp33_ASAP7_75t_L g1549 ( 
.A(n_1494),
.B(n_1457),
.C(n_1409),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1505),
.B(n_1418),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1480),
.A2(n_1463),
.B1(n_1406),
.B2(n_1407),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1496),
.B(n_1455),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1496),
.B(n_1455),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1486),
.B(n_1456),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1537),
.B(n_1468),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1544),
.B(n_1543),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1542),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1537),
.Y(n_1558)
);

INVxp67_ASAP7_75t_SL g1559 ( 
.A(n_1525),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1541),
.B(n_1473),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1536),
.B(n_1493),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1525),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1525),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1550),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1511),
.B(n_1473),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1550),
.Y(n_1566)
);

INVx4_ASAP7_75t_L g1567 ( 
.A(n_1540),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1511),
.B(n_1474),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1512),
.B(n_1474),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1536),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1542),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1552),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1512),
.B(n_1527),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1542),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1553),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1554),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1530),
.B(n_1474),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1530),
.B(n_1468),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1520),
.B(n_1493),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1533),
.B(n_1468),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1531),
.Y(n_1581)
);

INVx2_ASAP7_75t_SL g1582 ( 
.A(n_1540),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1521),
.B(n_1499),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_SL g1584 ( 
.A(n_1528),
.B(n_1490),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1531),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1517),
.B(n_1492),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1549),
.B(n_1492),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1538),
.Y(n_1588)
);

NOR2xp67_ASAP7_75t_L g1589 ( 
.A(n_1523),
.B(n_1484),
.Y(n_1589)
);

OR2x6_ASAP7_75t_L g1590 ( 
.A(n_1539),
.B(n_1489),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1540),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1519),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1545),
.Y(n_1593)
);

INVxp67_ASAP7_75t_SL g1594 ( 
.A(n_1515),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1562),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1562),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1563),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1563),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1587),
.B(n_1526),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1594),
.B(n_1516),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1557),
.Y(n_1601)
);

INVxp33_ASAP7_75t_L g1602 ( 
.A(n_1584),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1557),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1594),
.B(n_1518),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1587),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1558),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1558),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1593),
.B(n_1522),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1566),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1591),
.B(n_1547),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1566),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1590),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1555),
.B(n_1513),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1566),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1559),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1593),
.B(n_1588),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1588),
.B(n_1484),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1567),
.B(n_1534),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1591),
.B(n_1567),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1591),
.B(n_1529),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1559),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1564),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1567),
.B(n_1479),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1567),
.B(n_1479),
.Y(n_1624)
);

NAND3xp33_ASAP7_75t_L g1625 ( 
.A(n_1584),
.B(n_1507),
.C(n_1510),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1555),
.B(n_1477),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1560),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1564),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1586),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1580),
.B(n_1477),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1565),
.B(n_1479),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1586),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1565),
.B(n_1489),
.Y(n_1633)
);

INVxp67_ASAP7_75t_SL g1634 ( 
.A(n_1589),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1604),
.B(n_1580),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1608),
.B(n_1592),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1604),
.B(n_1556),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1595),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1627),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1595),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1620),
.B(n_1582),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1620),
.B(n_1582),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1596),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1629),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1608),
.B(n_1616),
.Y(n_1645)
);

AO22x1_ASAP7_75t_L g1646 ( 
.A1(n_1602),
.A2(n_1582),
.B1(n_1524),
.B2(n_1532),
.Y(n_1646)
);

AOI32xp33_ASAP7_75t_L g1647 ( 
.A1(n_1634),
.A2(n_1524),
.A3(n_1506),
.B1(n_1514),
.B2(n_1577),
.Y(n_1647)
);

AND2x2_ASAP7_75t_SL g1648 ( 
.A(n_1600),
.B(n_1498),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1612),
.B(n_1573),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1601),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1596),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1625),
.B(n_1556),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1616),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1612),
.B(n_1573),
.Y(n_1654)
);

INVx1_ASAP7_75t_SL g1655 ( 
.A(n_1600),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1599),
.B(n_1592),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1597),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1605),
.B(n_1583),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1597),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1599),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1598),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1625),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1598),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1622),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1622),
.Y(n_1665)
);

NOR2x1p5_ASAP7_75t_L g1666 ( 
.A(n_1613),
.B(n_1332),
.Y(n_1666)
);

NAND3xp33_ASAP7_75t_L g1667 ( 
.A(n_1605),
.B(n_1589),
.C(n_1509),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1628),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1613),
.A2(n_1508),
.B1(n_1590),
.B2(n_1535),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1628),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1605),
.B(n_1629),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1619),
.B(n_1565),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1632),
.B(n_1583),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1632),
.B(n_1576),
.Y(n_1674)
);

O2A1O1Ixp5_ASAP7_75t_L g1675 ( 
.A1(n_1618),
.A2(n_1534),
.B(n_1535),
.C(n_1490),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1610),
.B(n_1576),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1610),
.B(n_1572),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1638),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1650),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1652),
.B(n_1633),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1648),
.B(n_1618),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1662),
.A2(n_1590),
.B1(n_1618),
.B2(n_1619),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1648),
.B(n_1618),
.Y(n_1683)
);

NAND2x1p5_ASAP7_75t_L g1684 ( 
.A(n_1666),
.B(n_1601),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1641),
.B(n_1623),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1655),
.B(n_1630),
.Y(n_1686)
);

INVxp67_ASAP7_75t_L g1687 ( 
.A(n_1652),
.Y(n_1687)
);

OAI221xp5_ASAP7_75t_L g1688 ( 
.A1(n_1662),
.A2(n_1647),
.B1(n_1667),
.B2(n_1660),
.C(n_1669),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1640),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1641),
.B(n_1623),
.Y(n_1690)
);

INVx1_ASAP7_75t_SL g1691 ( 
.A(n_1650),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1642),
.B(n_1624),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1644),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1643),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1653),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1645),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1636),
.B(n_1332),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1651),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1656),
.B(n_1633),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1642),
.B(n_1649),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1649),
.B(n_1624),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1646),
.A2(n_1590),
.B(n_1617),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1637),
.B(n_1630),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1654),
.A2(n_1502),
.B1(n_1546),
.B2(n_1590),
.Y(n_1704)
);

CKINVDCx16_ASAP7_75t_R g1705 ( 
.A(n_1654),
.Y(n_1705)
);

OR2x6_ASAP7_75t_L g1706 ( 
.A(n_1671),
.B(n_1590),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1672),
.B(n_1627),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_SL g1708 ( 
.A1(n_1672),
.A2(n_1603),
.B1(n_1601),
.B2(n_1627),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1657),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1639),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1639),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1671),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1676),
.B(n_1631),
.Y(n_1713)
);

XOR2x2_ASAP7_75t_L g1714 ( 
.A(n_1688),
.B(n_1330),
.Y(n_1714)
);

OAI21xp33_ASAP7_75t_L g1715 ( 
.A1(n_1687),
.A2(n_1635),
.B(n_1677),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1693),
.Y(n_1716)
);

A2O1A1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1702),
.A2(n_1675),
.B(n_1635),
.C(n_1621),
.Y(n_1717)
);

OAI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1684),
.A2(n_1658),
.B1(n_1674),
.B2(n_1673),
.C(n_1663),
.Y(n_1718)
);

OAI322xp33_ASAP7_75t_L g1719 ( 
.A1(n_1696),
.A2(n_1615),
.A3(n_1621),
.B1(n_1658),
.B2(n_1673),
.C1(n_1661),
.C2(n_1659),
.Y(n_1719)
);

OAI22xp33_ASAP7_75t_SL g1720 ( 
.A1(n_1705),
.A2(n_1603),
.B1(n_1615),
.B2(n_1668),
.Y(n_1720)
);

NAND4xp25_ASAP7_75t_L g1721 ( 
.A(n_1695),
.B(n_1670),
.C(n_1665),
.D(n_1664),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1705),
.B(n_1631),
.Y(n_1722)
);

CKINVDCx20_ASAP7_75t_R g1723 ( 
.A(n_1697),
.Y(n_1723)
);

A2O1A1Ixp33_ASAP7_75t_L g1724 ( 
.A1(n_1704),
.A2(n_1626),
.B(n_1603),
.C(n_1617),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1712),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1712),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1712),
.Y(n_1727)
);

INVx1_ASAP7_75t_SL g1728 ( 
.A(n_1695),
.Y(n_1728)
);

OAI21xp33_ASAP7_75t_L g1729 ( 
.A1(n_1680),
.A2(n_1626),
.B(n_1611),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1679),
.B(n_1609),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1700),
.B(n_1578),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1712),
.Y(n_1732)
);

OAI21xp33_ASAP7_75t_L g1733 ( 
.A1(n_1704),
.A2(n_1611),
.B(n_1609),
.Y(n_1733)
);

OAI322xp33_ASAP7_75t_L g1734 ( 
.A1(n_1691),
.A2(n_1607),
.A3(n_1606),
.B1(n_1609),
.B2(n_1614),
.C1(n_1611),
.C2(n_1561),
.Y(n_1734)
);

OAI21xp5_ASAP7_75t_SL g1735 ( 
.A1(n_1684),
.A2(n_1548),
.B(n_1551),
.Y(n_1735)
);

NAND3xp33_ASAP7_75t_SL g1736 ( 
.A(n_1684),
.B(n_1708),
.C(n_1691),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_SL g1737 ( 
.A(n_1681),
.B(n_1579),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1681),
.A2(n_1498),
.B1(n_1501),
.B2(n_1481),
.Y(n_1738)
);

NAND3xp33_ASAP7_75t_L g1739 ( 
.A(n_1679),
.B(n_1614),
.C(n_1607),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1728),
.B(n_1700),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1725),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1722),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1723),
.B(n_1699),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1716),
.B(n_1713),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1726),
.Y(n_1745)
);

NAND3xp33_ASAP7_75t_L g1746 ( 
.A(n_1717),
.B(n_1682),
.C(n_1678),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1727),
.Y(n_1747)
);

OAI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1735),
.A2(n_1683),
.B1(n_1701),
.B2(n_1685),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1732),
.Y(n_1749)
);

INVx2_ASAP7_75t_SL g1750 ( 
.A(n_1730),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1721),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1737),
.B(n_1685),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1730),
.B(n_1690),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1715),
.B(n_1713),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1736),
.A2(n_1683),
.B1(n_1690),
.B2(n_1692),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1721),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1738),
.B(n_1692),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1739),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1720),
.Y(n_1759)
);

NAND3xp33_ASAP7_75t_SL g1760 ( 
.A(n_1755),
.B(n_1718),
.C(n_1724),
.Y(n_1760)
);

AOI21xp33_ASAP7_75t_SL g1761 ( 
.A1(n_1759),
.A2(n_1733),
.B(n_1714),
.Y(n_1761)
);

AOI221xp5_ASAP7_75t_L g1762 ( 
.A1(n_1756),
.A2(n_1719),
.B1(n_1734),
.B2(n_1729),
.C(n_1698),
.Y(n_1762)
);

AO22x2_ASAP7_75t_L g1763 ( 
.A1(n_1756),
.A2(n_1698),
.B1(n_1689),
.B2(n_1694),
.Y(n_1763)
);

OAI221xp5_ASAP7_75t_L g1764 ( 
.A1(n_1746),
.A2(n_1706),
.B1(n_1686),
.B2(n_1731),
.C(n_1709),
.Y(n_1764)
);

NAND4xp75_ASAP7_75t_L g1765 ( 
.A(n_1751),
.B(n_1678),
.C(n_1709),
.D(n_1689),
.Y(n_1765)
);

AOI211xp5_ASAP7_75t_SL g1766 ( 
.A1(n_1758),
.A2(n_1686),
.B(n_1694),
.C(n_1703),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1741),
.Y(n_1767)
);

NOR3xp33_ASAP7_75t_L g1768 ( 
.A(n_1743),
.B(n_1403),
.C(n_1395),
.Y(n_1768)
);

NOR3xp33_ASAP7_75t_L g1769 ( 
.A(n_1740),
.B(n_1711),
.C(n_1710),
.Y(n_1769)
);

AOI211xp5_ASAP7_75t_SL g1770 ( 
.A1(n_1748),
.A2(n_1703),
.B(n_1701),
.C(n_1710),
.Y(n_1770)
);

O2A1O1Ixp33_ASAP7_75t_L g1771 ( 
.A1(n_1754),
.A2(n_1706),
.B(n_1710),
.C(n_1711),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1763),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1766),
.B(n_1742),
.Y(n_1773)
);

NOR2x1_ASAP7_75t_L g1774 ( 
.A(n_1765),
.B(n_1741),
.Y(n_1774)
);

AOI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1761),
.A2(n_1742),
.B1(n_1744),
.B2(n_1747),
.C(n_1749),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1764),
.B(n_1752),
.Y(n_1776)
);

AOI211xp5_ASAP7_75t_L g1777 ( 
.A1(n_1760),
.A2(n_1752),
.B(n_1750),
.C(n_1745),
.Y(n_1777)
);

AO22x2_ASAP7_75t_L g1778 ( 
.A1(n_1767),
.A2(n_1745),
.B1(n_1750),
.B2(n_1763),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1770),
.B(n_1753),
.Y(n_1779)
);

INVx2_ASAP7_75t_SL g1780 ( 
.A(n_1768),
.Y(n_1780)
);

NAND3xp33_ASAP7_75t_SL g1781 ( 
.A(n_1762),
.B(n_1753),
.C(n_1757),
.Y(n_1781)
);

NAND4xp25_ASAP7_75t_L g1782 ( 
.A(n_1771),
.B(n_1757),
.C(n_1711),
.D(n_1707),
.Y(n_1782)
);

AOI211x1_ASAP7_75t_L g1783 ( 
.A1(n_1781),
.A2(n_1707),
.B(n_1769),
.C(n_1606),
.Y(n_1783)
);

NOR4xp25_ASAP7_75t_L g1784 ( 
.A(n_1772),
.B(n_1614),
.C(n_1706),
.D(n_1571),
.Y(n_1784)
);

NAND3x1_ASAP7_75t_L g1785 ( 
.A(n_1774),
.B(n_1388),
.C(n_1290),
.Y(n_1785)
);

AOI221xp5_ASAP7_75t_L g1786 ( 
.A1(n_1778),
.A2(n_1572),
.B1(n_1575),
.B2(n_1290),
.C(n_1388),
.Y(n_1786)
);

NAND3xp33_ASAP7_75t_L g1787 ( 
.A(n_1777),
.B(n_1706),
.C(n_1380),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1776),
.B(n_1706),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1773),
.B(n_1280),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1785),
.A2(n_1779),
.B1(n_1778),
.B2(n_1780),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1783),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1789),
.A2(n_1775),
.B1(n_1782),
.B2(n_1571),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1788),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1787),
.Y(n_1794)
);

AOI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1786),
.A2(n_1574),
.B1(n_1571),
.B2(n_1569),
.Y(n_1795)
);

AOI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1784),
.A2(n_1574),
.B1(n_1568),
.B2(n_1569),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1791),
.Y(n_1797)
);

BUFx12f_ASAP7_75t_L g1798 ( 
.A(n_1793),
.Y(n_1798)
);

AND2x4_ASAP7_75t_L g1799 ( 
.A(n_1794),
.B(n_1574),
.Y(n_1799)
);

NAND2x1p5_ASAP7_75t_L g1800 ( 
.A(n_1792),
.B(n_1280),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1790),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1800),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1798),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1801),
.B(n_1795),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1803),
.Y(n_1805)
);

OAI321xp33_ASAP7_75t_L g1806 ( 
.A1(n_1805),
.A2(n_1797),
.A3(n_1802),
.B1(n_1804),
.B2(n_1796),
.C(n_1799),
.Y(n_1806)
);

OAI21x1_ASAP7_75t_L g1807 ( 
.A1(n_1806),
.A2(n_1797),
.B(n_1579),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1806),
.Y(n_1808)
);

NAND3xp33_ASAP7_75t_SL g1809 ( 
.A(n_1808),
.B(n_1561),
.C(n_1371),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1807),
.Y(n_1810)
);

OAI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1810),
.A2(n_1808),
.B1(n_1575),
.B2(n_1570),
.Y(n_1811)
);

OAI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1809),
.A2(n_1581),
.B1(n_1585),
.B2(n_1382),
.Y(n_1812)
);

XNOR2x1_ASAP7_75t_L g1813 ( 
.A(n_1811),
.B(n_1382),
.Y(n_1813)
);

AOI322xp5_ASAP7_75t_L g1814 ( 
.A1(n_1813),
.A2(n_1812),
.A3(n_1568),
.B1(n_1569),
.B2(n_1577),
.C1(n_1581),
.C2(n_1585),
.Y(n_1814)
);

OAI221xp5_ASAP7_75t_R g1815 ( 
.A1(n_1814),
.A2(n_1404),
.B1(n_1502),
.B2(n_1568),
.C(n_1577),
.Y(n_1815)
);

AOI211xp5_ASAP7_75t_L g1816 ( 
.A1(n_1815),
.A2(n_1382),
.B(n_1390),
.C(n_1308),
.Y(n_1816)
);


endmodule