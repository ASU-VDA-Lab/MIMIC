module fake_jpeg_31573_n_136 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_136);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_26),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_25),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_2),
.B(n_5),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx11_ASAP7_75t_SL g56 ( 
.A(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_6),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_0),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_56),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_1),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_18),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_49),
.Y(n_81)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_74),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_44),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_70),
.A2(n_73),
.B1(n_60),
.B2(n_59),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_86),
.B1(n_3),
.B2(n_4),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_59),
.B1(n_60),
.B2(n_44),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_80),
.B1(n_48),
.B2(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_64),
.B1(n_56),
.B2(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_84),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_63),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_65),
.B1(n_64),
.B2(n_45),
.Y(n_86)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_98),
.B(n_16),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_86),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_99),
.Y(n_105)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_77),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_100),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_57),
.B1(n_47),
.B2(n_51),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_101)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_97),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_21),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_1),
.B(n_3),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_81),
.B(n_4),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_101),
.A2(n_105),
.B1(n_109),
.B2(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_27),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_28),
.B(n_12),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_107),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_89),
.C(n_22),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_14),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_35),
.B1(n_36),
.B2(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_40),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_15),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_112),
.C(n_29),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_114),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_118),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_34),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_121),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_104),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_115),
.B1(n_121),
.B2(n_120),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_129),
.B(n_124),
.C(n_112),
.Y(n_130)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_128),
.B(n_125),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_131),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_127),
.C(n_126),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_133),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_118),
.Y(n_135)
);

BUFx24_ASAP7_75t_SL g136 ( 
.A(n_135),
.Y(n_136)
);


endmodule