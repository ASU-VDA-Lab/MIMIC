module fake_jpeg_8123_n_313 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx2_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_7),
.B(n_1),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_7),
.Y(n_55)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_39),
.Y(n_53)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_30),
.B1(n_35),
.B2(n_33),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_59),
.B1(n_67),
.B2(n_20),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_30),
.B1(n_22),
.B2(n_33),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_62),
.B1(n_20),
.B2(n_34),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_53),
.Y(n_91)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_52),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

NOR3xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_18),
.C(n_23),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_26),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_23),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_60),
.B(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_37),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_22),
.B1(n_33),
.B2(n_27),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_27),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_34),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_33),
.B1(n_22),
.B2(n_32),
.Y(n_62)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_66),
.Y(n_73)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_22),
.B1(n_31),
.B2(n_25),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_82),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_55),
.B(n_52),
.C(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_71),
.B(n_80),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_72),
.A2(n_90),
.B1(n_103),
.B2(n_66),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_37),
.B1(n_43),
.B2(n_40),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_74),
.A2(n_85),
.B1(n_101),
.B2(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_75),
.B(n_76),
.Y(n_124)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_20),
.B1(n_34),
.B2(n_17),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_77),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

CKINVDCx10_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_95),
.B1(n_92),
.B2(n_76),
.Y(n_106)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_86),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_25),
.B1(n_17),
.B2(n_31),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_88),
.Y(n_123)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_89),
.B(n_96),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_46),
.A2(n_31),
.B1(n_25),
.B2(n_17),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_92),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_18),
.Y(n_93)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_18),
.Y(n_94)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_42),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_26),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_99),
.B(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_42),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_24),
.C(n_63),
.Y(n_114)
);

AO22x2_ASAP7_75t_SL g101 ( 
.A1(n_64),
.A2(n_38),
.B1(n_43),
.B2(n_40),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_64),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_63),
.A2(n_43),
.B1(n_21),
.B2(n_32),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_105),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_106),
.A2(n_100),
.B1(n_74),
.B2(n_85),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_109),
.B(n_114),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_97),
.A2(n_24),
.B1(n_63),
.B2(n_43),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_79),
.B(n_73),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_99),
.B1(n_96),
.B2(n_88),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_75),
.A2(n_48),
.B1(n_1),
.B2(n_2),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_14),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_119),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_101),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_104),
.Y(n_133)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_127),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_71),
.A2(n_48),
.B1(n_32),
.B2(n_28),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_82),
.B1(n_89),
.B2(n_81),
.Y(n_158)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_83),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_133),
.A2(n_144),
.B(n_162),
.Y(n_170)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_137),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_70),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_140),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_139),
.A2(n_149),
.B1(n_110),
.B2(n_128),
.Y(n_175)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_70),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_141),
.B(n_143),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_158),
.B1(n_160),
.B2(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_150),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_102),
.Y(n_148)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_80),
.Y(n_151)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_91),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_153),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_91),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_95),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_154),
.A2(n_131),
.B(n_111),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_118),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_119),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_127),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_156),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_115),
.Y(n_157)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_91),
.C(n_38),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_114),
.C(n_128),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_106),
.A2(n_38),
.B1(n_32),
.B2(n_28),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_38),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_132),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_171),
.B(n_172),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_144),
.A2(n_131),
.B(n_108),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_182),
.C(n_184),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_175),
.A2(n_186),
.B(n_188),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_162),
.A2(n_125),
.B1(n_120),
.B2(n_105),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_176),
.A2(n_177),
.B1(n_180),
.B2(n_191),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_151),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_145),
.A2(n_105),
.B1(n_112),
.B2(n_111),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_152),
.C(n_153),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_112),
.C(n_109),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_137),
.B(n_129),
.C(n_19),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_192),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_19),
.B(n_28),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_0),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_135),
.A2(n_28),
.B1(n_21),
.B2(n_19),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_21),
.C(n_0),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_145),
.A2(n_21),
.B1(n_0),
.B2(n_3),
.Y(n_193)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_142),
.B(n_2),
.C(n_3),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_195),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_3),
.C(n_4),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_136),
.A2(n_4),
.B1(n_5),
.B2(n_10),
.Y(n_196)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_197),
.Y(n_238)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_169),
.Y(n_200)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_161),
.Y(n_202)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_167),
.Y(n_204)
);

INVxp67_ASAP7_75t_SL g237 ( 
.A(n_204),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_182),
.B(n_164),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_205),
.B(n_191),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_154),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_208),
.Y(n_227)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_180),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_220),
.B1(n_221),
.B2(n_134),
.Y(n_228)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_213),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_170),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_218),
.Y(n_239)
);

BUFx12_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_188),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_188),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_222),
.A2(n_170),
.B(n_186),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_205),
.C(n_174),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_225),
.C(n_231),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_135),
.B1(n_160),
.B2(n_177),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_224),
.A2(n_218),
.B1(n_201),
.B2(n_206),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_172),
.C(n_184),
.Y(n_225)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_214),
.A2(n_147),
.B1(n_143),
.B2(n_187),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_229),
.A2(n_243),
.B1(n_199),
.B2(n_222),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_150),
.B(n_181),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_230),
.A2(n_201),
.B(n_212),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_185),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_192),
.C(n_164),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_241),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_203),
.A2(n_194),
.B1(n_155),
.B2(n_195),
.Y(n_236)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_163),
.C(n_166),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_203),
.A2(n_133),
.B1(n_178),
.B2(n_196),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_226),
.Y(n_249)
);

NOR2x1_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_207),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_245),
.A2(n_252),
.B1(n_258),
.B2(n_259),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_249),
.B(n_244),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_251),
.A2(n_229),
.B1(n_243),
.B2(n_242),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_232),
.B(n_215),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_254),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_239),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_240),
.B(n_215),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_256),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_235),
.B(n_210),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_257),
.A2(n_261),
.B(n_262),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_239),
.A2(n_206),
.B1(n_208),
.B2(n_221),
.Y(n_258)
);

OA22x2_ASAP7_75t_L g259 ( 
.A1(n_224),
.A2(n_212),
.B1(n_191),
.B2(n_197),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_233),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_270),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_223),
.C(n_225),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_268),
.C(n_276),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_231),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_271),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_241),
.C(n_234),
.Y(n_268)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_227),
.Y(n_270)
);

BUFx24_ASAP7_75t_SL g271 ( 
.A(n_260),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_237),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_274),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_238),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_219),
.C(n_235),
.Y(n_276)
);

NOR2x1_ASAP7_75t_SL g277 ( 
.A(n_263),
.B(n_245),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_5),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_254),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_13),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_247),
.B(n_254),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_283),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_261),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_282),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_275),
.A2(n_257),
.B(n_259),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_287),
.C(n_288),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_264),
.A2(n_259),
.B(n_219),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_259),
.C(n_191),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_279),
.A2(n_268),
.B1(n_10),
.B2(n_12),
.Y(n_290)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

OAI21x1_ASAP7_75t_L g293 ( 
.A1(n_277),
.A2(n_5),
.B(n_12),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_294),
.B(n_286),
.Y(n_301)
);

NOR2xp67_ASAP7_75t_SL g294 ( 
.A(n_288),
.B(n_12),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_296),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_13),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_14),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_301),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_283),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_302),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_305),
.Y(n_310)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_304),
.A2(n_291),
.A3(n_296),
.B1(n_287),
.B2(n_281),
.C1(n_285),
.C2(n_15),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_307),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_281),
.B(n_285),
.Y(n_307)
);

NOR2xp67_ASAP7_75t_SL g311 ( 
.A(n_309),
.B(n_308),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_310),
.C(n_299),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_298),
.C(n_16),
.Y(n_313)
);


endmodule