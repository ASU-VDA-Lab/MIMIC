module fake_aes_7284_n_35 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_7), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_3), .Y(n_12) );
AOI22xp5_ASAP7_75t_SL g13 ( .A1(n_9), .A2(n_6), .B1(n_10), .B2(n_8), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_0), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_4), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_6), .Y(n_17) );
AOI21xp5_ASAP7_75t_L g18 ( .A1(n_14), .A2(n_0), .B(n_1), .Y(n_18) );
A2O1A1Ixp33_ASAP7_75t_L g19 ( .A1(n_13), .A2(n_1), .B(n_2), .C(n_3), .Y(n_19) );
O2A1O1Ixp33_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_2), .B(n_4), .C(n_5), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_17), .B(n_5), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_11), .B(n_7), .Y(n_22) );
AND2x4_ASAP7_75t_L g23 ( .A(n_21), .B(n_14), .Y(n_23) );
BUFx2_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
CKINVDCx5p33_ASAP7_75t_R g25 ( .A(n_22), .Y(n_25) );
OR2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_19), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
NAND2x1p5_ASAP7_75t_L g28 ( .A(n_24), .B(n_13), .Y(n_28) );
INVx1_ASAP7_75t_SL g29 ( .A(n_27), .Y(n_29) );
OAI221xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_28), .B1(n_26), .B2(n_24), .C(n_20), .Y(n_30) );
OAI221xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_24), .B1(n_12), .B2(n_18), .C(n_16), .Y(n_31) );
BUFx2_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
CKINVDCx20_ASAP7_75t_R g33 ( .A(n_30), .Y(n_33) );
AOI31xp33_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_15), .A3(n_16), .B(n_23), .Y(n_34) );
AOI22xp33_ASAP7_75t_SL g35 ( .A1(n_34), .A2(n_33), .B1(n_32), .B2(n_23), .Y(n_35) );
endmodule