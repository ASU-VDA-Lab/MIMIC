module fake_jpeg_8418_n_119 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_119);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_31),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

BUFx2_ASAP7_75t_SL g87 ( 
.A(n_59),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_54),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_63),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_66),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_58),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_1),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_66),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_71),
.Y(n_89)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_68),
.A2(n_49),
.B1(n_55),
.B2(n_41),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_72),
.A2(n_76),
.B1(n_80),
.B2(n_88),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_51),
.B1(n_39),
.B2(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

OR2x2_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_62),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_85),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_46),
.B1(n_51),
.B2(n_53),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_61),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_86),
.B(n_84),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_56),
.B1(n_44),
.B2(n_3),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_40),
.Y(n_91)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_1),
.C(n_2),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_10),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_16),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_97),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_102),
.B1(n_89),
.B2(n_101),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_89),
.B1(n_95),
.B2(n_103),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_99),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_92),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_103),
.B1(n_83),
.B2(n_97),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_93),
.B(n_100),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_98),
.C(n_96),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_111),
.B(n_94),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_94),
.B(n_73),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_87),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_114),
.A2(n_17),
.B(n_18),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

AOI21x1_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_24),
.B(n_26),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_29),
.B(n_30),
.Y(n_119)
);


endmodule