module fake_netlist_5_1596_n_2028 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_2028);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2028;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_877;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_314;
wire n_604;
wire n_368;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1982;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1184;
wire n_1011;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_102),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_165),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_112),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_162),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_28),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_153),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_22),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_130),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_51),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_129),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_54),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_54),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_49),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_134),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_187),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_176),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_157),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_126),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_55),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_128),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_160),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_85),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_191),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_69),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_38),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_189),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_119),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_56),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_193),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_169),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_95),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_184),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_11),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_136),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_166),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_16),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_71),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_51),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_168),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_145),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_199),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_3),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_137),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_196),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_99),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_197),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_143),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_52),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_82),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_200),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_120),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_111),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_18),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_35),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_60),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_110),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_79),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_32),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_97),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_92),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_201),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_3),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_52),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_149),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_74),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_116),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_73),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_155),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_198),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_32),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_138),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_180),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_174),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_58),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_27),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_29),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_170),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_75),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_103),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_118),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_106),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_158),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_182),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_55),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_28),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_105),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_87),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_94),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_68),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_81),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_186),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_139),
.Y(n_299)
);

INVxp33_ASAP7_75t_R g300 ( 
.A(n_17),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_150),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_8),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_195),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_70),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_190),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_19),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_183),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_83),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_60),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_175),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_62),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_91),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_13),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_21),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_115),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_72),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_45),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_8),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_31),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_47),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_36),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_4),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_67),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_43),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_133),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_4),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_161),
.Y(n_327)
);

BUFx10_ASAP7_75t_L g328 ( 
.A(n_1),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_148),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_19),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_142),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_84),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_36),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_188),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_47),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_80),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_104),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_56),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_57),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_11),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_163),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_123),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_147),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_88),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_96),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_15),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_37),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_63),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_66),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_23),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_49),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_203),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_44),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_9),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_141),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_38),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_41),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_40),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_204),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_100),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_46),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_194),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_113),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_131),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_192),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_90),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_127),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_1),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_93),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_0),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_181),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_2),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_53),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_65),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_14),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_6),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_151),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_57),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_154),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_14),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_25),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_20),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_21),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_44),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_24),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_22),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_5),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_101),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_6),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_135),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_125),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_202),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_40),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_61),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_12),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_114),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_144),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_107),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_98),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_179),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_27),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_53),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_108),
.Y(n_403)
);

BUFx10_ASAP7_75t_L g404 ( 
.A(n_146),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_167),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_13),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_33),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_42),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_50),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_86),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_34),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_121),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_359),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_226),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_282),
.Y(n_415)
);

BUFx2_ASAP7_75t_SL g416 ( 
.A(n_359),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_376),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_380),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_218),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_239),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_226),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_226),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_282),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_211),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_213),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_208),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_226),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_302),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_257),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_296),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_226),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_304),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_277),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_243),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_277),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_208),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_277),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_302),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_277),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_236),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_247),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_249),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_273),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_277),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_317),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_275),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_317),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_288),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_209),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_317),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_339),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_317),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_260),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_339),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_317),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_402),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_212),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_402),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_402),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_402),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_402),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_408),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_218),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_261),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_408),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_408),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_408),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_408),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_215),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_217),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_232),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_235),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_245),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_326),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_326),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_302),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_216),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_255),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_248),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_262),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_292),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_306),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_313),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_319),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_250),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_354),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_253),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_340),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_254),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_265),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_340),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_361),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_328),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_361),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_370),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_375),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_269),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_311),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_291),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_385),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_394),
.Y(n_501)
);

INVxp33_ASAP7_75t_SL g502 ( 
.A(n_311),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_401),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_409),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_411),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_205),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_206),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_208),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_328),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_256),
.Y(n_510)
);

INVxp33_ASAP7_75t_L g511 ( 
.A(n_300),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_258),
.Y(n_512)
);

BUFx2_ASAP7_75t_SL g513 ( 
.A(n_266),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_240),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_214),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_240),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_309),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_393),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_246),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_448),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_421),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_413),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_421),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_414),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_427),
.Y(n_525)
);

INVx5_ASAP7_75t_L g526 ( 
.A(n_448),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_509),
.B(n_283),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_414),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_513),
.B(n_266),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_448),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_415),
.B(n_214),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_427),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_422),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_431),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_422),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_431),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_465),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_465),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_448),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_423),
.B(n_214),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_433),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_448),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_451),
.B(n_346),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_433),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_435),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_435),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_437),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_440),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_437),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_430),
.A2(n_283),
.B1(n_383),
.B2(n_351),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_439),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_439),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_444),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_444),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_445),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_445),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_443),
.B(n_316),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_447),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_447),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_450),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_506),
.B(n_273),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_450),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_502),
.A2(n_383),
.B1(n_407),
.B2(n_351),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_513),
.B(n_441),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_507),
.B(n_316),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_452),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_452),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_466),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_466),
.B(n_273),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_455),
.B(n_220),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_456),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_458),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_419),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_449),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_459),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_460),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_461),
.B(n_220),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_462),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_418),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_467),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_451),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_468),
.B(n_221),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_519),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_519),
.B(n_221),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_454),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_474),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_418),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_474),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_492),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_492),
.B(n_246),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_475),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_495),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_475),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_457),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_477),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_488),
.B(n_303),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_416),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_488),
.B(n_303),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_479),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_491),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_491),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_495),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_514),
.B(n_259),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_496),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_530),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_521),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_L g607 ( 
.A(n_557),
.B(n_288),
.Y(n_607)
);

OAI22xp33_ASAP7_75t_L g608 ( 
.A1(n_527),
.A2(n_381),
.B1(n_358),
.B2(n_318),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_557),
.A2(n_502),
.B1(n_348),
.B2(n_498),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_574),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_581),
.B(n_494),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_524),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_521),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_529),
.B(n_446),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_564),
.B(n_417),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_570),
.B(n_417),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_530),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_543),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_561),
.B(n_469),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_561),
.A2(n_348),
.B1(n_518),
.B2(n_463),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_527),
.Y(n_621)
);

NAND2x1p5_ASAP7_75t_L g622 ( 
.A(n_590),
.B(n_207),
.Y(n_622)
);

BUFx6f_ASAP7_75t_SL g623 ( 
.A(n_581),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_524),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_523),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_581),
.B(n_485),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_524),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_528),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_597),
.B(n_476),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_528),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_547),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_528),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_597),
.B(n_424),
.Y(n_633)
);

AOI21x1_ASAP7_75t_L g634 ( 
.A1(n_569),
.A2(n_238),
.B(n_225),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_533),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_543),
.B(n_424),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_533),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_533),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_535),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_523),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_573),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_525),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_530),
.Y(n_643)
);

OR2x6_ASAP7_75t_L g644 ( 
.A(n_603),
.B(n_416),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_535),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_L g646 ( 
.A(n_570),
.B(n_288),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_603),
.B(n_270),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_561),
.B(n_585),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_530),
.Y(n_649)
);

NAND2xp33_ASAP7_75t_L g650 ( 
.A(n_577),
.B(n_288),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_573),
.B(n_487),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_561),
.B(n_470),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_535),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_537),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_525),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_537),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_537),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_531),
.B(n_425),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_532),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_590),
.A2(n_472),
.B1(n_473),
.B2(n_471),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_531),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_577),
.B(n_425),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_532),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_582),
.B(n_428),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_538),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_534),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_L g667 ( 
.A1(n_550),
.A2(n_314),
.B1(n_321),
.B2(n_320),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_534),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_540),
.Y(n_669)
);

AND3x2_ASAP7_75t_L g670 ( 
.A(n_579),
.B(n_281),
.C(n_219),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_538),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_582),
.B(n_438),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_536),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_536),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_579),
.Y(n_675)
);

OR2x6_ASAP7_75t_L g676 ( 
.A(n_540),
.B(n_514),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_584),
.B(n_489),
.Y(n_677)
);

BUFx10_ASAP7_75t_L g678 ( 
.A(n_587),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_520),
.B(n_434),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_520),
.B(n_434),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_538),
.Y(n_681)
);

OAI22xp33_ASAP7_75t_L g682 ( 
.A1(n_550),
.A2(n_324),
.B1(n_330),
.B2(n_322),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_544),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_541),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_544),
.Y(n_685)
);

AND2x6_ASAP7_75t_L g686 ( 
.A(n_569),
.B(n_288),
.Y(n_686)
);

AND2x6_ASAP7_75t_L g687 ( 
.A(n_569),
.B(n_293),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_584),
.B(n_442),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_544),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_585),
.B(n_442),
.Y(n_690)
);

AND3x1_ASAP7_75t_L g691 ( 
.A(n_565),
.B(n_516),
.C(n_480),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_541),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_585),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_565),
.B(n_493),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_563),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_592),
.B(n_494),
.Y(n_696)
);

INVxp67_ASAP7_75t_R g697 ( 
.A(n_563),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_520),
.B(n_453),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_551),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_520),
.B(n_453),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_595),
.Y(n_701)
);

OAI22xp33_ASAP7_75t_L g702 ( 
.A1(n_592),
.A2(n_335),
.B1(n_338),
.B2(n_333),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_551),
.Y(n_703)
);

BUFx8_ASAP7_75t_SL g704 ( 
.A(n_548),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_552),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_569),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_546),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_552),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_553),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_602),
.B(n_516),
.Y(n_710)
);

AOI21x1_ASAP7_75t_L g711 ( 
.A1(n_553),
.A2(n_242),
.B(n_241),
.Y(n_711)
);

NAND3xp33_ASAP7_75t_L g712 ( 
.A(n_602),
.B(n_490),
.C(n_464),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_546),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_590),
.Y(n_714)
);

OAI22x1_ASAP7_75t_L g715 ( 
.A1(n_604),
.A2(n_395),
.B1(n_393),
.B2(n_464),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_542),
.Y(n_716)
);

AO21x2_ASAP7_75t_L g717 ( 
.A1(n_539),
.A2(n_251),
.B(n_244),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_590),
.A2(n_510),
.B1(n_512),
.B2(n_420),
.Y(n_718)
);

CKINVDCx11_ASAP7_75t_R g719 ( 
.A(n_522),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_546),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_549),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_549),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_556),
.B(n_490),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_596),
.B(n_497),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_549),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_555),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_555),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_555),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_560),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_556),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_559),
.Y(n_731)
);

BUFx4f_ASAP7_75t_L g732 ( 
.A(n_547),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_559),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_560),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_562),
.B(n_497),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_596),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_562),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_596),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_596),
.B(n_500),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_598),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_594),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_560),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_542),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_572),
.B(n_499),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_572),
.B(n_499),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_598),
.B(n_517),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_598),
.B(n_517),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_567),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_566),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_598),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_575),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_542),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_567),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_567),
.Y(n_754)
);

OR2x6_ASAP7_75t_L g755 ( 
.A(n_644),
.B(n_426),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_714),
.B(n_545),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_714),
.B(n_736),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_612),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_693),
.B(n_478),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_706),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_706),
.Y(n_761)
);

BUFx5_ASAP7_75t_L g762 ( 
.A(n_686),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_612),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_SL g764 ( 
.A(n_618),
.B(n_599),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_736),
.B(n_545),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_738),
.B(n_545),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_738),
.B(n_545),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_624),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_624),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_661),
.B(n_429),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_740),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_740),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_627),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_618),
.B(n_511),
.Y(n_774)
);

OAI22xp33_ASAP7_75t_L g775 ( 
.A1(n_664),
.A2(n_432),
.B1(n_436),
.B2(n_426),
.Y(n_775)
);

AND2x2_ASAP7_75t_SL g776 ( 
.A(n_675),
.B(n_263),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_641),
.B(n_611),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_627),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_628),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_SL g780 ( 
.A(n_626),
.B(n_407),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_661),
.B(n_222),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_L g782 ( 
.A(n_669),
.B(n_267),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_611),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_750),
.B(n_558),
.Y(n_784)
);

BUFx5_ASAP7_75t_L g785 ( 
.A(n_686),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_SL g786 ( 
.A(n_610),
.B(n_259),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_696),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_750),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_694),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_628),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_630),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_662),
.B(n_436),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_751),
.B(n_566),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_751),
.B(n_568),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_641),
.B(n_508),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_677),
.B(n_508),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_669),
.B(n_568),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_648),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_693),
.B(n_481),
.Y(n_799)
);

AND2x6_ASAP7_75t_L g800 ( 
.A(n_648),
.B(n_619),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_606),
.B(n_593),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_704),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_644),
.B(n_515),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_664),
.B(n_222),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_606),
.B(n_593),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_613),
.B(n_593),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_613),
.B(n_593),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_619),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_675),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_625),
.B(n_558),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_632),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_694),
.B(n_515),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_739),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_672),
.B(n_223),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_625),
.B(n_558),
.Y(n_815)
);

INVx8_ASAP7_75t_L g816 ( 
.A(n_623),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_672),
.B(n_223),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_635),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_640),
.B(n_558),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_615),
.B(n_224),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_614),
.A2(n_349),
.B1(n_210),
.B2(n_233),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_616),
.B(n_224),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_723),
.B(n_227),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_635),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_735),
.B(n_227),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_739),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_640),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_642),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_655),
.B(n_571),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_670),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_655),
.B(n_571),
.Y(n_831)
);

AOI211xp5_ASAP7_75t_L g832 ( 
.A1(n_608),
.A2(n_486),
.B(n_482),
.C(n_483),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_719),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_659),
.B(n_571),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_659),
.B(n_571),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_619),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_688),
.A2(n_252),
.B1(n_334),
.B2(n_284),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_744),
.B(n_328),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_663),
.B(n_601),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_745),
.B(n_228),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_633),
.B(n_228),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_L g842 ( 
.A(n_679),
.B(n_268),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_676),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_637),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_636),
.B(n_229),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_663),
.B(n_601),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_651),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_637),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_666),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_666),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_668),
.B(n_601),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_668),
.Y(n_852)
);

NOR2x1p5_ASAP7_75t_L g853 ( 
.A(n_712),
.B(n_395),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_724),
.A2(n_301),
.B1(n_278),
.B2(n_276),
.Y(n_854)
);

AND2x6_ASAP7_75t_SL g855 ( 
.A(n_644),
.B(n_484),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_673),
.B(n_601),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_676),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_673),
.B(n_575),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_674),
.B(n_684),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_676),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_638),
.Y(n_861)
);

INVx8_ASAP7_75t_L g862 ( 
.A(n_623),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_652),
.A2(n_299),
.B(n_264),
.C(n_271),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_638),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_692),
.B(n_576),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_692),
.B(n_576),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_741),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_639),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_699),
.B(n_578),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_609),
.B(n_229),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_620),
.B(n_230),
.Y(n_871)
);

NAND3xp33_ASAP7_75t_L g872 ( 
.A(n_658),
.B(n_350),
.C(n_347),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_746),
.A2(n_305),
.B1(n_294),
.B2(n_290),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_639),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_676),
.B(n_503),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_703),
.B(n_578),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_647),
.B(n_504),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_747),
.B(n_230),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_703),
.B(n_705),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_652),
.A2(n_379),
.B(n_295),
.C(n_327),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_680),
.B(n_231),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_705),
.B(n_580),
.Y(n_882)
);

INVx8_ASAP7_75t_L g883 ( 
.A(n_623),
.Y(n_883)
);

NAND2xp33_ASAP7_75t_SL g884 ( 
.A(n_629),
.B(n_353),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_644),
.B(n_505),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_708),
.B(n_580),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_645),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_708),
.B(n_583),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_645),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_709),
.B(n_730),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_698),
.B(n_231),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_691),
.Y(n_892)
);

NAND2xp33_ASAP7_75t_L g893 ( 
.A(n_700),
.B(n_272),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_741),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_652),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_709),
.B(n_730),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_718),
.B(n_702),
.Y(n_897)
);

OAI22xp33_ASAP7_75t_L g898 ( 
.A1(n_647),
.A2(n_289),
.B1(n_367),
.B2(n_363),
.Y(n_898)
);

INVxp33_ASAP7_75t_SL g899 ( 
.A(n_610),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_731),
.B(n_583),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_731),
.B(n_583),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_653),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_647),
.A2(n_352),
.B1(n_274),
.B2(n_279),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_667),
.B(n_682),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_733),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_737),
.A2(n_329),
.B1(n_360),
.B2(n_390),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_737),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_690),
.B(n_234),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_647),
.A2(n_287),
.B1(n_280),
.B2(n_285),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_749),
.B(n_717),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_749),
.Y(n_911)
);

OR2x2_ASAP7_75t_L g912 ( 
.A(n_621),
.B(n_500),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_710),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_710),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_717),
.B(n_547),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_678),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_717),
.B(n_547),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_798),
.Y(n_918)
);

BUFx10_ASAP7_75t_L g919 ( 
.A(n_796),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_809),
.Y(n_920)
);

INVx4_ASAP7_75t_L g921 ( 
.A(n_808),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_783),
.B(n_622),
.Y(n_922)
);

AND2x6_ASAP7_75t_SL g923 ( 
.A(n_845),
.B(n_501),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_758),
.Y(n_924)
);

OR2x6_ASAP7_75t_SL g925 ( 
.A(n_774),
.B(n_701),
.Y(n_925)
);

O2A1O1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_904),
.A2(n_607),
.B(n_646),
.C(n_650),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_827),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_761),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_795),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_859),
.B(n_622),
.Y(n_930)
);

BUFx4f_ASAP7_75t_L g931 ( 
.A(n_816),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_859),
.B(n_622),
.Y(n_932)
);

BUFx2_ASAP7_75t_SL g933 ( 
.A(n_867),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_912),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_777),
.Y(n_935)
);

AND2x4_ASAP7_75t_SL g936 ( 
.A(n_808),
.B(n_678),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_763),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_828),
.Y(n_938)
);

NAND2xp33_ASAP7_75t_L g939 ( 
.A(n_800),
.B(n_686),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_892),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_879),
.B(n_617),
.Y(n_941)
);

BUFx2_ASAP7_75t_SL g942 ( 
.A(n_833),
.Y(n_942)
);

AND2x6_ASAP7_75t_L g943 ( 
.A(n_910),
.B(n_293),
.Y(n_943)
);

AND2x6_ASAP7_75t_L g944 ( 
.A(n_910),
.B(n_915),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_812),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_879),
.B(n_617),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_768),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_769),
.Y(n_948)
);

AND2x6_ASAP7_75t_SL g949 ( 
.A(n_841),
.B(n_501),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_816),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_890),
.B(n_617),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_773),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_849),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_808),
.B(n_678),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_836),
.B(n_761),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_896),
.B(n_792),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_850),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_852),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_789),
.B(n_838),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_778),
.Y(n_960)
);

NAND2x1p5_ASAP7_75t_L g961 ( 
.A(n_836),
.B(n_631),
.Y(n_961)
);

NAND3xp33_ASAP7_75t_SL g962 ( 
.A(n_780),
.B(n_701),
.C(n_695),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_905),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_907),
.B(n_911),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_800),
.A2(n_650),
.B1(n_646),
.B2(n_686),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_761),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_779),
.Y(n_967)
);

NOR2xp67_ASAP7_75t_L g968 ( 
.A(n_847),
.B(n_715),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_914),
.B(n_356),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_881),
.B(n_649),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_790),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_891),
.B(n_788),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_791),
.Y(n_973)
);

NAND3xp33_ASAP7_75t_L g974 ( 
.A(n_821),
.B(n_660),
.C(n_607),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_800),
.A2(n_686),
.B1(n_687),
.B2(n_715),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_800),
.Y(n_976)
);

BUFx2_ASAP7_75t_SL g977 ( 
.A(n_802),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_877),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_888),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_888),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_762),
.B(n_732),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_811),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_800),
.A2(n_686),
.B1(n_687),
.B2(n_377),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_787),
.B(n_649),
.Y(n_984)
);

AND2x6_ASAP7_75t_SL g985 ( 
.A(n_755),
.B(n_697),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_757),
.A2(n_405),
.B1(n_341),
.B2(n_345),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_SL g987 ( 
.A1(n_786),
.A2(n_697),
.B1(n_366),
.B2(n_259),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_900),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_900),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_897),
.B(n_357),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_R g991 ( 
.A(n_764),
.B(n_634),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_894),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_776),
.B(n_368),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_804),
.B(n_814),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_762),
.B(n_732),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_901),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_817),
.B(n_372),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_818),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_759),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_816),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_901),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_757),
.A2(n_337),
.B1(n_410),
.B2(n_331),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_813),
.B(n_716),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_826),
.A2(n_687),
.B1(n_686),
.B2(n_332),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_899),
.Y(n_1005)
);

CKINVDCx20_ASAP7_75t_R g1006 ( 
.A(n_862),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_913),
.B(n_373),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_793),
.B(n_716),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_794),
.B(n_797),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_760),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_895),
.A2(n_687),
.B1(n_743),
.B2(n_716),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_762),
.B(n_732),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_843),
.B(n_586),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_SL g1014 ( 
.A(n_862),
.B(n_366),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_824),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_857),
.B(n_586),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_870),
.A2(n_687),
.B1(n_310),
.B2(n_293),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_770),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_860),
.B(n_588),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_875),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_771),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_862),
.Y(n_1022)
);

BUFx12f_ASAP7_75t_L g1023 ( 
.A(n_855),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_858),
.B(n_743),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_772),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_SL g1026 ( 
.A1(n_839),
.A2(n_754),
.B(n_753),
.C(n_748),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_846),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_846),
.A2(n_687),
.B1(n_310),
.B2(n_293),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_851),
.Y(n_1029)
);

NOR3xp33_ASAP7_75t_SL g1030 ( 
.A(n_898),
.B(n_382),
.C(n_378),
.Y(n_1030)
);

NOR2x1p5_ASAP7_75t_L g1031 ( 
.A(n_872),
.B(n_384),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_858),
.B(n_743),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_759),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_851),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_844),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_848),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_840),
.B(n_386),
.Y(n_1037)
);

INVx2_ASAP7_75t_SL g1038 ( 
.A(n_799),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_762),
.B(n_643),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_799),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_762),
.B(n_785),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_883),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_856),
.Y(n_1043)
);

NAND2xp33_ASAP7_75t_L g1044 ( 
.A(n_762),
.B(n_687),
.Y(n_1044)
);

INVx5_ASAP7_75t_L g1045 ( 
.A(n_883),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_861),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_864),
.Y(n_1047)
);

INVxp67_ASAP7_75t_L g1048 ( 
.A(n_885),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_853),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_865),
.B(n_683),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_868),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_883),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_916),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_830),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_865),
.B(n_683),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_785),
.B(n_643),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_874),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_781),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_866),
.B(n_685),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_856),
.A2(n_310),
.B1(n_293),
.B2(n_748),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_755),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_803),
.B(n_588),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_887),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_866),
.B(n_685),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_803),
.Y(n_1065)
);

BUFx12f_ASAP7_75t_L g1066 ( 
.A(n_803),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_810),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_810),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_889),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_902),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_815),
.Y(n_1071)
);

NAND2xp33_ASAP7_75t_L g1072 ( 
.A(n_785),
.B(n_643),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_SL g1073 ( 
.A1(n_878),
.A2(n_869),
.B(n_882),
.C(n_876),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_820),
.A2(n_631),
.B1(n_297),
.B2(n_298),
.Y(n_1074)
);

NOR2xp67_ASAP7_75t_L g1075 ( 
.A(n_837),
.B(n_634),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_822),
.B(n_387),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_815),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_908),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_819),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_819),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_SL g1081 ( 
.A(n_775),
.B(n_366),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_829),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_829),
.Y(n_1083)
);

BUFx12f_ASAP7_75t_L g1084 ( 
.A(n_832),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_869),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_876),
.B(n_689),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_823),
.B(n_389),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_756),
.A2(n_234),
.B1(n_237),
.B2(n_396),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_785),
.B(n_643),
.Y(n_1089)
);

AO22x1_ASAP7_75t_L g1090 ( 
.A1(n_882),
.A2(n_406),
.B1(n_396),
.B2(n_397),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_831),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_871),
.B(n_237),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_884),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_842),
.A2(n_893),
.B1(n_825),
.B2(n_782),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_886),
.B(n_689),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_831),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_SL g1097 ( 
.A1(n_903),
.A2(n_397),
.B1(n_398),
.B2(n_399),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_944),
.B(n_979),
.Y(n_1098)
);

OAI22x1_ASAP7_75t_L g1099 ( 
.A1(n_993),
.A2(n_909),
.B1(n_873),
.B2(n_854),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_920),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_L g1101 ( 
.A(n_993),
.B(n_906),
.C(n_880),
.Y(n_1101)
);

NOR3xp33_ASAP7_75t_L g1102 ( 
.A(n_962),
.B(n_863),
.C(n_886),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1072),
.A2(n_917),
.B(n_915),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_920),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_924),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_992),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1048),
.B(n_956),
.Y(n_1107)
);

NOR2x1_ASAP7_75t_L g1108 ( 
.A(n_933),
.B(n_801),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_1005),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_966),
.Y(n_1110)
);

NOR3xp33_ASAP7_75t_L g1111 ( 
.A(n_987),
.B(n_399),
.C(n_398),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_990),
.A2(n_805),
.B(n_806),
.C(n_807),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1048),
.B(n_834),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_930),
.A2(n_917),
.B(n_756),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_927),
.Y(n_1115)
);

OAI22x1_ASAP7_75t_L g1116 ( 
.A1(n_994),
.A2(n_400),
.B1(n_412),
.B2(n_403),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_944),
.B(n_834),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_977),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1020),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_980),
.A2(n_835),
.B1(n_784),
.B2(n_767),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_1020),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_990),
.A2(n_784),
.B(n_767),
.C(n_766),
.Y(n_1122)
);

NOR2xp67_ASAP7_75t_L g1123 ( 
.A(n_1045),
.B(n_835),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_994),
.A2(n_766),
.B(n_765),
.C(n_400),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_SL g1125 ( 
.A1(n_987),
.A2(n_286),
.B1(n_307),
.B2(n_308),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1062),
.B(n_765),
.Y(n_1126)
);

INVx1_ASAP7_75t_SL g1127 ( 
.A(n_940),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_932),
.A2(n_631),
.B(n_752),
.Y(n_1128)
);

BUFx12f_ASAP7_75t_L g1129 ( 
.A(n_985),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_1037),
.A2(n_365),
.B(n_344),
.C(n_343),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_945),
.A2(n_729),
.B(n_754),
.C(n_753),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_959),
.B(n_785),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_988),
.A2(n_310),
.B1(n_711),
.B2(n_742),
.Y(n_1133)
);

NAND2x1_ASAP7_75t_L g1134 ( 
.A(n_921),
.B(n_643),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1085),
.B(n_707),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1009),
.B(n_713),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_945),
.A2(n_729),
.B(n_734),
.C(n_728),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_989),
.A2(n_310),
.B1(n_711),
.B2(n_742),
.Y(n_1138)
);

O2A1O1Ixp5_ASAP7_75t_L g1139 ( 
.A1(n_972),
.A2(n_720),
.B(n_721),
.C(n_734),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_950),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_1037),
.B(n_392),
.C(n_391),
.Y(n_1141)
);

BUFx12f_ASAP7_75t_L g1142 ( 
.A(n_1066),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_937),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_929),
.B(n_785),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_996),
.A2(n_1001),
.B1(n_1077),
.B2(n_1082),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_974),
.A2(n_404),
.B1(n_362),
.B2(n_388),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_948),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_R g1148 ( 
.A(n_1042),
.B(n_312),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_919),
.B(n_315),
.Y(n_1149)
);

INVx1_ASAP7_75t_SL g1150 ( 
.A(n_1018),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_919),
.B(n_323),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_966),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_950),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_935),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_966),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_938),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_941),
.A2(n_752),
.B(n_605),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_935),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_997),
.A2(n_728),
.B(n_727),
.C(n_726),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1077),
.B(n_722),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_934),
.B(n_325),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1082),
.B(n_1091),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1062),
.B(n_589),
.Y(n_1163)
);

INVx5_ASAP7_75t_L g1164 ( 
.A(n_976),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1091),
.A2(n_727),
.B1(n_726),
.B2(n_725),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_997),
.A2(n_336),
.B(n_371),
.C(n_369),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1027),
.B(n_725),
.Y(n_1167)
);

AOI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1075),
.A2(n_656),
.B(n_681),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1073),
.A2(n_589),
.B(n_681),
.C(n_654),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1058),
.B(n_342),
.Y(n_1170)
);

AND3x1_ASAP7_75t_L g1171 ( 
.A(n_1081),
.B(n_600),
.C(n_591),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1029),
.B(n_653),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1083),
.B(n_654),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1061),
.B(n_591),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1073),
.A2(n_656),
.B(n_665),
.C(n_657),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_953),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_978),
.B(n_591),
.Y(n_1177)
);

NOR3xp33_ASAP7_75t_SL g1178 ( 
.A(n_1093),
.B(n_355),
.C(n_364),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1061),
.B(n_600),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_946),
.A2(n_752),
.B(n_605),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_951),
.A2(n_752),
.B(n_605),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_SL g1182 ( 
.A(n_942),
.B(n_404),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_1000),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_957),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1040),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_999),
.B(n_374),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1040),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1092),
.A2(n_657),
.B(n_665),
.C(n_671),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_958),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_963),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1054),
.Y(n_1191)
);

INVx3_ASAP7_75t_SL g1192 ( 
.A(n_1053),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1096),
.B(n_1034),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_1000),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1060),
.A2(n_600),
.B1(n_671),
.B2(n_539),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_918),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1033),
.B(n_404),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1038),
.B(n_542),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_966),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1043),
.A2(n_539),
.B(n_605),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1067),
.B(n_547),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1068),
.B(n_547),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_921),
.B(n_542),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1060),
.A2(n_554),
.B1(n_2),
.B2(n_5),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_952),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_964),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1071),
.B(n_554),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1084),
.B(n_0),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1045),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1092),
.A2(n_926),
.B(n_1079),
.C(n_1080),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_969),
.A2(n_554),
.B(n_9),
.C(n_10),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_952),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_969),
.B(n_554),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_960),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1024),
.A2(n_526),
.B(n_178),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1088),
.A2(n_7),
.B(n_10),
.C(n_12),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1050),
.B(n_7),
.Y(n_1217)
);

NOR3xp33_ASAP7_75t_L g1218 ( 
.A(n_1097),
.B(n_15),
.C(n_16),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_SL g1219 ( 
.A1(n_1094),
.A2(n_177),
.B(n_173),
.C(n_164),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_981),
.A2(n_526),
.B(n_159),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1055),
.B(n_17),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1028),
.A2(n_18),
.B1(n_20),
.B2(n_23),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_923),
.B(n_24),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1059),
.B(n_156),
.Y(n_1224)
);

NAND3xp33_ASAP7_75t_SL g1225 ( 
.A(n_1014),
.B(n_25),
.C(n_26),
.Y(n_1225)
);

INVxp67_ASAP7_75t_SL g1226 ( 
.A(n_961),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1064),
.B(n_152),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1086),
.B(n_140),
.Y(n_1228)
);

OAI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_968),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1095),
.B(n_30),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1028),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1010),
.B(n_35),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1045),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1078),
.B(n_37),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_973),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1010),
.B(n_39),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_973),
.Y(n_1237)
);

NOR3xp33_ASAP7_75t_SL g1238 ( 
.A(n_954),
.B(n_39),
.C(n_41),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_1049),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_995),
.A2(n_526),
.B(n_78),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1032),
.B(n_42),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1045),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_949),
.B(n_43),
.Y(n_1243)
);

NAND3xp33_ASAP7_75t_L g1244 ( 
.A(n_1102),
.B(n_1030),
.C(n_1090),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1107),
.B(n_1007),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1150),
.B(n_1087),
.Y(n_1246)
);

AOI21xp33_ASAP7_75t_L g1247 ( 
.A1(n_1099),
.A2(n_1076),
.B(n_986),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1103),
.A2(n_970),
.B(n_939),
.Y(n_1248)
);

OA21x2_ASAP7_75t_L g1249 ( 
.A1(n_1215),
.A2(n_1210),
.B(n_1200),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1114),
.A2(n_995),
.B(n_1012),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1168),
.A2(n_1128),
.B(n_1175),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1106),
.Y(n_1252)
);

NAND3xp33_ASAP7_75t_L g1253 ( 
.A(n_1111),
.B(n_1030),
.C(n_1002),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1104),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1154),
.B(n_1013),
.Y(n_1255)
);

BUFx10_ASAP7_75t_L g1256 ( 
.A(n_1109),
.Y(n_1256)
);

AOI221x1_ASAP7_75t_L g1257 ( 
.A1(n_1218),
.A2(n_1025),
.B1(n_1021),
.B2(n_1008),
.C(n_922),
.Y(n_1257)
);

AND3x4_ASAP7_75t_L g1258 ( 
.A(n_1140),
.B(n_1022),
.C(n_925),
.Y(n_1258)
);

AO22x2_ASAP7_75t_L g1259 ( 
.A1(n_1225),
.A2(n_954),
.B1(n_955),
.B2(n_1013),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1122),
.A2(n_1012),
.B(n_1044),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1112),
.A2(n_1041),
.B(n_961),
.Y(n_1261)
);

OAI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1182),
.A2(n_1065),
.B1(n_1023),
.B2(n_931),
.Y(n_1262)
);

CKINVDCx11_ASAP7_75t_R g1263 ( 
.A(n_1192),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_1100),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1115),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1136),
.A2(n_1041),
.B(n_1056),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1213),
.A2(n_1089),
.B(n_1039),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_SL g1268 ( 
.A1(n_1215),
.A2(n_976),
.B(n_965),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1101),
.A2(n_975),
.B(n_936),
.C(n_1031),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1156),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1117),
.A2(n_1026),
.B(n_943),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1206),
.B(n_1016),
.Y(n_1272)
);

INVx4_ASAP7_75t_L g1273 ( 
.A(n_1209),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1127),
.B(n_936),
.Y(n_1274)
);

NOR3xp33_ASAP7_75t_L g1275 ( 
.A(n_1197),
.B(n_955),
.C(n_1052),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1224),
.A2(n_1056),
.B(n_1026),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1176),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1224),
.A2(n_1003),
.B(n_984),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1121),
.B(n_1016),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1184),
.Y(n_1280)
);

NAND3x1_ASAP7_75t_L g1281 ( 
.A(n_1223),
.B(n_1006),
.C(n_928),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1113),
.B(n_1019),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1227),
.A2(n_983),
.B(n_1070),
.Y(n_1283)
);

OAI22x1_ASAP7_75t_L g1284 ( 
.A1(n_1243),
.A2(n_1019),
.B1(n_1052),
.B2(n_1011),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1189),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1157),
.A2(n_982),
.B(n_1070),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1180),
.A2(n_982),
.B(n_998),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1222),
.A2(n_1017),
.B(n_1074),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1193),
.B(n_971),
.Y(n_1289)
);

A2O1A1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1124),
.A2(n_1017),
.B(n_931),
.C(n_947),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1181),
.A2(n_998),
.B(n_1015),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1162),
.B(n_967),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1117),
.A2(n_943),
.B(n_1015),
.Y(n_1293)
);

O2A1O1Ixp5_ASAP7_75t_L g1294 ( 
.A1(n_1133),
.A2(n_1047),
.B(n_1063),
.C(n_1057),
.Y(n_1294)
);

OAI21xp33_ASAP7_75t_L g1295 ( 
.A1(n_1234),
.A2(n_991),
.B(n_1022),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1162),
.A2(n_1069),
.B1(n_1063),
.B2(n_1057),
.Y(n_1296)
);

BUFx12f_ASAP7_75t_L g1297 ( 
.A(n_1118),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1141),
.A2(n_1051),
.B(n_1069),
.C(n_1046),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1126),
.B(n_1047),
.Y(n_1299)
);

O2A1O1Ixp5_ASAP7_75t_L g1300 ( 
.A1(n_1133),
.A2(n_1036),
.B(n_1035),
.C(n_1046),
.Y(n_1300)
);

AO32x2_ASAP7_75t_L g1301 ( 
.A1(n_1138),
.A2(n_943),
.A3(n_991),
.B1(n_1035),
.B2(n_1036),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1126),
.B(n_943),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1098),
.A2(n_943),
.B(n_1004),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1228),
.A2(n_77),
.B(n_132),
.Y(n_1304)
);

BUFx10_ASAP7_75t_L g1305 ( 
.A(n_1149),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1158),
.B(n_45),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1145),
.B(n_46),
.Y(n_1307)
);

NOR2xp67_ASAP7_75t_L g1308 ( 
.A(n_1164),
.B(n_76),
.Y(n_1308)
);

AO21x2_ASAP7_75t_L g1309 ( 
.A1(n_1200),
.A2(n_89),
.B(n_124),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1145),
.B(n_48),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1228),
.A2(n_64),
.B(n_122),
.Y(n_1311)
);

INVx4_ASAP7_75t_L g1312 ( 
.A(n_1209),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1196),
.B(n_48),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1153),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1142),
.Y(n_1315)
);

OA22x2_ASAP7_75t_L g1316 ( 
.A1(n_1222),
.A2(n_50),
.B1(n_58),
.B2(n_59),
.Y(n_1316)
);

AO22x2_ASAP7_75t_L g1317 ( 
.A1(n_1231),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1190),
.B(n_1217),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1174),
.B(n_109),
.Y(n_1319)
);

AOI221x1_ASAP7_75t_L g1320 ( 
.A1(n_1211),
.A2(n_1138),
.B1(n_1204),
.B2(n_1116),
.C(n_1231),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1120),
.A2(n_1098),
.B(n_1226),
.Y(n_1321)
);

AOI221x1_ASAP7_75t_L g1322 ( 
.A1(n_1204),
.A2(n_117),
.B1(n_1241),
.B2(n_1120),
.C(n_1230),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1165),
.A2(n_1195),
.A3(n_1221),
.B(n_1201),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1169),
.A2(n_1165),
.B(n_1139),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1174),
.B(n_1179),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1214),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1164),
.Y(n_1327)
);

O2A1O1Ixp5_ASAP7_75t_SL g1328 ( 
.A1(n_1132),
.A2(n_1198),
.B(n_1151),
.C(n_1203),
.Y(n_1328)
);

AO31x2_ASAP7_75t_L g1329 ( 
.A1(n_1195),
.A2(n_1207),
.A3(n_1202),
.B(n_1236),
.Y(n_1329)
);

O2A1O1Ixp33_ASAP7_75t_SL g1330 ( 
.A1(n_1219),
.A2(n_1144),
.B(n_1130),
.C(n_1166),
.Y(n_1330)
);

AND2x2_ASAP7_75t_SL g1331 ( 
.A(n_1171),
.B(n_1146),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1183),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1119),
.B(n_1163),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1160),
.B(n_1167),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1229),
.A2(n_1216),
.B(n_1170),
.C(n_1238),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1163),
.B(n_1161),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1185),
.B(n_1187),
.Y(n_1337)
);

AO32x2_ASAP7_75t_L g1338 ( 
.A1(n_1125),
.A2(n_1239),
.A3(n_1232),
.B1(n_1188),
.B2(n_1159),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_SL g1339 ( 
.A1(n_1233),
.A2(n_1242),
.B(n_1135),
.Y(n_1339)
);

AOI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1123),
.A2(n_1172),
.B(n_1173),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1131),
.A2(n_1137),
.B(n_1108),
.C(n_1220),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1177),
.B(n_1179),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1172),
.A2(n_1240),
.B(n_1134),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1191),
.B(n_1148),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1143),
.A2(n_1205),
.B(n_1237),
.Y(n_1345)
);

AOI221xp5_ASAP7_75t_SL g1346 ( 
.A1(n_1147),
.A2(n_1212),
.B1(n_1235),
.B2(n_1186),
.C(n_1155),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1110),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1194),
.Y(n_1348)
);

A2O1A1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1178),
.A2(n_1208),
.B(n_1164),
.C(n_1242),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1233),
.A2(n_1110),
.B(n_1152),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1110),
.B(n_1152),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1129),
.Y(n_1352)
);

NOR2x1_ASAP7_75t_SL g1353 ( 
.A(n_1155),
.B(n_1199),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1199),
.B(n_1107),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1115),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1103),
.A2(n_1114),
.B(n_1072),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1150),
.B(n_618),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1107),
.B(n_1206),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1133),
.A2(n_1138),
.A3(n_1210),
.B(n_1120),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1101),
.A2(n_990),
.B(n_994),
.C(n_1037),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1105),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1115),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1115),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1168),
.A2(n_1128),
.B(n_1175),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1107),
.B(n_1206),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1150),
.B(n_618),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1103),
.A2(n_1114),
.B(n_1072),
.Y(n_1367)
);

OAI22x1_ASAP7_75t_L g1368 ( 
.A1(n_1107),
.A2(n_550),
.B1(n_904),
.B2(n_993),
.Y(n_1368)
);

AO31x2_ASAP7_75t_L g1369 ( 
.A1(n_1133),
.A2(n_1138),
.A3(n_1210),
.B(n_1120),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_SL g1370 ( 
.A(n_1150),
.B(n_597),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_R g1371 ( 
.A(n_1118),
.B(n_741),
.Y(n_1371)
);

INVx1_ASAP7_75t_SL g1372 ( 
.A(n_1106),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1107),
.B(n_777),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1107),
.B(n_777),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1168),
.A2(n_1128),
.B(n_1175),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1206),
.A2(n_1193),
.B1(n_956),
.B2(n_1107),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1107),
.B(n_1206),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1115),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1103),
.A2(n_1114),
.B(n_1072),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1107),
.B(n_777),
.Y(n_1380)
);

AO31x2_ASAP7_75t_L g1381 ( 
.A1(n_1133),
.A2(n_1138),
.A3(n_1210),
.B(n_1120),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1210),
.A2(n_1122),
.B(n_1114),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1115),
.Y(n_1383)
);

NOR2xp67_ASAP7_75t_L g1384 ( 
.A(n_1141),
.B(n_1094),
.Y(n_1384)
);

INVx8_ASAP7_75t_L g1385 ( 
.A(n_1164),
.Y(n_1385)
);

O2A1O1Ixp33_ASAP7_75t_SL g1386 ( 
.A1(n_1210),
.A2(n_904),
.B(n_1124),
.C(n_1211),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_SL g1387 ( 
.A1(n_1210),
.A2(n_1122),
.B(n_932),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1103),
.A2(n_1114),
.B(n_1072),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1115),
.Y(n_1389)
);

NOR2x1_ASAP7_75t_SL g1390 ( 
.A(n_1209),
.B(n_1233),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1210),
.A2(n_1122),
.B(n_1114),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1115),
.Y(n_1392)
);

NOR2xp67_ASAP7_75t_SL g1393 ( 
.A(n_1118),
.B(n_933),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1107),
.B(n_1206),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1103),
.A2(n_1114),
.B(n_1072),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1168),
.A2(n_1128),
.B(n_1175),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1360),
.A2(n_1245),
.B(n_1244),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1265),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1373),
.B(n_1374),
.Y(n_1399)
);

AOI222xp33_ASAP7_75t_L g1400 ( 
.A1(n_1368),
.A2(n_1317),
.B1(n_1380),
.B2(n_1365),
.C1(n_1394),
.C2(n_1358),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1332),
.Y(n_1401)
);

OAI21xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1316),
.A2(n_1331),
.B(n_1247),
.Y(n_1402)
);

CKINVDCx6p67_ASAP7_75t_R g1403 ( 
.A(n_1263),
.Y(n_1403)
);

OR2x6_ASAP7_75t_L g1404 ( 
.A(n_1268),
.B(n_1385),
.Y(n_1404)
);

OAI21xp33_ASAP7_75t_SL g1405 ( 
.A1(n_1247),
.A2(n_1377),
.B(n_1310),
.Y(n_1405)
);

O2A1O1Ixp33_ASAP7_75t_SL g1406 ( 
.A1(n_1269),
.A2(n_1310),
.B(n_1307),
.C(n_1288),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_SL g1407 ( 
.A1(n_1307),
.A2(n_1318),
.B(n_1335),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1325),
.B(n_1319),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1396),
.A2(n_1287),
.B(n_1286),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1354),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1256),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1345),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1246),
.A2(n_1376),
.B1(n_1336),
.B2(n_1282),
.Y(n_1413)
);

OAI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1244),
.A2(n_1384),
.B(n_1376),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1272),
.B(n_1289),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1270),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1254),
.Y(n_1417)
);

INVx1_ASAP7_75t_SL g1418 ( 
.A(n_1372),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1356),
.A2(n_1379),
.B(n_1367),
.Y(n_1419)
);

O2A1O1Ixp33_ASAP7_75t_SL g1420 ( 
.A1(n_1288),
.A2(n_1290),
.B(n_1341),
.C(n_1253),
.Y(n_1420)
);

O2A1O1Ixp5_ASAP7_75t_L g1421 ( 
.A1(n_1382),
.A2(n_1391),
.B(n_1293),
.C(n_1388),
.Y(n_1421)
);

OAI211xp5_ASAP7_75t_L g1422 ( 
.A1(n_1257),
.A2(n_1320),
.B(n_1322),
.C(n_1253),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1372),
.B(n_1354),
.Y(n_1423)
);

OAI21xp33_ASAP7_75t_SL g1424 ( 
.A1(n_1384),
.A2(n_1328),
.B(n_1308),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1317),
.A2(n_1259),
.B1(n_1391),
.B2(n_1382),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1385),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1342),
.B(n_1279),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1337),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1395),
.A2(n_1387),
.B(n_1248),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1324),
.A2(n_1293),
.B(n_1300),
.Y(n_1430)
);

NAND2x1p5_ASAP7_75t_L g1431 ( 
.A(n_1327),
.B(n_1393),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1277),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1291),
.A2(n_1250),
.B(n_1343),
.Y(n_1433)
);

OR2x6_ASAP7_75t_L g1434 ( 
.A(n_1339),
.B(n_1284),
.Y(n_1434)
);

O2A1O1Ixp33_ASAP7_75t_SL g1435 ( 
.A1(n_1349),
.A2(n_1302),
.B(n_1303),
.C(n_1298),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1321),
.A2(n_1283),
.B(n_1386),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1261),
.A2(n_1278),
.B(n_1260),
.Y(n_1437)
);

OA21x2_ASAP7_75t_L g1438 ( 
.A1(n_1294),
.A2(n_1271),
.B(n_1276),
.Y(n_1438)
);

AOI22x1_ASAP7_75t_L g1439 ( 
.A1(n_1259),
.A2(n_1304),
.B1(n_1311),
.B2(n_1389),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1295),
.A2(n_1266),
.B(n_1267),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1305),
.A2(n_1295),
.B1(n_1313),
.B2(n_1249),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1357),
.A2(n_1366),
.B1(n_1370),
.B2(n_1255),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1271),
.A2(n_1340),
.B(n_1303),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1333),
.B(n_1252),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_SL g1445 ( 
.A1(n_1305),
.A2(n_1249),
.B1(n_1371),
.B2(n_1319),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1299),
.B(n_1325),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1306),
.B(n_1392),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1275),
.A2(n_1378),
.B1(n_1355),
.B2(n_1362),
.Y(n_1448)
);

BUFx3_ASAP7_75t_L g1449 ( 
.A(n_1314),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1334),
.A2(n_1350),
.B(n_1296),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1292),
.B(n_1274),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1280),
.Y(n_1452)
);

AO21x2_ASAP7_75t_L g1453 ( 
.A1(n_1330),
.A2(n_1309),
.B(n_1383),
.Y(n_1453)
);

NOR2x1_ASAP7_75t_R g1454 ( 
.A(n_1297),
.B(n_1315),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1258),
.A2(n_1281),
.B1(n_1262),
.B2(n_1344),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1285),
.B(n_1363),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1346),
.A2(n_1301),
.B(n_1359),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1361),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1346),
.A2(n_1264),
.B(n_1351),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1347),
.A2(n_1329),
.B(n_1323),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1353),
.Y(n_1461)
);

NAND2x1p5_ASAP7_75t_L g1462 ( 
.A(n_1273),
.B(n_1312),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1329),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1256),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1329),
.A2(n_1323),
.B(n_1309),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1301),
.A2(n_1381),
.B(n_1369),
.Y(n_1466)
);

CKINVDCx11_ASAP7_75t_R g1467 ( 
.A(n_1352),
.Y(n_1467)
);

O2A1O1Ixp33_ASAP7_75t_SL g1468 ( 
.A1(n_1301),
.A2(n_1338),
.B(n_1381),
.C(n_1369),
.Y(n_1468)
);

AOI21xp33_ASAP7_75t_L g1469 ( 
.A1(n_1273),
.A2(n_1312),
.B(n_1338),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1323),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1359),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1390),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1359),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1348),
.A2(n_1338),
.B1(n_1369),
.B2(n_1381),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1360),
.B(n_847),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1345),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1263),
.Y(n_1477)
);

AO31x2_ASAP7_75t_L g1478 ( 
.A1(n_1322),
.A2(n_1320),
.A3(n_1360),
.B(n_1276),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1345),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1345),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_1332),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1332),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1265),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1251),
.A2(n_1375),
.B(n_1364),
.Y(n_1484)
);

INVx6_ASAP7_75t_SL g1485 ( 
.A(n_1256),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1325),
.B(n_1319),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1251),
.A2(n_1375),
.B(n_1364),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1245),
.B(n_1358),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1345),
.Y(n_1489)
);

CKINVDCx16_ASAP7_75t_R g1490 ( 
.A(n_1371),
.Y(n_1490)
);

AO31x2_ASAP7_75t_L g1491 ( 
.A1(n_1322),
.A2(n_1320),
.A3(n_1360),
.B(n_1276),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_SL g1492 ( 
.A1(n_1307),
.A2(n_1310),
.B(n_1318),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1382),
.A2(n_1391),
.B(n_1324),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1368),
.A2(n_1218),
.B1(n_1317),
.B2(n_780),
.Y(n_1494)
);

BUFx2_ASAP7_75t_SL g1495 ( 
.A(n_1332),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1251),
.A2(n_1375),
.B(n_1364),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1252),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1265),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1368),
.A2(n_1218),
.B1(n_1317),
.B2(n_780),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1332),
.Y(n_1500)
);

OAI221xp5_ASAP7_75t_SL g1501 ( 
.A1(n_1360),
.A2(n_550),
.B1(n_847),
.B2(n_987),
.C(n_1218),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1251),
.A2(n_1375),
.B(n_1364),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_1263),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1385),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1251),
.A2(n_1375),
.B(n_1364),
.Y(n_1505)
);

AOI21xp33_ASAP7_75t_SL g1506 ( 
.A1(n_1368),
.A2(n_899),
.B(n_701),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1373),
.B(n_1374),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1251),
.A2(n_1375),
.B(n_1364),
.Y(n_1508)
);

BUFx8_ASAP7_75t_SL g1509 ( 
.A(n_1315),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1368),
.A2(n_1218),
.B1(n_1317),
.B2(n_780),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1345),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1382),
.A2(n_1391),
.B(n_1324),
.Y(n_1512)
);

BUFx5_ASAP7_75t_L g1513 ( 
.A(n_1326),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1385),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1325),
.B(n_1319),
.Y(n_1515)
);

AO21x2_ASAP7_75t_L g1516 ( 
.A1(n_1382),
.A2(n_1391),
.B(n_1293),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1332),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1345),
.Y(n_1518)
);

O2A1O1Ixp33_ASAP7_75t_SL g1519 ( 
.A1(n_1360),
.A2(n_1269),
.B(n_1211),
.C(n_1247),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1385),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1332),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1372),
.Y(n_1522)
);

BUFx3_ASAP7_75t_L g1523 ( 
.A(n_1332),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1373),
.B(n_1374),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1360),
.B(n_847),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1382),
.A2(n_1391),
.B(n_1324),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1373),
.B(n_1374),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1265),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1385),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1368),
.A2(n_1218),
.B1(n_1317),
.B2(n_780),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1251),
.A2(n_1375),
.B(n_1364),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1265),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1251),
.A2(n_1375),
.B(n_1364),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1263),
.Y(n_1534)
);

BUFx8_ASAP7_75t_L g1535 ( 
.A(n_1254),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1358),
.A2(n_1365),
.B1(n_1394),
.B2(n_1377),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1325),
.B(n_1319),
.Y(n_1537)
);

OAI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1360),
.A2(n_796),
.B(n_677),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1251),
.A2(n_1375),
.B(n_1364),
.Y(n_1539)
);

INVxp67_ASAP7_75t_SL g1540 ( 
.A(n_1334),
.Y(n_1540)
);

OAI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1251),
.A2(n_1375),
.B(n_1364),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1385),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1345),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1373),
.B(n_1374),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1345),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1358),
.A2(n_1365),
.B1(n_1394),
.B2(n_1377),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1265),
.Y(n_1547)
);

BUFx2_ASAP7_75t_R g1548 ( 
.A(n_1315),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1251),
.A2(n_1375),
.B(n_1364),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1345),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1265),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1251),
.A2(n_1375),
.B(n_1364),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1345),
.Y(n_1553)
);

CKINVDCx6p67_ASAP7_75t_R g1554 ( 
.A(n_1263),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1373),
.B(n_1374),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1399),
.B(n_1507),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1509),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_SL g1558 ( 
.A1(n_1538),
.A2(n_1546),
.B(n_1536),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1509),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1501),
.A2(n_1494),
.B1(n_1510),
.B2(n_1499),
.Y(n_1560)
);

O2A1O1Ixp33_ASAP7_75t_L g1561 ( 
.A1(n_1475),
.A2(n_1525),
.B(n_1506),
.C(n_1414),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1540),
.B(n_1410),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1494),
.A2(n_1499),
.B1(n_1510),
.B2(n_1530),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1398),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1530),
.A2(n_1425),
.B1(n_1488),
.B2(n_1540),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1428),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1416),
.Y(n_1567)
);

O2A1O1Ixp5_ASAP7_75t_L g1568 ( 
.A1(n_1422),
.A2(n_1525),
.B(n_1475),
.C(n_1440),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1408),
.B(n_1486),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1425),
.A2(n_1555),
.B1(n_1544),
.B2(n_1527),
.Y(n_1570)
);

INVx3_ASAP7_75t_SL g1571 ( 
.A(n_1477),
.Y(n_1571)
);

BUFx12f_ASAP7_75t_L g1572 ( 
.A(n_1467),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1405),
.B(n_1397),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1524),
.B(n_1447),
.Y(n_1574)
);

O2A1O1Ixp33_ASAP7_75t_L g1575 ( 
.A1(n_1413),
.A2(n_1420),
.B(n_1519),
.C(n_1407),
.Y(n_1575)
);

OA21x2_ASAP7_75t_L g1576 ( 
.A1(n_1421),
.A2(n_1437),
.B(n_1409),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1428),
.B(n_1444),
.Y(n_1577)
);

AOI211xp5_ASAP7_75t_L g1578 ( 
.A1(n_1455),
.A2(n_1420),
.B(n_1402),
.C(n_1519),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1423),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1446),
.B(n_1423),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1492),
.B(n_1415),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1458),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1429),
.A2(n_1516),
.B(n_1419),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1442),
.B(n_1427),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1406),
.A2(n_1404),
.B(n_1526),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1400),
.B(n_1441),
.Y(n_1586)
);

OAI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1441),
.A2(n_1439),
.B1(n_1451),
.B2(n_1448),
.C(n_1424),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1446),
.B(n_1515),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1474),
.B(n_1448),
.Y(n_1589)
);

O2A1O1Ixp33_ASAP7_75t_L g1590 ( 
.A1(n_1435),
.A2(n_1459),
.B(n_1469),
.C(n_1522),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1401),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1493),
.A2(n_1512),
.B(n_1526),
.Y(n_1592)
);

OR2x2_ASAP7_75t_SL g1593 ( 
.A(n_1490),
.B(n_1426),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1497),
.B(n_1418),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1432),
.B(n_1452),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1483),
.B(n_1498),
.Y(n_1596)
);

AOI21x1_ASAP7_75t_SL g1597 ( 
.A1(n_1471),
.A2(n_1515),
.B(n_1537),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1513),
.B(n_1456),
.Y(n_1598)
);

AOI21x1_ASAP7_75t_SL g1599 ( 
.A1(n_1471),
.A2(n_1515),
.B(n_1537),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1456),
.B(n_1417),
.Y(n_1600)
);

O2A1O1Ixp5_ASAP7_75t_L g1601 ( 
.A1(n_1470),
.A2(n_1473),
.B(n_1463),
.C(n_1472),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1528),
.Y(n_1602)
);

A2O1A1Ixp33_ASAP7_75t_SL g1603 ( 
.A1(n_1463),
.A2(n_1461),
.B(n_1470),
.C(n_1514),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1532),
.B(n_1547),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1551),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1493),
.A2(n_1512),
.B(n_1526),
.Y(n_1606)
);

BUFx3_ASAP7_75t_L g1607 ( 
.A(n_1401),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1445),
.B(n_1431),
.Y(n_1608)
);

AOI21x1_ASAP7_75t_SL g1609 ( 
.A1(n_1485),
.A2(n_1491),
.B(n_1478),
.Y(n_1609)
);

AOI221x1_ASAP7_75t_SL g1610 ( 
.A1(n_1478),
.A2(n_1491),
.B1(n_1468),
.B2(n_1485),
.C(n_1535),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_SL g1611 ( 
.A1(n_1404),
.A2(n_1464),
.B(n_1411),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1434),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1404),
.A2(n_1434),
.B1(n_1457),
.B2(n_1466),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1493),
.A2(n_1512),
.B(n_1435),
.Y(n_1614)
);

O2A1O1Ixp33_ASAP7_75t_L g1615 ( 
.A1(n_1434),
.A2(n_1500),
.B(n_1521),
.C(n_1481),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1478),
.B(n_1491),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1449),
.B(n_1462),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1457),
.A2(n_1466),
.B1(n_1485),
.B2(n_1495),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1513),
.B(n_1491),
.Y(n_1619)
);

O2A1O1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1468),
.A2(n_1517),
.B(n_1482),
.C(n_1523),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1513),
.B(n_1453),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1460),
.B(n_1517),
.Y(n_1622)
);

NOR2x1_ASAP7_75t_SL g1623 ( 
.A(n_1453),
.B(n_1542),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_SL g1624 ( 
.A1(n_1504),
.A2(n_1520),
.B(n_1542),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1482),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1535),
.Y(n_1626)
);

BUFx2_ASAP7_75t_SL g1627 ( 
.A(n_1503),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1462),
.B(n_1523),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1450),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1457),
.A2(n_1466),
.B1(n_1503),
.B2(n_1554),
.Y(n_1630)
);

O2A1O1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1412),
.A2(n_1476),
.B(n_1489),
.C(n_1550),
.Y(n_1631)
);

O2A1O1Ixp33_ASAP7_75t_L g1632 ( 
.A1(n_1479),
.A2(n_1511),
.B(n_1550),
.C(n_1545),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1438),
.B(n_1543),
.Y(n_1633)
);

O2A1O1Ixp33_ASAP7_75t_L g1634 ( 
.A1(n_1480),
.A2(n_1543),
.B(n_1518),
.C(n_1489),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1529),
.B(n_1553),
.Y(n_1635)
);

AOI21xp5_ASAP7_75t_SL g1636 ( 
.A1(n_1529),
.A2(n_1454),
.B(n_1477),
.Y(n_1636)
);

BUFx12f_ASAP7_75t_L g1637 ( 
.A(n_1534),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1529),
.B(n_1403),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1430),
.B(n_1529),
.Y(n_1639)
);

OA21x2_ASAP7_75t_L g1640 ( 
.A1(n_1502),
.A2(n_1539),
.B(n_1533),
.Y(n_1640)
);

CKINVDCx20_ASAP7_75t_R g1641 ( 
.A(n_1534),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1548),
.B(n_1430),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1535),
.A2(n_1552),
.B1(n_1549),
.B2(n_1484),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1487),
.A2(n_1496),
.B1(n_1508),
.B2(n_1531),
.Y(n_1644)
);

AOI221xp5_ASAP7_75t_L g1645 ( 
.A1(n_1541),
.A2(n_1501),
.B1(n_1368),
.B2(n_1499),
.C(n_1494),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_1505),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_SL g1647 ( 
.A1(n_1505),
.A2(n_1360),
.B(n_1538),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1433),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_SL g1649 ( 
.A1(n_1538),
.A2(n_1360),
.B(n_1376),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1410),
.B(n_1524),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1399),
.B(n_1507),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1399),
.B(n_1507),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1399),
.B(n_1507),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1408),
.B(n_1486),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1410),
.B(n_1524),
.Y(n_1655)
);

BUFx6f_ASAP7_75t_L g1656 ( 
.A(n_1401),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1399),
.B(n_1507),
.Y(n_1657)
);

CKINVDCx11_ASAP7_75t_R g1658 ( 
.A(n_1503),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1410),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1399),
.B(n_1507),
.Y(n_1660)
);

INVx5_ASAP7_75t_L g1661 ( 
.A(n_1404),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1540),
.B(n_1410),
.Y(n_1662)
);

O2A1O1Ixp33_ASAP7_75t_L g1663 ( 
.A1(n_1501),
.A2(n_1360),
.B(n_1538),
.C(n_904),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1410),
.B(n_1524),
.Y(n_1664)
);

AO21x1_ASAP7_75t_L g1665 ( 
.A1(n_1538),
.A2(n_1525),
.B(n_1475),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1501),
.A2(n_1499),
.B1(n_1510),
.B2(n_1494),
.Y(n_1666)
);

INVx1_ASAP7_75t_SL g1667 ( 
.A(n_1410),
.Y(n_1667)
);

BUFx6f_ASAP7_75t_L g1668 ( 
.A(n_1401),
.Y(n_1668)
);

OA21x2_ASAP7_75t_L g1669 ( 
.A1(n_1436),
.A2(n_1465),
.B(n_1443),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1399),
.B(n_1507),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1593),
.Y(n_1671)
);

INVx2_ASAP7_75t_SL g1672 ( 
.A(n_1622),
.Y(n_1672)
);

AO21x2_ASAP7_75t_L g1673 ( 
.A1(n_1583),
.A2(n_1606),
.B(n_1592),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1665),
.A2(n_1666),
.B1(n_1560),
.B2(n_1563),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_SL g1675 ( 
.A1(n_1575),
.A2(n_1663),
.B(n_1561),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1619),
.B(n_1616),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_1661),
.Y(n_1677)
);

INVx3_ASAP7_75t_L g1678 ( 
.A(n_1635),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1560),
.A2(n_1666),
.B1(n_1563),
.B2(n_1578),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1601),
.Y(n_1680)
);

OAI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1558),
.A2(n_1568),
.B(n_1649),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1642),
.B(n_1564),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1562),
.B(n_1662),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1567),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1573),
.A2(n_1587),
.B(n_1647),
.Y(n_1685)
);

INVx3_ASAP7_75t_L g1686 ( 
.A(n_1635),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1562),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1605),
.B(n_1580),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1662),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1659),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1619),
.B(n_1589),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1598),
.B(n_1604),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1598),
.B(n_1667),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1602),
.Y(n_1694)
);

OA21x2_ASAP7_75t_L g1695 ( 
.A1(n_1614),
.A2(n_1621),
.B(n_1629),
.Y(n_1695)
);

OR2x6_ASAP7_75t_L g1696 ( 
.A(n_1585),
.B(n_1611),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1633),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1667),
.B(n_1630),
.Y(n_1698)
);

BUFx2_ASAP7_75t_L g1699 ( 
.A(n_1612),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1573),
.B(n_1566),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1595),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1639),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1596),
.Y(n_1703)
);

OR2x6_ASAP7_75t_L g1704 ( 
.A(n_1643),
.B(n_1613),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1639),
.Y(n_1705)
);

AO21x1_ASAP7_75t_SL g1706 ( 
.A1(n_1586),
.A2(n_1589),
.B(n_1581),
.Y(n_1706)
);

OA21x2_ASAP7_75t_L g1707 ( 
.A1(n_1587),
.A2(n_1586),
.B(n_1645),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1631),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1646),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1630),
.B(n_1574),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1618),
.Y(n_1711)
);

OR2x6_ASAP7_75t_L g1712 ( 
.A(n_1643),
.B(n_1615),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1632),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1634),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1579),
.B(n_1600),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1618),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1577),
.B(n_1650),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1582),
.Y(n_1718)
);

BUFx4f_ASAP7_75t_SL g1719 ( 
.A(n_1637),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1655),
.B(n_1664),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1640),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1640),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1581),
.B(n_1565),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1623),
.B(n_1648),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1584),
.B(n_1556),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1565),
.B(n_1570),
.Y(n_1726)
);

NAND2x1_ASAP7_75t_L g1727 ( 
.A(n_1624),
.B(n_1669),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1588),
.B(n_1670),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1610),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1610),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1576),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1651),
.B(n_1657),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1570),
.B(n_1590),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1576),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1652),
.B(n_1653),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1660),
.B(n_1645),
.Y(n_1736)
);

OAI21x1_ASAP7_75t_L g1737 ( 
.A1(n_1731),
.A2(n_1644),
.B(n_1609),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1702),
.B(n_1644),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1676),
.B(n_1608),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1727),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1702),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1705),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1684),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1684),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1705),
.B(n_1594),
.Y(n_1745)
);

OAI211xp5_ASAP7_75t_L g1746 ( 
.A1(n_1674),
.A2(n_1620),
.B(n_1658),
.C(n_1636),
.Y(n_1746)
);

BUFx2_ASAP7_75t_L g1747 ( 
.A(n_1724),
.Y(n_1747)
);

AOI222xp33_ASAP7_75t_L g1748 ( 
.A1(n_1679),
.A2(n_1572),
.B1(n_1626),
.B2(n_1571),
.C1(n_1638),
.C2(n_1625),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1687),
.B(n_1603),
.Y(n_1749)
);

AO21x2_ASAP7_75t_L g1750 ( 
.A1(n_1673),
.A2(n_1599),
.B(n_1597),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1697),
.B(n_1654),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1687),
.Y(n_1752)
);

NAND2x1p5_ASAP7_75t_L g1753 ( 
.A(n_1727),
.B(n_1617),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1695),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1689),
.Y(n_1755)
);

NAND2x1_ASAP7_75t_L g1756 ( 
.A(n_1696),
.B(n_1569),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1689),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1700),
.B(n_1628),
.Y(n_1758)
);

NOR2x1_ASAP7_75t_L g1759 ( 
.A(n_1681),
.B(n_1696),
.Y(n_1759)
);

BUFx2_ASAP7_75t_L g1760 ( 
.A(n_1724),
.Y(n_1760)
);

AND2x4_ASAP7_75t_SL g1761 ( 
.A(n_1677),
.B(n_1668),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1711),
.B(n_1607),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1700),
.B(n_1668),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1678),
.B(n_1686),
.Y(n_1764)
);

AOI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1679),
.A2(n_1627),
.B1(n_1591),
.B2(n_1668),
.C(n_1656),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1711),
.B(n_1656),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1692),
.B(n_1695),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1692),
.B(n_1569),
.Y(n_1768)
);

BUFx3_ASAP7_75t_L g1769 ( 
.A(n_1677),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1745),
.B(n_1717),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1746),
.A2(n_1681),
.B1(n_1733),
.B2(n_1726),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1748),
.A2(n_1707),
.B1(n_1726),
.B2(n_1733),
.Y(n_1772)
);

OA21x2_ASAP7_75t_L g1773 ( 
.A1(n_1737),
.A2(n_1722),
.B(n_1721),
.Y(n_1773)
);

AND2x4_ASAP7_75t_L g1774 ( 
.A(n_1747),
.B(n_1672),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_1761),
.Y(n_1775)
);

OAI332xp33_ASAP7_75t_L g1776 ( 
.A1(n_1749),
.A2(n_1723),
.A3(n_1729),
.B1(n_1730),
.B2(n_1691),
.B3(n_1680),
.C1(n_1694),
.C2(n_1675),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1746),
.A2(n_1675),
.B1(n_1671),
.B2(n_1685),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1765),
.A2(n_1671),
.B1(n_1759),
.B2(n_1685),
.Y(n_1778)
);

BUFx2_ASAP7_75t_L g1779 ( 
.A(n_1769),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_SL g1780 ( 
.A1(n_1739),
.A2(n_1707),
.B1(n_1671),
.B2(n_1723),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1741),
.Y(n_1781)
);

AOI222xp33_ASAP7_75t_SL g1782 ( 
.A1(n_1752),
.A2(n_1729),
.B1(n_1730),
.B2(n_1716),
.C1(n_1694),
.C2(n_1701),
.Y(n_1782)
);

NOR2x2_ASAP7_75t_L g1783 ( 
.A(n_1748),
.B(n_1712),
.Y(n_1783)
);

OAI221xp5_ASAP7_75t_L g1784 ( 
.A1(n_1759),
.A2(n_1707),
.B1(n_1712),
.B2(n_1696),
.C(n_1716),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_R g1785 ( 
.A(n_1762),
.B(n_1557),
.Y(n_1785)
);

OAI221xp5_ASAP7_75t_L g1786 ( 
.A1(n_1765),
.A2(n_1753),
.B1(n_1756),
.B2(n_1707),
.C(n_1712),
.Y(n_1786)
);

INVx2_ASAP7_75t_SL g1787 ( 
.A(n_1764),
.Y(n_1787)
);

INVx5_ASAP7_75t_L g1788 ( 
.A(n_1740),
.Y(n_1788)
);

INVxp67_ASAP7_75t_SL g1789 ( 
.A(n_1741),
.Y(n_1789)
);

OAI31xp33_ASAP7_75t_SL g1790 ( 
.A1(n_1739),
.A2(n_1710),
.A3(n_1736),
.B(n_1698),
.Y(n_1790)
);

OAI332xp33_ASAP7_75t_L g1791 ( 
.A1(n_1749),
.A2(n_1691),
.A3(n_1680),
.B1(n_1683),
.B2(n_1708),
.B3(n_1713),
.C1(n_1714),
.C2(n_1725),
.Y(n_1791)
);

AOI221xp5_ASAP7_75t_L g1792 ( 
.A1(n_1758),
.A2(n_1736),
.B1(n_1710),
.B2(n_1732),
.C(n_1683),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1743),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1743),
.Y(n_1794)
);

OAI33xp33_ASAP7_75t_L g1795 ( 
.A1(n_1752),
.A2(n_1703),
.A3(n_1701),
.B1(n_1690),
.B2(n_1717),
.B3(n_1718),
.Y(n_1795)
);

AOI221xp5_ASAP7_75t_L g1796 ( 
.A1(n_1758),
.A2(n_1698),
.B1(n_1703),
.B2(n_1682),
.C(n_1699),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1768),
.B(n_1751),
.Y(n_1797)
);

INVx3_ASAP7_75t_L g1798 ( 
.A(n_1764),
.Y(n_1798)
);

NAND4xp25_ASAP7_75t_L g1799 ( 
.A(n_1762),
.B(n_1699),
.C(n_1682),
.D(n_1688),
.Y(n_1799)
);

NAND4xp25_ASAP7_75t_L g1800 ( 
.A(n_1762),
.B(n_1688),
.C(n_1693),
.D(n_1715),
.Y(n_1800)
);

AOI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1763),
.A2(n_1715),
.B1(n_1735),
.B2(n_1728),
.C(n_1693),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1763),
.A2(n_1707),
.B1(n_1696),
.B2(n_1712),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1747),
.B(n_1760),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1744),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1766),
.A2(n_1709),
.B1(n_1696),
.B2(n_1712),
.Y(n_1805)
);

INVx1_ASAP7_75t_SL g1806 ( 
.A(n_1745),
.Y(n_1806)
);

AOI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1755),
.A2(n_1735),
.B1(n_1728),
.B2(n_1720),
.C(n_1672),
.Y(n_1807)
);

CKINVDCx16_ASAP7_75t_R g1808 ( 
.A(n_1751),
.Y(n_1808)
);

INVxp67_ASAP7_75t_L g1809 ( 
.A(n_1745),
.Y(n_1809)
);

INVx2_ASAP7_75t_SL g1810 ( 
.A(n_1788),
.Y(n_1810)
);

BUFx8_ASAP7_75t_L g1811 ( 
.A(n_1779),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1788),
.B(n_1740),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1788),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_L g1814 ( 
.A(n_1791),
.B(n_1776),
.Y(n_1814)
);

BUFx2_ASAP7_75t_L g1815 ( 
.A(n_1788),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1793),
.Y(n_1816)
);

OA21x2_ASAP7_75t_L g1817 ( 
.A1(n_1802),
.A2(n_1737),
.B(n_1734),
.Y(n_1817)
);

INVx4_ASAP7_75t_L g1818 ( 
.A(n_1775),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1794),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1804),
.Y(n_1820)
);

INVxp67_ASAP7_75t_SL g1821 ( 
.A(n_1781),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1789),
.Y(n_1822)
);

INVx2_ASAP7_75t_SL g1823 ( 
.A(n_1803),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1806),
.B(n_1767),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1809),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1803),
.B(n_1767),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1784),
.A2(n_1756),
.B(n_1750),
.Y(n_1827)
);

OAI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1772),
.A2(n_1753),
.B(n_1766),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1803),
.B(n_1740),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1770),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1792),
.B(n_1767),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1798),
.B(n_1740),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1773),
.Y(n_1833)
);

INVx4_ASAP7_75t_L g1834 ( 
.A(n_1775),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1785),
.B(n_1740),
.Y(n_1835)
);

INVxp67_ASAP7_75t_L g1836 ( 
.A(n_1782),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1833),
.Y(n_1837)
);

AOI221xp5_ASAP7_75t_L g1838 ( 
.A1(n_1814),
.A2(n_1771),
.B1(n_1772),
.B2(n_1777),
.C(n_1778),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1831),
.B(n_1800),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1818),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1823),
.B(n_1787),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1816),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1831),
.B(n_1757),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1814),
.A2(n_1786),
.B(n_1795),
.Y(n_1844)
);

OAI21xp33_ASAP7_75t_L g1845 ( 
.A1(n_1836),
.A2(n_1828),
.B(n_1780),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1825),
.B(n_1799),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1816),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1818),
.B(n_1719),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1818),
.B(n_1719),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1819),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1823),
.B(n_1808),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1829),
.B(n_1813),
.Y(n_1852)
);

BUFx3_ASAP7_75t_L g1853 ( 
.A(n_1813),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1836),
.B(n_1790),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1825),
.B(n_1742),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1829),
.B(n_1797),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1830),
.B(n_1807),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1833),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1833),
.Y(n_1859)
);

BUFx2_ASAP7_75t_L g1860 ( 
.A(n_1811),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1830),
.B(n_1796),
.Y(n_1861)
);

AND2x4_ASAP7_75t_SL g1862 ( 
.A(n_1818),
.B(n_1774),
.Y(n_1862)
);

AOI21xp5_ASAP7_75t_SL g1863 ( 
.A1(n_1835),
.A2(n_1783),
.B(n_1805),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1828),
.A2(n_1706),
.B1(n_1704),
.B2(n_1740),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1810),
.B(n_1740),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1829),
.B(n_1813),
.Y(n_1866)
);

NAND3xp33_ASAP7_75t_L g1867 ( 
.A(n_1827),
.B(n_1754),
.C(n_1740),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1815),
.B(n_1826),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1815),
.B(n_1760),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1818),
.B(n_1801),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1810),
.B(n_1774),
.Y(n_1871)
);

INVx1_ASAP7_75t_SL g1872 ( 
.A(n_1835),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1815),
.B(n_1774),
.Y(n_1873)
);

OR2x2_ASAP7_75t_SL g1874 ( 
.A(n_1822),
.B(n_1783),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1819),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1834),
.B(n_1766),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1822),
.B(n_1738),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1851),
.B(n_1810),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1843),
.B(n_1821),
.Y(n_1879)
);

NOR3xp33_ASAP7_75t_L g1880 ( 
.A(n_1838),
.B(n_1827),
.C(n_1834),
.Y(n_1880)
);

OAI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1839),
.A2(n_1834),
.B1(n_1704),
.B2(n_1756),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1851),
.B(n_1826),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_SL g1883 ( 
.A(n_1840),
.B(n_1785),
.Y(n_1883)
);

INVx1_ASAP7_75t_SL g1884 ( 
.A(n_1860),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1853),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1843),
.B(n_1821),
.Y(n_1886)
);

NOR2x1p5_ASAP7_75t_L g1887 ( 
.A(n_1840),
.B(n_1834),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1839),
.B(n_1855),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1855),
.B(n_1824),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1860),
.B(n_1812),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1868),
.B(n_1812),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1842),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1842),
.Y(n_1893)
);

XNOR2x1_ASAP7_75t_L g1894 ( 
.A(n_1854),
.B(n_1559),
.Y(n_1894)
);

INVxp67_ASAP7_75t_L g1895 ( 
.A(n_1870),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1853),
.Y(n_1896)
);

AND2x4_ASAP7_75t_SL g1897 ( 
.A(n_1871),
.B(n_1812),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1868),
.B(n_1812),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1847),
.Y(n_1899)
);

AND2x4_ASAP7_75t_L g1900 ( 
.A(n_1853),
.B(n_1812),
.Y(n_1900)
);

HB1xp67_ASAP7_75t_L g1901 ( 
.A(n_1852),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1847),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1877),
.B(n_1824),
.Y(n_1903)
);

INVx2_ASAP7_75t_SL g1904 ( 
.A(n_1862),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1852),
.B(n_1866),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1844),
.B(n_1820),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1850),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1866),
.B(n_1832),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1845),
.B(n_1820),
.Y(n_1909)
);

INVx1_ASAP7_75t_SL g1910 ( 
.A(n_1862),
.Y(n_1910)
);

OAI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1845),
.A2(n_1817),
.B(n_1753),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1850),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1856),
.B(n_1832),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1856),
.B(n_1832),
.Y(n_1914)
);

INVx1_ASAP7_75t_SL g1915 ( 
.A(n_1894),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1892),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1884),
.B(n_1872),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1901),
.Y(n_1918)
);

AOI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1880),
.A2(n_1861),
.B1(n_1857),
.B2(n_1864),
.Y(n_1919)
);

AOI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1894),
.A2(n_1863),
.B(n_1867),
.Y(n_1920)
);

BUFx3_ASAP7_75t_L g1921 ( 
.A(n_1885),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1892),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1893),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1888),
.B(n_1874),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1888),
.B(n_1874),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1878),
.B(n_1873),
.Y(n_1926)
);

INVx1_ASAP7_75t_SL g1927 ( 
.A(n_1897),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1878),
.B(n_1873),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1891),
.B(n_1871),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1893),
.Y(n_1930)
);

BUFx4f_ASAP7_75t_SL g1931 ( 
.A(n_1883),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1900),
.Y(n_1932)
);

INVx1_ASAP7_75t_SL g1933 ( 
.A(n_1897),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1899),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1899),
.Y(n_1935)
);

INVx2_ASAP7_75t_SL g1936 ( 
.A(n_1900),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1879),
.B(n_1846),
.Y(n_1937)
);

AND2x4_ASAP7_75t_L g1938 ( 
.A(n_1900),
.B(n_1871),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1902),
.Y(n_1939)
);

OR2x2_ASAP7_75t_L g1940 ( 
.A(n_1879),
.B(n_1846),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1886),
.B(n_1877),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1905),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1918),
.Y(n_1943)
);

OAI221xp5_ASAP7_75t_SL g1944 ( 
.A1(n_1919),
.A2(n_1895),
.B1(n_1906),
.B2(n_1863),
.C(n_1909),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1938),
.Y(n_1945)
);

OAI21xp33_ASAP7_75t_L g1946 ( 
.A1(n_1920),
.A2(n_1890),
.B(n_1911),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1921),
.B(n_1905),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1915),
.A2(n_1910),
.B1(n_1904),
.B2(n_1890),
.Y(n_1948)
);

OAI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1924),
.A2(n_1867),
.B1(n_1904),
.B2(n_1886),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1923),
.Y(n_1950)
);

AND2x4_ASAP7_75t_L g1951 ( 
.A(n_1936),
.B(n_1887),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1924),
.B(n_1885),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1923),
.Y(n_1953)
);

AND2x4_ASAP7_75t_L g1954 ( 
.A(n_1936),
.B(n_1887),
.Y(n_1954)
);

OAI31xp33_ASAP7_75t_L g1955 ( 
.A1(n_1925),
.A2(n_1881),
.A3(n_1848),
.B(n_1849),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1942),
.Y(n_1956)
);

NOR2xp33_ASAP7_75t_L g1957 ( 
.A(n_1931),
.B(n_1641),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1938),
.Y(n_1958)
);

INVxp67_ASAP7_75t_SL g1959 ( 
.A(n_1925),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_SL g1960 ( 
.A(n_1938),
.B(n_1891),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1942),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1937),
.B(n_1896),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1916),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1922),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1921),
.B(n_1896),
.Y(n_1965)
);

INVx1_ASAP7_75t_SL g1966 ( 
.A(n_1952),
.Y(n_1966)
);

INVxp67_ASAP7_75t_SL g1967 ( 
.A(n_1957),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1959),
.B(n_1932),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1945),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1948),
.B(n_1932),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1962),
.Y(n_1971)
);

NOR2x1_ASAP7_75t_L g1972 ( 
.A(n_1965),
.B(n_1943),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1958),
.B(n_1926),
.Y(n_1973)
);

INVx4_ASAP7_75t_L g1974 ( 
.A(n_1951),
.Y(n_1974)
);

INVx1_ASAP7_75t_SL g1975 ( 
.A(n_1947),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_R g1976 ( 
.A(n_1965),
.B(n_1917),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1956),
.B(n_1937),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1951),
.B(n_1926),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1955),
.B(n_1927),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_SL g1980 ( 
.A(n_1974),
.B(n_1933),
.Y(n_1980)
);

OAI22xp5_ASAP7_75t_R g1981 ( 
.A1(n_1967),
.A2(n_1961),
.B1(n_1964),
.B2(n_1963),
.Y(n_1981)
);

OAI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1970),
.A2(n_1944),
.B1(n_1946),
.B2(n_1940),
.Y(n_1982)
);

OAI21xp33_ASAP7_75t_L g1983 ( 
.A1(n_1979),
.A2(n_1960),
.B(n_1928),
.Y(n_1983)
);

O2A1O1Ixp33_ASAP7_75t_L g1984 ( 
.A1(n_1972),
.A2(n_1949),
.B(n_1955),
.C(n_1953),
.Y(n_1984)
);

AOI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1978),
.A2(n_1954),
.B1(n_1928),
.B2(n_1949),
.Y(n_1985)
);

OAI211xp5_ASAP7_75t_L g1986 ( 
.A1(n_1976),
.A2(n_1940),
.B(n_1950),
.C(n_1939),
.Y(n_1986)
);

AOI221xp5_ASAP7_75t_L g1987 ( 
.A1(n_1966),
.A2(n_1954),
.B1(n_1935),
.B2(n_1934),
.C(n_1930),
.Y(n_1987)
);

OAI21xp5_ASAP7_75t_SL g1988 ( 
.A1(n_1975),
.A2(n_1971),
.B(n_1978),
.Y(n_1988)
);

NAND4xp25_ASAP7_75t_L g1989 ( 
.A(n_1973),
.B(n_1929),
.C(n_1941),
.D(n_1898),
.Y(n_1989)
);

O2A1O1Ixp5_ASAP7_75t_L g1990 ( 
.A1(n_1974),
.A2(n_1941),
.B(n_1929),
.C(n_1898),
.Y(n_1990)
);

AOI22xp5_ASAP7_75t_L g1991 ( 
.A1(n_1980),
.A2(n_1969),
.B1(n_1968),
.B2(n_1977),
.Y(n_1991)
);

AOI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1983),
.A2(n_1908),
.B1(n_1882),
.B2(n_1865),
.Y(n_1992)
);

AOI221xp5_ASAP7_75t_SL g1993 ( 
.A1(n_1984),
.A2(n_1907),
.B1(n_1902),
.B2(n_1912),
.C(n_1908),
.Y(n_1993)
);

INVxp67_ASAP7_75t_L g1994 ( 
.A(n_1985),
.Y(n_1994)
);

A2O1A1Ixp33_ASAP7_75t_L g1995 ( 
.A1(n_1990),
.A2(n_1865),
.B(n_1912),
.C(n_1907),
.Y(n_1995)
);

NOR2x1_ASAP7_75t_L g1996 ( 
.A(n_1988),
.B(n_1865),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1986),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1996),
.B(n_1991),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1997),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1994),
.B(n_1987),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1993),
.B(n_1982),
.Y(n_2001)
);

NOR3xp33_ASAP7_75t_L g2002 ( 
.A(n_1995),
.B(n_1989),
.C(n_1981),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1992),
.B(n_1882),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1991),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1996),
.Y(n_2005)
);

INVx1_ASAP7_75t_SL g2006 ( 
.A(n_1998),
.Y(n_2006)
);

INVxp67_ASAP7_75t_SL g2007 ( 
.A(n_2005),
.Y(n_2007)
);

INVx1_ASAP7_75t_SL g2008 ( 
.A(n_2003),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_2004),
.B(n_1913),
.Y(n_2009)
);

OAI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_2000),
.A2(n_1876),
.B1(n_1903),
.B2(n_1889),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1999),
.Y(n_2011)
);

OR2x2_ASAP7_75t_L g2012 ( 
.A(n_2006),
.B(n_2001),
.Y(n_2012)
);

NAND4xp25_ASAP7_75t_L g2013 ( 
.A(n_2008),
.B(n_2002),
.C(n_1914),
.D(n_1913),
.Y(n_2013)
);

OAI21xp5_ASAP7_75t_L g2014 ( 
.A1(n_2007),
.A2(n_1903),
.B(n_1914),
.Y(n_2014)
);

NOR3xp33_ASAP7_75t_L g2015 ( 
.A(n_2013),
.B(n_2011),
.C(n_2009),
.Y(n_2015)
);

OAI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_2015),
.A2(n_2012),
.B1(n_2009),
.B2(n_2014),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_2016),
.Y(n_2017)
);

NOR2x1p5_ASAP7_75t_L g2018 ( 
.A(n_2016),
.B(n_2010),
.Y(n_2018)
);

INVx2_ASAP7_75t_SL g2019 ( 
.A(n_2018),
.Y(n_2019)
);

OAI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_2017),
.A2(n_1889),
.B1(n_1859),
.B2(n_1837),
.Y(n_2020)
);

AOI22xp33_ASAP7_75t_L g2021 ( 
.A1(n_2019),
.A2(n_1859),
.B1(n_1858),
.B2(n_1837),
.Y(n_2021)
);

CKINVDCx20_ASAP7_75t_R g2022 ( 
.A(n_2020),
.Y(n_2022)
);

OAI22xp5_ASAP7_75t_SL g2023 ( 
.A1(n_2022),
.A2(n_1865),
.B1(n_1858),
.B2(n_1871),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_2023),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_2024),
.B(n_2021),
.Y(n_2025)
);

INVxp67_ASAP7_75t_L g2026 ( 
.A(n_2025),
.Y(n_2026)
);

OA22x2_ASAP7_75t_L g2027 ( 
.A1(n_2026),
.A2(n_1869),
.B1(n_1875),
.B2(n_1841),
.Y(n_2027)
);

AOI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_2027),
.A2(n_1869),
.B1(n_1875),
.B2(n_1841),
.Y(n_2028)
);


endmodule