module fake_jpeg_1555_n_221 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_221);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_221;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_13),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_18),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_27),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_6),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_0),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_23),
.C(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_87),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_0),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_76),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_70),
.B1(n_77),
.B2(n_79),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_101),
.B1(n_84),
.B2(n_85),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_58),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_70),
.B1(n_77),
.B2(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_95),
.B(n_63),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_107),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_82),
.B1(n_83),
.B2(n_88),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_109),
.B1(n_113),
.B2(n_55),
.Y(n_129)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_97),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_111),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_82),
.B1(n_88),
.B2(n_81),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_110),
.A2(n_73),
.B1(n_69),
.B2(n_57),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_63),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_74),
.B1(n_71),
.B2(n_60),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_92),
.A2(n_71),
.B1(n_74),
.B2(n_85),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_73),
.B1(n_69),
.B2(n_57),
.Y(n_127)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_66),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_118),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_64),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_122),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_67),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_8),
.Y(n_145)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_102),
.B1(n_78),
.B2(n_75),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_126),
.B1(n_127),
.B2(n_138),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_72),
.C(n_84),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_34),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_122),
.Y(n_125)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_129),
.A2(n_37),
.B1(n_51),
.B2(n_50),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_106),
.B(n_68),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

OA22x2_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_68),
.B1(n_55),
.B2(n_24),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_134),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_1),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_140),
.B(n_144),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_112),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_142),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_8),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_145),
.B(n_15),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_149),
.Y(n_172)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_153),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_162),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_123),
.B1(n_134),
.B2(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_167),
.Y(n_176)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_136),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_163),
.B1(n_168),
.B2(n_15),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_12),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_158),
.B(n_164),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_145),
.B1(n_142),
.B2(n_132),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_124),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_14),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_169),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_133),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_161),
.A2(n_33),
.B(n_49),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_179),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_154),
.B1(n_19),
.B2(n_20),
.Y(n_196)
);

AND2x6_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_35),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_16),
.B(n_17),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_187),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_53),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_185),
.B(n_16),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_32),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_31),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_189),
.Y(n_204)
);

OAI322xp33_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_170),
.A3(n_162),
.B1(n_152),
.B2(n_148),
.C1(n_150),
.C2(n_157),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_198),
.C(n_183),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_172),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_193),
.A2(n_186),
.B(n_178),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_185),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_180),
.B1(n_187),
.B2(n_182),
.Y(n_202)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_154),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_191),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_203),
.C(n_205),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_188),
.C(n_173),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_176),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_181),
.C(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_207),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_200),
.A2(n_191),
.B(n_192),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_209),
.A2(n_210),
.B(n_204),
.Y(n_214)
);

O2A1O1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_211),
.A2(n_200),
.B(n_179),
.C(n_184),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_213),
.A2(n_214),
.B(n_195),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_212),
.B(n_208),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_42),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_217),
.A2(n_38),
.B(n_45),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_28),
.C(n_43),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_44),
.C(n_46),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_17),
.Y(n_221)
);


endmodule