module fake_jpeg_11209_n_119 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_119);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_26),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_5),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_57),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_48),
.B1(n_45),
.B2(n_8),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_1),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_3),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_5),
.Y(n_67)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_62),
.B(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_41),
.B1(n_48),
.B2(n_45),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_71),
.B1(n_74),
.B2(n_50),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_41),
.B1(n_38),
.B2(n_46),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_48),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_79),
.C(n_10),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_77),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_83),
.Y(n_91)
);

MAJx2_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_58),
.C(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_40),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_85),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_56),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_89),
.Y(n_94)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_23),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_6),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_7),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_24),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_96),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_100),
.B1(n_27),
.B2(n_30),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_9),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_98),
.B(n_101),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_99),
.A2(n_104),
.B(n_103),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_75),
.C(n_84),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_15),
.B(n_20),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_102),
.B(n_103),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_22),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_25),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_94),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_93),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_110),
.Y(n_111)
);

BUFx24_ASAP7_75t_SL g114 ( 
.A(n_112),
.Y(n_114)
);

AOI321xp33_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_108),
.A3(n_113),
.B1(n_106),
.B2(n_91),
.C(n_109),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_105),
.Y(n_116)
);

AOI21x1_ASAP7_75t_SL g117 ( 
.A1(n_116),
.A2(n_92),
.B(n_111),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_35),
.B(n_36),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_37),
.Y(n_119)
);


endmodule