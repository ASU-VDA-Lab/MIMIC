module fake_jpeg_14764_n_117 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_117);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_117;

wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx8_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx4f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_26),
.A2(n_14),
.B1(n_19),
.B2(n_18),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_29),
.A2(n_28),
.B1(n_25),
.B2(n_22),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_1),
.B(n_2),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_31),
.B1(n_13),
.B2(n_15),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_19),
.B1(n_18),
.B2(n_17),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_19),
.C(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_27),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_44),
.B1(n_49),
.B2(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_13),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_39),
.B1(n_23),
.B2(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_17),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_51),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_22),
.B1(n_23),
.B2(n_16),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_12),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_38),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_59),
.B(n_44),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_56),
.A2(n_40),
.B1(n_43),
.B2(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_16),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_60),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_42),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_71),
.B1(n_52),
.B2(n_44),
.Y(n_83)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_63),
.B(n_59),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_32),
.C(n_31),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_73),
.C(n_56),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_32),
.C(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_81),
.B(n_76),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_82),
.C(n_11),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_59),
.B(n_60),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_66),
.B1(n_42),
.B2(n_20),
.Y(n_92)
);

NOR4xp25_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_55),
.C(n_58),
.D(n_53),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_53),
.C(n_55),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_83),
.B(n_65),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_52),
.B(n_44),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_71),
.B(n_69),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_91),
.B1(n_2),
.B2(n_4),
.Y(n_98)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_93),
.C(n_11),
.Y(n_96)
);

AOI322xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_42),
.A3(n_38),
.B1(n_36),
.B2(n_11),
.C1(n_7),
.C2(n_8),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_90),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_75),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_20),
.Y(n_97)
);

AOI31xp33_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_92),
.A3(n_11),
.B(n_12),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_1),
.C(n_2),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_95),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_103),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_99),
.B(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_4),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_102),
.A2(n_97),
.B1(n_96),
.B2(n_105),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_109),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_100),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_32),
.C(n_11),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_112),
.Y(n_113)
);

AOI322xp5_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_36),
.A3(n_5),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_4),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_110),
.A2(n_107),
.B(n_7),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_114),
.B(n_5),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_SL g115 ( 
.A1(n_113),
.A2(n_5),
.A3(n_8),
.B1(n_9),
.B2(n_108),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_116),
.Y(n_117)
);


endmodule