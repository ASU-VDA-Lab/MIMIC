module real_jpeg_5430_n_32 (n_17, n_8, n_0, n_21, n_2, n_188, n_185, n_29, n_191, n_10, n_31, n_9, n_186, n_12, n_24, n_189, n_187, n_6, n_190, n_28, n_183, n_192, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_184, n_30, n_16, n_15, n_13, n_32);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_188;
input n_185;
input n_29;
input n_191;
input n_10;
input n_31;
input n_9;
input n_186;
input n_12;
input n_24;
input n_189;
input n_187;
input n_6;
input n_190;
input n_28;
input n_183;
input n_192;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_184;
input n_30;
input n_16;
input n_15;
input n_13;

output n_32;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_56;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_0),
.Y(n_154)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_1),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_1),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_2),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_2),
.B(n_164),
.Y(n_172)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_3),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_4),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_4),
.B(n_167),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_5),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_5),
.B(n_126),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_6),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_7),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_7),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_7),
.B(n_53),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_7),
.A2(n_50),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_8),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_10),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_10),
.B(n_78),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_11),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_13),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_14),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_15),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_15),
.B(n_88),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_16),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_17),
.Y(n_151)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_18),
.Y(n_110)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_19),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_20),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_20),
.B(n_73),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_21),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_21),
.B(n_150),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_22),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_22),
.B(n_91),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_23),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_24),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_24),
.B(n_140),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_25),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_25),
.B(n_113),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_26),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_26),
.B(n_70),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_27),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_28),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_28),
.B(n_64),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_29),
.B(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_31),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_178),
.Y(n_32)
);

AO21x1_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_42),
.B(n_176),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_36),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_38),
.B(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_38),
.B(n_151),
.Y(n_150)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_41),
.Y(n_147)
);

AO21x1_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_51),
.B(n_175),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_50),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_44),
.B(n_50),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_46),
.B(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_49),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_49),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_49),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_50),
.B(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_59),
.B(n_174),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_55),
.B(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_55),
.B(n_165),
.Y(n_164)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_89),
.Y(n_88)
);

BUFx8_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_162),
.B(n_171),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_142),
.B(n_156),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_83),
.B(n_130),
.C(n_139),
.Y(n_61)
);

NOR4xp25_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_69),
.C(n_72),
.D(n_77),
.Y(n_62)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_72),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21x1_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_125),
.B(n_129),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_120),
.B(n_124),
.Y(n_84)
);

AO221x1_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_95),
.B1(n_117),
.B2(n_118),
.C(n_119),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_141),
.Y(n_140)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_101),
.B(n_116),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_100),
.Y(n_116)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_112),
.B(n_115),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_106),
.B(n_111),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_110),
.Y(n_111)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_123),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B(n_136),
.C(n_137),
.D(n_138),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_148),
.C(n_152),
.Y(n_142)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_152),
.B(n_157),
.C(n_160),
.D(n_161),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_145),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_155),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_183),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_184),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_185),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_186),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_187),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_188),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_189),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_190),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_191),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_192),
.Y(n_127)
);


endmodule