module fake_aes_9800_n_635 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_635);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_635;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g74 ( .A(n_57), .Y(n_74) );
CKINVDCx5p33_ASAP7_75t_R g75 ( .A(n_5), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_6), .Y(n_76) );
CKINVDCx20_ASAP7_75t_R g77 ( .A(n_62), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_63), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_36), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_27), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_9), .Y(n_81) );
BUFx8_ASAP7_75t_SL g82 ( .A(n_18), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_38), .Y(n_83) );
INVxp33_ASAP7_75t_SL g84 ( .A(n_16), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_6), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_40), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_49), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_70), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_58), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_32), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_41), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_5), .Y(n_92) );
INVxp67_ASAP7_75t_L g93 ( .A(n_19), .Y(n_93) );
INVx1_ASAP7_75t_SL g94 ( .A(n_56), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_67), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_26), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_71), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_69), .Y(n_98) );
INVxp33_ASAP7_75t_SL g99 ( .A(n_8), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_48), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_43), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_16), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_3), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_0), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_54), .Y(n_105) );
CKINVDCx14_ASAP7_75t_R g106 ( .A(n_34), .Y(n_106) );
INVx2_ASAP7_75t_SL g107 ( .A(n_39), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_25), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_33), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_29), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_20), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_35), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_50), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_7), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_42), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_13), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_68), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_75), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_82), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_87), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_75), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_118), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_86), .Y(n_124) );
NOR2xp33_ASAP7_75t_SL g125 ( .A(n_78), .B(n_73), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_87), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_102), .Y(n_127) );
BUFx3_ASAP7_75t_L g128 ( .A(n_107), .Y(n_128) );
AND2x2_ASAP7_75t_SL g129 ( .A(n_108), .B(n_28), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_88), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_88), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_81), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_86), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_101), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_101), .Y(n_135) );
NAND2xp33_ASAP7_75t_R g136 ( .A(n_78), .B(n_24), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_96), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_96), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_118), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_106), .B(n_85), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_74), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_90), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_91), .Y(n_143) );
AND2x6_ASAP7_75t_L g144 ( .A(n_95), .B(n_30), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_107), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_98), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_85), .B(n_0), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_117), .B(n_1), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_117), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_102), .B(n_1), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_100), .Y(n_151) );
OAI21x1_ASAP7_75t_L g152 ( .A1(n_105), .A2(n_31), .B(n_66), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_109), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_77), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_80), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_111), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_113), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_147), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_135), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_147), .Y(n_160) );
BUFx6f_ASAP7_75t_SL g161 ( .A(n_129), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_154), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_135), .Y(n_163) );
INVx2_ASAP7_75t_SL g164 ( .A(n_140), .Y(n_164) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_152), .A2(n_116), .B(n_97), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_140), .B(n_79), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_128), .B(n_115), .Y(n_167) );
INVx5_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_155), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_119), .B(n_112), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_128), .B(n_76), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_147), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_129), .B(n_79), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_135), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_119), .B(n_83), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_135), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_135), .Y(n_177) );
INVx5_ASAP7_75t_L g178 ( .A(n_144), .Y(n_178) );
OR2x2_ASAP7_75t_L g179 ( .A(n_127), .B(n_114), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_135), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_147), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_149), .Y(n_182) );
INVx2_ASAP7_75t_SL g183 ( .A(n_128), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_151), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_141), .B(n_93), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_149), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_149), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_149), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_152), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_145), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_152), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_127), .B(n_112), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_151), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_145), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_151), .Y(n_195) );
AND2x6_ASAP7_75t_L g196 ( .A(n_123), .B(n_104), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_145), .Y(n_197) );
NOR2x1p5_ASAP7_75t_L g198 ( .A(n_120), .B(n_103), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_123), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_121), .B(n_92), .Y(n_200) );
INVx8_ASAP7_75t_L g201 ( .A(n_144), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_122), .B(n_89), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_151), .Y(n_203) );
INVx4_ASAP7_75t_L g204 ( .A(n_144), .Y(n_204) );
OR2x2_ASAP7_75t_L g205 ( .A(n_150), .B(n_83), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g206 ( .A(n_132), .Y(n_206) );
INVx4_ASAP7_75t_L g207 ( .A(n_144), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_141), .B(n_89), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_151), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_142), .B(n_99), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_166), .B(n_130), .Y(n_211) );
BUFx6f_ASAP7_75t_SL g212 ( .A(n_167), .Y(n_212) );
INVxp67_ASAP7_75t_SL g213 ( .A(n_158), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_204), .Y(n_214) );
BUFx8_ASAP7_75t_L g215 ( .A(n_161), .Y(n_215) );
OR2x2_ASAP7_75t_L g216 ( .A(n_179), .B(n_150), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_166), .B(n_130), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_161), .A2(n_129), .B1(n_110), .B2(n_99), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_208), .B(n_137), .Y(n_219) );
INVx2_ASAP7_75t_SL g220 ( .A(n_205), .Y(n_220) );
NOR3xp33_ASAP7_75t_SL g221 ( .A(n_173), .B(n_136), .C(n_148), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_164), .B(n_137), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_187), .Y(n_223) );
INVx5_ASAP7_75t_L g224 ( .A(n_196), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_164), .B(n_157), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_187), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_187), .Y(n_227) );
BUFx2_ASAP7_75t_L g228 ( .A(n_192), .Y(n_228) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_192), .Y(n_229) );
BUFx2_ASAP7_75t_L g230 ( .A(n_205), .Y(n_230) );
BUFx2_ASAP7_75t_L g231 ( .A(n_202), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_167), .B(n_131), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_167), .B(n_131), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_190), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_194), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_202), .Y(n_236) );
CKINVDCx11_ASAP7_75t_R g237 ( .A(n_206), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_161), .A2(n_121), .B1(n_126), .B2(n_139), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_171), .B(n_139), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_181), .Y(n_240) );
BUFx3_ASAP7_75t_L g241 ( .A(n_196), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_160), .A2(n_126), .B(n_157), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_197), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_171), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_171), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_200), .B(n_156), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_182), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_186), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_204), .B(n_207), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_210), .B(n_156), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_200), .B(n_153), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_170), .B(n_153), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_188), .Y(n_253) );
INVx1_ASAP7_75t_SL g254 ( .A(n_175), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_200), .B(n_185), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_179), .B(n_142), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_172), .B(n_143), .Y(n_257) );
INVx2_ASAP7_75t_SL g258 ( .A(n_198), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_204), .B(n_125), .Y(n_259) );
INVx4_ASAP7_75t_L g260 ( .A(n_196), .Y(n_260) );
AOI22xp33_ASAP7_75t_SL g261 ( .A1(n_162), .A2(n_84), .B1(n_125), .B2(n_148), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_199), .Y(n_262) );
NAND2x1_ASAP7_75t_L g263 ( .A(n_196), .B(n_144), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_181), .B(n_143), .Y(n_264) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_196), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_181), .B(n_146), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_260), .B(n_183), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_224), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_249), .A2(n_201), .B(n_207), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_244), .Y(n_270) );
BUFx8_ASAP7_75t_L g271 ( .A(n_212), .Y(n_271) );
AOI222xp33_ASAP7_75t_L g272 ( .A1(n_256), .A2(n_162), .B1(n_169), .B2(n_84), .C1(n_146), .C2(n_138), .Y(n_272) );
NAND2x1p5_ASAP7_75t_L g273 ( .A(n_260), .B(n_207), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_240), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_240), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_247), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_245), .Y(n_277) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_214), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_252), .B(n_196), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_252), .B(n_183), .Y(n_280) );
INVx4_ASAP7_75t_L g281 ( .A(n_224), .Y(n_281) );
INVx2_ASAP7_75t_SL g282 ( .A(n_224), .Y(n_282) );
NOR2x1_ASAP7_75t_R g283 ( .A(n_237), .B(n_169), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_214), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_254), .B(n_201), .Y(n_285) );
INVx6_ASAP7_75t_L g286 ( .A(n_224), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_220), .A2(n_201), .B1(n_144), .B2(n_191), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_225), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_230), .Y(n_289) );
OAI21xp5_ASAP7_75t_L g290 ( .A1(n_242), .A2(n_168), .B(n_178), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_229), .B(n_123), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_248), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_214), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_250), .B(n_201), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_225), .Y(n_295) );
BUFx8_ASAP7_75t_SL g296 ( .A(n_212), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_234), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_241), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_250), .B(n_123), .Y(n_299) );
INVx3_ASAP7_75t_SL g300 ( .A(n_216), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_253), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_211), .B(n_217), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_262), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_214), .Y(n_304) );
BUFx2_ASAP7_75t_L g305 ( .A(n_265), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_229), .B(n_138), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_228), .A2(n_144), .B1(n_189), .B2(n_191), .Y(n_307) );
AO32x1_ASAP7_75t_L g308 ( .A1(n_218), .A2(n_124), .A3(n_133), .B1(n_134), .B2(n_138), .Y(n_308) );
INVx3_ASAP7_75t_L g309 ( .A(n_263), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_249), .A2(n_168), .B(n_178), .Y(n_310) );
OAI21x1_ASAP7_75t_L g311 ( .A1(n_307), .A2(n_259), .B(n_238), .Y(n_311) );
INVx8_ASAP7_75t_L g312 ( .A(n_296), .Y(n_312) );
OAI21x1_ASAP7_75t_L g313 ( .A1(n_290), .A2(n_259), .B(n_238), .Y(n_313) );
OAI21xp33_ASAP7_75t_SL g314 ( .A1(n_280), .A2(n_213), .B(n_264), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_276), .Y(n_315) );
AO31x2_ASAP7_75t_L g316 ( .A1(n_276), .A2(n_134), .A3(n_133), .B(n_124), .Y(n_316) );
AOI21xp33_ASAP7_75t_SL g317 ( .A1(n_300), .A2(n_258), .B(n_236), .Y(n_317) );
OAI21x1_ASAP7_75t_L g318 ( .A1(n_309), .A2(n_219), .B(n_233), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_292), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_278), .Y(n_320) );
NOR2x1_ASAP7_75t_SL g321 ( .A(n_281), .B(n_235), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_300), .A2(n_231), .B1(n_215), .B2(n_261), .Y(n_322) );
AOI21x1_ASAP7_75t_L g323 ( .A1(n_292), .A2(n_193), .B(n_184), .Y(n_323) );
BUFx12f_ASAP7_75t_L g324 ( .A(n_271), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_272), .A2(n_213), .B1(n_264), .B2(n_257), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_303), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_271), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_281), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_302), .A2(n_255), .B(n_222), .C(n_251), .Y(n_329) );
CKINVDCx11_ASAP7_75t_R g330 ( .A(n_283), .Y(n_330) );
OAI21x1_ASAP7_75t_L g331 ( .A1(n_309), .A2(n_232), .B(n_239), .Y(n_331) );
INVx1_ASAP7_75t_SL g332 ( .A(n_289), .Y(n_332) );
CKINVDCx11_ASAP7_75t_R g333 ( .A(n_289), .Y(n_333) );
INVx1_ASAP7_75t_SL g334 ( .A(n_296), .Y(n_334) );
OR2x6_ASAP7_75t_L g335 ( .A(n_305), .B(n_246), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_303), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_301), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_271), .Y(n_338) );
AO21x2_ASAP7_75t_L g339 ( .A1(n_287), .A2(n_165), .B(n_221), .Y(n_339) );
OAI221xp5_ASAP7_75t_L g340 ( .A1(n_325), .A2(n_288), .B1(n_295), .B2(n_299), .C(n_221), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_337), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_315), .Y(n_342) );
OA21x2_ASAP7_75t_L g343 ( .A1(n_313), .A2(n_318), .B(n_311), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_325), .A2(n_215), .B1(n_306), .B2(n_291), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g345 ( .A1(n_329), .A2(n_291), .B1(n_306), .B2(n_257), .C(n_270), .Y(n_345) );
AOI222xp33_ASAP7_75t_L g346 ( .A1(n_322), .A2(n_277), .B1(n_266), .B2(n_243), .C1(n_146), .C2(n_279), .Y(n_346) );
AO21x1_ASAP7_75t_L g347 ( .A1(n_318), .A2(n_308), .B(n_297), .Y(n_347) );
OAI211xp5_ASAP7_75t_L g348 ( .A1(n_317), .A2(n_266), .B(n_133), .C(n_134), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_315), .B(n_297), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g350 ( .A1(n_317), .A2(n_124), .B1(n_151), .B2(n_227), .C(n_226), .Y(n_350) );
OAI221xp5_ASAP7_75t_L g351 ( .A1(n_314), .A2(n_294), .B1(n_285), .B2(n_275), .C(n_274), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_319), .B(n_274), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_314), .A2(n_308), .B(n_310), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_319), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g355 ( .A1(n_332), .A2(n_223), .B1(n_275), .B2(n_309), .C(n_191), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_326), .Y(n_356) );
OA21x2_ASAP7_75t_L g357 ( .A1(n_313), .A2(n_193), .B(n_184), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g358 ( .A1(n_337), .A2(n_305), .B1(n_265), .B2(n_304), .C(n_298), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_335), .A2(n_267), .B1(n_273), .B2(n_293), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_326), .Y(n_360) );
BUFx6f_ASAP7_75t_SL g361 ( .A(n_327), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_333), .A2(n_267), .B1(n_304), .B2(n_298), .Y(n_362) );
A2O1A1Ixp33_ASAP7_75t_L g363 ( .A1(n_336), .A2(n_267), .B(n_304), .C(n_298), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_336), .Y(n_364) );
INVxp67_ASAP7_75t_L g365 ( .A(n_361), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_349), .B(n_316), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_360), .B(n_335), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_342), .Y(n_368) );
AOI21xp5_ASAP7_75t_SL g369 ( .A1(n_359), .A2(n_321), .B(n_335), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_360), .B(n_321), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_342), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_349), .B(n_316), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_361), .B(n_338), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_354), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_361), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_357), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_354), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_356), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_352), .B(n_316), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_341), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_356), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_364), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_352), .B(n_316), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_364), .B(n_316), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_363), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_344), .B(n_335), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_357), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_340), .B(n_335), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_345), .B(n_331), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_353), .B(n_320), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_358), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_343), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_357), .Y(n_393) );
AND2x4_ASAP7_75t_L g394 ( .A(n_362), .B(n_320), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_343), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_347), .Y(n_396) );
AO31x2_ASAP7_75t_L g397 ( .A1(n_347), .A2(n_308), .A3(n_339), .B(n_177), .Y(n_397) );
OAI31xp33_ASAP7_75t_L g398 ( .A1(n_386), .A2(n_348), .A3(n_327), .B(n_351), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_368), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_366), .B(n_343), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_368), .Y(n_401) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_380), .A2(n_350), .B1(n_334), .B2(n_312), .C(n_94), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_370), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_366), .B(n_339), .Y(n_404) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_391), .A2(n_346), .B1(n_355), .B2(n_328), .C(n_282), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_371), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_388), .A2(n_328), .B1(n_282), .B2(n_191), .C(n_189), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_396), .A2(n_312), .B1(n_339), .B2(n_189), .C(n_191), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_371), .B(n_331), .Y(n_409) );
AOI322xp5_ASAP7_75t_L g410 ( .A1(n_375), .A2(n_324), .A3(n_312), .B1(n_330), .B2(n_7), .C1(n_8), .C2(n_9), .Y(n_410) );
OR2x6_ASAP7_75t_L g411 ( .A(n_369), .B(n_370), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_372), .B(n_165), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_386), .A2(n_324), .B1(n_328), .B2(n_312), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_370), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_370), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_395), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_377), .Y(n_417) );
OA211x2_ASAP7_75t_L g418 ( .A1(n_365), .A2(n_312), .B(n_308), .C(n_4), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_395), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_390), .B(n_328), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_395), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_367), .Y(n_422) );
AND2x2_ASAP7_75t_SL g423 ( .A(n_369), .B(n_189), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_372), .B(n_165), .Y(n_424) );
AO21x2_ASAP7_75t_L g425 ( .A1(n_396), .A2(n_311), .B(n_323), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_377), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_376), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_378), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_373), .B(n_2), .Y(n_429) );
NOR2xp67_ASAP7_75t_L g430 ( .A(n_376), .B(n_323), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_378), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_388), .B(n_2), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_376), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_374), .Y(n_434) );
OAI221xp5_ASAP7_75t_SL g435 ( .A1(n_385), .A2(n_209), .B1(n_195), .B2(n_203), .C(n_177), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_379), .B(n_3), .Y(n_436) );
BUFx2_ASAP7_75t_L g437 ( .A(n_367), .Y(n_437) );
OAI322xp33_ASAP7_75t_L g438 ( .A1(n_374), .A2(n_209), .A3(n_195), .B1(n_203), .B2(n_176), .C1(n_180), .C2(n_14), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_381), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_379), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_381), .Y(n_441) );
INVxp67_ASAP7_75t_SL g442 ( .A(n_383), .Y(n_442) );
NAND3xp33_ASAP7_75t_L g443 ( .A(n_384), .B(n_159), .C(n_163), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_382), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_399), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_404), .B(n_442), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_436), .B(n_383), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_436), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_440), .Y(n_449) );
BUFx2_ASAP7_75t_L g450 ( .A(n_411), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_415), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_404), .B(n_384), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_399), .B(n_382), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_401), .B(n_389), .Y(n_454) );
OAI211xp5_ASAP7_75t_SL g455 ( .A1(n_410), .A2(n_176), .B(n_180), .C(n_387), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_401), .B(n_389), .Y(n_456) );
INVx2_ASAP7_75t_SL g457 ( .A(n_403), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_406), .Y(n_458) );
NOR2xp67_ASAP7_75t_L g459 ( .A(n_443), .B(n_387), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_406), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_417), .B(n_394), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_417), .Y(n_462) );
NOR3xp33_ASAP7_75t_SL g463 ( .A(n_432), .B(n_4), .C(n_10), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_400), .B(n_392), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_400), .B(n_392), .Y(n_465) );
NAND2xp33_ASAP7_75t_R g466 ( .A(n_429), .B(n_10), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_426), .Y(n_467) );
BUFx2_ASAP7_75t_L g468 ( .A(n_411), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_422), .B(n_390), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_412), .B(n_390), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_426), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_412), .B(n_424), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_428), .B(n_394), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_424), .B(n_390), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_428), .Y(n_475) );
INVx5_ASAP7_75t_SL g476 ( .A(n_411), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_411), .B(n_394), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_431), .B(n_394), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_439), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_411), .B(n_393), .Y(n_480) );
INVx1_ASAP7_75t_SL g481 ( .A(n_403), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_431), .B(n_393), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_444), .B(n_385), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_414), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_422), .B(n_397), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_420), .B(n_393), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_416), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_439), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_420), .B(n_434), .Y(n_489) );
NOR3xp33_ASAP7_75t_L g490 ( .A(n_402), .B(n_281), .C(n_12), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_441), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_420), .B(n_393), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_441), .B(n_397), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_420), .B(n_393), .Y(n_494) );
AND2x2_ASAP7_75t_SL g495 ( .A(n_423), .B(n_393), .Y(n_495) );
NAND3xp33_ASAP7_75t_L g496 ( .A(n_410), .B(n_159), .C(n_163), .Y(n_496) );
AND2x4_ASAP7_75t_SL g497 ( .A(n_413), .B(n_293), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_434), .B(n_397), .Y(n_498) );
AND2x6_ASAP7_75t_SL g499 ( .A(n_466), .B(n_409), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_449), .B(n_437), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_452), .B(n_414), .Y(n_501) );
NOR3xp33_ASAP7_75t_L g502 ( .A(n_496), .B(n_405), .C(n_438), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_448), .B(n_437), .Y(n_503) );
NAND2x1p5_ASAP7_75t_L g504 ( .A(n_495), .B(n_423), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_445), .Y(n_505) );
INVxp67_ASAP7_75t_SL g506 ( .A(n_479), .Y(n_506) );
INVx1_ASAP7_75t_SL g507 ( .A(n_481), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_458), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_447), .B(n_444), .Y(n_509) );
INVxp67_ASAP7_75t_L g510 ( .A(n_451), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_472), .B(n_433), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_472), .B(n_433), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_460), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_452), .B(n_427), .Y(n_514) );
NAND2x1p5_ASAP7_75t_L g515 ( .A(n_495), .B(n_423), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_487), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_462), .Y(n_517) );
OAI322xp33_ASAP7_75t_L g518 ( .A1(n_464), .A2(n_407), .A3(n_427), .B1(n_421), .B2(n_416), .C1(n_419), .C2(n_11), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_487), .Y(n_519) );
OAI31xp33_ASAP7_75t_L g520 ( .A1(n_455), .A2(n_398), .A3(n_435), .B(n_419), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_446), .B(n_421), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_464), .B(n_425), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_467), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_490), .A2(n_408), .B(n_430), .C(n_418), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_471), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_483), .B(n_11), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_475), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_476), .A2(n_418), .B1(n_425), .B2(n_430), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_446), .B(n_425), .Y(n_529) );
NOR2x1_ASAP7_75t_L g530 ( .A(n_459), .B(n_12), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_470), .B(n_397), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_465), .B(n_397), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_488), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_491), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_453), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_465), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_482), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_470), .B(n_397), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_474), .B(n_13), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_482), .Y(n_540) );
NAND2x1p5_ASAP7_75t_L g541 ( .A(n_457), .B(n_293), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_469), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_454), .B(n_15), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_456), .B(n_15), .Y(n_544) );
INVx1_ASAP7_75t_SL g545 ( .A(n_457), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_474), .B(n_17), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_463), .A2(n_189), .B1(n_293), .B2(n_284), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_542), .Y(n_548) );
OAI32xp33_ASAP7_75t_L g549 ( .A1(n_507), .A2(n_469), .A3(n_485), .B1(n_484), .B2(n_473), .Y(n_549) );
INVx2_ASAP7_75t_SL g550 ( .A(n_545), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_542), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g552 ( .A(n_510), .B(n_493), .C(n_485), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_505), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_508), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_513), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_519), .Y(n_556) );
NAND2xp33_ASAP7_75t_L g557 ( .A(n_530), .B(n_484), .Y(n_557) );
AOI21xp5_ASAP7_75t_SL g558 ( .A1(n_506), .A2(n_518), .B(n_524), .Y(n_558) );
AOI221x1_ASAP7_75t_L g559 ( .A1(n_502), .A2(n_477), .B1(n_461), .B2(n_478), .C(n_480), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_502), .A2(n_477), .B1(n_468), .B2(n_450), .Y(n_560) );
OAI21xp33_ASAP7_75t_L g561 ( .A1(n_510), .A2(n_511), .B(n_512), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_536), .B(n_498), .Y(n_562) );
OAI21xp5_ASAP7_75t_L g563 ( .A1(n_524), .A2(n_450), .B(n_468), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_499), .B(n_497), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_516), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_526), .A2(n_477), .B1(n_476), .B2(n_480), .Y(n_566) );
OAI321xp33_ASAP7_75t_L g567 ( .A1(n_504), .A2(n_489), .A3(n_486), .B1(n_494), .B2(n_492), .C(n_498), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_517), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_501), .B(n_489), .Y(n_569) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_519), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g571 ( .A(n_526), .B(n_480), .C(n_494), .D(n_492), .Y(n_571) );
OAI211xp5_ASAP7_75t_L g572 ( .A1(n_547), .A2(n_486), .B(n_497), .C(n_476), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_514), .Y(n_573) );
INVx3_ASAP7_75t_L g574 ( .A(n_504), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_520), .A2(n_476), .B(n_293), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_506), .Y(n_576) );
NAND4xp75_ASAP7_75t_L g577 ( .A(n_539), .B(n_269), .C(n_22), .D(n_23), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_535), .B(n_174), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_500), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_531), .B(n_174), .Y(n_580) );
OAI22xp33_ASAP7_75t_L g581 ( .A1(n_515), .A2(n_284), .B1(n_278), .B2(n_268), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_569), .B(n_538), .Y(n_582) );
XNOR2x1_ASAP7_75t_L g583 ( .A(n_563), .B(n_515), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_571), .A2(n_532), .B1(n_546), .B2(n_529), .Y(n_584) );
AOI32xp33_ASAP7_75t_L g585 ( .A1(n_564), .A2(n_503), .A3(n_528), .B1(n_521), .B2(n_537), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g586 ( .A1(n_558), .A2(n_544), .B1(n_543), .B2(n_523), .C(n_527), .Y(n_586) );
NAND3xp33_ASAP7_75t_L g587 ( .A(n_557), .B(n_528), .C(n_534), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_548), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_573), .B(n_540), .Y(n_589) );
AND2x4_ASAP7_75t_SL g590 ( .A(n_550), .B(n_533), .Y(n_590) );
NOR3xp33_ASAP7_75t_L g591 ( .A(n_575), .B(n_525), .C(n_522), .Y(n_591) );
AOI221x1_ASAP7_75t_SL g592 ( .A1(n_564), .A2(n_516), .B1(n_509), .B2(n_541), .C(n_45), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_551), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_560), .A2(n_566), .B1(n_579), .B2(n_561), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_553), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_576), .B(n_541), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_566), .A2(n_159), .B1(n_163), .B2(n_174), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_554), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_555), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_549), .A2(n_174), .B1(n_163), .B2(n_159), .C(n_284), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_552), .B(n_174), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_574), .A2(n_159), .B1(n_163), .B2(n_278), .Y(n_602) );
AOI21xp33_ASAP7_75t_SL g603 ( .A1(n_583), .A2(n_574), .B(n_581), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_586), .A2(n_572), .B1(n_562), .B2(n_568), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_584), .B(n_570), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_590), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_585), .B(n_567), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_594), .B(n_570), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_587), .A2(n_559), .B(n_581), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_588), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_587), .A2(n_580), .B1(n_556), .B2(n_565), .Y(n_611) );
INVxp67_ASAP7_75t_L g612 ( .A(n_595), .Y(n_612) );
NOR2xp33_ASAP7_75t_R g613 ( .A(n_596), .B(n_592), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_591), .A2(n_556), .B1(n_565), .B2(n_577), .Y(n_614) );
NOR3xp33_ASAP7_75t_L g615 ( .A(n_601), .B(n_578), .C(n_268), .Y(n_615) );
AOI211x1_ASAP7_75t_SL g616 ( .A1(n_607), .A2(n_592), .B(n_600), .C(n_593), .Y(n_616) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_603), .A2(n_599), .B1(n_598), .B2(n_589), .C(n_582), .Y(n_617) );
AOI211xp5_ASAP7_75t_L g618 ( .A1(n_609), .A2(n_597), .B(n_602), .C(n_284), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_612), .B(n_21), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_608), .A2(n_284), .B1(n_278), .B2(n_46), .C(n_47), .Y(n_620) );
NAND5xp2_ASAP7_75t_SL g621 ( .A(n_611), .B(n_37), .C(n_44), .D(n_51), .E(n_52), .Y(n_621) );
NAND4xp25_ASAP7_75t_L g622 ( .A(n_614), .B(n_53), .C(n_55), .D(n_59), .Y(n_622) );
AND2x4_ASAP7_75t_L g623 ( .A(n_619), .B(n_606), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_617), .A2(n_605), .B(n_604), .Y(n_624) );
OAI22xp33_ASAP7_75t_SL g625 ( .A1(n_616), .A2(n_610), .B1(n_613), .B2(n_615), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_618), .Y(n_626) );
OR4x2_ASAP7_75t_L g627 ( .A(n_625), .B(n_622), .C(n_621), .D(n_620), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_626), .B(n_278), .C(n_168), .Y(n_628) );
XNOR2xp5_ASAP7_75t_L g629 ( .A(n_627), .B(n_623), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_628), .A2(n_624), .B1(n_286), .B2(n_168), .Y(n_630) );
XNOR2xp5_ASAP7_75t_L g631 ( .A(n_629), .B(n_60), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_631), .B(n_630), .Y(n_632) );
AOI222xp33_ASAP7_75t_L g633 ( .A1(n_632), .A2(n_286), .B1(n_168), .B2(n_178), .C1(n_72), .C2(n_64), .Y(n_633) );
AOI22x1_ASAP7_75t_L g634 ( .A1(n_633), .A2(n_273), .B1(n_65), .B2(n_61), .Y(n_634) );
OAI321xp33_ASAP7_75t_L g635 ( .A1(n_634), .A2(n_178), .A3(n_273), .B1(n_286), .B2(n_632), .C(n_630), .Y(n_635) );
endmodule