module real_aes_1587_n_239 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_239);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_239;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_503;
wire n_635;
wire n_287;
wire n_357;
wire n_673;
wire n_386;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_527;
wire n_434;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_653;
wire n_365;
wire n_290;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_0), .A2(n_85), .B1(n_330), .B2(n_569), .Y(n_568) );
XNOR2x1_ASAP7_75t_L g495 ( .A(n_1), .B(n_496), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_2), .A2(n_214), .B1(n_354), .B2(n_355), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_3), .A2(n_183), .B1(n_286), .B2(n_291), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_4), .A2(n_131), .B1(n_499), .B2(n_500), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_5), .A2(n_66), .B1(n_541), .B2(n_624), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_6), .A2(n_128), .B1(n_354), .B2(n_355), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_7), .A2(n_194), .B1(n_697), .B2(n_698), .Y(n_696) );
AO22x2_ASAP7_75t_L g266 ( .A1(n_8), .A2(n_171), .B1(n_267), .B2(n_268), .Y(n_266) );
INVx1_ASAP7_75t_L g671 ( .A(n_8), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_9), .A2(n_215), .B1(n_286), .B2(n_347), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_10), .A2(n_58), .B1(n_592), .B2(n_593), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_11), .A2(n_59), .B1(n_618), .B2(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_12), .A2(n_155), .B1(n_384), .B2(n_414), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g610 ( .A1(n_13), .A2(n_187), .B1(n_263), .B2(n_562), .Y(n_610) );
AO22x2_ASAP7_75t_L g270 ( .A1(n_14), .A2(n_48), .B1(n_267), .B2(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_14), .B(n_670), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_15), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_16), .A2(n_65), .B1(n_349), .B2(n_396), .Y(n_478) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_17), .A2(n_159), .B1(n_503), .B2(n_556), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_18), .A2(n_127), .B1(n_263), .B2(n_280), .Y(n_466) );
AO222x2_ASAP7_75t_SL g340 ( .A1(n_19), .A2(n_35), .B1(n_136), .B2(n_341), .C1(n_342), .C2(n_343), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_20), .A2(n_170), .B1(n_429), .B2(n_430), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_21), .A2(n_63), .B1(n_359), .B2(n_384), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_22), .A2(n_236), .B1(n_294), .B2(n_296), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_23), .A2(n_141), .B1(n_361), .B2(n_362), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_24), .A2(n_132), .B1(n_346), .B2(n_347), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_25), .B(n_302), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_26), .A2(n_106), .B1(n_571), .B2(n_596), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_27), .A2(n_211), .B1(n_349), .B2(n_350), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_28), .A2(n_225), .B1(n_655), .B2(n_656), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_29), .A2(n_105), .B1(n_280), .B2(n_560), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_30), .A2(n_116), .B1(n_426), .B2(n_516), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_31), .A2(n_165), .B1(n_263), .B2(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_32), .A2(n_186), .B1(n_286), .B2(n_291), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_33), .A2(n_111), .B1(n_263), .B2(n_280), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_34), .A2(n_117), .B1(n_325), .B2(n_382), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_36), .A2(n_158), .B1(n_325), .B2(n_382), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_37), .A2(n_168), .B1(n_545), .B2(n_546), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_38), .A2(n_130), .B1(n_545), .B2(n_626), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_39), .A2(n_52), .B1(n_417), .B2(n_419), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_40), .A2(n_200), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_41), .A2(n_222), .B1(n_617), .B2(n_618), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_42), .A2(n_69), .B1(n_349), .B2(n_350), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_43), .A2(n_216), .B1(n_538), .B2(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_SL g608 ( .A1(n_44), .A2(n_238), .B1(n_435), .B2(n_558), .Y(n_608) );
AOI22xp33_ASAP7_75t_SL g590 ( .A1(n_45), .A2(n_207), .B1(n_320), .B2(n_539), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_46), .A2(n_91), .B1(n_560), .B2(n_562), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_47), .A2(n_232), .B1(n_327), .B2(n_330), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_49), .A2(n_180), .B1(n_341), .B2(n_342), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_50), .A2(n_53), .B1(n_571), .B2(n_572), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_51), .A2(n_226), .B1(n_426), .B2(n_565), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_54), .A2(n_126), .B1(n_327), .B2(n_421), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_55), .A2(n_135), .B1(n_543), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_56), .A2(n_93), .B1(n_317), .B2(n_320), .Y(n_316) );
INVx3_ASAP7_75t_L g267 ( .A(n_57), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_60), .A2(n_124), .B1(n_324), .B2(n_325), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_61), .A2(n_221), .B1(n_341), .B2(n_342), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_62), .A2(n_109), .B1(n_652), .B2(n_653), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_64), .A2(n_89), .B1(n_679), .B2(n_681), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_67), .A2(n_75), .B1(n_359), .B2(n_384), .Y(n_458) );
INVx1_ASAP7_75t_SL g275 ( .A(n_68), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_68), .B(n_108), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_70), .A2(n_94), .B1(n_291), .B2(n_346), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_71), .A2(n_112), .B1(n_505), .B2(n_506), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_72), .A2(n_237), .B1(n_418), .B2(n_513), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_73), .A2(n_151), .B1(n_502), .B2(n_503), .Y(n_501) );
INVx2_ASAP7_75t_L g246 ( .A(n_74), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_76), .A2(n_217), .B1(n_419), .B2(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_77), .B(n_374), .Y(n_373) );
XOR2x2_ASAP7_75t_L g519 ( .A(n_78), .B(n_520), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_79), .A2(n_122), .B1(n_411), .B2(n_414), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_80), .A2(n_115), .B1(n_341), .B2(n_393), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_81), .A2(n_129), .B1(n_324), .B2(n_325), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_82), .A2(n_201), .B1(n_312), .B2(n_565), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_83), .A2(n_172), .B1(n_411), .B2(n_414), .Y(n_410) );
AOI22xp33_ASAP7_75t_SL g482 ( .A1(n_84), .A2(n_162), .B1(n_354), .B2(n_355), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_86), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_87), .A2(n_99), .B1(n_542), .B2(n_644), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_88), .A2(n_208), .B1(n_294), .B2(n_435), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_90), .B(n_440), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_92), .A2(n_173), .B1(n_311), .B2(n_359), .Y(n_379) );
XNOR2x1_ASAP7_75t_SL g603 ( .A(n_95), .B(n_604), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_96), .A2(n_119), .B1(n_421), .B2(n_641), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_97), .A2(n_198), .B1(n_442), .B2(n_444), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_98), .A2(n_228), .B1(n_535), .B2(n_536), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_100), .A2(n_163), .B1(n_433), .B2(n_436), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_101), .A2(n_147), .B1(n_317), .B2(n_567), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_102), .A2(n_230), .B1(n_527), .B2(n_528), .Y(n_526) );
AOI22xp33_ASAP7_75t_SL g400 ( .A1(n_103), .A2(n_154), .B1(n_354), .B2(n_355), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_104), .A2(n_174), .B1(n_541), .B2(n_543), .Y(n_540) );
OA21x2_ASAP7_75t_L g630 ( .A1(n_107), .A2(n_631), .B(n_657), .Y(n_630) );
INVx1_ASAP7_75t_L g659 ( .A(n_107), .Y(n_659) );
AO22x2_ASAP7_75t_L g278 ( .A1(n_108), .A2(n_182), .B1(n_267), .B2(n_279), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_110), .A2(n_133), .B1(n_528), .B2(n_638), .Y(n_692) );
INVx1_ASAP7_75t_L g708 ( .A(n_113), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_114), .A2(n_220), .B1(n_435), .B2(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g634 ( .A(n_118), .B(n_635), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_120), .A2(n_235), .B1(n_309), .B2(n_312), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_121), .A2(n_193), .B1(n_311), .B2(n_359), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_123), .A2(n_229), .B1(n_423), .B2(n_425), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_125), .A2(n_140), .B1(n_286), .B2(n_347), .Y(n_376) );
INVx1_ASAP7_75t_L g276 ( .A(n_134), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_137), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_138), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_139), .B(n_374), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_142), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_143), .A2(n_164), .B1(n_296), .B2(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_144), .A2(n_218), .B1(n_421), .B2(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_145), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_146), .A2(n_196), .B1(n_523), .B2(n_524), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_148), .B(n_391), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_149), .A2(n_150), .B1(n_324), .B2(n_325), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_152), .B(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_153), .A2(n_224), .B1(n_694), .B2(n_695), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_156), .A2(n_167), .B1(n_320), .B2(n_647), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_157), .A2(n_177), .B1(n_324), .B2(n_325), .Y(n_323) );
AO22x1_ASAP7_75t_L g637 ( .A1(n_160), .A2(n_210), .B1(n_433), .B2(n_638), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_161), .A2(n_675), .B1(n_700), .B2(n_701), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_161), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_166), .A2(n_209), .B1(n_361), .B2(n_362), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_169), .A2(n_223), .B1(n_418), .B2(n_457), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_175), .A2(n_190), .B1(n_314), .B2(n_460), .Y(n_459) );
AOI22xp33_ASAP7_75t_SL g395 ( .A1(n_176), .A2(n_184), .B1(n_349), .B2(n_396), .Y(n_395) );
OA22x2_ASAP7_75t_L g259 ( .A1(n_178), .A2(n_260), .B1(n_333), .B2(n_334), .Y(n_259) );
INVx1_ASAP7_75t_L g333 ( .A(n_178), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_179), .A2(n_203), .B1(n_311), .B2(n_359), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_181), .B(n_374), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_185), .A2(n_219), .B1(n_503), .B2(n_556), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_188), .A2(n_205), .B1(n_320), .B2(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_189), .B(n_440), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_191), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g667 ( .A(n_191), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_192), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_195), .A2(n_202), .B1(n_384), .B2(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g243 ( .A(n_197), .Y(n_243) );
AND2x2_ASAP7_75t_R g705 ( .A(n_197), .B(n_667), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g239 ( .A1(n_199), .A2(n_240), .B1(n_249), .B2(n_663), .C(n_673), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_204), .A2(n_234), .B1(n_311), .B2(n_405), .Y(n_404) );
INVxp67_ASAP7_75t_L g248 ( .A(n_206), .Y(n_248) );
AOI22x1_ASAP7_75t_SL g550 ( .A1(n_212), .A2(n_551), .B1(n_552), .B2(n_573), .Y(n_550) );
INVx1_ASAP7_75t_L g573 ( .A(n_212), .Y(n_573) );
XNOR2xp5_ASAP7_75t_L g407 ( .A(n_213), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_227), .B(n_391), .Y(n_390) );
XOR2x2_ASAP7_75t_L g577 ( .A(n_231), .B(n_578), .Y(n_577) );
XNOR2xp5_ASAP7_75t_L g470 ( .A(n_233), .B(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NOR2x1_ASAP7_75t_R g241 ( .A(n_242), .B(n_244), .Y(n_241) );
OR2x2_ASAP7_75t_L g714 ( .A(n_242), .B(n_245), .Y(n_714) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_243), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_489), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AOI21xp33_ASAP7_75t_L g663 ( .A1(n_251), .A2(n_490), .B(n_664), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_467), .B1(n_487), .B2(n_488), .Y(n_251) );
INVx1_ASAP7_75t_L g488 ( .A(n_252), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B1(n_450), .B2(n_451), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AO22x2_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_366), .B1(n_448), .B2(n_449), .Y(n_254) );
INVx1_ASAP7_75t_L g448 ( .A(n_255), .Y(n_448) );
OAI22xp5_ASAP7_75t_SL g255 ( .A1(n_256), .A2(n_335), .B1(n_364), .B2(n_365), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_259), .Y(n_364) );
INVx1_ASAP7_75t_L g334 ( .A(n_260), .Y(n_334) );
NOR2x1_ASAP7_75t_L g260 ( .A(n_261), .B(n_307), .Y(n_260) );
NAND4xp25_ASAP7_75t_L g261 ( .A(n_262), .B(n_285), .C(n_293), .D(n_301), .Y(n_261) );
BUFx6f_ASAP7_75t_SL g429 ( .A(n_263), .Y(n_429) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_264), .Y(n_505) );
INVx3_ASAP7_75t_L g561 ( .A(n_264), .Y(n_561) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_272), .Y(n_264) );
AND2x2_ASAP7_75t_L g319 ( .A(n_265), .B(n_287), .Y(n_319) );
AND2x4_ASAP7_75t_L g332 ( .A(n_265), .B(n_315), .Y(n_332) );
AND2x4_ASAP7_75t_L g349 ( .A(n_265), .B(n_272), .Y(n_349) );
AND2x2_ASAP7_75t_SL g354 ( .A(n_265), .B(n_287), .Y(n_354) );
AND2x6_ASAP7_75t_L g359 ( .A(n_265), .B(n_315), .Y(n_359) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_269), .Y(n_265) );
INVx2_ASAP7_75t_L g290 ( .A(n_266), .Y(n_290) );
AND2x2_ASAP7_75t_L g299 ( .A(n_266), .B(n_270), .Y(n_299) );
INVx1_ASAP7_75t_L g268 ( .A(n_267), .Y(n_268) );
INVx2_ASAP7_75t_L g271 ( .A(n_267), .Y(n_271) );
OAI22x1_ASAP7_75t_L g273 ( .A1(n_267), .A2(n_274), .B1(n_275), .B2(n_276), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_267), .Y(n_274) );
INVx1_ASAP7_75t_L g279 ( .A(n_267), .Y(n_279) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_269), .Y(n_284) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g289 ( .A(n_270), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g306 ( .A(n_270), .Y(n_306) );
AND2x2_ASAP7_75t_L g295 ( .A(n_272), .B(n_289), .Y(n_295) );
AND2x2_ASAP7_75t_L g324 ( .A(n_272), .B(n_305), .Y(n_324) );
AND2x4_ASAP7_75t_L g341 ( .A(n_272), .B(n_289), .Y(n_341) );
AND2x2_ASAP7_75t_L g382 ( .A(n_272), .B(n_305), .Y(n_382) );
AND2x4_ASAP7_75t_L g413 ( .A(n_272), .B(n_305), .Y(n_413) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_277), .Y(n_272) );
AND2x2_ASAP7_75t_L g282 ( .A(n_273), .B(n_278), .Y(n_282) );
INVx2_ASAP7_75t_L g288 ( .A(n_273), .Y(n_288) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_273), .Y(n_300) );
AND2x4_ASAP7_75t_L g315 ( .A(n_277), .B(n_288), .Y(n_315) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g287 ( .A(n_278), .B(n_288), .Y(n_287) );
BUFx2_ASAP7_75t_L g322 ( .A(n_278), .Y(n_322) );
BUFx2_ASAP7_75t_SL g656 ( .A(n_280), .Y(n_656) );
BUFx6f_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g431 ( .A(n_281), .Y(n_431) );
BUFx3_ASAP7_75t_L g506 ( .A(n_281), .Y(n_506) );
BUFx4f_ASAP7_75t_L g562 ( .A(n_281), .Y(n_562) );
INVx1_ASAP7_75t_L g699 ( .A(n_281), .Y(n_699) );
AND2x4_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g291 ( .A(n_282), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g304 ( .A(n_282), .B(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_L g343 ( .A(n_282), .B(n_305), .Y(n_343) );
AND2x2_ASAP7_75t_L g347 ( .A(n_282), .B(n_292), .Y(n_347) );
AND2x2_ASAP7_75t_L g350 ( .A(n_282), .B(n_283), .Y(n_350) );
AND2x2_ASAP7_75t_L g396 ( .A(n_282), .B(n_283), .Y(n_396) );
AND2x4_ASAP7_75t_L g446 ( .A(n_282), .B(n_292), .Y(n_446) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
AND2x6_ASAP7_75t_L g311 ( .A(n_287), .B(n_305), .Y(n_311) );
AND2x2_ASAP7_75t_L g346 ( .A(n_287), .B(n_289), .Y(n_346) );
AND2x2_ASAP7_75t_L g424 ( .A(n_287), .B(n_305), .Y(n_424) );
AND2x4_ASAP7_75t_L g443 ( .A(n_287), .B(n_289), .Y(n_443) );
AND2x4_ASAP7_75t_L g314 ( .A(n_289), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g362 ( .A(n_289), .B(n_315), .Y(n_362) );
INVxp67_ASAP7_75t_L g292 ( .A(n_290), .Y(n_292) );
AND2x4_ASAP7_75t_L g305 ( .A(n_290), .B(n_306), .Y(n_305) );
BUFx6f_ASAP7_75t_SL g527 ( .A(n_294), .Y(n_527) );
BUFx3_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g438 ( .A(n_295), .Y(n_438) );
BUFx5_ASAP7_75t_L g558 ( .A(n_295), .Y(n_558) );
BUFx3_ASAP7_75t_L g584 ( .A(n_295), .Y(n_584) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g500 ( .A(n_297), .Y(n_500) );
INVx3_ASAP7_75t_L g529 ( .A(n_297), .Y(n_529) );
INVx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx12f_ASAP7_75t_L g435 ( .A(n_298), .Y(n_435) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AND2x4_ASAP7_75t_L g321 ( .A(n_299), .B(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g325 ( .A(n_299), .B(n_315), .Y(n_325) );
AND2x2_ASAP7_75t_SL g342 ( .A(n_299), .B(n_300), .Y(n_342) );
AND2x4_ASAP7_75t_L g355 ( .A(n_299), .B(n_322), .Y(n_355) );
AND2x2_ASAP7_75t_SL g393 ( .A(n_299), .B(n_300), .Y(n_393) );
AND2x4_ASAP7_75t_L g415 ( .A(n_299), .B(n_315), .Y(n_415) );
INVx3_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
INVx4_ASAP7_75t_SL g374 ( .A(n_303), .Y(n_374) );
INVx4_ASAP7_75t_SL g391 ( .A(n_303), .Y(n_391) );
INVx3_ASAP7_75t_L g636 ( .A(n_303), .Y(n_636) );
BUFx2_ASAP7_75t_L g691 ( .A(n_303), .Y(n_691) );
INVx6_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x4_ASAP7_75t_L g329 ( .A(n_305), .B(n_315), .Y(n_329) );
AND2x2_ASAP7_75t_L g361 ( .A(n_305), .B(n_315), .Y(n_361) );
NAND4xp25_ASAP7_75t_L g307 ( .A(n_308), .B(n_316), .C(n_323), .D(n_326), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g460 ( .A(n_310), .Y(n_460) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g405 ( .A(n_313), .Y(n_405) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_314), .Y(n_385) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_314), .Y(n_426) );
BUFx3_ASAP7_75t_L g624 ( .A(n_314), .Y(n_624) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g539 ( .A(n_318), .Y(n_539) );
INVx2_ASAP7_75t_L g621 ( .A(n_318), .Y(n_621) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_319), .Y(n_418) );
BUFx3_ASAP7_75t_L g648 ( .A(n_319), .Y(n_648) );
BUFx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g419 ( .A(n_321), .Y(n_419) );
BUFx3_ASAP7_75t_L g457 ( .A(n_321), .Y(n_457) );
INVx5_ASAP7_75t_SL g514 ( .A(n_321), .Y(n_514) );
INVx3_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx3_ASAP7_75t_L g384 ( .A(n_328), .Y(n_384) );
INVx4_ASAP7_75t_L g542 ( .A(n_328), .Y(n_542) );
INVx2_ASAP7_75t_SL g565 ( .A(n_328), .Y(n_565) );
INVx2_ASAP7_75t_L g685 ( .A(n_328), .Y(n_685) );
INVx8_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g421 ( .A(n_331), .Y(n_421) );
INVx2_ASAP7_75t_L g546 ( .A(n_331), .Y(n_546) );
INVx2_ASAP7_75t_L g593 ( .A(n_331), .Y(n_593) );
INVx2_ASAP7_75t_SL g626 ( .A(n_331), .Y(n_626) );
INVx2_ASAP7_75t_L g681 ( .A(n_331), .Y(n_681) );
INVx8_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g365 ( .A(n_336), .Y(n_365) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
XOR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_363), .Y(n_337) );
NAND2x1_ASAP7_75t_L g338 ( .A(n_339), .B(n_351), .Y(n_338) );
NOR2x1_ASAP7_75t_L g339 ( .A(n_340), .B(n_344), .Y(n_339) );
INVx2_ASAP7_75t_SL g474 ( .A(n_343), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_348), .Y(n_344) );
NOR2x1_ASAP7_75t_L g351 ( .A(n_352), .B(n_357), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_356), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
INVx2_ASAP7_75t_L g449 ( .A(n_366), .Y(n_449) );
OA22x2_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_407), .B2(n_447), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
XNOR2x1_ASAP7_75t_L g368 ( .A(n_369), .B(n_386), .Y(n_368) );
XNOR2x1_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
NOR2x1_ASAP7_75t_L g371 ( .A(n_372), .B(n_378), .Y(n_371) );
NAND4xp25_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .C(n_376), .D(n_377), .Y(n_372) );
INVx1_ASAP7_75t_SL g581 ( .A(n_374), .Y(n_581) );
NAND4xp25_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .C(n_381), .D(n_383), .Y(n_378) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_385), .Y(n_543) );
INVx2_ASAP7_75t_L g645 ( .A(n_385), .Y(n_645) );
XOR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_406), .Y(n_386) );
NAND2x1_ASAP7_75t_L g387 ( .A(n_388), .B(n_398), .Y(n_387) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_389), .B(n_394), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
BUFx2_ASAP7_75t_L g440 ( .A(n_391), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_397), .Y(n_394) );
NOR2x1_ASAP7_75t_L g398 ( .A(n_399), .B(n_402), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx2_ASAP7_75t_SL g447 ( .A(n_407), .Y(n_447) );
NOR2xp67_ASAP7_75t_L g408 ( .A(n_409), .B(n_427), .Y(n_408) );
NAND4xp25_ASAP7_75t_L g409 ( .A(n_410), .B(n_416), .C(n_420), .D(n_422), .Y(n_409) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx3_ASAP7_75t_L g516 ( .A(n_412), .Y(n_516) );
INVx2_ASAP7_75t_L g535 ( .A(n_412), .Y(n_535) );
INVx2_ASAP7_75t_L g617 ( .A(n_412), .Y(n_617) );
INVx1_ASAP7_75t_SL g687 ( .A(n_412), .Y(n_687) );
INVx6_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx3_ASAP7_75t_L g571 ( .A(n_413), .Y(n_571) );
BUFx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx2_ASAP7_75t_SL g536 ( .A(n_415), .Y(n_536) );
BUFx3_ASAP7_75t_L g572 ( .A(n_415), .Y(n_572) );
INVx2_ASAP7_75t_L g597 ( .A(n_415), .Y(n_597) );
BUFx2_ASAP7_75t_SL g618 ( .A(n_415), .Y(n_618) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx3_ASAP7_75t_L g511 ( .A(n_424), .Y(n_511) );
BUFx2_ASAP7_75t_L g569 ( .A(n_424), .Y(n_569) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NAND4xp25_ASAP7_75t_L g427 ( .A(n_428), .B(n_432), .C(n_439), .D(n_441), .Y(n_427) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g532 ( .A(n_431), .Y(n_532) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g499 ( .A(n_438), .Y(n_499) );
BUFx2_ASAP7_75t_L g523 ( .A(n_442), .Y(n_523) );
BUFx4f_ASAP7_75t_SL g612 ( .A(n_442), .Y(n_612) );
BUFx2_ASAP7_75t_L g694 ( .A(n_442), .Y(n_694) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx3_ASAP7_75t_L g502 ( .A(n_443), .Y(n_502) );
BUFx2_ASAP7_75t_L g556 ( .A(n_443), .Y(n_556) );
BUFx2_ASAP7_75t_L g652 ( .A(n_443), .Y(n_652) );
INVx2_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g503 ( .A(n_445), .Y(n_503) );
INVx2_ASAP7_75t_L g524 ( .A(n_445), .Y(n_524) );
INVx2_ASAP7_75t_L g613 ( .A(n_445), .Y(n_613) );
INVx2_ASAP7_75t_SL g653 ( .A(n_445), .Y(n_653) );
INVx2_ASAP7_75t_L g695 ( .A(n_445), .Y(n_695) );
INVx6_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
XNOR2x1_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_462), .Y(n_454) );
NAND4xp25_ASAP7_75t_L g455 ( .A(n_456), .B(n_458), .C(n_459), .D(n_461), .Y(n_455) );
NAND4xp25_ASAP7_75t_SL g462 ( .A(n_463), .B(n_464), .C(n_465), .D(n_466), .Y(n_462) );
INVx1_ASAP7_75t_L g487 ( .A(n_467), .Y(n_487) );
INVx1_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_472), .B(n_480), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_477), .Y(n_472) );
OAI21xp5_ASAP7_75t_SL g473 ( .A1(n_474), .A2(n_475), .B(n_476), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_484), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
XNOR2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_601), .Y(n_490) );
OAI22xp5_ASAP7_75t_SL g491 ( .A1(n_492), .A2(n_547), .B1(n_548), .B2(n_600), .Y(n_491) );
INVx1_ASAP7_75t_L g600 ( .A(n_492), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B1(n_518), .B2(n_519), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
OR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_508), .Y(n_496) );
NAND4xp25_ASAP7_75t_L g497 ( .A(n_498), .B(n_501), .C(n_504), .D(n_507), .Y(n_497) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_505), .Y(n_655) );
NAND4xp25_ASAP7_75t_L g508 ( .A(n_509), .B(n_512), .C(n_515), .D(n_517), .Y(n_508) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_SL g545 ( .A(n_511), .Y(n_545) );
INVx2_ASAP7_75t_L g592 ( .A(n_511), .Y(n_592) );
INVx2_ASAP7_75t_L g642 ( .A(n_511), .Y(n_642) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g567 ( .A(n_514), .Y(n_567) );
INVx2_ASAP7_75t_L g683 ( .A(n_514), .Y(n_683) );
INVx5_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NOR2x1_ASAP7_75t_L g520 ( .A(n_521), .B(n_533), .Y(n_520) );
NAND4xp25_ASAP7_75t_L g521 ( .A(n_522), .B(n_525), .C(n_526), .D(n_530), .Y(n_521) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND4xp25_ASAP7_75t_L g533 ( .A(n_534), .B(n_537), .C(n_540), .D(n_544), .Y(n_533) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_574), .B1(n_575), .B2(n_599), .Y(n_548) );
INVx1_ASAP7_75t_L g599 ( .A(n_549), .Y(n_599) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_563), .Y(n_552) );
NAND4xp25_ASAP7_75t_SL g553 ( .A(n_554), .B(n_555), .C(n_557), .D(n_559), .Y(n_553) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx4_ASAP7_75t_L g697 ( .A(n_561), .Y(n_697) );
NAND4xp25_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .C(n_568), .D(n_570), .Y(n_563) );
INVx2_ASAP7_75t_L g680 ( .A(n_569), .Y(n_680) );
INVx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2x1_ASAP7_75t_L g578 ( .A(n_579), .B(n_588), .Y(n_578) );
NOR2x1_ASAP7_75t_L g579 ( .A(n_580), .B(n_585), .Y(n_579) );
OAI21xp5_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_582), .B(n_583), .Y(n_580) );
OAI21xp33_ASAP7_75t_L g606 ( .A1(n_581), .A2(n_607), .B(n_608), .Y(n_606) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_584), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
NOR2x1_ASAP7_75t_L g588 ( .A(n_589), .B(n_594), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_598), .Y(n_594) );
INVx2_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_627), .B1(n_660), .B2(n_661), .Y(n_601) );
INVx1_ASAP7_75t_L g660 ( .A(n_602), .Y(n_660) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_614), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_609), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_622), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_619), .Y(n_615) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g662 ( .A(n_630), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_631), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_650), .Y(n_632) );
NOR3xp33_ASAP7_75t_SL g633 ( .A(n_634), .B(n_637), .C(n_639), .Y(n_633) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND4xp25_ASAP7_75t_L g639 ( .A(n_640), .B(n_643), .C(n_646), .D(n_649), .Y(n_639) );
BUFx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_654), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_666), .B(n_669), .Y(n_711) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
OAI222xp33_ASAP7_75t_R g673 ( .A1(n_674), .A2(n_702), .B1(n_706), .B2(n_708), .C1(n_709), .C2(n_712), .Y(n_673) );
CKINVDCx16_ASAP7_75t_R g701 ( .A(n_675), .Y(n_701) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
XOR2x2_ASAP7_75t_L g707 ( .A(n_676), .B(n_708), .Y(n_707) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_677), .B(n_688), .Y(n_676) );
NAND4xp25_ASAP7_75t_L g677 ( .A(n_678), .B(n_682), .C(n_684), .D(n_686), .Y(n_677) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND4xp25_ASAP7_75t_L g688 ( .A(n_689), .B(n_692), .C(n_693), .D(n_696), .Y(n_688) );
INVx2_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
CKINVDCx6p67_ASAP7_75t_R g710 ( .A(n_711), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_714), .Y(n_713) );
endmodule