module fake_jpeg_7763_n_80 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_80);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_80;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_20),
.B(n_29),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_52),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_5),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_6),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_8),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_9),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

OR2x2_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_48),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_56),
.A2(n_37),
.B1(n_46),
.B2(n_45),
.Y(n_63)
);

AO22x2_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_43),
.B1(n_11),
.B2(n_14),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_42),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_61),
.C(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_72),
.B(n_70),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_69),
.C(n_68),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_64),
.C(n_62),
.Y(n_75)
);

NOR4xp25_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_10),
.C(n_17),
.D(n_22),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_25),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_26),
.C(n_27),
.Y(n_79)
);

AOI221xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.C(n_34),
.Y(n_80)
);


endmodule