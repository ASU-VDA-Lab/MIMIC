module fake_netlist_1_7337_n_1234 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1234);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1234;
wire n_963;
wire n_1034;
wire n_949;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_271;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_265;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_677;
wire n_283;
wire n_756;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_272;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_451;
wire n_487;
wire n_748;
wire n_258;
wire n_253;
wire n_266;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_280;
wire n_395;
wire n_257;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_252;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_275;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_251;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_795;
wire n_267;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_791;
wire n_707;
wire n_603;
wire n_885;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_366;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_1024;
wire n_321;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_710;
wire n_270;
wire n_1178;
wire n_259;
wire n_546;
wire n_412;
wire n_664;
wire n_788;
wire n_403;
wire n_516;
wire n_254;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_260;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_416;
wire n_536;
wire n_956;
wire n_264;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_269;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_998;
wire n_604;
wire n_755;
wire n_848;
wire n_1031;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_255;
wire n_844;
wire n_1160;
wire n_274;
wire n_1195;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_256;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_262;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_276;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_263;
wire n_1221;
wire n_428;
wire n_794;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_261;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
INVx1_ASAP7_75t_L g251 ( .A(n_166), .Y(n_251) );
BUFx5_ASAP7_75t_L g252 ( .A(n_109), .Y(n_252) );
INVxp67_ASAP7_75t_L g253 ( .A(n_55), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_119), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_49), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_33), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_132), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_157), .Y(n_258) );
BUFx2_ASAP7_75t_L g259 ( .A(n_110), .Y(n_259) );
INVx1_ASAP7_75t_SL g260 ( .A(n_8), .Y(n_260) );
INVxp67_ASAP7_75t_SL g261 ( .A(n_142), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_160), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_231), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_67), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_148), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_177), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_45), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_117), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_221), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_181), .Y(n_270) );
CKINVDCx16_ASAP7_75t_R g271 ( .A(n_90), .Y(n_271) );
INVx4_ASAP7_75t_R g272 ( .A(n_167), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_143), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_46), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_128), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_152), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_139), .Y(n_277) );
BUFx2_ASAP7_75t_SL g278 ( .A(n_20), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_222), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_145), .Y(n_280) );
INVxp33_ASAP7_75t_SL g281 ( .A(n_53), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_201), .Y(n_282) );
INVxp67_ASAP7_75t_L g283 ( .A(n_168), .Y(n_283) );
INVxp33_ASAP7_75t_L g284 ( .A(n_112), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_213), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_144), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_215), .Y(n_287) );
CKINVDCx16_ASAP7_75t_R g288 ( .A(n_208), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_103), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_18), .Y(n_290) );
INVxp67_ASAP7_75t_SL g291 ( .A(n_133), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_210), .Y(n_292) );
CKINVDCx14_ASAP7_75t_R g293 ( .A(n_238), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_11), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_178), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_150), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_48), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_105), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_31), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_114), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_55), .Y(n_301) );
INVxp33_ASAP7_75t_L g302 ( .A(n_106), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_248), .Y(n_303) );
BUFx5_ASAP7_75t_L g304 ( .A(n_16), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_102), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_237), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_224), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_57), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_171), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_88), .Y(n_310) );
INVxp67_ASAP7_75t_SL g311 ( .A(n_37), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_7), .Y(n_312) );
INVxp67_ASAP7_75t_L g313 ( .A(n_81), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_129), .Y(n_314) );
INVxp33_ASAP7_75t_SL g315 ( .A(n_60), .Y(n_315) );
INVxp33_ASAP7_75t_L g316 ( .A(n_218), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_140), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_241), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_11), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_230), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_29), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_47), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_205), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_61), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_63), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_229), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_170), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_233), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_53), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_84), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_15), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_43), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_39), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_52), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_249), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_6), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_89), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_183), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_85), .B(n_29), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_220), .Y(n_340) );
CKINVDCx14_ASAP7_75t_R g341 ( .A(n_159), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_158), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_87), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_169), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_52), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_138), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_153), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_226), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_71), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_56), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_36), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_239), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_172), .Y(n_353) );
CKINVDCx20_ASAP7_75t_R g354 ( .A(n_111), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_19), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_163), .Y(n_356) );
INVx1_ASAP7_75t_SL g357 ( .A(n_250), .Y(n_357) );
CKINVDCx16_ASAP7_75t_R g358 ( .A(n_27), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_58), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_20), .Y(n_360) );
INVx1_ASAP7_75t_SL g361 ( .A(n_120), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_204), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_113), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_187), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_79), .B(n_58), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_41), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_51), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_44), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_182), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_49), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_194), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_16), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_70), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_228), .Y(n_374) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_235), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_173), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_123), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_207), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_165), .Y(n_379) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_98), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_219), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_14), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_69), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_244), .B(n_36), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_324), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_304), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_331), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_252), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_304), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_269), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_331), .B(n_0), .Y(n_391) );
INVx3_ASAP7_75t_L g392 ( .A(n_304), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_266), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_358), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_304), .Y(n_395) );
BUFx8_ASAP7_75t_L g396 ( .A(n_259), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_252), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_304), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_284), .B(n_0), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_284), .B(n_1), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_263), .B(n_1), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_252), .Y(n_402) );
OAI21x1_ASAP7_75t_L g403 ( .A1(n_263), .A2(n_64), .B(n_62), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_252), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_345), .B(n_2), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_252), .Y(n_406) );
OA21x2_ASAP7_75t_L g407 ( .A1(n_279), .A2(n_66), .B(n_65), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_304), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_345), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_252), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_324), .Y(n_411) );
CKINVDCx16_ASAP7_75t_R g412 ( .A(n_271), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_273), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_324), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_253), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_256), .B(n_3), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_390), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_391), .A2(n_274), .B1(n_294), .B2(n_290), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_385), .Y(n_419) );
INVx4_ASAP7_75t_L g420 ( .A(n_392), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_387), .B(n_260), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_392), .Y(n_422) );
INVx3_ASAP7_75t_L g423 ( .A(n_405), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_392), .Y(n_424) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_385), .Y(n_425) );
INVx4_ASAP7_75t_L g426 ( .A(n_392), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_396), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_395), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_412), .B(n_302), .Y(n_429) );
INVxp67_ASAP7_75t_L g430 ( .A(n_415), .Y(n_430) );
AND2x4_ASAP7_75t_SL g431 ( .A(n_399), .B(n_300), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_396), .B(n_288), .Y(n_432) );
INVx2_ASAP7_75t_SL g433 ( .A(n_399), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_385), .Y(n_434) );
AND2x2_ASAP7_75t_SL g435 ( .A(n_405), .B(n_279), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_395), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_396), .B(n_316), .Y(n_437) );
INVx6_ASAP7_75t_L g438 ( .A(n_405), .Y(n_438) );
INVx3_ASAP7_75t_L g439 ( .A(n_405), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_396), .B(n_316), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_412), .B(n_255), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_415), .A2(n_315), .B1(n_281), .B2(n_306), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_395), .Y(n_443) );
INVx3_ASAP7_75t_L g444 ( .A(n_405), .Y(n_444) );
AO22x2_ASAP7_75t_L g445 ( .A1(n_391), .A2(n_278), .B1(n_311), .B2(n_299), .Y(n_445) );
INVx4_ASAP7_75t_L g446 ( .A(n_407), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_388), .Y(n_447) );
NAND2x1p5_ASAP7_75t_L g448 ( .A(n_400), .B(n_251), .Y(n_448) );
BUFx3_ASAP7_75t_L g449 ( .A(n_390), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_409), .B(n_283), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_388), .Y(n_451) );
BUFx2_ASAP7_75t_L g452 ( .A(n_400), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_388), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_391), .B(n_293), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_390), .B(n_293), .Y(n_455) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_385), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_397), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_397), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_452), .A2(n_330), .B1(n_354), .B2(n_393), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_417), .Y(n_460) );
INVx2_ASAP7_75t_SL g461 ( .A(n_454), .Y(n_461) );
NOR2x1_ASAP7_75t_L g462 ( .A(n_421), .B(n_401), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_423), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_433), .A2(n_333), .B1(n_334), .B2(n_301), .Y(n_464) );
BUFx3_ASAP7_75t_L g465 ( .A(n_427), .Y(n_465) );
AOI221xp5_ASAP7_75t_L g466 ( .A1(n_445), .A2(n_416), .B1(n_409), .B2(n_308), .C(n_319), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_427), .B(n_403), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_452), .B(n_416), .Y(n_468) );
AO22x1_ASAP7_75t_L g469 ( .A1(n_442), .A2(n_413), .B1(n_351), .B2(n_360), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_417), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_433), .A2(n_366), .B1(n_368), .B2(n_350), .Y(n_471) );
OAI221xp5_ASAP7_75t_L g472 ( .A1(n_418), .A2(n_297), .B1(n_322), .B2(n_321), .C(n_312), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_438), .Y(n_473) );
BUFx8_ASAP7_75t_L g474 ( .A(n_441), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_423), .Y(n_475) );
BUFx2_ASAP7_75t_L g476 ( .A(n_430), .Y(n_476) );
INVxp67_ASAP7_75t_SL g477 ( .A(n_448), .Y(n_477) );
BUFx8_ASAP7_75t_L g478 ( .A(n_441), .Y(n_478) );
INVx4_ASAP7_75t_L g479 ( .A(n_420), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_423), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_437), .B(n_403), .Y(n_481) );
BUFx2_ASAP7_75t_L g482 ( .A(n_421), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_448), .B(n_341), .Y(n_483) );
BUFx3_ASAP7_75t_L g484 ( .A(n_448), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_438), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_423), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_438), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_440), .B(n_432), .Y(n_488) );
INVx2_ASAP7_75t_SL g489 ( .A(n_431), .Y(n_489) );
OR2x4_ASAP7_75t_L g490 ( .A(n_429), .B(n_394), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_435), .B(n_386), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_435), .B(n_257), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_445), .A2(n_398), .B1(n_408), .B2(n_389), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_445), .A2(n_408), .B1(n_398), .B2(n_329), .Y(n_494) );
INVx4_ASAP7_75t_L g495 ( .A(n_420), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_439), .Y(n_496) );
OR2x6_ASAP7_75t_L g497 ( .A(n_445), .B(n_336), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_439), .B(n_359), .Y(n_498) );
OR2x6_ASAP7_75t_L g499 ( .A(n_431), .B(n_370), .Y(n_499) );
INVx4_ASAP7_75t_L g500 ( .A(n_420), .Y(n_500) );
NAND2x1p5_ASAP7_75t_L g501 ( .A(n_439), .B(n_372), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_449), .Y(n_502) );
AND2x2_ASAP7_75t_SL g503 ( .A(n_439), .B(n_407), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_449), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_444), .A2(n_402), .B1(n_404), .B2(n_397), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_444), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_444), .Y(n_507) );
BUFx3_ASAP7_75t_L g508 ( .A(n_458), .Y(n_508) );
INVxp67_ASAP7_75t_L g509 ( .A(n_450), .Y(n_509) );
NOR2x1p5_ASAP7_75t_L g510 ( .A(n_444), .B(n_267), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_451), .Y(n_511) );
INVx2_ASAP7_75t_SL g512 ( .A(n_455), .Y(n_512) );
INVx5_ASAP7_75t_L g513 ( .A(n_420), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_426), .B(n_275), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_446), .B(n_382), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_426), .B(n_285), .Y(n_516) );
BUFx3_ASAP7_75t_L g517 ( .A(n_458), .Y(n_517) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_446), .Y(n_518) );
AND2x6_ASAP7_75t_L g519 ( .A(n_447), .B(n_269), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_447), .A2(n_404), .B(n_406), .C(n_402), .Y(n_520) );
BUFx12f_ASAP7_75t_SL g521 ( .A(n_446), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_422), .B(n_287), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_453), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_453), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_446), .B(n_261), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_457), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_424), .Y(n_527) );
INVx4_ASAP7_75t_L g528 ( .A(n_428), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_424), .B(n_309), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_443), .B(n_291), .Y(n_530) );
OR2x6_ASAP7_75t_L g531 ( .A(n_428), .B(n_332), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_436), .B(n_404), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_472), .A2(n_406), .B(n_410), .C(n_443), .Y(n_533) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_508), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_517), .Y(n_535) );
INVx3_ASAP7_75t_L g536 ( .A(n_479), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_482), .B(n_355), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_476), .Y(n_538) );
INVx4_ASAP7_75t_L g539 ( .A(n_513), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_477), .Y(n_540) );
AOI222xp33_ASAP7_75t_L g541 ( .A1(n_466), .A2(n_469), .B1(n_474), .B2(n_478), .C1(n_468), .C2(n_459), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_518), .Y(n_542) );
AND2x2_ASAP7_75t_SL g543 ( .A(n_494), .B(n_407), .Y(n_543) );
INVx4_ASAP7_75t_L g544 ( .A(n_513), .Y(n_544) );
AOI22xp33_ASAP7_75t_SL g545 ( .A1(n_497), .A2(n_365), .B1(n_384), .B2(n_339), .Y(n_545) );
CKINVDCx14_ASAP7_75t_R g546 ( .A(n_531), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_518), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_507), .Y(n_548) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_513), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_503), .A2(n_407), .B(n_410), .Y(n_550) );
AND2x4_ASAP7_75t_L g551 ( .A(n_465), .B(n_313), .Y(n_551) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_493), .A2(n_365), .B(n_384), .C(n_339), .Y(n_552) );
INVxp67_ASAP7_75t_L g553 ( .A(n_531), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_484), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_499), .B(n_3), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_467), .A2(n_407), .B(n_262), .Y(n_556) );
BUFx2_ASAP7_75t_L g557 ( .A(n_499), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_498), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_497), .A2(n_264), .B1(n_265), .B2(n_254), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_523), .A2(n_268), .B1(n_276), .B2(n_270), .Y(n_560) );
CKINVDCx6p67_ASAP7_75t_R g561 ( .A(n_488), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_489), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_463), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_462), .B(n_367), .Y(n_564) );
BUFx12f_ASAP7_75t_L g565 ( .A(n_474), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_478), .Y(n_566) );
INVx2_ASAP7_75t_SL g567 ( .A(n_488), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_479), .B(n_310), .Y(n_568) );
INVx3_ASAP7_75t_L g569 ( .A(n_495), .Y(n_569) );
BUFx2_ASAP7_75t_L g570 ( .A(n_501), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_510), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_461), .B(n_320), .Y(n_572) );
OAI21xp33_ASAP7_75t_SL g573 ( .A1(n_523), .A2(n_282), .B(n_277), .Y(n_573) );
INVx3_ASAP7_75t_L g574 ( .A(n_495), .Y(n_574) );
NAND2xp33_ASAP7_75t_L g575 ( .A(n_519), .B(n_326), .Y(n_575) );
OAI22xp5_ASAP7_75t_SL g576 ( .A1(n_490), .A2(n_367), .B1(n_289), .B2(n_295), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_467), .A2(n_296), .B(n_286), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_509), .B(n_335), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_528), .Y(n_579) );
A2O1A1Ixp33_ASAP7_75t_L g580 ( .A1(n_515), .A2(n_305), .B(n_307), .C(n_298), .Y(n_580) );
AND2x4_ASAP7_75t_L g581 ( .A(n_512), .B(n_314), .Y(n_581) );
AND2x4_ASAP7_75t_L g582 ( .A(n_530), .B(n_318), .Y(n_582) );
BUFx3_ASAP7_75t_L g583 ( .A(n_515), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_530), .B(n_352), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_464), .B(n_292), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_524), .A2(n_327), .B1(n_328), .B2(n_323), .Y(n_586) );
NAND2x1_ASAP7_75t_L g587 ( .A(n_500), .B(n_272), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_471), .B(n_357), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_483), .B(n_356), .Y(n_589) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_528), .Y(n_590) );
A2O1A1Ixp33_ASAP7_75t_L g591 ( .A1(n_481), .A2(n_338), .B(n_342), .C(n_337), .Y(n_591) );
INVx3_ASAP7_75t_L g592 ( .A(n_485), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_463), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_491), .A2(n_367), .B1(n_344), .B2(n_346), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_475), .Y(n_595) );
AO21x2_ASAP7_75t_L g596 ( .A1(n_481), .A2(n_347), .B(n_343), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_525), .A2(n_475), .B1(n_486), .B2(n_480), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_480), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_486), .Y(n_599) );
INVx4_ASAP7_75t_L g600 ( .A(n_519), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_514), .B(n_363), .Y(n_601) );
A2O1A1Ixp33_ASAP7_75t_L g602 ( .A1(n_506), .A2(n_349), .B(n_353), .C(n_348), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_506), .Y(n_603) );
BUFx2_ASAP7_75t_R g604 ( .A(n_492), .Y(n_604) );
INVx3_ASAP7_75t_L g605 ( .A(n_485), .Y(n_605) );
A2O1A1Ixp33_ASAP7_75t_L g606 ( .A1(n_526), .A2(n_364), .B(n_371), .C(n_362), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_L g607 ( .A1(n_526), .A2(n_378), .B(n_379), .C(n_376), .Y(n_607) );
AO21x2_ASAP7_75t_L g608 ( .A1(n_520), .A2(n_383), .B(n_381), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_532), .B(n_4), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_525), .A2(n_340), .B1(n_373), .B2(n_303), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_496), .A2(n_280), .B1(n_377), .B2(n_374), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_527), .A2(n_377), .B(n_317), .Y(n_612) );
NOR2x1_ASAP7_75t_L g613 ( .A(n_522), .B(n_258), .Y(n_613) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_521), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_473), .A2(n_303), .B1(n_340), .B2(n_373), .Y(n_615) );
AND2x4_ASAP7_75t_L g616 ( .A(n_487), .B(n_4), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_511), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_505), .A2(n_369), .B1(n_361), .B2(n_411), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_529), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_460), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_516), .A2(n_414), .B(n_419), .Y(n_621) );
BUFx2_ASAP7_75t_SL g622 ( .A(n_519), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_470), .Y(n_623) );
INVx1_ASAP7_75t_SL g624 ( .A(n_519), .Y(n_624) );
INVx3_ASAP7_75t_L g625 ( .A(n_502), .Y(n_625) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_504), .Y(n_626) );
AND2x4_ASAP7_75t_L g627 ( .A(n_465), .B(n_5), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_477), .Y(n_628) );
BUFx2_ASAP7_75t_SL g629 ( .A(n_484), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_497), .A2(n_325), .B1(n_375), .B2(n_380), .Y(n_630) );
BUFx3_ASAP7_75t_L g631 ( .A(n_474), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_482), .B(n_6), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_482), .B(n_8), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_508), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_482), .B(n_9), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_497), .A2(n_325), .B1(n_375), .B2(n_380), .Y(n_636) );
INVx3_ASAP7_75t_SL g637 ( .A(n_531), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_465), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_550), .A2(n_425), .B(n_419), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_563), .Y(n_640) );
AOI22xp33_ASAP7_75t_SL g641 ( .A1(n_546), .A2(n_325), .B1(n_375), .B2(n_380), .Y(n_641) );
INVx8_ASAP7_75t_L g642 ( .A(n_565), .Y(n_642) );
OAI21xp5_ASAP7_75t_L g643 ( .A1(n_556), .A2(n_385), .B(n_375), .Y(n_643) );
INVx2_ASAP7_75t_SL g644 ( .A(n_631), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_566), .Y(n_645) );
OAI21xp5_ASAP7_75t_L g646 ( .A1(n_577), .A2(n_385), .B(n_380), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_593), .Y(n_647) );
INVx3_ASAP7_75t_L g648 ( .A(n_539), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_590), .Y(n_649) );
OAI21x1_ASAP7_75t_L g650 ( .A1(n_621), .A2(n_325), .B(n_385), .Y(n_650) );
OAI21x1_ASAP7_75t_SL g651 ( .A1(n_600), .A2(n_9), .B(n_10), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_540), .A2(n_10), .B1(n_12), .B2(n_13), .Y(n_652) );
BUFx3_ASAP7_75t_L g653 ( .A(n_538), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_590), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_553), .B(n_12), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_559), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_656) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_549), .Y(n_657) );
OAI21x1_ASAP7_75t_SL g658 ( .A1(n_600), .A2(n_17), .B(n_18), .Y(n_658) );
AO21x2_ASAP7_75t_L g659 ( .A1(n_596), .A2(n_456), .B(n_434), .Y(n_659) );
NAND2x1p5_ASAP7_75t_L g660 ( .A(n_570), .B(n_17), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_595), .Y(n_661) );
AND2x6_ASAP7_75t_L g662 ( .A(n_616), .B(n_21), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_557), .B(n_21), .Y(n_663) );
NOR2xp67_ASAP7_75t_L g664 ( .A(n_539), .B(n_68), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_598), .Y(n_665) );
INVx3_ASAP7_75t_L g666 ( .A(n_544), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_541), .B(n_456), .C(n_434), .Y(n_667) );
AND2x4_ASAP7_75t_L g668 ( .A(n_628), .B(n_22), .Y(n_668) );
OR2x2_ASAP7_75t_L g669 ( .A(n_537), .B(n_22), .Y(n_669) );
OAI21x1_ASAP7_75t_SL g670 ( .A1(n_559), .A2(n_23), .B(n_24), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_599), .Y(n_671) );
OR2x6_ASAP7_75t_L g672 ( .A(n_629), .B(n_23), .Y(n_672) );
BUFx3_ASAP7_75t_L g673 ( .A(n_637), .Y(n_673) );
BUFx3_ASAP7_75t_L g674 ( .A(n_554), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_590), .Y(n_675) );
AND2x6_ASAP7_75t_L g676 ( .A(n_616), .B(n_24), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_548), .Y(n_677) );
CKINVDCx14_ASAP7_75t_R g678 ( .A(n_576), .Y(n_678) );
INVx4_ASAP7_75t_SL g679 ( .A(n_627), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_581), .B(n_25), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_561), .B(n_25), .Y(n_681) );
CKINVDCx11_ASAP7_75t_R g682 ( .A(n_627), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_603), .Y(n_683) );
BUFx4f_ASAP7_75t_L g684 ( .A(n_555), .Y(n_684) );
OAI21x1_ASAP7_75t_L g685 ( .A1(n_612), .A2(n_73), .B(n_72), .Y(n_685) );
NAND2x1p5_ASAP7_75t_L g686 ( .A(n_638), .B(n_26), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_581), .B(n_26), .Y(n_687) );
AOI22x1_ASAP7_75t_L g688 ( .A1(n_542), .A2(n_136), .B1(n_246), .B2(n_245), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_534), .B(n_27), .Y(n_689) );
OAI22xp33_ASAP7_75t_L g690 ( .A1(n_632), .A2(n_28), .B1(n_30), .B2(n_31), .Y(n_690) );
INVx2_ASAP7_75t_SL g691 ( .A(n_614), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_541), .A2(n_28), .B1(n_30), .B2(n_32), .Y(n_692) );
A2O1A1Ixp33_ASAP7_75t_L g693 ( .A1(n_619), .A2(n_32), .B(n_33), .C(n_34), .Y(n_693) );
AO21x2_ASAP7_75t_L g694 ( .A1(n_596), .A2(n_75), .B(n_74), .Y(n_694) );
CKINVDCx6p67_ASAP7_75t_R g695 ( .A(n_551), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_609), .A2(n_34), .B1(n_35), .B2(n_37), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_633), .B(n_35), .Y(n_697) );
AO32x2_ASAP7_75t_L g698 ( .A1(n_560), .A2(n_38), .A3(n_39), .B1(n_40), .B2(n_41), .Y(n_698) );
INVx4_ASAP7_75t_L g699 ( .A(n_534), .Y(n_699) );
OAI21x1_ASAP7_75t_L g700 ( .A1(n_547), .A2(n_141), .B(n_243), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_576), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_560), .A2(n_38), .B1(n_40), .B2(n_42), .C(n_43), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_617), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_551), .B(n_42), .Y(n_704) );
AOI22xp33_ASAP7_75t_SL g705 ( .A1(n_571), .A2(n_44), .B1(n_45), .B2(n_46), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_635), .B(n_582), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_597), .Y(n_707) );
O2A1O1Ixp33_ASAP7_75t_L g708 ( .A1(n_552), .A2(n_47), .B(n_48), .C(n_50), .Y(n_708) );
OAI21x1_ASAP7_75t_L g709 ( .A1(n_625), .A2(n_149), .B(n_242), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_549), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_549), .Y(n_711) );
OAI21x1_ASAP7_75t_L g712 ( .A1(n_625), .A2(n_147), .B(n_240), .Y(n_712) );
OAI22xp33_ASAP7_75t_L g713 ( .A1(n_636), .A2(n_50), .B1(n_51), .B2(n_54), .Y(n_713) );
AND2x4_ASAP7_75t_SL g714 ( .A(n_534), .B(n_54), .Y(n_714) );
AO21x2_ASAP7_75t_L g715 ( .A1(n_608), .A2(n_146), .B(n_236), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_567), .A2(n_56), .B1(n_57), .B2(n_59), .Y(n_716) );
NAND2x1p5_ASAP7_75t_L g717 ( .A(n_544), .B(n_59), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_597), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_564), .Y(n_719) );
OAI221xp5_ASAP7_75t_L g720 ( .A1(n_585), .A2(n_60), .B1(n_76), .B2(n_77), .C(n_78), .Y(n_720) );
BUFx2_ASAP7_75t_L g721 ( .A(n_583), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_582), .A2(n_80), .B1(n_82), .B2(n_83), .Y(n_722) );
AO21x2_ASAP7_75t_L g723 ( .A1(n_608), .A2(n_86), .B(n_91), .Y(n_723) );
OR2x2_ASAP7_75t_L g724 ( .A(n_578), .B(n_92), .Y(n_724) );
AND2x4_ASAP7_75t_L g725 ( .A(n_558), .B(n_247), .Y(n_725) );
BUFx6f_ASAP7_75t_L g726 ( .A(n_536), .Y(n_726) );
CKINVDCx5p33_ASAP7_75t_R g727 ( .A(n_604), .Y(n_727) );
OAI21x1_ASAP7_75t_L g728 ( .A1(n_620), .A2(n_93), .B(n_94), .Y(n_728) );
OAI222xp33_ASAP7_75t_L g729 ( .A1(n_545), .A2(n_95), .B1(n_96), .B2(n_97), .C1(n_99), .C2(n_100), .Y(n_729) );
BUFx10_ASAP7_75t_L g730 ( .A(n_562), .Y(n_730) );
INVxp67_ASAP7_75t_SL g731 ( .A(n_630), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_623), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_586), .Y(n_733) );
INVx4_ASAP7_75t_L g734 ( .A(n_536), .Y(n_734) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_535), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_579), .Y(n_736) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_569), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_626), .Y(n_738) );
AO32x2_ASAP7_75t_L g739 ( .A1(n_586), .A2(n_101), .A3(n_104), .B1(n_107), .B2(n_108), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_533), .Y(n_740) );
AND2x4_ASAP7_75t_L g741 ( .A(n_634), .B(n_115), .Y(n_741) );
AND2x4_ASAP7_75t_L g742 ( .A(n_569), .B(n_234), .Y(n_742) );
OAI21x1_ASAP7_75t_L g743 ( .A1(n_587), .A2(n_116), .B(n_118), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_574), .Y(n_744) );
INVx2_ASAP7_75t_SL g745 ( .A(n_592), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_588), .B(n_121), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_574), .Y(n_747) );
OAI21x1_ASAP7_75t_L g748 ( .A1(n_613), .A2(n_122), .B(n_124), .Y(n_748) );
OAI22xp33_ASAP7_75t_L g749 ( .A1(n_636), .A2(n_125), .B1(n_126), .B2(n_127), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_626), .Y(n_750) );
BUFx2_ASAP7_75t_L g751 ( .A(n_573), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_584), .B(n_130), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_580), .B(n_131), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_573), .B(n_134), .Y(n_754) );
AND2x4_ASAP7_75t_L g755 ( .A(n_592), .B(n_135), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_611), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_703), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_639), .A2(n_643), .B(n_543), .Y(n_758) );
OR2x2_ASAP7_75t_L g759 ( .A(n_653), .B(n_572), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_703), .Y(n_760) );
AOI222xp33_ASAP7_75t_L g761 ( .A1(n_733), .A2(n_606), .B1(n_589), .B2(n_575), .C1(n_594), .C2(n_602), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_695), .B(n_605), .Y(n_762) );
AO31x2_ASAP7_75t_L g763 ( .A1(n_751), .A2(n_591), .A3(n_630), .B(n_611), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_668), .Y(n_764) );
INVx3_ASAP7_75t_L g765 ( .A(n_657), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_682), .B(n_605), .Y(n_766) );
AOI221xp5_ASAP7_75t_L g767 ( .A1(n_690), .A2(n_607), .B1(n_610), .B2(n_615), .C(n_601), .Y(n_767) );
OR2x2_ASAP7_75t_L g768 ( .A(n_669), .B(n_618), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_668), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_706), .B(n_618), .Y(n_770) );
AOI21xp33_ASAP7_75t_L g771 ( .A1(n_708), .A2(n_624), .B(n_626), .Y(n_771) );
INVxp67_ASAP7_75t_L g772 ( .A(n_672), .Y(n_772) );
OAI21xp5_ASAP7_75t_L g773 ( .A1(n_740), .A2(n_568), .B(n_622), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_684), .B(n_137), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_732), .Y(n_775) );
INVx4_ASAP7_75t_L g776 ( .A(n_642), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_640), .Y(n_777) );
AOI21xp5_ASAP7_75t_L g778 ( .A1(n_731), .A2(n_151), .B(n_154), .Y(n_778) );
OAI221xp5_ASAP7_75t_L g779 ( .A1(n_692), .A2(n_155), .B1(n_156), .B2(n_161), .C(n_162), .Y(n_779) );
INVx2_ASAP7_75t_SL g780 ( .A(n_642), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_707), .B(n_164), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_707), .A2(n_174), .B1(n_175), .B2(n_176), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_640), .Y(n_783) );
INVx3_ASAP7_75t_L g784 ( .A(n_657), .Y(n_784) );
BUFx12f_ASAP7_75t_L g785 ( .A(n_644), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_732), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_647), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_647), .Y(n_788) );
AOI221xp5_ASAP7_75t_L g789 ( .A1(n_756), .A2(n_179), .B1(n_180), .B2(n_184), .C(n_185), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_718), .B(n_186), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_756), .B(n_232), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_718), .B(n_188), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_678), .B(n_704), .Y(n_793) );
A2O1A1Ixp33_ASAP7_75t_L g794 ( .A1(n_746), .A2(n_189), .B(n_190), .C(n_191), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_656), .A2(n_192), .B1(n_193), .B2(n_195), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_662), .A2(n_196), .B1(n_197), .B2(n_198), .Y(n_796) );
OAI22xp33_ASAP7_75t_L g797 ( .A1(n_701), .A2(n_199), .B1(n_200), .B2(n_202), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_662), .A2(n_203), .B1(n_206), .B2(n_209), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_661), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_661), .B(n_211), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_665), .Y(n_801) );
AND2x2_ASAP7_75t_L g802 ( .A(n_679), .B(n_212), .Y(n_802) );
OAI211xp5_ASAP7_75t_L g803 ( .A1(n_656), .A2(n_214), .B(n_216), .C(n_217), .Y(n_803) );
AO31x2_ASAP7_75t_L g804 ( .A1(n_740), .A2(n_223), .A3(n_225), .B(n_227), .Y(n_804) );
CKINVDCx11_ASAP7_75t_R g805 ( .A(n_645), .Y(n_805) );
OAI21xp5_ASAP7_75t_L g806 ( .A1(n_754), .A2(n_646), .B(n_671), .Y(n_806) );
INVx3_ASAP7_75t_L g807 ( .A(n_657), .Y(n_807) );
OAI211xp5_ASAP7_75t_L g808 ( .A1(n_705), .A2(n_702), .B(n_641), .C(n_716), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_662), .A2(n_676), .B1(n_684), .B2(n_697), .Y(n_809) );
BUFx6f_ASAP7_75t_L g810 ( .A(n_699), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_662), .A2(n_676), .B1(n_719), .B2(n_655), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_665), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_676), .A2(n_719), .B1(n_672), .B2(n_687), .Y(n_813) );
AND2x2_ASAP7_75t_L g814 ( .A(n_679), .B(n_660), .Y(n_814) );
OR2x6_ASAP7_75t_L g815 ( .A(n_673), .B(n_717), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_671), .Y(n_816) );
A2O1A1Ixp33_ASAP7_75t_L g817 ( .A1(n_725), .A2(n_667), .B(n_753), .C(n_693), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_683), .Y(n_818) );
OAI22xp33_ASAP7_75t_L g819 ( .A1(n_686), .A2(n_727), .B1(n_680), .B2(n_696), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_683), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_735), .B(n_676), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_674), .B(n_721), .Y(n_822) );
AOI21xp33_ASAP7_75t_L g823 ( .A1(n_720), .A2(n_659), .B(n_713), .Y(n_823) );
OR2x6_ASAP7_75t_L g824 ( .A(n_725), .B(n_742), .Y(n_824) );
INVx3_ASAP7_75t_L g825 ( .A(n_699), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_730), .B(n_663), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_670), .A2(n_681), .B1(n_752), .B2(n_691), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_741), .A2(n_652), .B1(n_648), .B2(n_666), .Y(n_828) );
AO21x2_ASAP7_75t_L g829 ( .A1(n_715), .A2(n_723), .B(n_659), .Y(n_829) );
AND2x2_ASAP7_75t_L g830 ( .A(n_730), .B(n_714), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_677), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_741), .A2(n_648), .B1(n_666), .B2(n_744), .Y(n_832) );
INVx3_ASAP7_75t_L g833 ( .A(n_734), .Y(n_833) );
AOI221xp5_ASAP7_75t_L g834 ( .A1(n_689), .A2(n_729), .B1(n_651), .B2(n_658), .C(n_749), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_744), .A2(n_747), .B1(n_742), .B2(n_724), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_747), .A2(n_755), .B1(n_734), .B2(n_736), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_649), .Y(n_837) );
AND2x2_ASAP7_75t_L g838 ( .A(n_698), .B(n_745), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_698), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_654), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_698), .B(n_675), .Y(n_841) );
INVx3_ASAP7_75t_L g842 ( .A(n_726), .Y(n_842) );
OAI22xp33_ASAP7_75t_L g843 ( .A1(n_726), .A2(n_737), .B1(n_664), .B2(n_711), .Y(n_843) );
BUFx3_ASAP7_75t_L g844 ( .A(n_710), .Y(n_844) );
OAI221xp5_ASAP7_75t_SL g845 ( .A1(n_722), .A2(n_739), .B1(n_738), .B2(n_750), .C(n_694), .Y(n_845) );
INVx6_ASAP7_75t_L g846 ( .A(n_726), .Y(n_846) );
INVx3_ASAP7_75t_L g847 ( .A(n_737), .Y(n_847) );
OR2x2_ASAP7_75t_L g848 ( .A(n_737), .B(n_755), .Y(n_848) );
NAND3xp33_ASAP7_75t_L g849 ( .A(n_688), .B(n_739), .C(n_748), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_739), .A2(n_709), .B1(n_712), .B2(n_728), .Y(n_850) );
AOI222xp33_ASAP7_75t_L g851 ( .A1(n_743), .A2(n_733), .B1(n_576), .B2(n_701), .C1(n_682), .C2(n_466), .Y(n_851) );
AOI22xp5_ASAP7_75t_L g852 ( .A1(n_685), .A2(n_733), .B1(n_482), .B2(n_393), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_700), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_668), .Y(n_854) );
AOI21xp33_ASAP7_75t_L g855 ( .A1(n_708), .A2(n_740), .B(n_497), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_756), .B(n_452), .Y(n_856) );
AOI21xp5_ASAP7_75t_L g857 ( .A1(n_639), .A2(n_556), .B(n_643), .Y(n_857) );
AOI22x1_ASAP7_75t_SL g858 ( .A1(n_733), .A2(n_566), .B1(n_727), .B2(n_701), .Y(n_858) );
OA21x2_ASAP7_75t_L g859 ( .A1(n_643), .A2(n_639), .B(n_650), .Y(n_859) );
OR2x2_ASAP7_75t_L g860 ( .A(n_653), .B(n_482), .Y(n_860) );
BUFx12f_ASAP7_75t_L g861 ( .A(n_682), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_707), .B(n_718), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_733), .B(n_482), .Y(n_863) );
BUFx3_ASAP7_75t_L g864 ( .A(n_642), .Y(n_864) );
AOI221xp5_ASAP7_75t_L g865 ( .A1(n_690), .A2(n_445), .B1(n_576), .B2(n_472), .C(n_482), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_733), .A2(n_497), .B1(n_541), .B2(n_662), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_733), .A2(n_482), .B1(n_393), .B2(n_413), .Y(n_867) );
OAI22xp33_ASAP7_75t_L g868 ( .A1(n_733), .A2(n_497), .B1(n_531), .B2(n_637), .Y(n_868) );
NAND2xp5_ASAP7_75t_SL g869 ( .A(n_733), .B(n_679), .Y(n_869) );
OAI22xp33_ASAP7_75t_L g870 ( .A1(n_733), .A2(n_497), .B1(n_531), .B2(n_637), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_824), .B(n_757), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_824), .B(n_760), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_859), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_799), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_824), .B(n_777), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_783), .Y(n_876) );
INVx1_ASAP7_75t_SL g877 ( .A(n_805), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_787), .Y(n_878) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_860), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_788), .B(n_820), .Y(n_880) );
INVx2_ASAP7_75t_L g881 ( .A(n_829), .Y(n_881) );
AND2x2_ASAP7_75t_L g882 ( .A(n_801), .B(n_812), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_816), .B(n_818), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_775), .B(n_786), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_831), .B(n_862), .Y(n_885) );
INVx4_ASAP7_75t_L g886 ( .A(n_810), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_863), .B(n_770), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_862), .B(n_866), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_839), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_809), .B(n_851), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_838), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_841), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_804), .Y(n_893) );
INVx4_ASAP7_75t_L g894 ( .A(n_810), .Y(n_894) );
BUFx2_ASAP7_75t_L g895 ( .A(n_821), .Y(n_895) );
INVx3_ASAP7_75t_L g896 ( .A(n_810), .Y(n_896) );
HB1xp67_ASAP7_75t_L g897 ( .A(n_822), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_851), .B(n_764), .Y(n_898) );
BUFx3_ASAP7_75t_L g899 ( .A(n_833), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_865), .B(n_768), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_804), .Y(n_901) );
INVx3_ASAP7_75t_L g902 ( .A(n_833), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_804), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_769), .B(n_854), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_837), .B(n_840), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_800), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_800), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_781), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_868), .A2(n_870), .B1(n_819), .B2(n_761), .Y(n_909) );
HB1xp67_ASAP7_75t_L g910 ( .A(n_815), .Y(n_910) );
INVxp67_ASAP7_75t_L g911 ( .A(n_864), .Y(n_911) );
INVx2_ASAP7_75t_SL g912 ( .A(n_815), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_813), .B(n_811), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_781), .Y(n_914) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_815), .Y(n_915) );
BUFx2_ASAP7_75t_L g916 ( .A(n_848), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_790), .Y(n_917) );
OR2x2_ASAP7_75t_L g918 ( .A(n_856), .B(n_869), .Y(n_918) );
HB1xp67_ASAP7_75t_L g919 ( .A(n_759), .Y(n_919) );
HB1xp67_ASAP7_75t_L g920 ( .A(n_772), .Y(n_920) );
BUFx2_ASAP7_75t_L g921 ( .A(n_853), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_825), .B(n_847), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_790), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_792), .Y(n_924) );
INVxp67_ASAP7_75t_SL g925 ( .A(n_835), .Y(n_925) );
AND2x4_ASAP7_75t_L g926 ( .A(n_765), .B(n_807), .Y(n_926) );
BUFx2_ASAP7_75t_L g927 ( .A(n_765), .Y(n_927) );
INVxp67_ASAP7_75t_L g928 ( .A(n_867), .Y(n_928) );
HB1xp67_ASAP7_75t_L g929 ( .A(n_830), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_825), .B(n_842), .Y(n_930) );
OR2x2_ASAP7_75t_L g931 ( .A(n_827), .B(n_836), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_791), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_806), .Y(n_933) );
NOR2x1_ASAP7_75t_SL g934 ( .A(n_795), .B(n_782), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_806), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_793), .B(n_826), .Y(n_936) );
INVx2_ASAP7_75t_L g937 ( .A(n_784), .Y(n_937) );
HB1xp67_ASAP7_75t_L g938 ( .A(n_814), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_842), .B(n_847), .Y(n_939) );
INVx5_ASAP7_75t_SL g940 ( .A(n_776), .Y(n_940) );
INVx2_ASAP7_75t_SL g941 ( .A(n_846), .Y(n_941) );
INVx2_ASAP7_75t_L g942 ( .A(n_784), .Y(n_942) );
INVx2_ASAP7_75t_L g943 ( .A(n_807), .Y(n_943) );
BUFx2_ASAP7_75t_L g944 ( .A(n_844), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_802), .B(n_832), .Y(n_945) );
OAI21xp33_ASAP7_75t_L g946 ( .A1(n_795), .A2(n_852), .B(n_808), .Y(n_946) );
OR2x2_ASAP7_75t_L g947 ( .A(n_828), .B(n_763), .Y(n_947) );
AND2x2_ASAP7_75t_L g948 ( .A(n_763), .B(n_846), .Y(n_948) );
BUFx2_ASAP7_75t_L g949 ( .A(n_763), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_850), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_850), .Y(n_951) );
AND2x4_ASAP7_75t_L g952 ( .A(n_773), .B(n_758), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_849), .Y(n_953) );
OR2x2_ASAP7_75t_L g954 ( .A(n_845), .B(n_817), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_849), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_761), .A2(n_767), .B1(n_855), .B2(n_834), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_855), .B(n_773), .Y(n_957) );
AND2x4_ASAP7_75t_L g958 ( .A(n_857), .B(n_778), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_891), .B(n_823), .Y(n_959) );
INVx1_ASAP7_75t_SL g960 ( .A(n_879), .Y(n_960) );
INVx2_ASAP7_75t_L g961 ( .A(n_873), .Y(n_961) );
INVx2_ASAP7_75t_SL g962 ( .A(n_899), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_891), .B(n_823), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_882), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_882), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_885), .B(n_766), .Y(n_966) );
NOR3xp33_ASAP7_75t_L g967 ( .A(n_928), .B(n_776), .C(n_774), .Y(n_967) );
AND2x4_ASAP7_75t_L g968 ( .A(n_948), .B(n_798), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_892), .B(n_782), .Y(n_969) );
AND2x4_ASAP7_75t_L g970 ( .A(n_948), .B(n_796), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_889), .Y(n_971) );
INVx3_ASAP7_75t_L g972 ( .A(n_886), .Y(n_972) );
OAI211xp5_ASAP7_75t_L g973 ( .A1(n_909), .A2(n_762), .B(n_803), .C(n_771), .Y(n_973) );
NAND2x1_ASAP7_75t_L g974 ( .A(n_902), .B(n_843), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_883), .Y(n_975) );
INVx2_ASAP7_75t_SL g976 ( .A(n_899), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_956), .A2(n_797), .B1(n_779), .B2(n_789), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_885), .B(n_780), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_883), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_898), .B(n_858), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_898), .B(n_785), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_884), .Y(n_982) );
INVx1_ASAP7_75t_SL g983 ( .A(n_938), .Y(n_983) );
INVx2_ASAP7_75t_L g984 ( .A(n_873), .Y(n_984) );
AND2x4_ASAP7_75t_L g985 ( .A(n_892), .B(n_794), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_900), .B(n_771), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_884), .B(n_861), .Y(n_987) );
INVx2_ASAP7_75t_L g988 ( .A(n_873), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_876), .B(n_888), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_889), .Y(n_990) );
AND2x2_ASAP7_75t_L g991 ( .A(n_876), .B(n_888), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_874), .Y(n_992) );
AOI221xp5_ASAP7_75t_L g993 ( .A1(n_890), .A2(n_946), .B1(n_887), .B2(n_925), .C(n_919), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_876), .B(n_874), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_949), .B(n_880), .Y(n_995) );
AND2x4_ASAP7_75t_L g996 ( .A(n_886), .B(n_894), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_949), .B(n_880), .Y(n_997) );
NOR2xp33_ASAP7_75t_SL g998 ( .A(n_877), .B(n_912), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_878), .B(n_957), .Y(n_999) );
INVx5_ASAP7_75t_L g1000 ( .A(n_940), .Y(n_1000) );
BUFx8_ASAP7_75t_L g1001 ( .A(n_912), .Y(n_1001) );
INVx2_ASAP7_75t_SL g1002 ( .A(n_899), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_878), .B(n_957), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_947), .B(n_905), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_947), .B(n_905), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_890), .B(n_897), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_904), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_950), .B(n_951), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_950), .B(n_951), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_904), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_918), .Y(n_1011) );
AO22x1_ASAP7_75t_L g1012 ( .A1(n_921), .A2(n_913), .B1(n_895), .B2(n_915), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_921), .B(n_913), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_918), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_952), .B(n_871), .Y(n_1015) );
AOI22xp5_ASAP7_75t_L g1016 ( .A1(n_946), .A2(n_931), .B1(n_872), .B2(n_875), .Y(n_1016) );
OR2x2_ASAP7_75t_L g1017 ( .A(n_895), .B(n_931), .Y(n_1017) );
AND2x4_ASAP7_75t_SL g1018 ( .A(n_910), .B(n_886), .Y(n_1018) );
AND2x4_ASAP7_75t_L g1019 ( .A(n_886), .B(n_894), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_893), .Y(n_1020) );
INVx3_ASAP7_75t_L g1021 ( .A(n_894), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_871), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_872), .B(n_875), .Y(n_1023) );
INVx3_ASAP7_75t_L g1024 ( .A(n_894), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_952), .B(n_933), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_916), .B(n_920), .Y(n_1026) );
HB1xp67_ASAP7_75t_L g1027 ( .A(n_944), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_916), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_952), .B(n_933), .Y(n_1029) );
INVx2_ASAP7_75t_SL g1030 ( .A(n_896), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_929), .B(n_944), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_952), .B(n_935), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_935), .B(n_917), .Y(n_1033) );
OAI21xp33_ASAP7_75t_L g1034 ( .A1(n_993), .A2(n_954), .B(n_936), .Y(n_1034) );
NOR3xp33_ASAP7_75t_SL g1035 ( .A(n_973), .B(n_940), .C(n_901), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_1013), .B(n_945), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_964), .B(n_945), .Y(n_1037) );
OR2x2_ASAP7_75t_L g1038 ( .A(n_960), .B(n_927), .Y(n_1038) );
AND2x2_ASAP7_75t_SL g1039 ( .A(n_1018), .B(n_954), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_1025), .B(n_955), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_992), .Y(n_1041) );
NAND2xp5_ASAP7_75t_SL g1042 ( .A(n_962), .B(n_902), .Y(n_1042) );
NAND4xp25_ASAP7_75t_L g1043 ( .A(n_1006), .B(n_911), .C(n_932), .D(n_930), .Y(n_1043) );
AND2x4_ASAP7_75t_L g1044 ( .A(n_1015), .B(n_881), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_1013), .B(n_927), .Y(n_1045) );
HB1xp67_ASAP7_75t_L g1046 ( .A(n_1027), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_965), .B(n_930), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_975), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_979), .B(n_923), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_982), .Y(n_1050) );
INVxp67_ASAP7_75t_SL g1051 ( .A(n_961), .Y(n_1051) );
AND2x4_ASAP7_75t_L g1052 ( .A(n_1015), .B(n_881), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_966), .B(n_922), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_971), .Y(n_1054) );
OR2x2_ASAP7_75t_L g1055 ( .A(n_983), .B(n_896), .Y(n_1055) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_984), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_1023), .B(n_922), .Y(n_1057) );
AND2x4_ASAP7_75t_L g1058 ( .A(n_1025), .B(n_881), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_971), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_1004), .B(n_896), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_1007), .B(n_923), .Y(n_1061) );
INVx2_ASAP7_75t_SL g1062 ( .A(n_1018), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_990), .Y(n_1063) );
XNOR2x2_ASAP7_75t_L g1064 ( .A(n_1031), .B(n_903), .Y(n_1064) );
INVx4_ASAP7_75t_L g1065 ( .A(n_1000), .Y(n_1065) );
OR2x6_ASAP7_75t_L g1066 ( .A(n_1012), .B(n_902), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1010), .B(n_914), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_990), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1026), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_1004), .B(n_896), .Y(n_1070) );
NOR2xp67_ASAP7_75t_SL g1071 ( .A(n_1000), .B(n_940), .Y(n_1071) );
NOR2xp33_ASAP7_75t_L g1072 ( .A(n_981), .B(n_932), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_1005), .B(n_939), .Y(n_1073) );
OR2x2_ASAP7_75t_L g1074 ( .A(n_1017), .B(n_902), .Y(n_1074) );
HB1xp67_ASAP7_75t_L g1075 ( .A(n_988), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_994), .Y(n_1076) );
NOR2xp33_ASAP7_75t_L g1077 ( .A(n_980), .B(n_934), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_1011), .B(n_908), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_994), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1014), .Y(n_1080) );
NOR2xp67_ASAP7_75t_L g1081 ( .A(n_1000), .B(n_955), .Y(n_1081) );
BUFx3_ASAP7_75t_L g1082 ( .A(n_1001), .Y(n_1082) );
CKINVDCx5p33_ASAP7_75t_R g1083 ( .A(n_1001), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1028), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_999), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_999), .Y(n_1086) );
OR2x2_ASAP7_75t_L g1087 ( .A(n_1017), .B(n_907), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1003), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_1003), .B(n_917), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_1005), .B(n_939), .Y(n_1090) );
NOR2xp67_ASAP7_75t_SL g1091 ( .A(n_1000), .B(n_940), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_995), .Y(n_1092) );
AND2x4_ASAP7_75t_SL g1093 ( .A(n_996), .B(n_926), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1029), .B(n_953), .Y(n_1094) );
OR2x2_ASAP7_75t_L g1095 ( .A(n_1085), .B(n_1029), .Y(n_1095) );
OR2x2_ASAP7_75t_L g1096 ( .A(n_1086), .B(n_1032), .Y(n_1096) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1056), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_1040), .B(n_1032), .Y(n_1098) );
INVx1_ASAP7_75t_SL g1099 ( .A(n_1083), .Y(n_1099) );
OR2x6_ASAP7_75t_L g1100 ( .A(n_1066), .B(n_1012), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1041), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1046), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g1103 ( .A(n_1046), .Y(n_1103) );
NAND2x1_ASAP7_75t_SL g1104 ( .A(n_1065), .B(n_972), .Y(n_1104) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_1069), .B(n_1088), .Y(n_1105) );
O2A1O1Ixp33_ASAP7_75t_L g1106 ( .A1(n_1034), .A2(n_967), .B(n_987), .C(n_978), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1054), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_1080), .B(n_1036), .Y(n_1108) );
OAI22xp5_ASAP7_75t_L g1109 ( .A1(n_1039), .A2(n_1000), .B1(n_1016), .B2(n_940), .Y(n_1109) );
INVx2_ASAP7_75t_L g1110 ( .A(n_1056), .Y(n_1110) );
AOI21xp5_ASAP7_75t_L g1111 ( .A1(n_1042), .A2(n_934), .B(n_974), .Y(n_1111) );
INVx2_ASAP7_75t_L g1112 ( .A(n_1075), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_1048), .B(n_989), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1059), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1040), .B(n_1008), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1050), .B(n_989), .Y(n_1116) );
INVx2_ASAP7_75t_L g1117 ( .A(n_1075), .Y(n_1117) );
BUFx2_ASAP7_75t_L g1118 ( .A(n_1062), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1063), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1094), .B(n_1008), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1068), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_1092), .B(n_991), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1084), .Y(n_1123) );
INVx6_ASAP7_75t_L g1124 ( .A(n_1065), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1076), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1094), .B(n_1009), .Y(n_1126) );
OR2x2_ASAP7_75t_L g1127 ( .A(n_1079), .B(n_997), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1047), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1044), .B(n_1009), .Y(n_1129) );
OR2x2_ASAP7_75t_L g1130 ( .A(n_1087), .B(n_995), .Y(n_1130) );
NAND3xp33_ASAP7_75t_SL g1131 ( .A(n_1083), .B(n_998), .C(n_974), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1044), .B(n_997), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1044), .B(n_959), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1072), .B(n_991), .Y(n_1134) );
HB1xp67_ASAP7_75t_L g1135 ( .A(n_1038), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_1072), .B(n_1033), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_1037), .B(n_1033), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1073), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1090), .Y(n_1139) );
OAI221xp5_ASAP7_75t_L g1140 ( .A1(n_1106), .A2(n_1043), .B1(n_1077), .B2(n_1082), .C(n_1035), .Y(n_1140) );
OAI21xp5_ASAP7_75t_L g1141 ( .A1(n_1131), .A2(n_1035), .B(n_1039), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1103), .Y(n_1142) );
O2A1O1Ixp5_ASAP7_75t_L g1143 ( .A1(n_1109), .A2(n_1065), .B(n_1091), .C(n_1071), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1101), .Y(n_1144) );
OAI21xp33_ASAP7_75t_L g1145 ( .A1(n_1133), .A2(n_1077), .B(n_1066), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1146 ( .A(n_1115), .B(n_1057), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_1135), .A2(n_970), .B1(n_968), .B2(n_1045), .Y(n_1147) );
AOI21xp5_ASAP7_75t_L g1148 ( .A1(n_1111), .A2(n_1042), .B(n_1066), .Y(n_1148) );
OAI21xp33_ASAP7_75t_L g1149 ( .A1(n_1133), .A2(n_1055), .B(n_1053), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1102), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1123), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1095), .Y(n_1152) );
AOI21xp33_ASAP7_75t_SL g1153 ( .A1(n_1100), .A2(n_1062), .B(n_1019), .Y(n_1153) );
OAI22xp33_ASAP7_75t_L g1154 ( .A1(n_1124), .A2(n_1082), .B1(n_1081), .B2(n_1002), .Y(n_1154) );
OAI22xp33_ASAP7_75t_L g1155 ( .A1(n_1124), .A2(n_962), .B1(n_1002), .B2(n_976), .Y(n_1155) );
NAND2x1_ASAP7_75t_L g1156 ( .A(n_1124), .B(n_972), .Y(n_1156) );
OAI21xp5_ASAP7_75t_SL g1157 ( .A1(n_1118), .A2(n_1093), .B(n_996), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1095), .Y(n_1158) );
OAI31xp33_ASAP7_75t_SL g1159 ( .A1(n_1099), .A2(n_996), .A3(n_1019), .B(n_1060), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1098), .B(n_1070), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1098), .B(n_1052), .Y(n_1161) );
OR2x2_ASAP7_75t_L g1162 ( .A(n_1130), .B(n_1089), .Y(n_1162) );
AOI21xp33_ASAP7_75t_L g1163 ( .A1(n_1100), .A2(n_1078), .B(n_1049), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1115), .B(n_1052), .Y(n_1164) );
XNOR2xp5_ASAP7_75t_L g1165 ( .A(n_1138), .B(n_1093), .Y(n_1165) );
NOR2xp33_ASAP7_75t_L g1166 ( .A(n_1128), .B(n_1001), .Y(n_1166) );
OAI21xp33_ASAP7_75t_L g1167 ( .A1(n_1100), .A2(n_1052), .B(n_963), .Y(n_1167) );
AND2x4_ASAP7_75t_L g1168 ( .A(n_1118), .B(n_1058), .Y(n_1168) );
INVxp67_ASAP7_75t_L g1169 ( .A(n_1097), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1142), .Y(n_1170) );
AOI21xp5_ASAP7_75t_L g1171 ( .A1(n_1159), .A2(n_1100), .B(n_1019), .Y(n_1171) );
OAI211xp5_ASAP7_75t_L g1172 ( .A1(n_1157), .A2(n_1104), .B(n_1105), .C(n_1136), .Y(n_1172) );
INVxp67_ASAP7_75t_SL g1173 ( .A(n_1169), .Y(n_1173) );
AOI21xp33_ASAP7_75t_L g1174 ( .A1(n_1140), .A2(n_1061), .B(n_1067), .Y(n_1174) );
INVxp67_ASAP7_75t_SL g1175 ( .A(n_1169), .Y(n_1175) );
NAND2xp5_ASAP7_75t_SL g1176 ( .A(n_1143), .B(n_1097), .Y(n_1176) );
A2O1A1Ixp33_ASAP7_75t_L g1177 ( .A1(n_1153), .A2(n_1104), .B(n_1130), .C(n_1134), .Y(n_1177) );
AOI222xp33_ASAP7_75t_L g1178 ( .A1(n_1140), .A2(n_1139), .B1(n_1125), .B2(n_1126), .C1(n_1120), .C2(n_1129), .Y(n_1178) );
OAI222xp33_ASAP7_75t_L g1179 ( .A1(n_1148), .A2(n_1127), .B1(n_1096), .B2(n_1108), .C1(n_1120), .C2(n_1126), .Y(n_1179) );
OAI21xp5_ASAP7_75t_L g1180 ( .A1(n_1143), .A2(n_977), .B(n_976), .Y(n_1180) );
OAI21xp5_ASAP7_75t_L g1181 ( .A1(n_1148), .A2(n_986), .B(n_1024), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1144), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1151), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1150), .Y(n_1184) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1152), .Y(n_1185) );
AOI21xp33_ASAP7_75t_L g1186 ( .A1(n_1167), .A2(n_1121), .B(n_1107), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1158), .Y(n_1187) );
OAI22xp5_ASAP7_75t_L g1188 ( .A1(n_1165), .A2(n_1124), .B1(n_1127), .B2(n_1096), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g1189 ( .A1(n_1141), .A2(n_1137), .B1(n_1122), .B2(n_1113), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1178), .B(n_1164), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1185), .Y(n_1191) );
OAI221xp5_ASAP7_75t_SL g1192 ( .A1(n_1172), .A2(n_1145), .B1(n_1147), .B2(n_1154), .C(n_1149), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1185), .Y(n_1193) );
OAI21xp33_ASAP7_75t_L g1194 ( .A1(n_1177), .A2(n_1163), .B(n_1168), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1182), .Y(n_1195) );
AOI221xp5_ASAP7_75t_L g1196 ( .A1(n_1179), .A2(n_1146), .B1(n_1166), .B2(n_1160), .C(n_1162), .Y(n_1196) );
AOI221xp5_ASAP7_75t_L g1197 ( .A1(n_1189), .A2(n_1168), .B1(n_1161), .B2(n_1155), .C(n_1114), .Y(n_1197) );
AOI21xp33_ASAP7_75t_L g1198 ( .A1(n_1180), .A2(n_1156), .B(n_1119), .Y(n_1198) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1183), .Y(n_1199) );
HB1xp67_ASAP7_75t_L g1200 ( .A(n_1173), .Y(n_1200) );
AOI21xp33_ASAP7_75t_L g1201 ( .A1(n_1181), .A2(n_941), .B(n_1030), .Y(n_1201) );
AOI21xp5_ASAP7_75t_L g1202 ( .A1(n_1171), .A2(n_1116), .B(n_1112), .Y(n_1202) );
INVx2_ASAP7_75t_SL g1203 ( .A(n_1200), .Y(n_1203) );
AOI221xp5_ASAP7_75t_L g1204 ( .A1(n_1192), .A2(n_1174), .B1(n_1188), .B2(n_1186), .C(n_1177), .Y(n_1204) );
AND2x2_ASAP7_75t_SL g1205 ( .A(n_1200), .B(n_1176), .Y(n_1205) );
AOI222xp33_ASAP7_75t_L g1206 ( .A1(n_1196), .A2(n_1176), .B1(n_1175), .B2(n_1170), .C1(n_1187), .C2(n_1184), .Y(n_1206) );
NAND3xp33_ASAP7_75t_L g1207 ( .A(n_1192), .B(n_1030), .C(n_901), .Y(n_1207) );
AOI221xp5_ASAP7_75t_L g1208 ( .A1(n_1197), .A2(n_1129), .B1(n_1132), .B2(n_1022), .C(n_1112), .Y(n_1208) );
A2O1A1Ixp33_ASAP7_75t_L g1209 ( .A1(n_1202), .A2(n_1132), .B(n_1024), .C(n_1021), .Y(n_1209) );
OAI321xp33_ASAP7_75t_L g1210 ( .A1(n_1194), .A2(n_1074), .A3(n_963), .B1(n_959), .B2(n_1117), .C(n_1110), .Y(n_1210) );
AOI211xp5_ASAP7_75t_L g1211 ( .A1(n_1198), .A2(n_969), .B(n_985), .C(n_970), .Y(n_1211) );
NAND5xp2_ASAP7_75t_L g1212 ( .A(n_1204), .B(n_1190), .C(n_1201), .D(n_969), .E(n_1195), .Y(n_1212) );
NAND2xp33_ASAP7_75t_R g1213 ( .A(n_1205), .B(n_1024), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1203), .B(n_1199), .Y(n_1214) );
NOR3xp33_ASAP7_75t_L g1215 ( .A(n_1207), .B(n_1193), .C(n_1191), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1209), .Y(n_1216) );
OAI221xp5_ASAP7_75t_L g1217 ( .A1(n_1206), .A2(n_1117), .B1(n_1110), .B2(n_972), .C(n_1021), .Y(n_1217) );
NAND3xp33_ASAP7_75t_SL g1218 ( .A(n_1216), .B(n_1208), .C(n_1211), .Y(n_1218) );
NAND3xp33_ASAP7_75t_L g1219 ( .A(n_1213), .B(n_1210), .C(n_941), .Y(n_1219) );
OAI221xp5_ASAP7_75t_SL g1220 ( .A1(n_1217), .A2(n_1021), .B1(n_1064), .B2(n_1020), .C(n_1051), .Y(n_1220) );
INVx2_ASAP7_75t_L g1221 ( .A(n_1214), .Y(n_1221) );
NOR2xp33_ASAP7_75t_L g1222 ( .A(n_1212), .B(n_1064), .Y(n_1222) );
OAI22xp5_ASAP7_75t_SL g1223 ( .A1(n_1222), .A2(n_1213), .B1(n_1215), .B2(n_985), .Y(n_1223) );
NAND3xp33_ASAP7_75t_L g1224 ( .A(n_1219), .B(n_926), .C(n_937), .Y(n_1224) );
OAI21xp5_ASAP7_75t_L g1225 ( .A1(n_1218), .A2(n_985), .B(n_958), .Y(n_1225) );
BUFx3_ASAP7_75t_L g1226 ( .A(n_1221), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1226), .Y(n_1227) );
OAI22xp5_ASAP7_75t_L g1228 ( .A1(n_1223), .A2(n_1220), .B1(n_1058), .B2(n_1020), .Y(n_1228) );
OAI22x1_ASAP7_75t_L g1229 ( .A1(n_1224), .A2(n_926), .B1(n_968), .B2(n_970), .Y(n_1229) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1227), .Y(n_1230) );
OAI21xp5_ASAP7_75t_L g1231 ( .A1(n_1228), .A2(n_1225), .B(n_1229), .Y(n_1231) );
OAI221xp5_ASAP7_75t_L g1232 ( .A1(n_1230), .A2(n_907), .B1(n_906), .B2(n_924), .C(n_908), .Y(n_1232) );
AO221x2_ASAP7_75t_L g1233 ( .A1(n_1232), .A2(n_1231), .B1(n_937), .B2(n_943), .C(n_942), .Y(n_1233) );
AOI21xp5_ASAP7_75t_L g1234 ( .A1(n_1233), .A2(n_943), .B(n_937), .Y(n_1234) );
endmodule