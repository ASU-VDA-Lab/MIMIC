module fake_jpeg_29784_n_549 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_549);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_549;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_15),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_55),
.B(n_85),
.Y(n_137)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_57),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_21),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_58),
.B(n_71),
.Y(n_117)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g167 ( 
.A(n_61),
.Y(n_167)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_63),
.Y(n_168)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_15),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_74),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_21),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_72),
.Y(n_141)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_22),
.B(n_15),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_75),
.B(n_77),
.Y(n_144)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_21),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_83),
.Y(n_148)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_22),
.B(n_14),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx11_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_88),
.Y(n_165)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_89),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_90),
.Y(n_164)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_27),
.B(n_14),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_93),
.B(n_105),
.C(n_26),
.Y(n_146)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_25),
.B(n_12),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_97),
.B(n_100),
.Y(n_147)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_18),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_18),
.Y(n_102)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_18),
.Y(n_103)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_18),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

HAxp5_ASAP7_75t_SL g105 ( 
.A(n_47),
.B(n_1),
.CON(n_105),
.SN(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_18),
.Y(n_107)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_18),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

BUFx10_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_53),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_119),
.B(n_128),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_127),
.B(n_134),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_53),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_68),
.B(n_25),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g205 ( 
.A1(n_129),
.A2(n_174),
.B(n_45),
.Y(n_205)
);

CKINVDCx9p33_ASAP7_75t_R g131 ( 
.A(n_94),
.Y(n_131)
);

CKINVDCx9p33_ASAP7_75t_R g208 ( 
.A(n_131),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_54),
.A2(n_51),
.B1(n_49),
.B2(n_31),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_135),
.A2(n_101),
.B1(n_96),
.B2(n_82),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_76),
.A2(n_47),
.B1(n_26),
.B2(n_20),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_145),
.A2(n_32),
.B(n_38),
.Y(n_210)
);

OR2x2_ASAP7_75t_SL g193 ( 
.A(n_146),
.B(n_42),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_104),
.B(n_20),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_156),
.B(n_169),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_110),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_104),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_171),
.B(n_175),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_92),
.Y(n_173)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_95),
.B(n_24),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_63),
.B(n_24),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_27),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_176),
.B(n_178),
.Y(n_245)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_177),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_40),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_117),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_179),
.B(n_180),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_40),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_40),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_181),
.B(n_192),
.Y(n_258)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_136),
.Y(n_183)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_183),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_139),
.A2(n_87),
.B1(n_62),
.B2(n_70),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_185),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_187),
.A2(n_200),
.B1(n_78),
.B2(n_57),
.Y(n_240)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_188),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_136),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_189),
.B(n_193),
.Y(n_238)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_190),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_191),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_118),
.B(n_44),
.Y(n_192)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_133),
.Y(n_194)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_194),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_124),
.Y(n_195)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_195),
.Y(n_259)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_196),
.Y(n_267)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_135),
.Y(n_197)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_197),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_198),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_123),
.A2(n_60),
.B1(n_48),
.B2(n_35),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_199),
.A2(n_207),
.B1(n_212),
.B2(n_214),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_113),
.A2(n_79),
.B1(n_67),
.B2(n_90),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_133),
.Y(n_201)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_201),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_219),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_123),
.A2(n_48),
.B1(n_45),
.B2(n_31),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_121),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_209),
.B(n_215),
.Y(n_268)
);

OA21x2_ASAP7_75t_L g266 ( 
.A1(n_210),
.A2(n_235),
.B(n_29),
.Y(n_266)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_157),
.Y(n_211)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_211),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_130),
.A2(n_49),
.B1(n_29),
.B2(n_19),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_213),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_140),
.A2(n_51),
.B1(n_49),
.B2(n_31),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_157),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_217),
.Y(n_243)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_218),
.B(n_220),
.Y(n_272)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_143),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_132),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_223),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_155),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_222),
.B(n_224),
.Y(n_275)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_149),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_111),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_225),
.A2(n_228),
.B1(n_233),
.B2(n_234),
.Y(n_281)
);

CKINVDCx12_ASAP7_75t_R g226 ( 
.A(n_122),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_226),
.B(n_227),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_143),
.Y(n_227)
);

INVx11_ASAP7_75t_L g228 ( 
.A(n_155),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_230),
.Y(n_256)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_163),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_167),
.A2(n_51),
.B(n_30),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_231),
.A2(n_167),
.B(n_19),
.Y(n_244)
);

XNOR2x1_ASAP7_75t_SL g232 ( 
.A(n_115),
.B(n_32),
.Y(n_232)
);

MAJx2_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_19),
.C(n_30),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_165),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_112),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_116),
.B(n_40),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_111),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_236),
.A2(n_111),
.B1(n_172),
.B2(n_168),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_237),
.B(n_274),
.C(n_284),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_262),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_197),
.A2(n_164),
.B1(n_160),
.B2(n_112),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_L g242 ( 
.A1(n_208),
.A2(n_164),
.B1(n_149),
.B2(n_151),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_244),
.B(n_265),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_210),
.A2(n_160),
.B1(n_81),
.B2(n_158),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_246),
.A2(n_195),
.B1(n_224),
.B2(n_191),
.Y(n_295)
);

OA22x2_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_102),
.B1(n_172),
.B2(n_141),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_253),
.Y(n_314)
);

AOI32xp33_ASAP7_75t_L g255 ( 
.A1(n_232),
.A2(n_141),
.A3(n_148),
.B1(n_154),
.B2(n_38),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g289 ( 
.A1(n_255),
.A2(n_204),
.B(n_203),
.C(n_219),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_193),
.A2(n_158),
.B1(n_152),
.B2(n_151),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_229),
.A2(n_148),
.B(n_165),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_195),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_230),
.A2(n_29),
.B(n_30),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_42),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_206),
.B(n_107),
.C(n_109),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_177),
.A2(n_152),
.B1(n_161),
.B2(n_126),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_276),
.A2(n_280),
.B1(n_183),
.B2(n_189),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_208),
.A2(n_196),
.B1(n_216),
.B2(n_234),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_206),
.B(n_161),
.C(n_103),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_277),
.Y(n_285)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_285),
.Y(n_331)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_277),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_287),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_289),
.B(n_309),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_278),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_290),
.B(n_293),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_291),
.Y(n_339)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_245),
.B(n_268),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_294),
.B(n_297),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_295),
.A2(n_312),
.B1(n_315),
.B2(n_320),
.Y(n_338)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_248),
.Y(n_296)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_296),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_244),
.B(n_182),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_271),
.A2(n_222),
.B1(n_194),
.B2(n_198),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_298),
.A2(n_259),
.B1(n_281),
.B2(n_261),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_299),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_270),
.Y(n_300)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_300),
.Y(n_346)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_270),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_301),
.B(n_303),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_256),
.B(n_213),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_302),
.B(n_313),
.Y(n_337)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_248),
.Y(n_304)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_304),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_249),
.A2(n_188),
.B1(n_185),
.B2(n_183),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_305),
.A2(n_323),
.B1(n_283),
.B2(n_257),
.Y(n_340)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_306),
.Y(n_351)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_273),
.Y(n_308)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_308),
.Y(n_359)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_250),
.Y(n_309)
);

AND2x6_ASAP7_75t_L g310 ( 
.A(n_255),
.B(n_223),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_310),
.B(n_262),
.Y(n_333)
);

INVx13_ASAP7_75t_L g311 ( 
.A(n_257),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_311),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_271),
.A2(n_190),
.B1(n_221),
.B2(n_154),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_256),
.B(n_211),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_264),
.A2(n_246),
.B1(n_249),
.B2(n_284),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_247),
.B(n_201),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_318),
.Y(n_348)
);

INVx2_ASAP7_75t_R g318 ( 
.A(n_266),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_247),
.B(n_217),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_259),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_253),
.A2(n_72),
.B1(n_125),
.B2(n_228),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_252),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_321),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_247),
.B(n_218),
.C(n_215),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_274),
.C(n_265),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_254),
.A2(n_202),
.B1(n_225),
.B2(n_125),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_266),
.B(n_251),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_324),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_326),
.B(n_332),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_288),
.A2(n_253),
.B(n_272),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_329),
.A2(n_335),
.B(n_312),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_314),
.A2(n_253),
.B1(n_238),
.B2(n_269),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_330),
.A2(n_344),
.B1(n_345),
.B2(n_354),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_238),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_303),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_288),
.A2(n_238),
.B(n_252),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_340),
.A2(n_286),
.B1(n_317),
.B2(n_285),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_294),
.B(n_258),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_341),
.B(n_307),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_315),
.A2(n_240),
.B1(n_242),
.B2(n_252),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_343),
.A2(n_356),
.B1(n_317),
.B2(n_299),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_297),
.A2(n_237),
.B1(n_275),
.B2(n_267),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_352),
.B(n_292),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_318),
.A2(n_267),
.B1(n_283),
.B2(n_243),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_318),
.A2(n_243),
.B1(n_263),
.B2(n_279),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_313),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_357),
.B(n_302),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_360),
.B(n_366),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_361),
.Y(n_405)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_328),
.Y(n_362)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_362),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_348),
.A2(n_319),
.B(n_316),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_363),
.A2(n_368),
.B(n_327),
.Y(n_412)
);

AND2x6_ASAP7_75t_L g364 ( 
.A(n_333),
.B(n_310),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_364),
.A2(n_388),
.B(n_389),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_365),
.A2(n_384),
.B1(n_354),
.B2(n_344),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_330),
.B(n_356),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_367),
.B(n_338),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_348),
.A2(n_322),
.B(n_289),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_331),
.Y(n_369)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_369),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_342),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_371),
.B(n_372),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_263),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_328),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_373),
.B(n_377),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_334),
.A2(n_320),
.B1(n_295),
.B2(n_286),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_374),
.A2(n_338),
.B1(n_343),
.B2(n_339),
.Y(n_413)
);

OR2x2_ASAP7_75t_SL g375 ( 
.A(n_335),
.B(n_287),
.Y(n_375)
);

AOI21xp33_ASAP7_75t_L g406 ( 
.A1(n_375),
.A2(n_345),
.B(n_327),
.Y(n_406)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_336),
.Y(n_376)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_376),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_353),
.B(n_301),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_346),
.Y(n_378)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_378),
.Y(n_411)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_350),
.Y(n_379)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_379),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_380),
.B(n_383),
.Y(n_393)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_346),
.Y(n_381)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_381),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_342),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_382),
.B(n_390),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_309),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_336),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_385),
.B(n_386),
.Y(n_397)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_387),
.B(n_391),
.Y(n_410)
);

AND2x6_ASAP7_75t_L g389 ( 
.A(n_349),
.B(n_311),
.Y(n_389)
);

INVx6_ASAP7_75t_L g390 ( 
.A(n_331),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_359),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_388),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_394),
.B(n_402),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_395),
.A2(n_355),
.B1(n_369),
.B2(n_390),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_367),
.A2(n_329),
.B(n_349),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_396),
.A2(n_422),
.B(n_125),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_332),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_401),
.B(n_414),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_383),
.B(n_347),
.Y(n_402)
);

AND2x2_ASAP7_75t_SL g450 ( 
.A(n_406),
.B(n_1),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_408),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_412),
.B(n_254),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_413),
.A2(n_387),
.B1(n_379),
.B2(n_355),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_326),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_361),
.B(n_357),
.Y(n_416)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_416),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_368),
.B(n_363),
.C(n_375),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_418),
.B(n_365),
.C(n_376),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_370),
.B(n_341),
.Y(n_420)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_420),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_380),
.B(n_337),
.Y(n_421)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_421),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_367),
.A2(n_347),
.B(n_358),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_370),
.B(n_352),
.Y(n_423)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_423),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_399),
.B(n_358),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_425),
.B(n_432),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_405),
.A2(n_374),
.B1(n_389),
.B2(n_364),
.Y(n_426)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_426),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_427),
.B(n_437),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_405),
.A2(n_325),
.B1(n_386),
.B2(n_385),
.Y(n_428)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_428),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_414),
.B(n_325),
.C(n_391),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_429),
.B(n_433),
.C(n_440),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_430),
.A2(n_431),
.B1(n_439),
.B2(n_441),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_419),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_351),
.C(n_359),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_407),
.B(n_308),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_434),
.B(n_435),
.Y(n_473)
);

FAx1_ASAP7_75t_SL g435 ( 
.A(n_416),
.B(n_306),
.CI(n_296),
.CON(n_435),
.SN(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_400),
.B(n_304),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_436),
.B(n_448),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_413),
.A2(n_260),
.B1(n_279),
.B2(n_282),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_418),
.B(n_282),
.C(n_202),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_408),
.A2(n_260),
.B1(n_126),
.B2(n_120),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_412),
.B(n_120),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_445),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_395),
.A2(n_12),
.B1(n_11),
.B2(n_44),
.Y(n_444)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_444),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_408),
.A2(n_11),
.B1(n_2),
.B2(n_4),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_450),
.B(n_422),
.Y(n_456)
);

INVxp33_ASAP7_75t_L g452 ( 
.A(n_446),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_452),
.B(n_456),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_402),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_454),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_447),
.B(n_438),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_424),
.B(n_409),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_466),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_424),
.B(n_409),
.C(n_394),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_463),
.B(n_464),
.C(n_462),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_433),
.B(n_396),
.C(n_423),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_393),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_437),
.B(n_393),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_467),
.B(n_468),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_440),
.B(n_397),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_449),
.B(n_421),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_469),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_450),
.B(n_397),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_472),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_442),
.B(n_410),
.Y(n_472)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_473),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_481),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_489),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_463),
.A2(n_445),
.B(n_443),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_479),
.A2(n_404),
.B1(n_441),
.B2(n_411),
.Y(n_505)
);

BUFx12f_ASAP7_75t_SL g480 ( 
.A(n_452),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_472),
.Y(n_497)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_458),
.Y(n_481)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_470),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_491),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_457),
.A2(n_451),
.B1(n_448),
.B2(n_430),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_484),
.A2(n_459),
.B1(n_431),
.B2(n_465),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_460),
.B(n_435),
.C(n_443),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_485),
.B(n_417),
.C(n_411),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_460),
.B(n_450),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_487),
.B(n_462),
.Y(n_494)
);

OAI21xp33_ASAP7_75t_L g489 ( 
.A1(n_465),
.A2(n_435),
.B(n_404),
.Y(n_489)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_461),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_474),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_492),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_494),
.B(n_502),
.Y(n_516)
);

CKINVDCx14_ASAP7_75t_R g518 ( 
.A(n_497),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_487),
.B(n_466),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_499),
.B(n_500),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_478),
.B(n_464),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_489),
.B(n_467),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_501),
.B(n_507),
.C(n_476),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_477),
.B(n_455),
.C(n_439),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_503),
.B(n_504),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_410),
.C(n_415),
.Y(n_504)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_505),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_482),
.B(n_417),
.Y(n_506)
);

BUFx24_ASAP7_75t_SL g511 ( 
.A(n_506),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_480),
.Y(n_508)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_508),
.Y(n_517)
);

AOI21xp33_ASAP7_75t_L g510 ( 
.A1(n_495),
.A2(n_488),
.B(n_490),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_510),
.A2(n_514),
.B(n_512),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_512),
.B(n_493),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_476),
.C(n_482),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_513),
.B(n_515),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_493),
.B(n_486),
.C(n_415),
.Y(n_515)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_508),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_519),
.B(n_521),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_498),
.A2(n_398),
.B1(n_486),
.B2(n_403),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_496),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_522),
.B(n_398),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_516),
.B(n_513),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_523),
.B(n_525),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_527),
.B(n_531),
.Y(n_538)
);

AOI21x1_ASAP7_75t_SL g528 ( 
.A1(n_518),
.A2(n_497),
.B(n_501),
.Y(n_528)
);

NAND3xp33_ASAP7_75t_SL g537 ( 
.A(n_528),
.B(n_529),
.C(n_530),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_517),
.A2(n_496),
.B(n_403),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_520),
.B(n_44),
.C(n_5),
.Y(n_531)
);

INVxp33_ASAP7_75t_L g532 ( 
.A(n_509),
.Y(n_532)
);

OAI21xp33_ASAP7_75t_L g533 ( 
.A1(n_532),
.A2(n_511),
.B(n_515),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_533),
.B(n_44),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_526),
.A2(n_516),
.B(n_44),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_535),
.B(n_538),
.C(n_528),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_524),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_536),
.B(n_532),
.Y(n_539)
);

AOI322xp5_ASAP7_75t_L g544 ( 
.A1(n_539),
.A2(n_540),
.A3(n_541),
.B1(n_542),
.B2(n_2),
.C1(n_7),
.C2(n_8),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_537),
.B(n_525),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_542),
.A2(n_534),
.B(n_5),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_543),
.A2(n_544),
.B(n_7),
.Y(n_545)
);

NAND3xp33_ASAP7_75t_L g546 ( 
.A(n_545),
.B(n_7),
.C(n_9),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_546),
.A2(n_7),
.B(n_9),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_9),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_548),
.Y(n_549)
);


endmodule