module fake_netlist_1_1286_n_1124 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_225, n_39, n_1124);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1124;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_963;
wire n_1092;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_667;
wire n_496;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_383;
wire n_288;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_476;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_345;
wire n_360;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_1097;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_955;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1025;
wire n_1011;
wire n_880;
wire n_1101;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_506;
wire n_533;
wire n_490;
wire n_393;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_1000;
wire n_893;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_950;
wire n_910;
wire n_460;
wire n_1046;
wire n_478;
wire n_482;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_1089;
wire n_1058;
wire n_370;
wire n_1050;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_363;
wire n_315;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_912;
wire n_947;
wire n_1043;
wire n_924;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_994;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
wire n_269;
INVx1_ASAP7_75t_L g261 ( .A(n_220), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_6), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_122), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_240), .Y(n_264) );
INVxp33_ASAP7_75t_SL g265 ( .A(n_243), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_141), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_129), .B(n_222), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_15), .Y(n_268) );
INVx1_ASAP7_75t_SL g269 ( .A(n_260), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_160), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_258), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_116), .Y(n_272) );
CKINVDCx16_ASAP7_75t_R g273 ( .A(n_86), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_201), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_72), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_139), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_217), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_177), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_68), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_98), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_249), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_230), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_219), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_114), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g285 ( .A(n_51), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_76), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_175), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_218), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_163), .B(n_107), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_192), .Y(n_290) );
BUFx2_ASAP7_75t_L g291 ( .A(n_44), .Y(n_291) );
NOR2xp67_ASAP7_75t_L g292 ( .A(n_128), .B(n_241), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_191), .Y(n_293) );
BUFx2_ASAP7_75t_L g294 ( .A(n_185), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_209), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_246), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_127), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_242), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_213), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_184), .Y(n_300) );
CKINVDCx20_ASAP7_75t_R g301 ( .A(n_195), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_196), .Y(n_302) );
BUFx10_ASAP7_75t_L g303 ( .A(n_215), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_77), .Y(n_304) );
CKINVDCx14_ASAP7_75t_R g305 ( .A(n_214), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_43), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_138), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_174), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_77), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_148), .Y(n_310) );
INVxp67_ASAP7_75t_L g311 ( .A(n_91), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_247), .Y(n_312) );
NOR2xp67_ASAP7_75t_L g313 ( .A(n_76), .B(n_131), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_169), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_221), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_178), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_118), .Y(n_317) );
CKINVDCx14_ASAP7_75t_R g318 ( .A(n_37), .Y(n_318) );
BUFx2_ASAP7_75t_SL g319 ( .A(n_216), .Y(n_319) );
INVxp67_ASAP7_75t_SL g320 ( .A(n_187), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_159), .Y(n_321) );
CKINVDCx20_ASAP7_75t_R g322 ( .A(n_135), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_223), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_147), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_170), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_37), .Y(n_326) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_182), .Y(n_327) );
CKINVDCx14_ASAP7_75t_R g328 ( .A(n_233), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_154), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_108), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_73), .Y(n_331) );
INVx3_ASAP7_75t_L g332 ( .A(n_144), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_237), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_115), .Y(n_334) );
INVxp67_ASAP7_75t_SL g335 ( .A(n_121), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_68), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_225), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_158), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_29), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_117), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_257), .Y(n_341) );
INVx1_ASAP7_75t_SL g342 ( .A(n_90), .Y(n_342) );
INVx1_ASAP7_75t_SL g343 ( .A(n_227), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_253), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_132), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_17), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_130), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_239), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_80), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_102), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_125), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_134), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_84), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_229), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_149), .Y(n_355) );
CKINVDCx16_ASAP7_75t_R g356 ( .A(n_207), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_124), .Y(n_357) );
CKINVDCx14_ASAP7_75t_R g358 ( .A(n_48), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_20), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_5), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_231), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_78), .Y(n_362) );
INVxp67_ASAP7_75t_L g363 ( .A(n_259), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_224), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_232), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_101), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_165), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_137), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_51), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_126), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_226), .Y(n_371) );
CKINVDCx20_ASAP7_75t_R g372 ( .A(n_146), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_69), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_156), .Y(n_374) );
BUFx10_ASAP7_75t_L g375 ( .A(n_142), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_4), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_244), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_53), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_50), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_143), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_133), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_48), .Y(n_382) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_189), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_18), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_25), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_136), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_250), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_86), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_254), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_120), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_183), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_248), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_145), .Y(n_393) );
INVxp67_ASAP7_75t_L g394 ( .A(n_78), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_236), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_55), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_59), .Y(n_397) );
INVxp67_ASAP7_75t_L g398 ( .A(n_152), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_123), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_59), .Y(n_400) );
INVx1_ASAP7_75t_SL g401 ( .A(n_61), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_23), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_212), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_171), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_155), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_119), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_45), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_45), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_66), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_34), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_318), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_333), .Y(n_412) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_333), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_287), .B(n_0), .Y(n_414) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_333), .Y(n_415) );
BUFx2_ASAP7_75t_L g416 ( .A(n_318), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_307), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_303), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_333), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_336), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_379), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_379), .Y(n_422) );
OAI22x1_ASAP7_75t_SL g423 ( .A1(n_285), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_294), .B(n_1), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_388), .Y(n_425) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_345), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_291), .Y(n_427) );
BUFx3_ASAP7_75t_L g428 ( .A(n_307), .Y(n_428) );
NAND2xp33_ASAP7_75t_L g429 ( .A(n_277), .B(n_109), .Y(n_429) );
OA21x2_ASAP7_75t_L g430 ( .A1(n_344), .A2(n_111), .B(n_110), .Y(n_430) );
BUFx8_ASAP7_75t_L g431 ( .A(n_314), .Y(n_431) );
BUFx2_ASAP7_75t_L g432 ( .A(n_358), .Y(n_432) );
BUFx2_ASAP7_75t_L g433 ( .A(n_358), .Y(n_433) );
OA21x2_ASAP7_75t_L g434 ( .A1(n_344), .A2(n_113), .B(n_112), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_388), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_282), .Y(n_436) );
INVx3_ASAP7_75t_L g437 ( .A(n_303), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_307), .B(n_2), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_261), .Y(n_439) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_345), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_332), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_303), .Y(n_442) );
INVx5_ASAP7_75t_L g443 ( .A(n_332), .Y(n_443) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_345), .Y(n_444) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_345), .Y(n_445) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_383), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_263), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_264), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_266), .Y(n_449) );
BUFx2_ASAP7_75t_L g450 ( .A(n_280), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_273), .B(n_4), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_270), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_438), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_436), .B(n_356), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_418), .B(n_297), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_438), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_418), .B(n_341), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_438), .A2(n_268), .B1(n_279), .B2(n_262), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_431), .Y(n_459) );
BUFx10_ASAP7_75t_L g460 ( .A(n_438), .Y(n_460) );
AND2x6_ASAP7_75t_L g461 ( .A(n_428), .B(n_332), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_439), .B(n_348), .Y(n_462) );
INVxp67_ASAP7_75t_SL g463 ( .A(n_411), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_450), .A2(n_265), .B1(n_397), .B2(n_280), .Y(n_464) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_412), .Y(n_465) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_412), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_439), .B(n_348), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_436), .B(n_404), .Y(n_468) );
BUFx2_ASAP7_75t_L g469 ( .A(n_411), .Y(n_469) );
BUFx4f_ASAP7_75t_L g470 ( .A(n_416), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_428), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_418), .B(n_397), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_437), .B(n_409), .Y(n_473) );
BUFx10_ASAP7_75t_L g474 ( .A(n_427), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_417), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_431), .Y(n_476) );
NAND2xp33_ASAP7_75t_L g477 ( .A(n_443), .B(n_383), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_432), .B(n_305), .Y(n_478) );
INVx8_ASAP7_75t_L g479 ( .A(n_437), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_432), .B(n_305), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_437), .B(n_409), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_447), .B(n_365), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_437), .B(n_410), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_447), .A2(n_286), .B1(n_306), .B2(n_304), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_417), .Y(n_485) );
AND2x6_ASAP7_75t_L g486 ( .A(n_441), .B(n_299), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_442), .B(n_363), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_448), .B(n_365), .Y(n_488) );
INVxp33_ASAP7_75t_L g489 ( .A(n_433), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_433), .A2(n_322), .B1(n_327), .B2(n_301), .Y(n_490) );
BUFx2_ASAP7_75t_L g491 ( .A(n_450), .Y(n_491) );
BUFx6f_ASAP7_75t_SL g492 ( .A(n_449), .Y(n_492) );
OR2x6_ASAP7_75t_L g493 ( .A(n_451), .B(n_319), .Y(n_493) );
OAI21xp33_ASAP7_75t_SL g494 ( .A1(n_449), .A2(n_339), .B(n_326), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_460), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_468), .B(n_442), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_489), .B(n_442), .Y(n_497) );
NAND2x1p5_ASAP7_75t_L g498 ( .A(n_470), .B(n_349), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_453), .B(n_452), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_456), .B(n_455), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_490), .B(n_454), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_475), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_456), .B(n_452), .Y(n_503) );
INVx8_ASAP7_75t_L g504 ( .A(n_479), .Y(n_504) );
NOR3xp33_ASAP7_75t_L g505 ( .A(n_494), .B(n_424), .C(n_414), .Y(n_505) );
NAND2xp33_ASAP7_75t_L g506 ( .A(n_461), .B(n_443), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_469), .B(n_414), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_485), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_455), .B(n_424), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_457), .B(n_443), .Y(n_510) );
AOI221xp5_ASAP7_75t_L g511 ( .A1(n_484), .A2(n_423), .B1(n_311), .B2(n_394), .C(n_420), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_474), .B(n_275), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_457), .B(n_443), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_489), .B(n_431), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_461), .B(n_443), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_462), .Y(n_516) );
INVx2_ASAP7_75t_SL g517 ( .A(n_474), .Y(n_517) );
INVx2_ASAP7_75t_SL g518 ( .A(n_478), .Y(n_518) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_484), .A2(n_423), .B1(n_421), .B2(n_422), .C(n_420), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_463), .Y(n_520) );
AND2x6_ASAP7_75t_L g521 ( .A(n_480), .B(n_441), .Y(n_521) );
NAND2x1_ASAP7_75t_L g522 ( .A(n_461), .B(n_430), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_461), .B(n_443), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_462), .Y(n_524) );
BUFx6f_ASAP7_75t_SL g525 ( .A(n_493), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_461), .B(n_429), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_458), .B(n_281), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_464), .B(n_342), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_493), .A2(n_322), .B1(n_327), .B2(n_301), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_472), .B(n_398), .Y(n_530) );
BUFx3_ASAP7_75t_L g531 ( .A(n_459), .Y(n_531) );
NAND2xp33_ASAP7_75t_SL g532 ( .A(n_492), .B(n_330), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_458), .B(n_281), .Y(n_533) );
INVx2_ASAP7_75t_SL g534 ( .A(n_479), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_473), .B(n_283), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_493), .B(n_401), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_471), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_481), .B(n_483), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_476), .B(n_309), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_479), .B(n_283), .Y(n_540) );
INVxp67_ASAP7_75t_SL g541 ( .A(n_487), .Y(n_541) );
BUFx3_ASAP7_75t_L g542 ( .A(n_486), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_467), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_482), .B(n_393), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_492), .A2(n_330), .B1(n_386), .B2(n_372), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_488), .B(n_393), .Y(n_546) );
INVx2_ASAP7_75t_SL g547 ( .A(n_486), .Y(n_547) );
OR2x6_ASAP7_75t_L g548 ( .A(n_486), .B(n_353), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_477), .A2(n_434), .B(n_430), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_477), .A2(n_328), .B1(n_373), .B2(n_359), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_465), .B(n_406), .Y(n_551) );
INVx3_ASAP7_75t_L g552 ( .A(n_465), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_466), .B(n_350), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_466), .A2(n_386), .B1(n_399), .B2(n_372), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_489), .B(n_375), .Y(n_555) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_461), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_454), .A2(n_399), .B1(n_366), .B2(n_384), .Y(n_557) );
INVxp33_ASAP7_75t_L g558 ( .A(n_491), .Y(n_558) );
AND2x6_ASAP7_75t_SL g559 ( .A(n_493), .B(n_376), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_468), .B(n_328), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_460), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_491), .Y(n_562) );
INVx8_ASAP7_75t_L g563 ( .A(n_479), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_468), .B(n_320), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_456), .A2(n_378), .B1(n_396), .B2(n_382), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_474), .B(n_360), .Y(n_566) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_461), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_456), .A2(n_400), .B1(n_407), .B2(n_402), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_454), .A2(n_385), .B1(n_408), .B2(n_346), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_503), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_522), .A2(n_434), .B(n_430), .Y(n_571) );
AO22x1_ASAP7_75t_L g572 ( .A1(n_545), .A2(n_285), .B1(n_362), .B2(n_346), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_509), .B(n_425), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_503), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_500), .A2(n_434), .B(n_430), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_500), .A2(n_513), .B(n_510), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_507), .B(n_362), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_558), .B(n_369), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_510), .A2(n_434), .B(n_430), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_504), .A2(n_369), .B1(n_335), .B2(n_425), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_501), .B(n_375), .Y(n_581) );
A2O1A1Ixp33_ASAP7_75t_L g582 ( .A1(n_538), .A2(n_313), .B(n_435), .C(n_272), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_513), .A2(n_434), .B(n_274), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_504), .A2(n_435), .B1(n_331), .B2(n_271), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_549), .A2(n_278), .B(n_276), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_509), .B(n_375), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_499), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_499), .A2(n_288), .B(n_284), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_508), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_517), .Y(n_590) );
A2O1A1Ixp33_ASAP7_75t_L g591 ( .A1(n_541), .A2(n_293), .B(n_296), .C(n_295), .Y(n_591) );
BUFx2_ASAP7_75t_L g592 ( .A(n_562), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_526), .A2(n_308), .B(n_298), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_514), .B(n_269), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_496), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_520), .B(n_316), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_504), .B(n_290), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_526), .A2(n_312), .B(n_310), .Y(n_598) );
O2A1O1Ixp33_ASAP7_75t_L g599 ( .A1(n_505), .A2(n_321), .B(n_323), .C(n_315), .Y(n_599) );
OAI21xp33_ASAP7_75t_L g600 ( .A1(n_569), .A2(n_302), .B(n_300), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_563), .A2(n_331), .B1(n_337), .B2(n_334), .Y(n_601) );
AOI21x1_ASAP7_75t_L g602 ( .A1(n_515), .A2(n_292), .B(n_338), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_521), .A2(n_331), .B1(n_347), .B2(n_340), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_560), .A2(n_354), .B(n_352), .Y(n_604) );
BUFx3_ASAP7_75t_L g605 ( .A(n_563), .Y(n_605) );
INVx3_ASAP7_75t_L g606 ( .A(n_563), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_515), .A2(n_361), .B(n_355), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_534), .B(n_317), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_523), .A2(n_370), .B(n_368), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_516), .A2(n_377), .B(n_374), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_524), .A2(n_381), .B(n_380), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_518), .B(n_343), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_498), .B(n_324), .Y(n_613) );
AO22x1_ASAP7_75t_L g614 ( .A1(n_531), .A2(n_329), .B1(n_351), .B2(n_325), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_543), .A2(n_390), .B(n_389), .Y(n_615) );
A2O1A1Ixp33_ASAP7_75t_L g616 ( .A1(n_530), .A2(n_392), .B(n_395), .C(n_391), .Y(n_616) );
INVx4_ASAP7_75t_L g617 ( .A(n_556), .Y(n_617) );
NOR2xp33_ASAP7_75t_SL g618 ( .A(n_567), .B(n_357), .Y(n_618) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_512), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_551), .A2(n_405), .B(n_403), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_566), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_551), .A2(n_267), .B(n_289), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_498), .B(n_364), .Y(n_623) );
NOR2xp33_ASAP7_75t_SL g624 ( .A(n_567), .B(n_367), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_536), .B(n_371), .Y(n_625) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_567), .Y(n_626) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_542), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_539), .B(n_387), .Y(n_628) );
AND2x2_ASAP7_75t_SL g629 ( .A(n_519), .B(n_383), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_537), .A2(n_446), .B(n_413), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_511), .A2(n_440), .B1(n_445), .B2(n_444), .C(n_426), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_564), .B(n_6), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_497), .A2(n_440), .B1(n_413), .B2(n_415), .Y(n_633) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_535), .A2(n_413), .B(n_415), .C(n_412), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_495), .A2(n_413), .B(n_412), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_527), .B(n_7), .Y(n_636) );
AO21x1_ASAP7_75t_L g637 ( .A1(n_506), .A2(n_553), .B(n_533), .Y(n_637) );
INVx3_ASAP7_75t_L g638 ( .A(n_561), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_527), .B(n_7), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_533), .A2(n_440), .B1(n_446), .B2(n_413), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_557), .B(n_8), .Y(n_641) );
NOR3xp33_ASAP7_75t_L g642 ( .A(n_532), .B(n_8), .C(n_9), .Y(n_642) );
NAND3xp33_ASAP7_75t_L g643 ( .A(n_565), .B(n_568), .C(n_550), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_540), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_540), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_528), .B(n_555), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_544), .B(n_10), .Y(n_647) );
BUFx2_ASAP7_75t_L g648 ( .A(n_559), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_525), .B(n_10), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_546), .B(n_11), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_547), .B(n_11), .Y(n_651) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_548), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_548), .B(n_12), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_552), .B(n_12), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_509), .B(n_13), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_504), .A2(n_426), .B1(n_444), .B2(n_419), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_504), .B(n_419), .Y(n_657) );
AND2x2_ASAP7_75t_SL g658 ( .A(n_554), .B(n_14), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_502), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_502), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_509), .B(n_16), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_509), .B(n_17), .Y(n_662) );
NOR2xp33_ASAP7_75t_SL g663 ( .A(n_504), .B(n_426), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_558), .B(n_18), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_509), .B(n_19), .Y(n_665) );
AO32x2_ASAP7_75t_L g666 ( .A1(n_547), .A2(n_445), .A3(n_444), .B1(n_446), .B2(n_22), .Y(n_666) );
AO21x1_ASAP7_75t_L g667 ( .A1(n_522), .A2(n_446), .B(n_445), .Y(n_667) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_522), .A2(n_445), .B(n_444), .Y(n_668) );
BUFx8_ASAP7_75t_L g669 ( .A(n_525), .Y(n_669) );
AOI22x1_ASAP7_75t_L g670 ( .A1(n_549), .A2(n_445), .B1(n_446), .B2(n_444), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_545), .B(n_21), .C(n_22), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_522), .A2(n_446), .B(n_445), .Y(n_672) );
O2A1O1Ixp33_ASAP7_75t_L g673 ( .A1(n_509), .A2(n_26), .B(n_24), .C(n_25), .Y(n_673) );
OR2x6_ASAP7_75t_L g674 ( .A(n_504), .B(n_24), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_629), .A2(n_28), .B1(n_26), .B2(n_27), .Y(n_675) );
O2A1O1Ixp33_ASAP7_75t_L g676 ( .A1(n_616), .A2(n_29), .B(n_27), .C(n_28), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_595), .B(n_30), .Y(n_677) );
INVx2_ASAP7_75t_SL g678 ( .A(n_605), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_587), .B(n_30), .Y(n_679) );
A2O1A1Ixp33_ASAP7_75t_L g680 ( .A1(n_599), .A2(n_33), .B(n_31), .C(n_32), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_589), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_577), .B(n_592), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_570), .B(n_32), .Y(n_683) );
AO31x2_ASAP7_75t_L g684 ( .A1(n_667), .A2(n_585), .A3(n_637), .B(n_583), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_621), .B(n_35), .Y(n_685) );
AOI21xp33_ASAP7_75t_L g686 ( .A1(n_628), .A2(n_36), .B(n_38), .Y(n_686) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_674), .Y(n_687) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_626), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_573), .Y(n_689) );
INVx1_ASAP7_75t_SL g690 ( .A(n_674), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_574), .B(n_39), .Y(n_691) );
AO32x2_ASAP7_75t_L g692 ( .A1(n_640), .A2(n_40), .A3(n_41), .B1(n_42), .B2(n_43), .Y(n_692) );
O2A1O1Ixp33_ASAP7_75t_L g693 ( .A1(n_591), .A2(n_40), .B(n_42), .C(n_44), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_646), .B(n_46), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_576), .A2(n_672), .B(n_668), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g696 ( .A1(n_604), .A2(n_46), .B(n_47), .C(n_49), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_644), .B(n_47), .Y(n_697) );
OR2x6_ASAP7_75t_L g698 ( .A(n_674), .B(n_49), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_659), .Y(n_699) );
O2A1O1Ixp33_ASAP7_75t_SL g700 ( .A1(n_634), .A2(n_157), .B(n_256), .C(n_255), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_655), .Y(n_701) );
A2O1A1Ixp33_ASAP7_75t_L g702 ( .A1(n_581), .A2(n_52), .B(n_53), .C(n_54), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_578), .B(n_54), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_645), .B(n_55), .Y(n_704) );
NAND2x1p5_ASAP7_75t_L g705 ( .A(n_606), .B(n_56), .Y(n_705) );
A2O1A1Ixp33_ASAP7_75t_L g706 ( .A1(n_593), .A2(n_57), .B(n_58), .C(n_60), .Y(n_706) );
BUFx6f_ASAP7_75t_L g707 ( .A(n_626), .Y(n_707) );
BUFx8_ASAP7_75t_L g708 ( .A(n_648), .Y(n_708) );
INVx3_ASAP7_75t_SL g709 ( .A(n_590), .Y(n_709) );
NOR2xp67_ASAP7_75t_SL g710 ( .A(n_606), .B(n_57), .Y(n_710) );
AO31x2_ASAP7_75t_L g711 ( .A1(n_582), .A2(n_58), .A3(n_61), .B(n_62), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_586), .B(n_62), .Y(n_712) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_598), .A2(n_63), .B(n_64), .C(n_65), .Y(n_713) );
AO31x2_ASAP7_75t_L g714 ( .A1(n_636), .A2(n_63), .A3(n_64), .B(n_65), .Y(n_714) );
AND2x4_ASAP7_75t_L g715 ( .A(n_638), .B(n_66), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_643), .B(n_67), .Y(n_716) );
BUFx8_ASAP7_75t_L g717 ( .A(n_652), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_643), .B(n_67), .Y(n_718) );
AO32x2_ASAP7_75t_L g719 ( .A1(n_584), .A2(n_69), .A3(n_70), .B1(n_71), .B2(n_72), .Y(n_719) );
INVxp67_ASAP7_75t_L g720 ( .A(n_619), .Y(n_720) );
AO31x2_ASAP7_75t_L g721 ( .A1(n_639), .A2(n_71), .A3(n_73), .B(n_74), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_661), .A2(n_74), .B1(n_75), .B2(n_79), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_662), .Y(n_723) );
BUFx12f_ASAP7_75t_L g724 ( .A(n_669), .Y(n_724) );
A2O1A1Ixp33_ASAP7_75t_L g725 ( .A1(n_620), .A2(n_79), .B(n_80), .C(n_81), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_660), .Y(n_726) );
O2A1O1Ixp33_ASAP7_75t_SL g727 ( .A1(n_665), .A2(n_179), .B(n_252), .C(n_251), .Y(n_727) );
INVx3_ASAP7_75t_L g728 ( .A(n_617), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_641), .B(n_81), .Y(n_729) );
OAI21xp5_ASAP7_75t_L g730 ( .A1(n_588), .A2(n_176), .B(n_245), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_658), .A2(n_82), .B1(n_83), .B2(n_84), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_580), .B(n_82), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_632), .Y(n_733) );
A2O1A1Ixp33_ASAP7_75t_L g734 ( .A1(n_607), .A2(n_85), .B(n_87), .C(n_88), .Y(n_734) );
NOR2x1_ASAP7_75t_SL g735 ( .A(n_626), .B(n_89), .Y(n_735) );
AO32x2_ASAP7_75t_L g736 ( .A1(n_601), .A2(n_90), .A3(n_91), .B1(n_92), .B2(n_93), .Y(n_736) );
AO21x1_ASAP7_75t_L g737 ( .A1(n_673), .A2(n_181), .B(n_238), .Y(n_737) );
A2O1A1Ixp33_ASAP7_75t_L g738 ( .A1(n_609), .A2(n_92), .B(n_93), .C(n_94), .Y(n_738) );
OAI21x1_ASAP7_75t_L g739 ( .A1(n_630), .A2(n_602), .B(n_635), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_603), .A2(n_95), .B1(n_96), .B2(n_97), .Y(n_740) );
O2A1O1Ixp5_ASAP7_75t_L g741 ( .A1(n_622), .A2(n_180), .B(n_235), .C(n_234), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_594), .A2(n_95), .B1(n_96), .B2(n_97), .Y(n_742) );
BUFx12f_ASAP7_75t_L g743 ( .A(n_669), .Y(n_743) );
NOR2x1_ASAP7_75t_L g744 ( .A(n_597), .B(n_98), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g745 ( .A1(n_610), .A2(n_173), .B(n_228), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g746 ( .A1(n_611), .A2(n_99), .B(n_100), .C(n_101), .Y(n_746) );
BUFx12f_ASAP7_75t_L g747 ( .A(n_627), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_596), .B(n_103), .Y(n_748) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_653), .Y(n_749) );
INVx4_ASAP7_75t_L g750 ( .A(n_617), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_625), .B(n_104), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_613), .B(n_104), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_647), .Y(n_753) );
INVx1_ASAP7_75t_SL g754 ( .A(n_650), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_623), .B(n_105), .Y(n_755) );
INVx2_ASAP7_75t_SL g756 ( .A(n_614), .Y(n_756) );
AOI221x1_ASAP7_75t_L g757 ( .A1(n_671), .A2(n_105), .B1(n_106), .B2(n_107), .C(n_140), .Y(n_757) );
NOR2x1_ASAP7_75t_L g758 ( .A(n_649), .B(n_106), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_642), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_666), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_654), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_664), .Y(n_762) );
AO31x2_ASAP7_75t_L g763 ( .A1(n_651), .A2(n_150), .A3(n_151), .B(n_153), .Y(n_763) );
AND2x4_ASAP7_75t_L g764 ( .A(n_608), .B(n_161), .Y(n_764) );
AO31x2_ASAP7_75t_L g765 ( .A1(n_656), .A2(n_162), .A3(n_164), .B(n_166), .Y(n_765) );
NOR3xp33_ASAP7_75t_L g766 ( .A(n_600), .B(n_167), .C(n_168), .Y(n_766) );
AOI21xp5_ASAP7_75t_SL g767 ( .A1(n_663), .A2(n_172), .B(n_186), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_615), .Y(n_768) );
AOI31xp67_ASAP7_75t_L g769 ( .A1(n_633), .A2(n_188), .A3(n_190), .B(n_193), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_666), .Y(n_770) );
INVx2_ASAP7_75t_SL g771 ( .A(n_657), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g772 ( .A1(n_663), .A2(n_194), .B(n_197), .Y(n_772) );
OA21x2_ASAP7_75t_L g773 ( .A1(n_631), .A2(n_198), .B(n_199), .Y(n_773) );
AO31x2_ASAP7_75t_L g774 ( .A1(n_666), .A2(n_200), .A3(n_202), .B(n_203), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_612), .Y(n_775) );
AO31x2_ASAP7_75t_L g776 ( .A1(n_618), .A2(n_204), .A3(n_205), .B(n_206), .Y(n_776) );
AO31x2_ASAP7_75t_L g777 ( .A1(n_618), .A2(n_208), .A3(n_210), .B(n_211), .Y(n_777) );
BUFx3_ASAP7_75t_L g778 ( .A(n_624), .Y(n_778) );
INVx1_ASAP7_75t_SL g779 ( .A(n_592), .Y(n_779) );
OAI21x1_ASAP7_75t_L g780 ( .A1(n_670), .A2(n_571), .B(n_672), .Y(n_780) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_592), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_589), .Y(n_782) );
NAND2x1p5_ASAP7_75t_L g783 ( .A(n_605), .B(n_606), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_621), .B(n_558), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_575), .A2(n_579), .B(n_571), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_595), .B(n_509), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_575), .A2(n_579), .B(n_571), .Y(n_787) );
O2A1O1Ixp33_ASAP7_75t_L g788 ( .A1(n_616), .A2(n_591), .B(n_599), .C(n_501), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_689), .B(n_786), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_698), .B(n_779), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_782), .Y(n_791) );
INVx3_ASAP7_75t_L g792 ( .A(n_717), .Y(n_792) );
AOI21xp5_ASAP7_75t_SL g793 ( .A1(n_675), .A2(n_778), .B(n_715), .Y(n_793) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_781), .Y(n_794) );
AO21x2_ASAP7_75t_L g795 ( .A1(n_760), .A2(n_770), .B(n_718), .Y(n_795) );
OR2x2_ASAP7_75t_L g796 ( .A(n_720), .B(n_709), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g797 ( .A1(n_701), .A2(n_723), .B(n_788), .Y(n_797) );
OR2x2_ASAP7_75t_L g798 ( .A(n_784), .B(n_690), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_733), .B(n_753), .Y(n_799) );
OA21x2_ASAP7_75t_L g800 ( .A1(n_739), .A2(n_741), .B(n_737), .Y(n_800) );
BUFx8_ASAP7_75t_L g801 ( .A(n_724), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_679), .Y(n_802) );
INVx3_ASAP7_75t_L g803 ( .A(n_747), .Y(n_803) );
AND2x2_ASAP7_75t_L g804 ( .A(n_775), .B(n_687), .Y(n_804) );
INVx3_ASAP7_75t_L g805 ( .A(n_750), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_759), .B(n_768), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g807 ( .A1(n_761), .A2(n_712), .B(n_751), .Y(n_807) );
OAI221xp5_ASAP7_75t_L g808 ( .A1(n_731), .A2(n_732), .B1(n_729), .B2(n_703), .C(n_694), .Y(n_808) );
OAI21x1_ASAP7_75t_SL g809 ( .A1(n_735), .A2(n_756), .B(n_772), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_715), .A2(n_705), .B1(n_691), .B2(n_683), .Y(n_810) );
OA21x2_ASAP7_75t_L g811 ( .A1(n_730), .A2(n_757), .B(n_745), .Y(n_811) );
INVx4_ASAP7_75t_SL g812 ( .A(n_776), .Y(n_812) );
AND2x4_ASAP7_75t_L g813 ( .A(n_750), .B(n_764), .Y(n_813) );
AOI21xp5_ASAP7_75t_L g814 ( .A1(n_700), .A2(n_677), .B(n_727), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_699), .B(n_726), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_697), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_762), .B(n_704), .Y(n_817) );
INVx3_ASAP7_75t_L g818 ( .A(n_728), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_749), .B(n_754), .Y(n_819) );
AO31x2_ASAP7_75t_L g820 ( .A1(n_735), .A2(n_713), .A3(n_706), .B(n_680), .Y(n_820) );
AOI21xp5_ASAP7_75t_L g821 ( .A1(n_748), .A2(n_755), .B(n_752), .Y(n_821) );
OAI21x1_ASAP7_75t_SL g822 ( .A1(n_693), .A2(n_773), .B(n_676), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_714), .Y(n_823) );
AOI22xp33_ASAP7_75t_SL g824 ( .A1(n_742), .A2(n_685), .B1(n_764), .B2(n_722), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_714), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_702), .A2(n_696), .B1(n_758), .B2(n_725), .Y(n_826) );
AOI21xp5_ASAP7_75t_L g827 ( .A1(n_767), .A2(n_734), .B(n_738), .Y(n_827) );
OA21x2_ASAP7_75t_L g828 ( .A1(n_766), .A2(n_746), .B(n_686), .Y(n_828) );
AND2x4_ASAP7_75t_L g829 ( .A(n_678), .B(n_728), .Y(n_829) );
OA21x2_ASAP7_75t_L g830 ( .A1(n_684), .A2(n_769), .B(n_774), .Y(n_830) );
BUFx10_ASAP7_75t_L g831 ( .A(n_771), .Y(n_831) );
OR2x2_ASAP7_75t_L g832 ( .A(n_783), .B(n_711), .Y(n_832) );
AO21x2_ASAP7_75t_L g833 ( .A1(n_684), .A2(n_740), .B(n_774), .Y(n_833) );
AOI21xp5_ASAP7_75t_L g834 ( .A1(n_688), .A2(n_707), .B(n_744), .Y(n_834) );
INVxp67_ASAP7_75t_L g835 ( .A(n_710), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_721), .Y(n_836) );
AND2x2_ASAP7_75t_L g837 ( .A(n_736), .B(n_719), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_736), .A2(n_692), .B1(n_719), .B2(n_711), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_763), .A2(n_765), .B(n_692), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_736), .B(n_719), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_692), .B(n_721), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_763), .B(n_765), .Y(n_842) );
OA21x2_ASAP7_75t_L g843 ( .A1(n_777), .A2(n_776), .B(n_708), .Y(n_843) );
AO31x2_ASAP7_75t_L g844 ( .A1(n_776), .A2(n_787), .A3(n_785), .B(n_770), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g845 ( .A(n_777), .B(n_529), .Y(n_845) );
INVx1_ASAP7_75t_SL g846 ( .A(n_777), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_689), .B(n_786), .Y(n_847) );
OA21x2_ASAP7_75t_L g848 ( .A1(n_785), .A2(n_787), .B(n_780), .Y(n_848) );
OAI21xp5_ASAP7_75t_L g849 ( .A1(n_716), .A2(n_576), .B(n_585), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_681), .Y(n_850) );
AOI21xp33_ASAP7_75t_SL g851 ( .A1(n_709), .A2(n_545), .B(n_572), .Y(n_851) );
INVx3_ASAP7_75t_SL g852 ( .A(n_709), .Y(n_852) );
BUFx8_ASAP7_75t_L g853 ( .A(n_724), .Y(n_853) );
AO31x2_ASAP7_75t_L g854 ( .A1(n_785), .A2(n_787), .A3(n_770), .B(n_760), .Y(n_854) );
INVx4_ASAP7_75t_L g855 ( .A(n_724), .Y(n_855) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_715), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_681), .Y(n_857) );
AOI21xp5_ASAP7_75t_L g858 ( .A1(n_785), .A2(n_787), .B(n_695), .Y(n_858) );
BUFx2_ASAP7_75t_L g859 ( .A(n_698), .Y(n_859) );
AO31x2_ASAP7_75t_L g860 ( .A1(n_785), .A2(n_787), .A3(n_770), .B(n_760), .Y(n_860) );
AND2x4_ASAP7_75t_L g861 ( .A(n_689), .B(n_786), .Y(n_861) );
OR3x4_ASAP7_75t_SL g862 ( .A(n_724), .B(n_743), .C(n_423), .Y(n_862) );
CKINVDCx5p33_ASAP7_75t_R g863 ( .A(n_724), .Y(n_863) );
BUFx2_ASAP7_75t_L g864 ( .A(n_698), .Y(n_864) );
OR2x6_ASAP7_75t_L g865 ( .A(n_698), .B(n_674), .Y(n_865) );
AOI21xp5_ASAP7_75t_L g866 ( .A1(n_785), .A2(n_787), .B(n_695), .Y(n_866) );
NOR2xp33_ASAP7_75t_L g867 ( .A(n_749), .B(n_529), .Y(n_867) );
INVx5_ASAP7_75t_L g868 ( .A(n_698), .Y(n_868) );
A2O1A1Ixp33_ASAP7_75t_L g869 ( .A1(n_788), .A2(n_689), .B(n_786), .C(n_629), .Y(n_869) );
AOI21xp5_ASAP7_75t_L g870 ( .A1(n_785), .A2(n_787), .B(n_695), .Y(n_870) );
OA21x2_ASAP7_75t_L g871 ( .A1(n_785), .A2(n_787), .B(n_780), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_698), .A2(n_629), .B1(n_658), .B2(n_646), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_681), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_682), .B(n_577), .Y(n_874) );
NAND2x1p5_ASAP7_75t_L g875 ( .A(n_750), .B(n_605), .Y(n_875) );
BUFx2_ASAP7_75t_L g876 ( .A(n_698), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_681), .Y(n_877) );
OAI221xp5_ASAP7_75t_SL g878 ( .A1(n_698), .A2(n_529), .B1(n_519), .B2(n_731), .C(n_511), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_806), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_806), .Y(n_880) );
INVx2_ASAP7_75t_SL g881 ( .A(n_875), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_823), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_825), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_861), .B(n_789), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_836), .Y(n_885) );
HB1xp67_ASAP7_75t_L g886 ( .A(n_794), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_789), .B(n_847), .Y(n_887) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_847), .Y(n_888) );
OR2x6_ASAP7_75t_L g889 ( .A(n_865), .B(n_793), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_791), .Y(n_890) );
BUFx2_ASAP7_75t_L g891 ( .A(n_865), .Y(n_891) );
INVxp67_ASAP7_75t_L g892 ( .A(n_859), .Y(n_892) );
OR2x6_ASAP7_75t_L g893 ( .A(n_865), .B(n_856), .Y(n_893) );
NAND2x1p5_ASAP7_75t_L g894 ( .A(n_868), .B(n_813), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_850), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_857), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_854), .Y(n_897) );
INVx2_ASAP7_75t_SL g898 ( .A(n_875), .Y(n_898) );
OA21x2_ASAP7_75t_L g899 ( .A1(n_858), .A2(n_870), .B(n_866), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_854), .Y(n_900) );
INVx2_ASAP7_75t_L g901 ( .A(n_854), .Y(n_901) );
INVx2_ASAP7_75t_L g902 ( .A(n_860), .Y(n_902) );
INVx2_ASAP7_75t_L g903 ( .A(n_860), .Y(n_903) );
OR2x2_ASAP7_75t_L g904 ( .A(n_815), .B(n_819), .Y(n_904) );
OR2x2_ASAP7_75t_L g905 ( .A(n_815), .B(n_819), .Y(n_905) );
BUFx2_ASAP7_75t_L g906 ( .A(n_813), .Y(n_906) );
INVx2_ASAP7_75t_L g907 ( .A(n_848), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_874), .B(n_867), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_873), .B(n_877), .Y(n_909) );
BUFx2_ASAP7_75t_SL g910 ( .A(n_868), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_799), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_804), .Y(n_912) );
BUFx2_ASAP7_75t_L g913 ( .A(n_832), .Y(n_913) );
AO21x2_ASAP7_75t_L g914 ( .A1(n_839), .A2(n_842), .B(n_866), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_797), .B(n_802), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_797), .B(n_816), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_817), .B(n_837), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_840), .B(n_841), .Y(n_918) );
HB1xp67_ASAP7_75t_L g919 ( .A(n_868), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_872), .A2(n_824), .B1(n_869), .B2(n_878), .Y(n_920) );
OR2x6_ASAP7_75t_L g921 ( .A(n_864), .B(n_876), .Y(n_921) );
CKINVDCx5p33_ASAP7_75t_R g922 ( .A(n_801), .Y(n_922) );
NOR2x1_ASAP7_75t_L g923 ( .A(n_792), .B(n_805), .Y(n_923) );
AND2x4_ASAP7_75t_L g924 ( .A(n_805), .B(n_818), .Y(n_924) );
AO21x2_ASAP7_75t_L g925 ( .A1(n_839), .A2(n_842), .B(n_858), .Y(n_925) );
INVx4_ASAP7_75t_SL g926 ( .A(n_820), .Y(n_926) );
OAI21xp5_ASAP7_75t_L g927 ( .A1(n_821), .A2(n_807), .B(n_808), .Y(n_927) );
OR2x6_ASAP7_75t_L g928 ( .A(n_810), .B(n_809), .Y(n_928) );
INVx4_ASAP7_75t_L g929 ( .A(n_792), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_829), .Y(n_930) );
OR2x6_ASAP7_75t_L g931 ( .A(n_810), .B(n_834), .Y(n_931) );
AND2x2_ASAP7_75t_L g932 ( .A(n_807), .B(n_845), .Y(n_932) );
INVxp33_ASAP7_75t_L g933 ( .A(n_796), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_831), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_820), .B(n_821), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_851), .B(n_790), .Y(n_936) );
INVx3_ASAP7_75t_L g937 ( .A(n_831), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_838), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_820), .B(n_838), .Y(n_939) );
AO21x2_ASAP7_75t_L g940 ( .A1(n_822), .A2(n_814), .B(n_833), .Y(n_940) );
OR2x2_ASAP7_75t_L g941 ( .A(n_913), .B(n_918), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_882), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_918), .B(n_833), .Y(n_943) );
HB1xp67_ASAP7_75t_L g944 ( .A(n_888), .Y(n_944) );
INVx2_ASAP7_75t_SL g945 ( .A(n_881), .Y(n_945) );
BUFx2_ASAP7_75t_L g946 ( .A(n_913), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_932), .B(n_844), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_882), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_932), .B(n_844), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_917), .B(n_844), .Y(n_950) );
AND2x2_ASAP7_75t_L g951 ( .A(n_917), .B(n_795), .Y(n_951) );
INVx2_ASAP7_75t_L g952 ( .A(n_907), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_939), .B(n_887), .Y(n_953) );
AND2x2_ASAP7_75t_L g954 ( .A(n_939), .B(n_795), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_883), .Y(n_955) );
INVxp67_ASAP7_75t_SL g956 ( .A(n_884), .Y(n_956) );
BUFx3_ASAP7_75t_L g957 ( .A(n_894), .Y(n_957) );
AND2x4_ASAP7_75t_L g958 ( .A(n_926), .B(n_812), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_935), .B(n_871), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_935), .B(n_830), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_938), .B(n_830), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_938), .B(n_843), .Y(n_962) );
BUFx3_ASAP7_75t_L g963 ( .A(n_894), .Y(n_963) );
AND2x2_ASAP7_75t_L g964 ( .A(n_915), .B(n_843), .Y(n_964) );
HB1xp67_ASAP7_75t_L g965 ( .A(n_886), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_885), .Y(n_966) );
AND2x4_ASAP7_75t_SL g967 ( .A(n_889), .B(n_803), .Y(n_967) );
OR2x2_ASAP7_75t_L g968 ( .A(n_904), .B(n_798), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_915), .B(n_846), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_916), .B(n_846), .Y(n_970) );
AND2x2_ASAP7_75t_L g971 ( .A(n_916), .B(n_927), .Y(n_971) );
OR2x2_ASAP7_75t_L g972 ( .A(n_905), .B(n_826), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_879), .B(n_849), .Y(n_973) );
BUFx2_ASAP7_75t_L g974 ( .A(n_928), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_911), .B(n_808), .Y(n_975) );
OR2x2_ASAP7_75t_L g976 ( .A(n_880), .B(n_852), .Y(n_976) );
OR2x2_ASAP7_75t_L g977 ( .A(n_880), .B(n_811), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_909), .B(n_800), .Y(n_978) );
BUFx3_ASAP7_75t_L g979 ( .A(n_894), .Y(n_979) );
OR2x2_ASAP7_75t_L g980 ( .A(n_912), .B(n_828), .Y(n_980) );
BUFx2_ASAP7_75t_L g981 ( .A(n_931), .Y(n_981) );
INVxp67_ASAP7_75t_L g982 ( .A(n_965), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_942), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_953), .B(n_914), .Y(n_984) );
OR2x2_ASAP7_75t_L g985 ( .A(n_941), .B(n_914), .Y(n_985) );
AND2x4_ASAP7_75t_L g986 ( .A(n_958), .B(n_931), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_953), .B(n_914), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_942), .Y(n_988) );
OR2x2_ASAP7_75t_L g989 ( .A(n_941), .B(n_925), .Y(n_989) );
BUFx3_ASAP7_75t_L g990 ( .A(n_957), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_948), .Y(n_991) );
NOR2xp33_ASAP7_75t_L g992 ( .A(n_976), .B(n_922), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_943), .B(n_925), .Y(n_993) );
INVx2_ASAP7_75t_L g994 ( .A(n_952), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_943), .B(n_925), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_955), .Y(n_996) );
BUFx2_ASAP7_75t_L g997 ( .A(n_946), .Y(n_997) );
HB1xp67_ASAP7_75t_L g998 ( .A(n_944), .Y(n_998) );
AND2x4_ASAP7_75t_L g999 ( .A(n_958), .B(n_931), .Y(n_999) );
CKINVDCx16_ASAP7_75t_R g1000 ( .A(n_957), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_950), .B(n_897), .Y(n_1001) );
OR2x2_ASAP7_75t_L g1002 ( .A(n_946), .B(n_936), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_950), .B(n_900), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_971), .B(n_901), .Y(n_1004) );
INVx2_ASAP7_75t_SL g1005 ( .A(n_945), .Y(n_1005) );
NAND2x1p5_ASAP7_75t_L g1006 ( .A(n_957), .B(n_891), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_971), .B(n_902), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_947), .B(n_902), .Y(n_1008) );
OR2x2_ASAP7_75t_L g1009 ( .A(n_980), .B(n_899), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_956), .B(n_968), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_949), .B(n_903), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_966), .Y(n_1012) );
OR2x2_ASAP7_75t_SL g1013 ( .A(n_972), .B(n_919), .Y(n_1013) );
OR2x2_ASAP7_75t_L g1014 ( .A(n_951), .B(n_899), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_951), .B(n_940), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_978), .B(n_940), .Y(n_1016) );
OR2x2_ASAP7_75t_L g1017 ( .A(n_985), .B(n_954), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_1010), .B(n_973), .Y(n_1018) );
INVx2_ASAP7_75t_L g1019 ( .A(n_994), .Y(n_1019) );
OR2x2_ASAP7_75t_L g1020 ( .A(n_989), .B(n_959), .Y(n_1020) );
INVxp67_ASAP7_75t_L g1021 ( .A(n_998), .Y(n_1021) );
OR2x2_ASAP7_75t_L g1022 ( .A(n_989), .B(n_959), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_984), .B(n_964), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_987), .B(n_962), .Y(n_1024) );
OR2x2_ASAP7_75t_L g1025 ( .A(n_1014), .B(n_977), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_1015), .B(n_962), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_1015), .B(n_960), .Y(n_1027) );
AND2x4_ASAP7_75t_L g1028 ( .A(n_986), .B(n_981), .Y(n_1028) );
NOR2xp33_ASAP7_75t_L g1029 ( .A(n_992), .B(n_933), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_983), .Y(n_1030) );
NAND4xp25_ASAP7_75t_L g1031 ( .A(n_1002), .B(n_920), .C(n_975), .D(n_908), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_993), .B(n_960), .Y(n_1032) );
INVx1_ASAP7_75t_SL g1033 ( .A(n_1000), .Y(n_1033) );
OR2x2_ASAP7_75t_L g1034 ( .A(n_1014), .B(n_978), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_983), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_988), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_993), .B(n_995), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_988), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_995), .B(n_969), .Y(n_1039) );
AND2x2_ASAP7_75t_SL g1040 ( .A(n_1000), .B(n_974), .Y(n_1040) );
INVx2_ASAP7_75t_L g1041 ( .A(n_994), .Y(n_1041) );
NOR2xp33_ASAP7_75t_L g1042 ( .A(n_982), .B(n_933), .Y(n_1042) );
HB1xp67_ASAP7_75t_L g1043 ( .A(n_997), .Y(n_1043) );
INVx2_ASAP7_75t_SL g1044 ( .A(n_1005), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_1016), .B(n_969), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_991), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_1016), .B(n_970), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_996), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_1001), .B(n_970), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_1001), .B(n_961), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1025), .Y(n_1051) );
INVx1_ASAP7_75t_SL g1052 ( .A(n_1033), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1030), .Y(n_1053) );
INVx2_ASAP7_75t_L g1054 ( .A(n_1019), .Y(n_1054) );
INVx2_ASAP7_75t_L g1055 ( .A(n_1019), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1025), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1057 ( .A(n_1037), .B(n_1004), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_1037), .B(n_1024), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1030), .Y(n_1059) );
OR2x2_ASAP7_75t_L g1060 ( .A(n_1034), .B(n_1002), .Y(n_1060) );
NOR2xp67_ASAP7_75t_L g1061 ( .A(n_1044), .B(n_1005), .Y(n_1061) );
OAI32xp33_ASAP7_75t_L g1062 ( .A1(n_1021), .A2(n_1006), .A3(n_979), .B1(n_963), .B2(n_990), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1026), .B(n_1007), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_1032), .B(n_1003), .Y(n_1064) );
HB1xp67_ASAP7_75t_L g1065 ( .A(n_1043), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_1032), .B(n_1003), .Y(n_1066) );
AOI32xp33_ASAP7_75t_L g1067 ( .A1(n_1029), .A2(n_967), .A3(n_997), .B1(n_929), .B2(n_963), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1027), .B(n_1008), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_1027), .B(n_1008), .Y(n_1069) );
INVx1_ASAP7_75t_SL g1070 ( .A(n_1040), .Y(n_1070) );
INVx2_ASAP7_75t_L g1071 ( .A(n_1041), .Y(n_1071) );
INVxp67_ASAP7_75t_L g1072 ( .A(n_1042), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1036), .Y(n_1073) );
INVx2_ASAP7_75t_L g1074 ( .A(n_1041), .Y(n_1074) );
OR2x2_ASAP7_75t_L g1075 ( .A(n_1034), .B(n_1009), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1036), .Y(n_1076) );
AOI22xp5_ASAP7_75t_L g1077 ( .A1(n_1070), .A2(n_1031), .B1(n_1018), .B2(n_1028), .Y(n_1077) );
INVx1_ASAP7_75t_SL g1078 ( .A(n_1052), .Y(n_1078) );
INVx1_ASAP7_75t_SL g1079 ( .A(n_1060), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1051), .Y(n_1080) );
NAND2xp5_ASAP7_75t_SL g1081 ( .A(n_1061), .B(n_1020), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1051), .Y(n_1082) );
INVx2_ASAP7_75t_L g1083 ( .A(n_1075), .Y(n_1083) );
NAND2xp5_ASAP7_75t_L g1084 ( .A(n_1056), .B(n_1064), .Y(n_1084) );
NOR3xp33_ASAP7_75t_SL g1085 ( .A(n_1062), .B(n_863), .C(n_862), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_1066), .B(n_1023), .Y(n_1086) );
NAND3xp33_ASAP7_75t_L g1087 ( .A(n_1065), .B(n_892), .C(n_934), .Y(n_1087) );
INVx5_ASAP7_75t_L g1088 ( .A(n_1062), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1060), .Y(n_1089) );
NOR2xp33_ASAP7_75t_L g1090 ( .A(n_1072), .B(n_855), .Y(n_1090) );
NAND3xp33_ASAP7_75t_L g1091 ( .A(n_1067), .B(n_923), .C(n_853), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1084), .Y(n_1092) );
AOI22xp5_ASAP7_75t_L g1093 ( .A1(n_1077), .A2(n_1085), .B1(n_1078), .B2(n_1081), .Y(n_1093) );
OR2x2_ASAP7_75t_L g1094 ( .A(n_1083), .B(n_1058), .Y(n_1094) );
AOI221xp5_ASAP7_75t_L g1095 ( .A1(n_1087), .A2(n_1068), .B1(n_1069), .B2(n_1057), .C(n_1063), .Y(n_1095) );
INVx1_ASAP7_75t_SL g1096 ( .A(n_1079), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1080), .Y(n_1097) );
NAND3xp33_ASAP7_75t_SL g1098 ( .A(n_1091), .B(n_1006), .C(n_906), .Y(n_1098) );
AOI221x1_ASAP7_75t_L g1099 ( .A1(n_1090), .A2(n_1053), .B1(n_1073), .B2(n_1076), .C(n_1059), .Y(n_1099) );
AOI22xp5_ASAP7_75t_L g1100 ( .A1(n_1089), .A2(n_1045), .B1(n_1047), .B2(n_1039), .Y(n_1100) );
AOI322xp5_ASAP7_75t_L g1101 ( .A1(n_1086), .A2(n_1039), .A3(n_1049), .B1(n_1050), .B2(n_1076), .C1(n_1059), .C2(n_1011), .Y(n_1101) );
NOR2x1_ASAP7_75t_L g1102 ( .A(n_1087), .B(n_910), .Y(n_1102) );
AOI31xp33_ASAP7_75t_L g1103 ( .A1(n_1088), .A2(n_898), .A3(n_1013), .B(n_1020), .Y(n_1103) );
AOI221xp5_ASAP7_75t_L g1104 ( .A1(n_1082), .A2(n_1049), .B1(n_1038), .B2(n_1048), .C(n_1035), .Y(n_1104) );
AOI221xp5_ASAP7_75t_L g1105 ( .A1(n_1077), .A2(n_1046), .B1(n_1017), .B2(n_1022), .C(n_1054), .Y(n_1105) );
AOI221xp5_ASAP7_75t_L g1106 ( .A1(n_1077), .A2(n_1074), .B1(n_1071), .B2(n_1055), .C(n_1012), .Y(n_1106) );
NOR2xp33_ASAP7_75t_L g1107 ( .A(n_1093), .B(n_1096), .Y(n_1107) );
NOR2xp33_ASAP7_75t_SL g1108 ( .A(n_1102), .B(n_1098), .Y(n_1108) );
NAND3xp33_ASAP7_75t_L g1109 ( .A(n_1099), .B(n_1105), .C(n_1106), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1110 ( .A(n_1095), .B(n_1101), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1092), .Y(n_1111) );
NOR2xp33_ASAP7_75t_L g1112 ( .A(n_1107), .B(n_1097), .Y(n_1112) );
NOR2x1_ASAP7_75t_L g1113 ( .A(n_1109), .B(n_1103), .Y(n_1113) );
NAND4xp25_ASAP7_75t_L g1114 ( .A(n_1113), .B(n_1110), .C(n_1108), .D(n_1111), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_1112), .A2(n_1100), .B1(n_1094), .B2(n_1104), .Y(n_1115) );
HB1xp67_ASAP7_75t_L g1116 ( .A(n_1114), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1115), .Y(n_1117) );
XNOR2xp5_ASAP7_75t_L g1118 ( .A(n_1116), .B(n_921), .Y(n_1118) );
OAI22x1_ASAP7_75t_L g1119 ( .A1(n_1117), .A2(n_937), .B1(n_835), .B2(n_930), .Y(n_1119) );
AOI21xp5_ASAP7_75t_L g1120 ( .A1(n_1118), .A2(n_921), .B(n_893), .Y(n_1120) );
OA22x2_ASAP7_75t_L g1121 ( .A1(n_1120), .A2(n_1119), .B1(n_893), .B2(n_895), .Y(n_1121) );
AO21x2_ASAP7_75t_L g1122 ( .A1(n_1121), .A2(n_896), .B(n_890), .Y(n_1122) );
AO21x2_ASAP7_75t_L g1123 ( .A1(n_1122), .A2(n_827), .B(n_814), .Y(n_1123) );
AOI22xp5_ASAP7_75t_L g1124 ( .A1(n_1123), .A2(n_999), .B1(n_906), .B2(n_924), .Y(n_1124) );
endmodule