module fake_jpeg_5742_n_164 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_2),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_0),
.B(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_1),
.B(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_17),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_35),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_34),
.Y(n_46)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_17),
.B(n_1),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_43),
.B1(n_20),
.B2(n_21),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_38),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_1),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_29),
.Y(n_60)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

OA22x2_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_20),
.B1(n_14),
.B2(n_26),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_44),
.A2(n_66),
.B1(n_69),
.B2(n_7),
.Y(n_94)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_49),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_30),
.B(n_22),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_26),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_56),
.C(n_39),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_61),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_25),
.B1(n_29),
.B2(n_22),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_59),
.A2(n_2),
.B1(n_8),
.B2(n_7),
.Y(n_93)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_40),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_35),
.B(n_15),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_15),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_21),
.B1(n_19),
.B2(n_16),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_39),
.A2(n_23),
.B1(n_16),
.B2(n_19),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_60),
.B1(n_44),
.B2(n_57),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_SL g68 ( 
.A(n_31),
.B(n_8),
.C(n_10),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g69 ( 
.A1(n_38),
.A2(n_23),
.A3(n_4),
.B1(n_5),
.B2(n_2),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_31),
.B(n_24),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_28),
.Y(n_87)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_79),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_75),
.Y(n_113)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_63),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_94),
.Y(n_108)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_93),
.B1(n_48),
.B2(n_56),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_44),
.A2(n_40),
.B1(n_31),
.B2(n_4),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_92),
.A2(n_83),
.B1(n_74),
.B2(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_72),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_69),
.B1(n_56),
.B2(n_57),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_78),
.B(n_80),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_102),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_84),
.B1(n_90),
.B2(n_107),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_73),
.B(n_54),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_112),
.B(n_102),
.Y(n_125)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_100),
.B(n_106),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_47),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_107),
.C(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_70),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_70),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_72),
.Y(n_111)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_88),
.B1(n_95),
.B2(n_86),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_115),
.B1(n_122),
.B2(n_108),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_108),
.A2(n_75),
.B1(n_81),
.B2(n_76),
.Y(n_115)
);

AO21x1_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_104),
.B(n_113),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_121),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_123),
.B(n_126),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_99),
.Y(n_136)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_127),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_131),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_105),
.C(n_108),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_138),
.C(n_117),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_115),
.B(n_103),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_132),
.B(n_135),
.Y(n_140)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_133),
.B(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_111),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_98),
.C(n_100),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_114),
.B1(n_116),
.B2(n_125),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_145),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_141),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_131),
.B(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_147),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_130),
.A2(n_117),
.B1(n_121),
.B2(n_138),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_146),
.A2(n_128),
.B(n_139),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_134),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_152),
.B(n_142),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_145),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_149),
.B(n_142),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_146),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_150),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_156),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_157),
.A2(n_151),
.B(n_152),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_154),
.B(n_151),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_158),
.B(n_159),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_160),
.B(n_140),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_161),
.Y(n_163)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_163),
.Y(n_164)
);


endmodule