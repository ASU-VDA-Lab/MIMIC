module fake_jpeg_11500_n_40 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_40);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_40;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

INVx4_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_10),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_19),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_23),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_1),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_26)
);

AO21x1_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_28),
.B(n_17),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_2),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_4),
.B(n_5),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_1),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_33),
.C(n_34),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_8),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_37),
.A2(n_9),
.B(n_13),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_3),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_35),
.Y(n_40)
);


endmodule