module fake_jpeg_18278_n_262 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_262);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_26),
.Y(n_60)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_20),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_1),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_28),
.Y(n_74)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_20),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_53),
.Y(n_84)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_37),
.Y(n_53)
);

OA22x2_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_36),
.B1(n_18),
.B2(n_21),
.Y(n_54)
);

AO22x1_ASAP7_75t_SL g103 ( 
.A1(n_54),
.A2(n_35),
.B1(n_19),
.B2(n_29),
.Y(n_103)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_26),
.B1(n_33),
.B2(n_31),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_56),
.A2(n_57),
.B1(n_64),
.B2(n_32),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_26),
.B1(n_33),
.B2(n_31),
.Y(n_57)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_59),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_65),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_33),
.B1(n_25),
.B2(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_30),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_66),
.B(n_73),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_43),
.B1(n_37),
.B2(n_22),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_67),
.A2(n_60),
.B1(n_77),
.B2(n_61),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_36),
.B(n_19),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_29),
.C(n_27),
.Y(n_113)
);

HAxp5_ASAP7_75t_SL g72 ( 
.A(n_44),
.B(n_36),
.CON(n_72),
.SN(n_72)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_72),
.A2(n_32),
.B1(n_31),
.B2(n_35),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_17),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_22),
.Y(n_101)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_79),
.Y(n_87)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_24),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_35),
.B1(n_19),
.B2(n_36),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_82),
.A2(n_103),
.B1(n_95),
.B2(n_100),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_24),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_88),
.B(n_91),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_34),
.B(n_36),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_89),
.A2(n_23),
.B(n_29),
.Y(n_132)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_30),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_97),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_98),
.A2(n_81),
.B1(n_51),
.B2(n_62),
.Y(n_127)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_101),
.B(n_106),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_68),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_110),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_23),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_103),
.B(n_82),
.C(n_105),
.Y(n_124)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_54),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_SL g141 ( 
.A(n_109),
.B(n_113),
.C(n_63),
.Y(n_141)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_63),
.Y(n_131)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_73),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_113),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_81),
.B1(n_78),
.B2(n_75),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_124),
.B1(n_127),
.B2(n_134),
.Y(n_148)
);

NAND2xp33_ASAP7_75t_SL g123 ( 
.A(n_82),
.B(n_54),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_112),
.C(n_2),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_84),
.B(n_59),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_125),
.B(n_138),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_58),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_128),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_58),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_29),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_129),
.B(n_136),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_131),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_6),
.B(n_7),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_89),
.A2(n_62),
.B1(n_27),
.B2(n_80),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_141),
.B1(n_104),
.B2(n_27),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_86),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_142),
.Y(n_150)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_82),
.A2(n_23),
.A3(n_27),
.B1(n_3),
.B2(n_4),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_83),
.B(n_1),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_166),
.B(n_138),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_90),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_121),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_129),
.A2(n_96),
.B1(n_94),
.B2(n_108),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_157),
.B1(n_163),
.B2(n_167),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_1),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_9),
.Y(n_178)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_136),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_110),
.C(n_112),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_146),
.C(n_161),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_124),
.A2(n_96),
.B1(n_94),
.B2(n_104),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_114),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_158),
.B(n_162),
.Y(n_191)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_160),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_161),
.A2(n_136),
.B(n_139),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_92),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_6),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_124),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_169),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_116),
.B(n_9),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_176),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_172),
.A2(n_181),
.B(n_188),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_173),
.B(n_177),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_141),
.B(n_139),
.Y(n_174)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_180),
.C(n_166),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_132),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_115),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_178),
.B(n_189),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_124),
.B1(n_122),
.B2(n_134),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_183),
.A2(n_148),
.B1(n_153),
.B2(n_163),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_135),
.Y(n_184)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_135),
.Y(n_186)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_SL g188 ( 
.A1(n_148),
.A2(n_119),
.B(n_117),
.C(n_140),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_151),
.B(n_140),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_165),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_155),
.C(n_165),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_172),
.C(n_173),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_201),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_185),
.B(n_11),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_207),
.B1(n_188),
.B2(n_179),
.Y(n_213)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_149),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_202),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_167),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_152),
.Y(n_220)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_205),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_147),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_206),
.A2(n_196),
.B(n_209),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_179),
.A2(n_158),
.B1(n_156),
.B2(n_154),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_221),
.C(n_201),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_217),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_180),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_220),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_197),
.A2(n_188),
.B1(n_189),
.B2(n_181),
.Y(n_215)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_199),
.A2(n_188),
.B1(n_170),
.B2(n_182),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_194),
.A2(n_188),
.B1(n_182),
.B2(n_156),
.Y(n_218)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_207),
.A2(n_175),
.B1(n_185),
.B2(n_160),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_219),
.A2(n_224),
.B(n_196),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_159),
.C(n_178),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_223),
.B(n_208),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_210),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_225),
.A2(n_231),
.B(n_233),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_193),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_214),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_206),
.B(n_203),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_236),
.C(n_221),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_224),
.A2(n_206),
.B(n_195),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_219),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_168),
.C(n_11),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_218),
.B1(n_216),
.B2(n_222),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_237),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_239),
.Y(n_245)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_231),
.C(n_230),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_212),
.C(n_223),
.Y(n_243)
);

OAI221xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_244),
.B1(n_229),
.B2(n_12),
.C(n_13),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_236),
.A2(n_213),
.B1(n_212),
.B2(n_13),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_247),
.B(n_10),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_235),
.B1(n_228),
.B2(n_226),
.Y(n_248)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_248),
.Y(n_254)
);

AO21x1_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_234),
.B(n_229),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_250),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_238),
.C(n_241),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_249),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_253),
.A2(n_10),
.B(n_13),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_257),
.C(n_252),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_251),
.B(n_246),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_256),
.Y(n_259)
);

OAI21x1_ASAP7_75t_L g260 ( 
.A1(n_258),
.A2(n_254),
.B(n_14),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_259),
.C(n_15),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_15),
.Y(n_262)
);


endmodule