module fake_jpeg_21043_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVxp33_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_19),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_40),
.Y(n_73)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_56),
.B(n_70),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_17),
.B1(n_21),
.B2(n_35),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_26),
.B1(n_31),
.B2(n_30),
.Y(n_92)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_17),
.B1(n_27),
.B2(n_33),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_26),
.B1(n_18),
.B2(n_33),
.Y(n_80)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g111 ( 
.A(n_65),
.Y(n_111)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_27),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_24),
.B(n_49),
.C(n_28),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_72),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_73),
.B(n_102),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_74),
.Y(n_122)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_49),
.B1(n_17),
.B2(n_50),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_75),
.A2(n_92),
.B1(n_63),
.B2(n_46),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_52),
.C(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_81),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_80),
.A2(n_25),
.B1(n_34),
.B2(n_20),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_50),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_82),
.B(n_91),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_42),
.B1(n_43),
.B2(n_18),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_86),
.B1(n_65),
.B2(n_58),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_43),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_88),
.Y(n_119)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_42),
.B1(n_30),
.B2(n_31),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_51),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_25),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_36),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_99),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_36),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_62),
.A2(n_24),
.B1(n_28),
.B2(n_22),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_25),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_53),
.B(n_40),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_105),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_36),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_107),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_36),
.C(n_46),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_67),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_109),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_53),
.B(n_24),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_58),
.B(n_15),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_112),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_130),
.B1(n_85),
.B2(n_110),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_63),
.B1(n_65),
.B2(n_24),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_123),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_146),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_131),
.B1(n_135),
.B2(n_83),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_63),
.B1(n_34),
.B2(n_20),
.Y(n_130)
);

OAI22x1_ASAP7_75t_SL g131 ( 
.A1(n_72),
.A2(n_22),
.B1(n_25),
.B2(n_23),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_34),
.B1(n_15),
.B2(n_14),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_144),
.A2(n_80),
.B1(n_81),
.B2(n_86),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_95),
.A2(n_14),
.B1(n_13),
.B2(n_23),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_145),
.A2(n_111),
.B1(n_90),
.B2(n_79),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_78),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_77),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_171),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_151),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_153),
.A2(n_157),
.B1(n_161),
.B2(n_114),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_94),
.C(n_73),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_116),
.C(n_139),
.Y(n_187)
);

AO21x2_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_75),
.B(n_82),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_133),
.B1(n_143),
.B2(n_138),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_75),
.B1(n_103),
.B2(n_88),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_164),
.B1(n_172),
.B2(n_144),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_94),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_178),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_122),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_160),
.B(n_165),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_93),
.B1(n_107),
.B2(n_106),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_129),
.A2(n_103),
.B(n_112),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_162),
.A2(n_117),
.B(n_5),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_163),
.A2(n_148),
.B1(n_114),
.B2(n_7),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_126),
.A2(n_111),
.B1(n_90),
.B2(n_79),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_132),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_131),
.A2(n_98),
.B1(n_89),
.B2(n_111),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_120),
.B(n_133),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_132),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_170),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_0),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_126),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_129),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_3),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_121),
.B(n_97),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_179),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_115),
.A2(n_122),
.B(n_121),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_176),
.A2(n_120),
.B(n_143),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_87),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_140),
.B(n_2),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_113),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_148),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_3),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_4),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_182),
.A2(n_193),
.B1(n_211),
.B2(n_156),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_125),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_183),
.B(n_190),
.Y(n_233)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_162),
.A2(n_125),
.B(n_137),
.C(n_116),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_184),
.B(n_200),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_118),
.B1(n_146),
.B2(n_147),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_195),
.B1(n_201),
.B2(n_205),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_191),
.C(n_178),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_188),
.A2(n_197),
.B(n_198),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_130),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_134),
.C(n_113),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_176),
.A2(n_152),
.B(n_168),
.Y(n_198)
);

XOR2x1_ASAP7_75t_SL g199 ( 
.A(n_156),
.B(n_158),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_199),
.A2(n_204),
.B(n_212),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_138),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_157),
.A2(n_148),
.B1(n_6),
.B2(n_7),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_207),
.A2(n_213),
.B1(n_164),
.B2(n_173),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_166),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_180),
.Y(n_238)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_209),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_172),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_177),
.A2(n_6),
.B(n_8),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_202),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_228),
.Y(n_244)
);

AOI22x1_ASAP7_75t_L g217 ( 
.A1(n_199),
.A2(n_156),
.B1(n_167),
.B2(n_151),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_217),
.A2(n_204),
.B1(n_190),
.B2(n_212),
.Y(n_250)
);

AND2x2_ASAP7_75t_SL g219 ( 
.A(n_197),
.B(n_168),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_219),
.A2(n_221),
.B(n_239),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_177),
.B(n_161),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_233),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_189),
.B1(n_194),
.B2(n_213),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_229),
.C(n_241),
.Y(n_243)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_183),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_230),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_185),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_227),
.B(n_234),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_191),
.C(n_187),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_173),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_206),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_156),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_217),
.Y(n_249)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_154),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_165),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_225),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_249),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_223),
.A2(n_201),
.B1(n_195),
.B2(n_207),
.Y(n_245)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_245),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_215),
.A2(n_182),
.B1(n_208),
.B2(n_189),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_253),
.B1(n_254),
.B2(n_228),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_248),
.B(n_229),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_235),
.A2(n_232),
.B1(n_217),
.B2(n_221),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_257),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_239),
.A2(n_196),
.B1(n_210),
.B2(n_169),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_214),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_231),
.Y(n_274)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_220),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_214),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_258),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_236),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_259),
.A2(n_219),
.B(n_230),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_218),
.B(n_8),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_261),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_251),
.B(n_218),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_264),
.B(n_277),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_274),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_224),
.C(n_233),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_248),
.C(n_260),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_241),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_280),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_271),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_245),
.B1(n_252),
.B2(n_244),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_255),
.A2(n_239),
.B1(n_240),
.B2(n_216),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_273),
.A2(n_276),
.B1(n_278),
.B2(n_249),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_243),
.A2(n_240),
.B1(n_231),
.B2(n_237),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_242),
.A2(n_219),
.B1(n_222),
.B2(n_11),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_9),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_254),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_287),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_286),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_281),
.A2(n_266),
.B1(n_244),
.B2(n_275),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_265),
.C(n_276),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_291),
.C(n_292),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_296),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_247),
.C(n_262),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_262),
.C(n_246),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_279),
.B(n_259),
.Y(n_293)
);

INVx11_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_267),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_246),
.C(n_263),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_300),
.C(n_291),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_278),
.C(n_257),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_266),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_300),
.Y(n_314)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_305),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_297),
.A2(n_285),
.B(n_290),
.Y(n_307)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_284),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_308),
.B(n_309),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_306),
.A2(n_289),
.B1(n_295),
.B2(n_292),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_310),
.B(n_311),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_282),
.C(n_11),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_10),
.B1(n_12),
.B2(n_298),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_312),
.B(n_314),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_305),
.Y(n_316)
);

OA21x2_ASAP7_75t_L g322 ( 
.A1(n_316),
.A2(n_302),
.B(n_297),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_311),
.B(n_301),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_317),
.B(n_310),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_322),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_304),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_320),
.B(n_315),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_324),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_325),
.B(n_319),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_321),
.B(n_316),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_304),
.B(n_10),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_12),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_12),
.Y(n_331)
);


endmodule