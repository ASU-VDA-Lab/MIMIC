module real_jpeg_13083_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_343, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_343;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_0),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_0),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_0),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_61),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_0),
.A2(n_44),
.B1(n_45),
.B2(n_61),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_3),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_62)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_3),
.A2(n_57),
.B1(n_58),
.B2(n_66),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g195 ( 
.A(n_3),
.B(n_64),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_4),
.A2(n_63),
.B1(n_64),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_4),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_4),
.A2(n_44),
.B1(n_45),
.B2(n_151),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_151),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_4),
.A2(n_57),
.B1(n_58),
.B2(n_151),
.Y(n_268)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_6),
.A2(n_43),
.B1(n_63),
.B2(n_64),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_6),
.A2(n_43),
.B1(n_57),
.B2(n_58),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_43),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_7),
.A2(n_63),
.B1(n_64),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_7),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_7),
.A2(n_57),
.B1(n_58),
.B2(n_83),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_83),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_83),
.Y(n_161)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_9),
.A2(n_57),
.B1(n_58),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_9),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_9),
.A2(n_63),
.B1(n_64),
.B2(n_73),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_73),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_73),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_10),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_10),
.A2(n_39),
.B1(n_63),
.B2(n_64),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_10),
.A2(n_39),
.B1(n_57),
.B2(n_58),
.Y(n_328)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_11),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_12),
.B(n_157),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_12),
.A2(n_63),
.B(n_80),
.C(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_12),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_12),
.B(n_57),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_171),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_12),
.B(n_34),
.C(n_48),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_12),
.B(n_81),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_12),
.A2(n_116),
.B(n_219),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_171),
.Y(n_245)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_13),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_14),
.A2(n_53),
.B1(n_63),
.B2(n_64),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_53),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_14),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_17),
.A2(n_57),
.B1(n_58),
.B2(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_17),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_17),
.A2(n_44),
.B1(n_45),
.B2(n_125),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_17),
.A2(n_63),
.B1(n_64),
.B2(n_125),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_17),
.A2(n_33),
.B1(n_34),
.B2(n_125),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_18),
.A2(n_20),
.B(n_339),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_18),
.B(n_340),
.Y(n_339)
);

AOI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_334),
.B(n_337),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_326),
.B(n_330),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_313),
.B(n_325),
.Y(n_22)
);

AO21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_141),
.B(n_310),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_128),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_103),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_26),
.B(n_103),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_26),
.Y(n_342)
);

FAx1_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_74),
.CI(n_89),
.CON(n_26),
.SN(n_26)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_27),
.B(n_74),
.C(n_89),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B(n_55),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_28),
.A2(n_29),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_40),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_30),
.A2(n_31),
.B1(n_55),
.B2(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_30),
.A2(n_31),
.B1(n_40),
.B2(n_41),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_36),
.B(n_37),
.Y(n_31)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_32),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_32),
.B(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_32),
.A2(n_36),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_32),
.A2(n_36),
.B1(n_115),
.B2(n_199),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_34),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_33),
.B(n_235),
.Y(n_234)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_36),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_36),
.B(n_174),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_38),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_46),
.B1(n_51),
.B2(n_54),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_42),
.A2(n_46),
.B1(n_54),
.B2(n_120),
.Y(n_119)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

AO22x1_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_45),
.B1(n_79),
.B2(n_80),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_44),
.B(n_209),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_45),
.A2(n_79),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_46),
.A2(n_54),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_46),
.B(n_166),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_46),
.A2(n_54),
.B1(n_164),
.B2(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_46),
.A2(n_54),
.B1(n_120),
.B2(n_187),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_50),
.A2(n_52),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_50),
.A2(n_186),
.B(n_188),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_50),
.A2(n_188),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_50),
.B(n_171),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_54),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_62),
.B(n_67),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_56),
.A2(n_62),
.B1(n_69),
.B2(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_58),
.A2(n_69),
.B(n_171),
.C(n_180),
.Y(n_179)
);

AOI32xp33_ASAP7_75t_L g194 ( 
.A1(n_58),
.A2(n_63),
.A3(n_66),
.B1(n_181),
.B2(n_195),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_62),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_62),
.B(n_72),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_62),
.A2(n_69),
.B1(n_101),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_62),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_62),
.A2(n_67),
.B(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_62),
.A2(n_69),
.B1(n_124),
.B2(n_268),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_64),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_68),
.A2(n_157),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_68),
.A2(n_157),
.B1(n_320),
.B2(n_328),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_68),
.A2(n_157),
.B(n_328),
.Y(n_336)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_69),
.A2(n_124),
.B(n_126),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_75),
.B(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_86),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_76),
.A2(n_82),
.B1(n_84),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_76),
.A2(n_84),
.B1(n_94),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_76),
.A2(n_84),
.B1(n_150),
.B2(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_76),
.A2(n_245),
.B(n_246),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_76),
.A2(n_184),
.B(n_246),
.Y(n_266)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_81),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_77),
.B(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_77),
.A2(n_81),
.B(n_317),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_81),
.B(n_153),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_84),
.A2(n_150),
.B(n_152),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_84),
.A2(n_122),
.B(n_152),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_87),
.A2(n_163),
.B(n_165),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_87),
.A2(n_165),
.B(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_SL g139 ( 
.A(n_91),
.B(n_96),
.C(n_100),
.Y(n_139)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_95),
.A2(n_96),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_96),
.B(n_133),
.C(n_137),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_100),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_100),
.B(n_132),
.C(n_139),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_109),
.C(n_110),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_104),
.A2(n_105),
.B1(n_109),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_109),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_110),
.B(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_121),
.C(n_123),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_111),
.A2(n_112),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_113),
.A2(n_118),
.B1(n_119),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_113),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_116),
.A2(n_117),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_116),
.A2(n_117),
.B1(n_161),
.B2(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_116),
.A2(n_218),
.B(n_219),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_117),
.A2(n_160),
.B(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_117),
.A2(n_173),
.B(n_224),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_117),
.B(n_171),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_121),
.B(n_123),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_127),
.B(n_179),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g310 ( 
.A1(n_128),
.A2(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_140),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_129),
.B(n_140),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_139),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_134),
.Y(n_319)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_138),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_304),
.B(n_309),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_292),
.B(n_303),
.Y(n_142)
);

OAI321xp33_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_260),
.A3(n_285),
.B1(n_290),
.B2(n_291),
.C(n_343),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_200),
.B(n_259),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_175),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_146),
.B(n_175),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_162),
.C(n_167),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_147),
.A2(n_148),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_154),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_155),
.C(n_159),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_162),
.A2(n_167),
.B1(n_168),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_162),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_169),
.B(n_172),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_190),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_176),
.B(n_191),
.C(n_192),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_182),
.B2(n_189),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_177),
.B(n_183),
.C(n_185),
.Y(n_274)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_193),
.B(n_197),
.Y(n_270)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_252),
.B(n_258),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_239),
.B(n_251),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_220),
.B(n_238),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_210),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_204),
.B(n_210),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_208),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_217),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_215),
.C(n_217),
.Y(n_240)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_216),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_218),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_228),
.B(n_237),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_222),
.B(n_226),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_232),
.B(n_236),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_230),
.B(n_231),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_240),
.B(n_241),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_247),
.C(n_250),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.Y(n_243)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_244),
.Y(n_250)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_253),
.B(n_254),
.Y(n_258)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_275),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_275),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_271),
.C(n_274),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_262),
.A2(n_263),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_270),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_269),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_269),
.C(n_270),
.Y(n_284)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_271),
.B(n_274),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_273),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_284),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_279),
.C(n_284),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_282),
.C(n_283),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_286),
.B(n_287),
.Y(n_290)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_302),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_302),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_297),
.C(n_298),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_306),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_324),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_324),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_323),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_318),
.B1(n_321),
.B2(n_322),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_316),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_318),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_321),
.C(n_323),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_327),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_335),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_329),
.Y(n_333)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_336),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_338),
.Y(n_337)
);


endmodule