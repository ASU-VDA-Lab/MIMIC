module fake_jpeg_15688_n_26 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_26);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_26;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

OAI22xp5_ASAP7_75t_SL g8 ( 
.A1(n_5),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_0),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_5),
.A2(n_6),
.B1(n_1),
.B2(n_0),
.Y(n_13)
);

HAxp5_ASAP7_75t_SL g14 ( 
.A(n_1),
.B(n_0),
.CON(n_14),
.SN(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_9),
.B(n_10),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_9),
.B(n_10),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_13),
.A2(n_12),
.B1(n_7),
.B2(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_11),
.C(n_14),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_7),
.A2(n_12),
.B(n_11),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_24),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_17),
.B(n_19),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_12),
.B1(n_22),
.B2(n_21),
.Y(n_26)
);


endmodule