module fake_jpeg_23858_n_132 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_28),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_15),
.A2(n_0),
.B(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_35),
.Y(n_42)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_0),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_56),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_19),
.B1(n_14),
.B2(n_13),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_20),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_31),
.A2(n_19),
.B1(n_14),
.B2(n_13),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_29),
.A2(n_26),
.B1(n_21),
.B2(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_30),
.B(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_24),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_37),
.B(n_38),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_61),
.B1(n_74),
.B2(n_77),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_R g92 ( 
.A(n_60),
.B(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_63),
.Y(n_79)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_73),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_33),
.C(n_34),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_57),
.C(n_55),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_24),
.B1(n_32),
.B2(n_27),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_20),
.B1(n_18),
.B2(n_21),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_50),
.B1(n_55),
.B2(n_40),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_3),
.Y(n_72)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_7),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_34),
.B(n_10),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_77),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_91),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_88),
.B1(n_76),
.B2(n_58),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_8),
.B1(n_11),
.B2(n_61),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_69),
.B(n_60),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_72),
.B1(n_60),
.B2(n_68),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_96),
.B(n_99),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_63),
.B1(n_64),
.B2(n_75),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_98),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_81),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_101),
.C(n_102),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_91),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_82),
.Y(n_102)
);

INVx4_ASAP7_75t_SL g103 ( 
.A(n_92),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_103),
.A2(n_84),
.B(n_87),
.Y(n_110)
);

OAI22x1_ASAP7_75t_SL g105 ( 
.A1(n_103),
.A2(n_83),
.B1(n_95),
.B2(n_82),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_84),
.B1(n_94),
.B2(n_78),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_83),
.B(n_85),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_110),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_100),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_112),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_115),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_114),
.A2(n_117),
.B1(n_107),
.B2(n_65),
.Y(n_121)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_107),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_104),
.A2(n_94),
.B1(n_90),
.B2(n_73),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_121),
.Y(n_127)
);

OR2x6_ASAP7_75t_SL g124 ( 
.A(n_119),
.B(n_113),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_126),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_120),
.A2(n_118),
.B(n_58),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_122),
.Y(n_129)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_129),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_128),
.B(n_125),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_123),
.Y(n_132)
);


endmodule