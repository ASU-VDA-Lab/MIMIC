module fake_jpeg_30162_n_116 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_116);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx12_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_20),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_6),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_56)
);

AO21x1_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_60),
.B(n_6),
.Y(n_67)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_44),
.B1(n_51),
.B2(n_53),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_40),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_47),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_57),
.B(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_73),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_48),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_69),
.B(n_15),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_7),
.B(n_8),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_71),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_29),
.B(n_37),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_44),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_52),
.B1(n_50),
.B2(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_74),
.B(n_80),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_30),
.C(n_31),
.Y(n_97)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_40),
.B1(n_9),
.B2(n_10),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

NOR3xp33_ASAP7_75t_SL g87 ( 
.A(n_84),
.B(n_18),
.C(n_21),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_87),
.B(n_89),
.Y(n_106)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_23),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_93),
.B(n_90),
.Y(n_105)
);

NOR3xp33_ASAP7_75t_SL g89 ( 
.A(n_77),
.B(n_24),
.C(n_25),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_26),
.C(n_28),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_38),
.C(n_75),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_99),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_96),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_32),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_34),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_100),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_36),
.Y(n_101)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_103),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_104),
.C(n_105),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_111),
.C(n_109),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_103),
.B(n_92),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_88),
.B(n_92),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_109),
.B1(n_87),
.B2(n_106),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_89),
.Y(n_115)
);

BUFx24_ASAP7_75t_SL g116 ( 
.A(n_115),
.Y(n_116)
);


endmodule