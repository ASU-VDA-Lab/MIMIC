module real_jpeg_9456_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_206;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_39),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_2),
.A2(n_56),
.B1(n_57),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_2),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_68),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_68),
.Y(n_172)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_3),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_4),
.A2(n_72),
.B1(n_79),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_4),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_4),
.A2(n_56),
.B1(n_57),
.B2(n_82),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_82),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_82),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_5),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_5),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_5),
.A2(n_59),
.B1(n_72),
.B2(n_79),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_59),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_59),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_6),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_6),
.A2(n_56),
.B1(n_57),
.B2(n_86),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_86),
.Y(n_165)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_SL g63 ( 
.A(n_10),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_12),
.A2(n_72),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_12),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_12),
.A2(n_57),
.B(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_12),
.B(n_83),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_12),
.A2(n_31),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_12),
.B(n_31),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_12),
.A2(n_46),
.B1(n_96),
.B2(n_149),
.Y(n_151)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_123),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_121),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_20),
.B(n_105),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_89),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_51),
.B1(n_52),
.B2(n_88),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_22),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_43),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_36),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_24),
.A2(n_28),
.B(n_31),
.C(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_24),
.B(n_38),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_24),
.A2(n_41),
.B1(n_137),
.B2(n_139),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_24),
.B(n_78),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_24),
.A2(n_41),
.B1(n_139),
.B2(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_24),
.A2(n_41),
.B1(n_162),
.B2(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_24),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_25),
.B(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_25),
.B(n_29),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_25),
.B(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_26),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_140)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_31),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_31),
.A2(n_32),
.B1(n_62),
.B2(n_63),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_31),
.B(n_62),
.Y(n_179)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_32),
.A2(n_64),
.B1(n_174),
.B2(n_179),
.Y(n_178)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_40),
.A2(n_85),
.B(n_87),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_41),
.A2(n_172),
.B(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_42),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_46),
.B(n_49),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_44),
.A2(n_46),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_46),
.A2(n_96),
.B1(n_131),
.B2(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_46),
.A2(n_133),
.B(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_46),
.A2(n_49),
.B(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_47),
.B(n_50),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_47),
.A2(n_48),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_50),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_48),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_48),
.B(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_69),
.C(n_84),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_53),
.A2(n_54),
.B1(n_84),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_66),
.B2(n_67),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_55),
.A2(n_60),
.B1(n_66),
.B2(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_57),
.B1(n_73),
.B2(n_74),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_62),
.B(n_64),
.C(n_65),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_62),
.Y(n_64)
);

HAxp5_ASAP7_75t_SL g174 ( 
.A(n_57),
.B(n_78),
.CON(n_174),
.SN(n_174)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_60),
.A2(n_67),
.B(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_61),
.A2(n_65),
.B1(n_116),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_66),
.B(n_78),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_77),
.B1(n_80),
.B2(n_83),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_76),
.B1(n_81),
.B2(n_100),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B(n_75),
.C(n_76),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_73),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_72),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_73),
.B(n_78),
.C(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_78),
.B(n_96),
.Y(n_153)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_85),
.B(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_97),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_94),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_96),
.B(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_101),
.B2(n_104),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_101),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.C(n_111),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_106),
.B(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_109),
.A2(n_111),
.B1(n_112),
.B2(n_205),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_109),
.Y(n_205)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.C(n_118),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_113),
.A2(n_114),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_117),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_201),
.B(n_206),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_184),
.B(n_200),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_167),
.B(n_183),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_156),
.B(n_166),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_145),
.B(n_155),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_134),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_129),
.B(n_134),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_140),
.B2(n_144),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_135),
.B(n_144),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_138),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_140),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_150),
.B(n_154),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_147),
.B(n_148),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_157),
.B(n_158),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_159),
.B(n_168),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_161),
.CI(n_163),
.CON(n_159),
.SN(n_159)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_165),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_177),
.B2(n_182),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_171),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_173),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_176),
.C(n_182),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_177),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_180),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_185),
.B(n_186),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_192),
.B2(n_193),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_195),
.C(n_198),
.Y(n_202)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_198),
.B2(n_199),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_194),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_195),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_202),
.B(n_203),
.Y(n_206)
);


endmodule