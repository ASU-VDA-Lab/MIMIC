module fake_jpeg_12054_n_148 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_148);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_32),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_1),
.C(n_2),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_18),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_38),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_21),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_23),
.B1(n_30),
.B2(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_54),
.Y(n_74)
);

AO22x2_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_23),
.B1(n_29),
.B2(n_20),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_60),
.B1(n_22),
.B2(n_37),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_32),
.A2(n_22),
.B1(n_29),
.B2(n_20),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_31),
.A2(n_28),
.B(n_27),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_19),
.Y(n_66)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_40),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_33),
.A2(n_20),
.B1(n_17),
.B2(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_62),
.B(n_64),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_46),
.B(n_24),
.Y(n_64)
);

AO21x1_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_68),
.B(n_77),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_69),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_24),
.B(n_16),
.C(n_37),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_49),
.A3(n_43),
.B1(n_53),
.B2(n_52),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_17),
.B1(n_25),
.B2(n_19),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_75),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_25),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_53),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_79),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_17),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_9),
.Y(n_79)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_82),
.A2(n_77),
.B(n_68),
.Y(n_109)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_49),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_93),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_57),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_92),
.C(n_71),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_61),
.B(n_52),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_74),
.B(n_77),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_59),
.C(n_3),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_109),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_74),
.B(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_98),
.B(n_95),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_100),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_67),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_103),
.C(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_65),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_77),
.C(n_65),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_110),
.C(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_108),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_80),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_81),
.B1(n_95),
.B2(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_111),
.B(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_94),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_115),
.A2(n_104),
.B(n_88),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_117),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_106),
.C(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_87),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_86),
.B1(n_81),
.B2(n_82),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_97),
.B1(n_109),
.B2(n_83),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_122),
.B(n_125),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_80),
.C(n_4),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_87),
.B(n_69),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_117),
.B(n_80),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_118),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_123),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_127),
.A2(n_118),
.B1(n_119),
.B2(n_2),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_135),
.B(n_126),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_128),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_137),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_124),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_122),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_132),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_141),
.A2(n_143),
.B(n_144),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_134),
.Y(n_143)
);

AOI322xp5_ASAP7_75t_L g146 ( 
.A1(n_143),
.A2(n_4),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_14),
.C2(n_142),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_11),
.C(n_14),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_145),
.Y(n_148)
);


endmodule