module fake_jpeg_28284_n_141 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_141);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_65),
.Y(n_77)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_66),
.B(n_41),
.Y(n_85)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_78),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_47),
.B1(n_56),
.B2(n_50),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_51),
.B1(n_40),
.B2(n_52),
.Y(n_88)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_42),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_58),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_0),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_91),
.Y(n_103)
);

AO22x1_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_54),
.B1(n_52),
.B2(n_40),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_88),
.Y(n_97)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_93),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_54),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_71),
.A2(n_55),
.B1(n_57),
.B2(n_45),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_19),
.B1(n_37),
.B2(n_36),
.Y(n_104)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_67),
.A2(n_73),
.B1(n_55),
.B2(n_68),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_46),
.B1(n_1),
.B2(n_2),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_66),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_96),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_101),
.B1(n_84),
.B2(n_94),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_3),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_100),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_109),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_81),
.B1(n_7),
.B2(n_8),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_112),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_113),
.B(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_102),
.A2(n_90),
.B(n_92),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_105),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_117),
.C(n_119),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_104),
.C(n_82),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_5),
.B(n_10),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_83),
.C(n_99),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_121),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_17),
.C(n_35),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_24),
.C(n_12),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_112),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_115),
.C(n_119),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_130),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_116),
.A2(n_26),
.B(n_13),
.Y(n_130)
);

XNOR2x1_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_127),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_133),
.A2(n_120),
.B(n_132),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_125),
.B(n_130),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_126),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_123),
.B(n_14),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_28),
.B(n_15),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_29),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_31),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_21),
.Y(n_141)
);


endmodule