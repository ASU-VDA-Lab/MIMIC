module fake_jpeg_8354_n_113 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_113);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_113;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_0),
.Y(n_13)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_27),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_34),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_15),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_19),
.B1(n_25),
.B2(n_23),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_49),
.B1(n_20),
.B2(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_23),
.C(n_18),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_17),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_28),
.A2(n_19),
.B1(n_18),
.B2(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_14),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_63),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_15),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_41),
.B1(n_37),
.B2(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_12),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_64),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_0),
.B(n_1),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_62),
.A2(n_5),
.B(n_6),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_3),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_63),
.B(n_64),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVxp33_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_5),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_76),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_51),
.C(n_52),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_84),
.C(n_86),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_83),
.B(n_71),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_42),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_66),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_53),
.B(n_50),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_82),
.B(n_72),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_88),
.B(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_85),
.B(n_69),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_86),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_93),
.Y(n_97)
);

MAJx2_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_92),
.C(n_79),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_84),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_94),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_98),
.A2(n_78),
.B1(n_83),
.B2(n_87),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_100),
.A2(n_97),
.B(n_96),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_102),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_SL g102 ( 
.A(n_95),
.B(n_74),
.C(n_37),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_8),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_102),
.A2(n_80),
.B1(n_8),
.B2(n_7),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_7),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_103),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_60),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_110),
.B(n_60),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

BUFx24_ASAP7_75t_SL g113 ( 
.A(n_112),
.Y(n_113)
);


endmodule