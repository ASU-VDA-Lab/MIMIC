module fake_jpeg_10899_n_472 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_472);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_472;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_13),
.B(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g127 ( 
.A(n_45),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_46),
.Y(n_122)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_48),
.Y(n_126)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_50),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_52),
.B(n_63),
.Y(n_133)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_54),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_58),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx6_ASAP7_75t_SL g123 ( 
.A(n_67),
.Y(n_123)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_22),
.B(n_29),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_91),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_16),
.Y(n_87)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_26),
.A2(n_15),
.B1(n_12),
.B2(n_10),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_88),
.A2(n_38),
.B1(n_30),
.B2(n_28),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_16),
.Y(n_90)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_32),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_45),
.A2(n_26),
.B1(n_41),
.B2(n_19),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_95),
.A2(n_117),
.B1(n_130),
.B2(n_137),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_46),
.A2(n_26),
.B1(n_33),
.B2(n_18),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_55),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_119),
.B(n_143),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_129),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_89),
.A2(n_21),
.B1(n_79),
.B2(n_88),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_58),
.A2(n_38),
.B1(n_33),
.B2(n_18),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_131),
.B(n_32),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_45),
.A2(n_41),
.B1(n_32),
.B2(n_16),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_51),
.A2(n_41),
.B1(n_32),
.B2(n_16),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_141),
.A2(n_30),
.B1(n_59),
.B2(n_28),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_57),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_83),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_146),
.B(n_165),
.Y(n_191)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_147),
.Y(n_198)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_151),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_152),
.B(n_163),
.Y(n_200)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

BUFx2_ASAP7_75t_SL g197 ( 
.A(n_153),
.Y(n_197)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_117),
.A2(n_71),
.B1(n_50),
.B2(n_54),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_155),
.A2(n_159),
.B1(n_185),
.B2(n_188),
.Y(n_210)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_99),
.B(n_83),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_158),
.A2(n_180),
.B(n_186),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_141),
.A2(n_65),
.B1(n_78),
.B2(n_75),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_99),
.A2(n_62),
.B1(n_48),
.B2(n_70),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_167),
.B1(n_120),
.B2(n_110),
.Y(n_194)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_164),
.B(n_169),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_104),
.B(n_81),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_166),
.A2(n_175),
.B1(n_181),
.B2(n_183),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_118),
.A2(n_74),
.B1(n_64),
.B2(n_60),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_172),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_106),
.B(n_57),
.C(n_67),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_184),
.C(n_158),
.Y(n_192)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_173),
.Y(n_220)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_176),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_114),
.A2(n_39),
.B1(n_86),
.B2(n_32),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

INVx4_ASAP7_75t_SL g177 ( 
.A(n_107),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_178),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_107),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_94),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_95),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_114),
.A2(n_39),
.B1(n_32),
.B2(n_42),
.Y(n_181)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

AOI32xp33_ASAP7_75t_L g184 ( 
.A1(n_137),
.A2(n_81),
.A3(n_66),
.B1(n_43),
.B2(n_42),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_139),
.B(n_66),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_190),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_110),
.A2(n_43),
.B1(n_22),
.B2(n_29),
.Y(n_188)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_189),
.A2(n_124),
.B1(n_132),
.B2(n_105),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_124),
.Y(n_190)
);

XNOR2x1_ASAP7_75t_L g249 ( 
.A(n_192),
.B(n_67),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_140),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_156),
.A2(n_145),
.B1(n_120),
.B2(n_100),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_196),
.A2(n_205),
.B1(n_214),
.B2(n_221),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_166),
.A2(n_93),
.B1(n_102),
.B2(n_96),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_155),
.A2(n_105),
.B1(n_132),
.B2(n_128),
.Y(n_207)
);

OA22x2_ASAP7_75t_L g245 ( 
.A1(n_207),
.A2(n_138),
.B1(n_168),
.B2(n_172),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_109),
.C(n_103),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_209),
.C(n_213),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_116),
.C(n_98),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_101),
.C(n_134),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_156),
.A2(n_128),
.B1(n_113),
.B2(n_140),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_182),
.A2(n_113),
.B1(n_138),
.B2(n_122),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_156),
.B(n_20),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_224),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_160),
.B(n_20),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_150),
.B(n_30),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_225),
.B(n_186),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_214),
.A2(n_148),
.B1(n_164),
.B2(n_161),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_226),
.Y(n_265)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_227),
.Y(n_261)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_157),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_230),
.B(n_235),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_231),
.A2(n_256),
.B1(n_194),
.B2(n_196),
.Y(n_272)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_176),
.C(n_173),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_248),
.C(n_205),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_191),
.B(n_37),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_236),
.Y(n_264)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_206),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_240),
.Y(n_271)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_242),
.Y(n_270)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_199),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_250),
.Y(n_277)
);

XNOR2x1_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_249),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_247),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_183),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_246),
.A2(n_215),
.B(n_204),
.Y(n_285)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_206),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_154),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_198),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_254),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_219),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_252),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_206),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_229),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_210),
.A2(n_149),
.B1(n_147),
.B2(n_100),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_213),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_257),
.B(n_275),
.C(n_193),
.Y(n_304)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_235),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_253),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_237),
.A2(n_210),
.B1(n_195),
.B2(n_207),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_267),
.A2(n_268),
.B1(n_282),
.B2(n_283),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_237),
.A2(n_221),
.B1(n_209),
.B2(n_225),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_228),
.A2(n_200),
.B(n_219),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_274),
.B(n_247),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_272),
.A2(n_276),
.B1(n_279),
.B2(n_197),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_201),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_273),
.B(n_177),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_228),
.A2(n_200),
.B(n_219),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_256),
.A2(n_218),
.B1(n_224),
.B2(n_201),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_231),
.A2(n_198),
.B1(n_202),
.B2(n_215),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_233),
.A2(n_220),
.B1(n_222),
.B2(n_198),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_254),
.A2(n_220),
.B1(n_216),
.B2(n_163),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_285),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_227),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_265),
.A2(n_255),
.B1(n_236),
.B2(n_240),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_287),
.A2(n_301),
.B1(n_307),
.B2(n_313),
.Y(n_324)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_261),
.Y(n_288)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_288),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_289),
.B(n_284),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_290),
.B(n_305),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_291),
.B(n_292),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_270),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_261),
.Y(n_293)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_293),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_272),
.A2(n_234),
.B1(n_250),
.B2(n_246),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_294),
.A2(n_298),
.B1(n_299),
.B2(n_303),
.Y(n_336)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_262),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_295),
.B(n_302),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_296),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_286),
.A2(n_253),
.B1(n_231),
.B2(n_244),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_275),
.A2(n_248),
.B1(n_239),
.B2(n_245),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_257),
.B(n_280),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_304),
.C(n_306),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_265),
.A2(n_232),
.B1(n_251),
.B2(n_238),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_243),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_265),
.A2(n_245),
.B1(n_216),
.B2(n_204),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_262),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_178),
.C(n_217),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_276),
.A2(n_245),
.B1(n_217),
.B2(n_241),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_278),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_310),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_273),
.B(n_282),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_271),
.C(n_264),
.Y(n_329)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_264),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_312),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_267),
.A2(n_242),
.B1(n_197),
.B2(n_171),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_266),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_317),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_271),
.A2(n_151),
.B1(n_153),
.B2(n_169),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_316),
.A2(n_274),
.B1(n_269),
.B2(n_281),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_284),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_320),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_291),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_322),
.B(n_333),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_302),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_325),
.B(n_327),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_316),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_330),
.C(n_331),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_271),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_300),
.B(n_277),
.Y(n_331)
);

OA21x2_ASAP7_75t_L g333 ( 
.A1(n_314),
.A2(n_259),
.B(n_268),
.Y(n_333)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_335),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_281),
.C(n_259),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_340),
.C(n_342),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_285),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_297),
.A2(n_314),
.B1(n_287),
.B2(n_292),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_341),
.A2(n_343),
.B1(n_344),
.B2(n_346),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_299),
.B(n_259),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_297),
.A2(n_263),
.B1(n_279),
.B2(n_266),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_289),
.A2(n_263),
.B1(n_270),
.B2(n_260),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_294),
.A2(n_260),
.B1(n_33),
.B2(n_174),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_328),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_347),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_321),
.A2(n_295),
.B1(n_310),
.B2(n_308),
.Y(n_348)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_348),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_328),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_349),
.A2(n_372),
.B1(n_326),
.B2(n_318),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_341),
.A2(n_303),
.B1(n_307),
.B2(n_313),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_350),
.A2(n_357),
.B1(n_365),
.B2(n_339),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_334),
.A2(n_288),
.B1(n_305),
.B2(n_293),
.Y(n_355)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_355),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_298),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_356),
.B(n_366),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_343),
.A2(n_306),
.B1(n_315),
.B2(n_179),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_337),
.Y(n_359)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_359),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_344),
.B(n_336),
.Y(n_360)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_360),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_322),
.A2(n_37),
.B(n_39),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_361),
.A2(n_40),
.B(n_9),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_336),
.A2(n_33),
.B1(n_15),
.B2(n_10),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_363),
.A2(n_371),
.B1(n_370),
.B2(n_368),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_10),
.Y(n_364)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_364),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_333),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_40),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_332),
.Y(n_367)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_367),
.Y(n_393)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_345),
.Y(n_368)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_368),
.Y(n_387)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_345),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_370),
.B(n_371),
.Y(n_379)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_326),
.Y(n_371)
);

NAND3xp33_ASAP7_75t_L g372 ( 
.A(n_320),
.B(n_10),
.C(n_9),
.Y(n_372)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_373),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_351),
.B(n_323),
.C(n_330),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_375),
.B(n_377),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_351),
.B(n_323),
.C(n_342),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_356),
.B(n_362),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_384),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_382),
.A2(n_394),
.B1(n_361),
.B2(n_367),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_369),
.A2(n_333),
.B(n_318),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_383),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_362),
.B(n_319),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_340),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_385),
.B(n_395),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_386),
.B(n_365),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_358),
.A2(n_324),
.B1(n_339),
.B2(n_346),
.Y(n_388)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_388),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_358),
.A2(n_335),
.B1(n_9),
.B2(n_2),
.Y(n_390)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_390),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_352),
.B(n_9),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_396),
.A2(n_409),
.B1(n_390),
.B2(n_389),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_375),
.B(n_380),
.C(n_377),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_399),
.B(n_403),
.Y(n_416)
);

XNOR2x1_ASAP7_75t_SL g401 ( 
.A(n_385),
.B(n_352),
.Y(n_401)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_401),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_354),
.C(n_369),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_379),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_405),
.B(n_406),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_376),
.B(n_354),
.C(n_366),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_350),
.C(n_353),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_408),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_391),
.B(n_393),
.C(n_381),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_378),
.B(n_363),
.C(n_1),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_410),
.B(n_411),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_392),
.B(n_0),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_374),
.B(n_0),
.C(n_1),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_413),
.B(n_0),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_383),
.C(n_386),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_415),
.B(n_420),
.Y(n_433)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_417),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_402),
.B(n_387),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_418),
.B(n_421),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_412),
.A2(n_379),
.B(n_387),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_388),
.C(n_382),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_400),
.B(n_395),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_422),
.B(n_424),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_396),
.B(n_394),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_412),
.A2(n_0),
.B(n_2),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_426),
.B(n_7),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_428),
.B(n_429),
.Y(n_436)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_397),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_2),
.C(n_3),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_430),
.B(n_7),
.C(n_4),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_415),
.A2(n_407),
.B(n_406),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_431),
.A2(n_434),
.B(n_419),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_417),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_432),
.B(n_438),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_416),
.A2(n_401),
.B(n_413),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_425),
.A2(n_414),
.B1(n_410),
.B2(n_398),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_398),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_439),
.B(n_440),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_441),
.B(n_427),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_424),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_442),
.B(n_444),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_3),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_446),
.B(n_437),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_447),
.A2(n_450),
.B(n_442),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_436),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_449),
.B(n_451),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_433),
.A2(n_419),
.B(n_430),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_435),
.B(n_422),
.C(n_424),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_422),
.Y(n_452)
);

AO21x1_ASAP7_75t_L g462 ( 
.A1(n_452),
.A2(n_453),
.B(n_455),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_426),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_443),
.B(n_3),
.Y(n_455)
);

AOI21x1_ASAP7_75t_L g464 ( 
.A1(n_456),
.A2(n_461),
.B(n_4),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_458),
.B(n_459),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_445),
.B(n_437),
.C(n_441),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_448),
.B(n_440),
.C(n_4),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_460),
.A2(n_4),
.B(n_5),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_3),
.Y(n_461)
);

OAI31xp33_ASAP7_75t_SL g463 ( 
.A1(n_462),
.A2(n_455),
.A3(n_454),
.B(n_6),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_463),
.A2(n_464),
.B(n_6),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_465),
.B(n_5),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_467),
.B(n_468),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_469),
.A2(n_457),
.B(n_466),
.Y(n_470)
);

AOI21x1_ASAP7_75t_L g471 ( 
.A1(n_470),
.A2(n_458),
.B(n_6),
.Y(n_471)
);

BUFx24_ASAP7_75t_SL g472 ( 
.A(n_471),
.Y(n_472)
);


endmodule