module real_aes_2658_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_785, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_785;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_769;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_733;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_691;
wire n_765;
wire n_498;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g159 ( .A(n_0), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_1), .B(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_2), .B(n_165), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_3), .B(n_162), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_4), .A2(n_43), .B1(n_435), .B2(n_436), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_4), .Y(n_435) );
INVx1_ASAP7_75t_L g125 ( .A(n_5), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_6), .B(n_165), .Y(n_187) );
NAND2xp33_ASAP7_75t_SL g145 ( .A(n_7), .B(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g116 ( .A(n_8), .Y(n_116) );
CKINVDCx16_ASAP7_75t_R g453 ( .A(n_9), .Y(n_453) );
AND2x2_ASAP7_75t_L g185 ( .A(n_10), .B(n_168), .Y(n_185) );
AND2x2_ASAP7_75t_L g488 ( .A(n_11), .B(n_141), .Y(n_488) );
AND2x2_ASAP7_75t_L g539 ( .A(n_12), .B(n_196), .Y(n_539) );
INVx2_ASAP7_75t_L g119 ( .A(n_13), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_14), .B(n_162), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_15), .Y(n_441) );
AOI221x1_ASAP7_75t_L g137 ( .A1(n_16), .A2(n_138), .B1(n_140), .B2(n_141), .C(n_144), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_17), .B(n_165), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_18), .B(n_165), .Y(n_544) );
INVx1_ASAP7_75t_L g445 ( .A(n_19), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_20), .A2(n_91), .B1(n_120), .B2(n_165), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_21), .A2(n_140), .B(n_189), .Y(n_188) );
AOI221xp5_ASAP7_75t_SL g232 ( .A1(n_22), .A2(n_35), .B1(n_140), .B2(n_165), .C(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_23), .B(n_160), .Y(n_190) );
OR2x2_ASAP7_75t_L g118 ( .A(n_24), .B(n_90), .Y(n_118) );
OA21x2_ASAP7_75t_L g143 ( .A1(n_24), .A2(n_90), .B(n_119), .Y(n_143) );
INVxp67_ASAP7_75t_L g136 ( .A(n_25), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_26), .B(n_162), .Y(n_227) );
AND2x2_ASAP7_75t_L g179 ( .A(n_27), .B(n_167), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_28), .A2(n_140), .B(n_158), .Y(n_157) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_29), .A2(n_141), .B(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_30), .B(n_162), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_31), .A2(n_140), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_32), .B(n_162), .Y(n_520) );
AND2x2_ASAP7_75t_L g127 ( .A(n_33), .B(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g131 ( .A(n_33), .Y(n_131) );
AND2x2_ASAP7_75t_L g146 ( .A(n_33), .B(n_125), .Y(n_146) );
OR2x6_ASAP7_75t_L g443 ( .A(n_34), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_36), .B(n_165), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_37), .A2(n_83), .B1(n_129), .B2(n_140), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_38), .B(n_162), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_39), .A2(n_48), .B1(n_767), .B2(n_768), .Y(n_766) );
INVx1_ASAP7_75t_L g768 ( .A(n_39), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_40), .B(n_165), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_41), .B(n_160), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_42), .A2(n_140), .B(n_484), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_43), .Y(n_436) );
AND2x2_ASAP7_75t_L g166 ( .A(n_44), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_45), .B(n_160), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_46), .B(n_167), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_47), .B(n_165), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_48), .Y(n_767) );
INVx1_ASAP7_75t_L g123 ( .A(n_49), .Y(n_123) );
INVx1_ASAP7_75t_L g150 ( .A(n_49), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_50), .B(n_162), .Y(n_486) );
AND2x2_ASAP7_75t_L g498 ( .A(n_51), .B(n_167), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_52), .B(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_53), .B(n_165), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_54), .B(n_160), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_55), .B(n_160), .Y(n_519) );
AND2x2_ASAP7_75t_L g208 ( .A(n_56), .B(n_167), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_57), .B(n_165), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_58), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_59), .B(n_165), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_60), .A2(n_140), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_61), .B(n_160), .Y(n_206) );
AND2x2_ASAP7_75t_SL g228 ( .A(n_62), .B(n_168), .Y(n_228) );
XNOR2xp5_ASAP7_75t_L g765 ( .A(n_63), .B(n_766), .Y(n_765) );
AOI221xp5_ASAP7_75t_L g103 ( .A1(n_64), .A2(n_104), .B1(n_450), .B2(n_455), .C(n_461), .Y(n_103) );
XNOR2x1_ASAP7_75t_SL g105 ( .A(n_64), .B(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g550 ( .A(n_64), .B(n_168), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_65), .A2(n_140), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_66), .B(n_162), .Y(n_191) );
AND2x2_ASAP7_75t_SL g200 ( .A(n_67), .B(n_196), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_68), .B(n_160), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_69), .B(n_160), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_70), .A2(n_93), .B1(n_129), .B2(n_140), .Y(n_493) );
XNOR2xp5_ASAP7_75t_L g764 ( .A(n_71), .B(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_SL g773 ( .A(n_72), .B(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_73), .B(n_162), .Y(n_547) );
INVx1_ASAP7_75t_L g128 ( .A(n_74), .Y(n_128) );
INVx1_ASAP7_75t_L g152 ( .A(n_74), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_75), .B(n_160), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_76), .A2(n_140), .B(n_502), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_77), .A2(n_140), .B(n_476), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_78), .A2(n_140), .B(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g522 ( .A(n_79), .B(n_168), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_80), .B(n_167), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_81), .A2(n_85), .B1(n_120), .B2(n_165), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_82), .B(n_165), .Y(n_207) );
INVx1_ASAP7_75t_L g446 ( .A(n_84), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_86), .B(n_160), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_87), .B(n_160), .Y(n_235) );
AND2x2_ASAP7_75t_L g479 ( .A(n_88), .B(n_196), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_89), .A2(n_140), .B(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_92), .B(n_162), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_94), .A2(n_140), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_95), .B(n_162), .Y(n_477) );
OAI22x1_ASAP7_75t_R g432 ( .A1(n_96), .A2(n_433), .B1(n_434), .B2(n_437), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_96), .Y(n_437) );
INVxp67_ASAP7_75t_L g139 ( .A(n_97), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_98), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_99), .B(n_162), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_100), .A2(n_140), .B(n_225), .Y(n_224) );
BUFx2_ASAP7_75t_L g549 ( .A(n_101), .Y(n_549) );
BUFx2_ASAP7_75t_L g454 ( .A(n_102), .Y(n_454) );
BUFx2_ASAP7_75t_SL g459 ( .A(n_102), .Y(n_459) );
OAI21xp33_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_438), .B(n_447), .Y(n_104) );
OAI22x1_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_108), .B1(n_431), .B2(n_432), .Y(n_106) );
OAI22x1_ASAP7_75t_L g463 ( .A1(n_107), .A2(n_464), .B1(n_466), .B2(n_761), .Y(n_463) );
INVx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OA22x2_ASAP7_75t_L g771 ( .A1(n_108), .A2(n_464), .B1(n_467), .B2(n_772), .Y(n_771) );
AND2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_308), .Y(n_108) );
NOR4xp25_ASAP7_75t_L g109 ( .A(n_110), .B(n_251), .C(n_290), .D(n_297), .Y(n_109) );
OAI221xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_169), .B1(n_209), .B2(n_218), .C(n_237), .Y(n_110) );
OR2x2_ASAP7_75t_L g381 ( .A(n_111), .B(n_243), .Y(n_381) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g296 ( .A(n_112), .B(n_221), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_112), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_SL g361 ( .A(n_112), .B(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_L g112 ( .A(n_113), .B(n_153), .Y(n_112) );
AND2x4_ASAP7_75t_SL g220 ( .A(n_113), .B(n_221), .Y(n_220) );
INVx3_ASAP7_75t_L g242 ( .A(n_113), .Y(n_242) );
AND2x2_ASAP7_75t_L g277 ( .A(n_113), .B(n_250), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_113), .B(n_154), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_113), .B(n_244), .Y(n_329) );
OR2x2_ASAP7_75t_L g407 ( .A(n_113), .B(n_221), .Y(n_407) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_137), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B1(n_129), .B2(n_135), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_117), .B(n_136), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_117), .B(n_139), .Y(n_138) );
NOR3xp33_ASAP7_75t_L g144 ( .A(n_117), .B(n_145), .C(n_147), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_117), .A2(n_187), .B(n_188), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_117), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_117), .A2(n_509), .B(n_510), .Y(n_508) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
AND2x2_ASAP7_75t_SL g168 ( .A(n_118), .B(n_119), .Y(n_168) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_126), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_124), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g134 ( .A(n_123), .B(n_125), .Y(n_134) );
AND2x4_ASAP7_75t_L g162 ( .A(n_123), .B(n_151), .Y(n_162) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x6_ASAP7_75t_L g140 ( .A(n_127), .B(n_134), .Y(n_140) );
INVx2_ASAP7_75t_L g133 ( .A(n_128), .Y(n_133) );
AND2x6_ASAP7_75t_L g160 ( .A(n_128), .B(n_149), .Y(n_160) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_134), .Y(n_129) );
NOR2x1p5_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx3_ASAP7_75t_L g515 ( .A(n_141), .Y(n_515) );
INVx4_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AOI21x1_ASAP7_75t_L g155 ( .A1(n_142), .A2(n_156), .B(n_166), .Y(n_155) );
AO21x2_ASAP7_75t_L g481 ( .A1(n_142), .A2(n_482), .B(n_488), .Y(n_481) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx4f_ASAP7_75t_L g196 ( .A(n_143), .Y(n_196) );
INVx5_ASAP7_75t_L g163 ( .A(n_146), .Y(n_163) );
AND2x4_ASAP7_75t_L g165 ( .A(n_146), .B(n_148), .Y(n_165) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g229 ( .A(n_154), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_154), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g255 ( .A(n_154), .Y(n_255) );
OR2x2_ASAP7_75t_L g260 ( .A(n_154), .B(n_244), .Y(n_260) );
AND2x2_ASAP7_75t_L g273 ( .A(n_154), .B(n_231), .Y(n_273) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_154), .Y(n_276) );
INVx1_ASAP7_75t_L g288 ( .A(n_154), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_154), .B(n_242), .Y(n_353) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_164), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_161), .B(n_163), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_160), .B(n_549), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_163), .A2(n_175), .B(n_176), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_163), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_163), .A2(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_163), .A2(n_226), .B(n_227), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_163), .A2(n_234), .B(n_235), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_163), .A2(n_477), .B(n_478), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_163), .A2(n_485), .B(n_486), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_163), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_163), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_163), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_163), .A2(n_536), .B(n_537), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_163), .A2(n_547), .B(n_548), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_167), .Y(n_178) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_167), .A2(n_232), .B(n_236), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_167), .A2(n_474), .B(n_475), .Y(n_473) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_167), .A2(n_492), .B(n_493), .Y(n_491) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_170), .B(n_180), .Y(n_169) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OR2x2_ASAP7_75t_L g217 ( .A(n_171), .B(n_201), .Y(n_217) );
AND2x4_ASAP7_75t_L g247 ( .A(n_171), .B(n_184), .Y(n_247) );
INVx2_ASAP7_75t_L g281 ( .A(n_171), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_171), .B(n_201), .Y(n_339) );
AND2x2_ASAP7_75t_L g386 ( .A(n_171), .B(n_215), .Y(n_386) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_178), .B(n_179), .Y(n_171) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_172), .A2(n_178), .B(n_179), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_177), .Y(n_172) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_178), .A2(n_202), .B(n_208), .Y(n_201) );
AOI21x1_ASAP7_75t_L g532 ( .A1(n_178), .A2(n_533), .B(n_539), .Y(n_532) );
AOI222xp33_ASAP7_75t_L g374 ( .A1(n_180), .A2(n_246), .B1(n_289), .B2(n_349), .C1(n_375), .C2(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_192), .Y(n_181) );
AND2x2_ASAP7_75t_L g293 ( .A(n_182), .B(n_213), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_182), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g422 ( .A(n_182), .B(n_262), .Y(n_422) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_183), .A2(n_253), .B(n_257), .Y(n_252) );
AND2x2_ASAP7_75t_L g333 ( .A(n_183), .B(n_216), .Y(n_333) );
OR2x2_ASAP7_75t_L g358 ( .A(n_183), .B(n_217), .Y(n_358) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx5_ASAP7_75t_L g212 ( .A(n_184), .Y(n_212) );
AND2x2_ASAP7_75t_L g299 ( .A(n_184), .B(n_281), .Y(n_299) );
AND2x2_ASAP7_75t_L g325 ( .A(n_184), .B(n_201), .Y(n_325) );
OR2x2_ASAP7_75t_L g328 ( .A(n_184), .B(n_215), .Y(n_328) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_184), .Y(n_346) );
AND2x4_ASAP7_75t_SL g403 ( .A(n_184), .B(n_280), .Y(n_403) );
OR2x2_ASAP7_75t_L g412 ( .A(n_184), .B(n_239), .Y(n_412) );
OR2x6_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
INVx1_ASAP7_75t_L g245 ( .A(n_192), .Y(n_245) );
AOI221xp5_ASAP7_75t_SL g363 ( .A1(n_192), .A2(n_247), .B1(n_364), .B2(n_366), .C(n_367), .Y(n_363) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_201), .Y(n_192) );
OR2x2_ASAP7_75t_L g302 ( .A(n_193), .B(n_272), .Y(n_302) );
OR2x2_ASAP7_75t_L g312 ( .A(n_193), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g338 ( .A(n_193), .B(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g344 ( .A(n_193), .B(n_263), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_193), .B(n_327), .Y(n_356) );
INVx2_ASAP7_75t_L g369 ( .A(n_193), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_193), .B(n_247), .Y(n_390) );
AND2x2_ASAP7_75t_L g394 ( .A(n_193), .B(n_216), .Y(n_394) );
AND2x2_ASAP7_75t_L g402 ( .A(n_193), .B(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g215 ( .A(n_194), .Y(n_215) );
AOI21x1_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_197), .B(n_200), .Y(n_194) );
INVx2_ASAP7_75t_SL g195 ( .A(n_196), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_196), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_196), .A2(n_544), .B(n_545), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_201), .B(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g246 ( .A(n_201), .B(n_215), .Y(n_246) );
INVx2_ASAP7_75t_L g263 ( .A(n_201), .Y(n_263) );
AND2x4_ASAP7_75t_L g280 ( .A(n_201), .B(n_281), .Y(n_280) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_201), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_207), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_213), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
OR2x2_ASAP7_75t_L g392 ( .A(n_211), .B(n_214), .Y(n_392) );
AND2x4_ASAP7_75t_L g238 ( .A(n_212), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g279 ( .A(n_212), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g306 ( .A(n_212), .B(n_246), .Y(n_306) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_216), .Y(n_213) );
AND2x2_ASAP7_75t_L g410 ( .A(n_214), .B(n_411), .Y(n_410) );
BUFx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g262 ( .A(n_215), .B(n_263), .Y(n_262) );
OAI21xp5_ASAP7_75t_SL g282 ( .A1(n_216), .A2(n_283), .B(n_289), .Y(n_282) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_229), .Y(n_219) );
INVx1_ASAP7_75t_SL g336 ( .A(n_220), .Y(n_336) );
AND2x2_ASAP7_75t_L g366 ( .A(n_220), .B(n_276), .Y(n_366) );
AND2x4_ASAP7_75t_L g377 ( .A(n_220), .B(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g243 ( .A(n_221), .B(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g250 ( .A(n_221), .Y(n_250) );
AND2x4_ASAP7_75t_L g256 ( .A(n_221), .B(n_242), .Y(n_256) );
INVx2_ASAP7_75t_L g267 ( .A(n_221), .Y(n_267) );
INVx1_ASAP7_75t_L g316 ( .A(n_221), .Y(n_316) );
OR2x2_ASAP7_75t_L g337 ( .A(n_221), .B(n_321), .Y(n_337) );
OR2x2_ASAP7_75t_L g351 ( .A(n_221), .B(n_231), .Y(n_351) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_221), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_221), .B(n_273), .Y(n_423) );
OR2x6_ASAP7_75t_L g221 ( .A(n_222), .B(n_228), .Y(n_221) );
INVx1_ASAP7_75t_L g268 ( .A(n_229), .Y(n_268) );
AND2x2_ASAP7_75t_L g401 ( .A(n_229), .B(n_267), .Y(n_401) );
AND2x2_ASAP7_75t_L g426 ( .A(n_229), .B(n_256), .Y(n_426) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g244 ( .A(n_231), .Y(n_244) );
BUFx3_ASAP7_75t_L g286 ( .A(n_231), .Y(n_286) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_231), .Y(n_313) );
INVx1_ASAP7_75t_L g322 ( .A(n_231), .Y(n_322) );
AOI33xp33_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_240), .A3(n_245), .B1(n_246), .B2(n_247), .B3(n_248), .Y(n_237) );
AOI21x1_ASAP7_75t_SL g340 ( .A1(n_238), .A2(n_262), .B(n_324), .Y(n_340) );
INVx2_ASAP7_75t_L g370 ( .A(n_238), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_238), .B(n_369), .Y(n_376) );
AND2x2_ASAP7_75t_L g324 ( .A(n_239), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
AND2x2_ASAP7_75t_L g287 ( .A(n_242), .B(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g388 ( .A(n_243), .Y(n_388) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_244), .Y(n_378) );
OAI32xp33_ASAP7_75t_L g427 ( .A1(n_245), .A2(n_247), .A3(n_423), .B1(n_428), .B2(n_430), .Y(n_427) );
AND2x2_ASAP7_75t_L g345 ( .A(n_246), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_SL g335 ( .A(n_247), .Y(n_335) );
AND2x2_ASAP7_75t_L g400 ( .A(n_247), .B(n_344), .Y(n_400) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OAI221xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_261), .B1(n_264), .B2(n_278), .C(n_282), .Y(n_251) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_255), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_256), .B(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_256), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_256), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g305 ( .A(n_260), .Y(n_305) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NOR3xp33_ASAP7_75t_L g264 ( .A(n_265), .B(n_269), .C(n_274), .Y(n_264) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
OAI22xp33_ASAP7_75t_L g367 ( .A1(n_266), .A2(n_328), .B1(n_368), .B2(n_371), .Y(n_367) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx1_ASAP7_75t_L g271 ( .A(n_267), .Y(n_271) );
NOR2x1p5_ASAP7_75t_L g285 ( .A(n_267), .B(n_286), .Y(n_285) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_267), .Y(n_307) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OAI322xp33_ASAP7_75t_L g334 ( .A1(n_270), .A2(n_312), .A3(n_335), .B1(n_336), .B2(n_337), .C1(n_338), .C2(n_340), .Y(n_334) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_272), .A2(n_291), .B(n_292), .C(n_294), .Y(n_290) );
OR2x2_ASAP7_75t_L g382 ( .A(n_272), .B(n_336), .Y(n_382) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g289 ( .A(n_273), .B(n_277), .Y(n_289) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g295 ( .A(n_279), .B(n_296), .Y(n_295) );
INVx3_ASAP7_75t_SL g327 ( .A(n_280), .Y(n_327) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_284), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx1_ASAP7_75t_SL g331 ( .A(n_287), .Y(n_331) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_288), .Y(n_373) );
OR2x6_ASAP7_75t_SL g428 ( .A(n_291), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVxp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AOI211xp5_ASAP7_75t_L g418 ( .A1(n_296), .A2(n_419), .B(n_420), .C(n_427), .Y(n_418) );
O2A1O1Ixp33_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_300), .B(n_303), .C(n_307), .Y(n_297) );
OAI211xp5_ASAP7_75t_SL g309 ( .A1(n_298), .A2(n_310), .B(n_317), .C(n_341), .Y(n_309) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVxp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
NOR3xp33_ASAP7_75t_L g308 ( .A(n_309), .B(n_354), .C(n_398), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_314), .Y(n_310) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_313), .Y(n_405) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g360 ( .A(n_316), .Y(n_360) );
NOR3xp33_ASAP7_75t_SL g317 ( .A(n_318), .B(n_330), .C(n_334), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_323), .B1(n_326), .B2(n_329), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g362 ( .A(n_322), .Y(n_362) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_322), .Y(n_429) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx1_ASAP7_75t_SL g415 ( .A(n_328), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
OR2x2_ASAP7_75t_L g365 ( .A(n_331), .B(n_351), .Y(n_365) );
OR2x2_ASAP7_75t_L g416 ( .A(n_331), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g414 ( .A(n_339), .Y(n_414) );
OR2x2_ASAP7_75t_L g430 ( .A(n_339), .B(n_369), .Y(n_430) );
OAI21xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_345), .B(n_347), .Y(n_341) );
OAI31xp33_ASAP7_75t_L g355 ( .A1(n_342), .A2(n_356), .A3(n_357), .B(n_359), .Y(n_355) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g387 ( .A(n_352), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND4xp25_ASAP7_75t_SL g354 ( .A(n_355), .B(n_363), .C(n_374), .D(n_379), .Y(n_354) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_362), .Y(n_397) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_383), .B1(n_387), .B2(n_389), .C(n_391), .Y(n_379) );
NAND2xp33_ASAP7_75t_SL g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_L g424 ( .A(n_383), .Y(n_424) );
AND2x2_ASAP7_75t_SL g383 ( .A(n_384), .B(n_386), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI21xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B(n_395), .Y(n_391) );
INVx1_ASAP7_75t_L g419 ( .A(n_393), .Y(n_419) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_399), .B(n_418), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_402), .B2(n_404), .C(n_408), .Y(n_399) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
AOI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_413), .B(n_416), .Y(n_408) );
INVxp33_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_423), .B1(n_424), .B2(n_425), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVxp33_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx2_ASAP7_75t_R g439 ( .A(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_L g449 ( .A(n_440), .Y(n_449) );
BUFx2_ASAP7_75t_L g783 ( .A(n_440), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
AND2x6_ASAP7_75t_SL g465 ( .A(n_441), .B(n_443), .Y(n_465) );
OR2x6_ASAP7_75t_SL g763 ( .A(n_441), .B(n_442), .Y(n_763) );
OR2x2_ASAP7_75t_L g777 ( .A(n_441), .B(n_443), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g460 ( .A(n_449), .Y(n_460) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_SL g451 ( .A(n_452), .B(n_454), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_452), .A2(n_457), .B(n_460), .Y(n_456) );
INVx2_ASAP7_75t_L g782 ( .A(n_452), .Y(n_782) );
NAND2xp5_ASAP7_75t_SL g781 ( .A(n_454), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
CKINVDCx11_ASAP7_75t_R g457 ( .A(n_458), .Y(n_457) );
CKINVDCx8_ASAP7_75t_R g458 ( .A(n_459), .Y(n_458) );
AOI31xp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_769), .A3(n_773), .B(n_778), .Y(n_461) );
NAND2xp33_ASAP7_75t_SL g462 ( .A(n_463), .B(n_764), .Y(n_462) );
CKINVDCx11_ASAP7_75t_R g464 ( .A(n_465), .Y(n_464) );
INVx3_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
AND2x4_ASAP7_75t_SL g467 ( .A(n_468), .B(n_657), .Y(n_467) );
NOR3xp33_ASAP7_75t_SL g468 ( .A(n_469), .B(n_566), .C(n_598), .Y(n_468) );
OAI221xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_494), .B1(n_523), .B2(n_540), .C(n_551), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_480), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g529 ( .A(n_472), .B(n_481), .Y(n_529) );
INVx4_ASAP7_75t_L g557 ( .A(n_472), .Y(n_557) );
AND2x4_ASAP7_75t_SL g597 ( .A(n_472), .B(n_531), .Y(n_597) );
BUFx2_ASAP7_75t_L g607 ( .A(n_472), .Y(n_607) );
NOR2x1_ASAP7_75t_L g673 ( .A(n_472), .B(n_612), .Y(n_673) );
AND2x2_ASAP7_75t_L g682 ( .A(n_472), .B(n_610), .Y(n_682) );
OR2x2_ASAP7_75t_L g690 ( .A(n_472), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g716 ( .A(n_472), .B(n_555), .Y(n_716) );
AND2x4_ASAP7_75t_L g735 ( .A(n_472), .B(n_736), .Y(n_735) );
OR2x6_ASAP7_75t_L g472 ( .A(n_473), .B(n_479), .Y(n_472) );
INVx2_ASAP7_75t_SL g648 ( .A(n_480), .Y(n_648) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_489), .Y(n_480) );
AND2x2_ASAP7_75t_L g555 ( .A(n_481), .B(n_532), .Y(n_555) );
INVx2_ASAP7_75t_L g582 ( .A(n_481), .Y(n_582) );
INVx2_ASAP7_75t_L g612 ( .A(n_481), .Y(n_612) );
AND2x2_ASAP7_75t_L g626 ( .A(n_481), .B(n_531), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_487), .Y(n_482) );
AND2x2_ASAP7_75t_L g556 ( .A(n_489), .B(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g579 ( .A(n_489), .Y(n_579) );
BUFx3_ASAP7_75t_L g593 ( .A(n_489), .Y(n_593) );
AND2x2_ASAP7_75t_L g622 ( .A(n_489), .B(n_623), .Y(n_622) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
AND2x4_ASAP7_75t_L g527 ( .A(n_490), .B(n_491), .Y(n_527) );
INVx1_ASAP7_75t_L g628 ( .A(n_494), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_505), .Y(n_494) );
OR2x2_ASAP7_75t_L g739 ( .A(n_495), .B(n_540), .Y(n_739) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g595 ( .A(n_496), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_496), .B(n_505), .Y(n_656) );
OR2x2_ASAP7_75t_L g754 ( .A(n_496), .B(n_676), .Y(n_754) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g565 ( .A(n_497), .B(n_541), .Y(n_565) );
OR2x2_ASAP7_75t_SL g575 ( .A(n_497), .B(n_576), .Y(n_575) );
INVx4_ASAP7_75t_L g586 ( .A(n_497), .Y(n_586) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_497), .Y(n_637) );
NAND2x1_ASAP7_75t_L g643 ( .A(n_497), .B(n_542), .Y(n_643) );
AND2x2_ASAP7_75t_L g668 ( .A(n_497), .B(n_507), .Y(n_668) );
OR2x2_ASAP7_75t_L g689 ( .A(n_497), .B(n_572), .Y(n_689) );
OR2x6_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g584 ( .A(n_505), .Y(n_584) );
O2A1O1Ixp33_ASAP7_75t_L g677 ( .A1(n_505), .A2(n_678), .B(n_681), .C(n_683), .Y(n_677) );
AND2x2_ASAP7_75t_L g750 ( .A(n_505), .B(n_526), .Y(n_750) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_514), .Y(n_505) );
INVx1_ASAP7_75t_L g617 ( .A(n_506), .Y(n_617) );
AND2x2_ASAP7_75t_L g687 ( .A(n_506), .B(n_542), .Y(n_687) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g561 ( .A(n_507), .Y(n_561) );
OR2x2_ASAP7_75t_L g576 ( .A(n_507), .B(n_542), .Y(n_576) );
INVx1_ASAP7_75t_L g592 ( .A(n_507), .Y(n_592) );
AND2x2_ASAP7_75t_L g604 ( .A(n_507), .B(n_514), .Y(n_604) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_507), .Y(n_710) );
NOR2x1_ASAP7_75t_SL g541 ( .A(n_514), .B(n_542), .Y(n_541) );
AO21x1_ASAP7_75t_SL g514 ( .A1(n_515), .A2(n_516), .B(n_522), .Y(n_514) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_515), .A2(n_516), .B(n_522), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_521), .Y(n_516) );
INVxp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_528), .Y(n_524) );
OR2x2_ASAP7_75t_L g674 ( .A(n_525), .B(n_609), .Y(n_674) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_526), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g756 ( .A(n_526), .B(n_653), .Y(n_756) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g601 ( .A(n_527), .B(n_582), .Y(n_601) );
AND2x2_ASAP7_75t_L g697 ( .A(n_527), .B(n_610), .Y(n_697) );
INVx1_ASAP7_75t_L g614 ( .A(n_528), .Y(n_614) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g664 ( .A(n_529), .Y(n_664) );
INVx2_ASAP7_75t_L g631 ( .A(n_530), .Y(n_631) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g581 ( .A(n_531), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g611 ( .A(n_531), .Y(n_611) );
INVx1_ASAP7_75t_L g736 ( .A(n_531), .Y(n_736) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_532), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_538), .Y(n_533) );
OR2x2_ASAP7_75t_L g707 ( .A(n_540), .B(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_SL g562 ( .A(n_542), .Y(n_562) );
OR2x2_ASAP7_75t_L g585 ( .A(n_542), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g596 ( .A(n_542), .B(n_572), .Y(n_596) );
AND2x2_ASAP7_75t_L g670 ( .A(n_542), .B(n_586), .Y(n_670) );
BUFx2_ASAP7_75t_L g753 ( .A(n_542), .Y(n_753) );
OR2x6_ASAP7_75t_L g542 ( .A(n_543), .B(n_550), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_558), .B(n_563), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
AND2x2_ASAP7_75t_L g705 ( .A(n_554), .B(n_627), .Y(n_705) );
BUFx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g564 ( .A(n_555), .B(n_557), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_556), .B(n_626), .Y(n_727) );
INVx1_ASAP7_75t_L g757 ( .A(n_556), .Y(n_757) );
NAND2x1p5_ASAP7_75t_L g653 ( .A(n_557), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_557), .B(n_693), .Y(n_730) );
INVxp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
AND2x4_ASAP7_75t_SL g594 ( .A(n_560), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_560), .B(n_588), .Y(n_741) );
INVx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_561), .B(n_643), .Y(n_699) );
AND2x2_ASAP7_75t_L g717 ( .A(n_561), .B(n_670), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_562), .B(n_604), .Y(n_620) );
A2O1A1Ixp33_ASAP7_75t_L g649 ( .A1(n_562), .A2(n_608), .B(n_650), .C(n_655), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_562), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g744 ( .A1(n_564), .A2(n_637), .B1(n_745), .B2(n_751), .C(n_755), .Y(n_744) );
INVx1_ASAP7_75t_SL g732 ( .A(n_565), .Y(n_732) );
OAI221xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_577), .B1(n_583), .B2(n_587), .C(n_785), .Y(n_566) );
INVx2_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
AND2x4_ASAP7_75t_L g568 ( .A(n_569), .B(n_574), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g642 ( .A(n_571), .Y(n_642) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g616 ( .A(n_572), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g647 ( .A(n_572), .B(n_592), .Y(n_647) );
INVx2_ASAP7_75t_L g680 ( .A(n_572), .Y(n_680) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI32xp33_ASAP7_75t_L g731 ( .A1(n_575), .A2(n_622), .A3(n_653), .B1(n_732), .B2(n_733), .Y(n_731) );
OR2x2_ASAP7_75t_L g702 ( .A(n_576), .B(n_689), .Y(n_702) );
INVx1_ASAP7_75t_L g712 ( .A(n_577), .Y(n_712) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
INVx2_ASAP7_75t_L g627 ( .A(n_578), .Y(n_627) );
AND2x2_ASAP7_75t_L g698 ( .A(n_578), .B(n_673), .Y(n_698) );
OR2x2_ASAP7_75t_L g729 ( .A(n_578), .B(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_579), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g623 ( .A(n_582), .Y(n_623) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx2_ASAP7_75t_SL g588 ( .A(n_585), .Y(n_588) );
OR2x2_ASAP7_75t_L g675 ( .A(n_585), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_586), .B(n_604), .Y(n_603) );
NOR2xp67_ASAP7_75t_L g709 ( .A(n_586), .B(n_710), .Y(n_709) );
BUFx2_ASAP7_75t_L g722 ( .A(n_586), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B(n_594), .C(n_597), .Y(n_587) );
AND2x2_ASAP7_75t_L g737 ( .A(n_589), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
BUFx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g663 ( .A(n_593), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_593), .B(n_597), .Y(n_684) );
AND2x2_ASAP7_75t_L g715 ( .A(n_593), .B(n_716), .Y(n_715) );
O2A1O1Ixp33_ASAP7_75t_L g725 ( .A1(n_595), .A2(n_726), .B(n_728), .C(n_731), .Y(n_725) );
AOI222xp33_ASAP7_75t_L g599 ( .A1(n_596), .A2(n_600), .B1(n_602), .B2(n_605), .C1(n_613), .C2(n_615), .Y(n_599) );
AND2x2_ASAP7_75t_L g667 ( .A(n_596), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g600 ( .A(n_597), .B(n_601), .Y(n_600) );
INVx2_ASAP7_75t_SL g621 ( .A(n_597), .Y(n_621) );
NAND4xp25_ASAP7_75t_L g598 ( .A(n_599), .B(n_618), .C(n_639), .D(n_649), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_601), .B(n_607), .Y(n_661) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g669 ( .A(n_604), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_SL g676 ( .A(n_604), .Y(n_676) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
A2O1A1Ixp33_ASAP7_75t_L g639 ( .A1(n_606), .A2(n_640), .B(n_644), .C(n_648), .Y(n_639) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_607), .B(n_622), .Y(n_743) );
OR2x2_ASAP7_75t_L g747 ( .A(n_607), .B(n_633), .Y(n_747) );
INVx1_ASAP7_75t_L g720 ( .A(n_608), .Y(n_720) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_SL g654 ( .A(n_611), .Y(n_654) );
INVx1_ASAP7_75t_L g634 ( .A(n_612), .Y(n_634) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_614), .B(n_651), .Y(n_650) );
BUFx2_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g638 ( .A(n_616), .Y(n_638) );
AOI322xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_621), .A3(n_622), .B1(n_624), .B2(n_628), .C1(n_629), .C2(n_635), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
O2A1O1Ixp33_ASAP7_75t_SL g700 ( .A1(n_621), .A2(n_701), .B(n_702), .C(n_703), .Y(n_700) );
INVx1_ASAP7_75t_L g723 ( .A(n_622), .Y(n_723) );
NOR2xp67_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g681 ( .A(n_627), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_633), .Y(n_703) );
INVx2_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
INVx3_ASAP7_75t_L g646 ( .A(n_643), .Y(n_646) );
OR2x2_ASAP7_75t_L g714 ( .A(n_643), .B(n_676), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_643), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx1_ASAP7_75t_SL g746 ( .A(n_647), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_648), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND3xp33_ASAP7_75t_SL g751 ( .A(n_656), .B(n_752), .C(n_754), .Y(n_751) );
NOR3xp33_ASAP7_75t_SL g657 ( .A(n_658), .B(n_695), .C(n_724), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_659), .B(n_677), .Y(n_658) );
O2A1O1Ixp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_662), .B(n_665), .C(n_671), .Y(n_659) );
OAI31xp33_ASAP7_75t_L g704 ( .A1(n_660), .A2(n_682), .A3(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
INVx2_ASAP7_75t_L g719 ( .A(n_667), .Y(n_719) );
INVx1_ASAP7_75t_L g694 ( .A(n_669), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_674), .B(n_675), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g721 ( .A(n_679), .B(n_722), .Y(n_721) );
INVxp67_ASAP7_75t_L g760 ( .A(n_680), .Y(n_760) );
OAI22xp33_ASAP7_75t_SL g683 ( .A1(n_684), .A2(n_685), .B1(n_690), .B2(n_694), .Y(n_683) );
INVx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x4_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_689), .Y(n_701) );
OR2x2_ASAP7_75t_L g752 ( .A(n_689), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND3xp33_ASAP7_75t_SL g695 ( .A(n_696), .B(n_704), .C(n_711), .Y(n_695) );
O2A1O1Ixp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B(n_699), .C(n_700), .Y(n_696) );
INVx2_ASAP7_75t_L g733 ( .A(n_697), .Y(n_733) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_713), .B1(n_715), .B2(n_717), .C(n_718), .Y(n_711) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI22xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .B1(n_721), .B2(n_723), .Y(n_718) );
NAND3xp33_ASAP7_75t_SL g724 ( .A(n_725), .B(n_734), .C(n_744), .Y(n_724) );
INVxp33_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_737), .B1(n_740), .B2(n_742), .Y(n_734) );
INVx2_ASAP7_75t_L g748 ( .A(n_735), .Y(n_748) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B1(n_748), .B2(n_749), .Y(n_745) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
OAI22xp33_ASAP7_75t_SL g755 ( .A1(n_754), .A2(n_756), .B1(n_757), .B2(n_758), .Y(n_755) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
BUFx4f_ASAP7_75t_SL g772 ( .A(n_761), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_762), .Y(n_761) );
CKINVDCx11_ASAP7_75t_R g762 ( .A(n_763), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_764), .B(n_771), .Y(n_770) );
INVxp33_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx2_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
INVx3_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_783), .Y(n_779) );
INVxp67_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
endmodule