module fake_jpeg_24911_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_10),
.B(n_12),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g64 ( 
.A(n_37),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_0),
.B(n_1),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_38),
.A2(n_44),
.B(n_0),
.Y(n_68)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NAND3xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_28),
.C(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_R g49 ( 
.A(n_44),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_71),
.Y(n_88)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_70),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_22),
.B1(n_19),
.B2(n_33),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_49),
.B1(n_59),
.B2(n_66),
.Y(n_76)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_59),
.B(n_34),
.Y(n_82)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_63),
.A2(n_65),
.B1(n_27),
.B2(n_17),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_12),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_21),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_23),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_74),
.B(n_81),
.Y(n_136)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_75),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_76),
.A2(n_103),
.B1(n_50),
.B2(n_60),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_39),
.B1(n_30),
.B2(n_29),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_78),
.A2(n_90),
.B1(n_95),
.B2(n_107),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_71),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_80),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_23),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_82),
.B(n_100),
.Y(n_118)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_32),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_84),
.B(n_93),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_34),
.B1(n_18),
.B2(n_20),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_85),
.A2(n_98),
.B1(n_99),
.B2(n_0),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_45),
.B(n_42),
.C(n_41),
.Y(n_87)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_89),
.A2(n_105),
.B1(n_113),
.B2(n_114),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_30),
.B1(n_17),
.B2(n_27),
.Y(n_90)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_32),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_53),
.A2(n_27),
.B1(n_29),
.B2(n_26),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_64),
.A2(n_45),
.B(n_42),
.C(n_29),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_62),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_62),
.A2(n_32),
.B(n_16),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_4),
.C(n_5),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_51),
.A2(n_16),
.B1(n_20),
.B2(n_26),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_52),
.B(n_32),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_106),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_62),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_72),
.B(n_16),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_28),
.B1(n_30),
.B2(n_56),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_73),
.A2(n_30),
.B1(n_14),
.B2(n_26),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_62),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_50),
.B(n_32),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_50),
.C(n_45),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_70),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_117),
.A2(n_120),
.B1(n_130),
.B2(n_132),
.Y(n_159)
);

NAND2xp33_ASAP7_75t_SL g119 ( 
.A(n_74),
.B(n_32),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_119),
.A2(n_125),
.B(n_144),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_76),
.A2(n_80),
.B1(n_99),
.B2(n_88),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_52),
.B1(n_29),
.B2(n_26),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_139),
.B1(n_106),
.B2(n_86),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_42),
.C(n_52),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_104),
.Y(n_157)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_96),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_88),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_88),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_137),
.B1(n_141),
.B2(n_143),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_90),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

AOI22x1_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_81),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_146),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_140),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_83),
.B(n_86),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_147),
.A2(n_152),
.B(n_166),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_82),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_157),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_149),
.Y(n_202)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_151),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

OA21x2_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_113),
.B(n_87),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_153),
.A2(n_164),
.B1(n_171),
.B2(n_173),
.Y(n_199)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_155),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_112),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_161),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g158 ( 
.A(n_136),
.B(n_93),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_158),
.A2(n_175),
.B(n_177),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_112),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_133),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_165),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_122),
.B1(n_123),
.B2(n_133),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_163),
.A2(n_156),
.B1(n_165),
.B2(n_147),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_123),
.A2(n_110),
.B1(n_114),
.B2(n_91),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_136),
.A2(n_92),
.B(n_105),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_137),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_172),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_97),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_170),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_120),
.B(n_103),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_139),
.A2(n_119),
.B1(n_115),
.B2(n_125),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_115),
.A2(n_144),
.B1(n_135),
.B2(n_142),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_135),
.B(n_134),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_77),
.Y(n_176)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_100),
.B(n_77),
.Y(n_177)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_193),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_167),
.A2(n_129),
.B1(n_111),
.B2(n_126),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_SL g233 ( 
.A1(n_181),
.A2(n_188),
.B(n_206),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_182),
.A2(n_160),
.B(n_154),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_95),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_196),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_129),
.B1(n_101),
.B2(n_91),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_189),
.B1(n_198),
.B2(n_153),
.Y(n_212)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_191),
.Y(n_214)
);

INVxp33_ASAP7_75t_SL g188 ( 
.A(n_149),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_150),
.A2(n_101),
.B1(n_87),
.B2(n_131),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_207),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_L g196 ( 
.A1(n_157),
.A2(n_111),
.A3(n_94),
.B1(n_131),
.B2(n_126),
.C1(n_79),
.C2(n_75),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_163),
.A2(n_126),
.B1(n_79),
.B2(n_7),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_155),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_201),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_94),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_173),
.C(n_148),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_SL g206 ( 
.A1(n_174),
.A2(n_94),
.B(n_6),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_152),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_176),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_209),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_163),
.B1(n_159),
.B2(n_146),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_211),
.A2(n_223),
.B1(n_237),
.B2(n_198),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_212),
.A2(n_226),
.B1(n_235),
.B2(n_236),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_158),
.B(n_175),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_213),
.A2(n_225),
.B(n_228),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_145),
.Y(n_218)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_219),
.B(n_229),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_158),
.Y(n_220)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_201),
.B(n_172),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_221),
.B(n_205),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_199),
.A2(n_159),
.B1(n_170),
.B2(n_168),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_187),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_224),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_158),
.B(n_171),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_231),
.C(n_200),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_190),
.A2(n_157),
.B(n_152),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_192),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_157),
.Y(n_230)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_179),
.C(n_194),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_152),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_179),
.B(n_160),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_204),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_182),
.A2(n_154),
.B1(n_7),
.B2(n_8),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_199),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_242),
.C(n_250),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_204),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_212),
.B1(n_236),
.B2(n_235),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_211),
.A2(n_184),
.B1(n_208),
.B2(n_185),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_244),
.A2(n_255),
.B1(n_232),
.B2(n_215),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_218),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_219),
.B(n_186),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_249),
.B(n_259),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_228),
.A2(n_197),
.B(n_195),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_213),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_200),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_254),
.C(n_258),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_189),
.C(n_202),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_202),
.B1(n_207),
.B2(n_181),
.Y(n_255)
);

NAND2x1_ASAP7_75t_SL g257 ( 
.A(n_210),
.B(n_183),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_257),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_180),
.C(n_8),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_221),
.B(n_7),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_265),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_269),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_243),
.A2(n_217),
.B1(n_222),
.B2(n_214),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_217),
.B1(n_222),
.B2(n_214),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_258),
.Y(n_265)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_251),
.B(n_229),
.Y(n_270)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_271),
.A2(n_252),
.B(n_246),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_220),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_272),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_251),
.A2(n_224),
.B1(n_237),
.B2(n_223),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_273),
.A2(n_257),
.B1(n_9),
.B2(n_11),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_216),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_278),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_248),
.A2(n_234),
.B1(n_216),
.B2(n_10),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_276),
.A2(n_239),
.B1(n_238),
.B2(n_248),
.Y(n_282)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_277),
.A2(n_260),
.B1(n_255),
.B2(n_256),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_8),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_254),
.C(n_240),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_283),
.C(n_286),
.Y(n_300)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_247),
.C(n_246),
.Y(n_283)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_285),
.A2(n_272),
.B(n_277),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_247),
.C(n_242),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_256),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_267),
.Y(n_295)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

OAI21x1_ASAP7_75t_L g293 ( 
.A1(n_261),
.A2(n_9),
.B(n_260),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_293),
.A2(n_266),
.B(n_278),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_294),
.A2(n_302),
.B(n_304),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_292),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_268),
.Y(n_297)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_282),
.A2(n_269),
.B1(n_265),
.B2(n_276),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_298),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_303),
.B1(n_287),
.B2(n_302),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

INVxp33_ASAP7_75t_SL g303 ( 
.A(n_290),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_285),
.A2(n_279),
.B(n_288),
.Y(n_304)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_279),
.Y(n_306)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_283),
.C(n_286),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_308),
.C(n_313),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_280),
.C(n_292),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_295),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_296),
.B(n_298),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_294),
.C(n_301),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_305),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_316),
.A2(n_318),
.B(n_315),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_319),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_308),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_313),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_310),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_323),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_321),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_321),
.B(n_317),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_324),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_327),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_315),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_314),
.Y(n_331)
);


endmodule