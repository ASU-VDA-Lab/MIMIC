module fake_jpeg_1648_n_144 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_144);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_19),
.B(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_38),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_57),
.B(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_58),
.Y(n_62)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_63),
.B(n_69),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_52),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_42),
.B1(n_53),
.B2(n_51),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_60),
.B1(n_47),
.B2(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_42),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_60),
.B1(n_56),
.B2(n_43),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_64),
.B1(n_76),
.B2(n_73),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_59),
.B(n_44),
.C(n_50),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_85),
.C(n_1),
.Y(n_97)
);

AO22x1_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_56),
.B1(n_54),
.B2(n_40),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_71),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_33),
.Y(n_93)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_44),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_84),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_49),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_36),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_48),
.B(n_71),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_98),
.B1(n_87),
.B2(n_8),
.Y(n_114)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_0),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_94),
.B(n_99),
.Y(n_115)
);

AOI32xp33_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_97),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_81),
.B(n_5),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_92),
.B(n_74),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_14),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_85),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_21),
.C(n_26),
.Y(n_123)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_89),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_109),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_85),
.B1(n_79),
.B2(n_7),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_12),
.B(n_13),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_5),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_6),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_112),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_6),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_87),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_114),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_102),
.B(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_119),
.Y(n_128)
);

AOI32xp33_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_11),
.B(n_12),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_123),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_18),
.C(n_24),
.Y(n_124)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_127),
.A2(n_111),
.B1(n_115),
.B2(n_114),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_123),
.C(n_122),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_118),
.B(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_131),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_135),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_130),
.B(n_132),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_132),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_137),
.B(n_117),
.Y(n_141)
);

AOI322xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_129),
.A3(n_126),
.B1(n_120),
.B2(n_100),
.C1(n_27),
.C2(n_23),
.Y(n_142)
);

AOI221xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_124),
.B1(n_129),
.B2(n_22),
.C(n_15),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_17),
.Y(n_144)
);


endmodule