module fake_jpeg_3396_n_217 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_217);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_217;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_2),
.B(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_36),
.B(n_38),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_7),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_14),
.B(n_7),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_51),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_6),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_20),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_8),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_33),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_62),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_13),
.B1(n_30),
.B2(n_31),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_67),
.A2(n_69),
.B1(n_83),
.B2(n_97),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_12),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_35),
.A2(n_13),
.B1(n_30),
.B2(n_31),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_20),
.C(n_32),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_70),
.B(n_73),
.C(n_94),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_24),
.C(n_32),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_42),
.A2(n_17),
.B1(n_29),
.B2(n_27),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_86),
.B1(n_52),
.B2(n_43),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_46),
.A2(n_30),
.B1(n_24),
.B2(n_29),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_34),
.B(n_33),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_68),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_37),
.A2(n_27),
.B1(n_25),
.B2(n_23),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_25),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_23),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_8),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_44),
.Y(n_96)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_101),
.B(n_99),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_62),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_105),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_40),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_123),
.C(n_72),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_61),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_47),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_112),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_78),
.A2(n_44),
.B1(n_43),
.B2(n_40),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_111),
.B1(n_71),
.B2(n_64),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_114),
.Y(n_143)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_65),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_0),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_98),
.A2(n_5),
.B1(n_11),
.B2(n_94),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_116),
.A2(n_71),
.B1(n_100),
.B2(n_91),
.Y(n_127)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_5),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_124),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_11),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_122),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_11),
.Y(n_122)
);

AOI32xp33_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_93),
.A3(n_91),
.B1(n_64),
.B2(n_82),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

BUFx24_ASAP7_75t_SL g128 ( 
.A(n_113),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_144),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_129),
.B(n_135),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_131),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_87),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_142),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_106),
.A2(n_87),
.B1(n_92),
.B2(n_75),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_137),
.A2(n_138),
.B1(n_140),
.B2(n_148),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_105),
.A2(n_75),
.B1(n_80),
.B2(n_66),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_80),
.A3(n_100),
.B1(n_66),
.B2(n_72),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_145),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_63),
.B1(n_77),
.B2(n_122),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_77),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_63),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_63),
.B(n_103),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_104),
.A2(n_112),
.B1(n_121),
.B2(n_114),
.Y(n_148)
);

NOR4xp25_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_114),
.C(n_117),
.D(n_111),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_150),
.B(n_159),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_110),
.B1(n_125),
.B2(n_108),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_162),
.Y(n_167)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_119),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_120),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_161),
.Y(n_166)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_148),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_165),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_137),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_135),
.B(n_129),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_142),
.C(n_131),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_175),
.C(n_177),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_126),
.B1(n_136),
.B2(n_143),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_162),
.B1(n_154),
.B2(n_156),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_160),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_172),
.B(n_174),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_138),
.C(n_141),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_143),
.C(n_130),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_147),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_182),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_158),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_158),
.B(n_149),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_186),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_158),
.B(n_149),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_168),
.C(n_175),
.Y(n_193)
);

XOR2x2_ASAP7_75t_SL g190 ( 
.A(n_182),
.B(n_170),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_193),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_191),
.A2(n_186),
.B(n_185),
.Y(n_201)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_179),
.C(n_184),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_201),
.Y(n_206)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_192),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_199),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_190),
.B(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_195),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_195),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_203),
.A2(n_187),
.B1(n_194),
.B2(n_191),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_196),
.A2(n_179),
.B(n_176),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_204),
.A2(n_196),
.B(n_177),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_157),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_205),
.B(n_151),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_210),
.C(n_206),
.Y(n_213)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_208),
.Y(n_211)
);

AOI31xp67_ASAP7_75t_SL g209 ( 
.A1(n_202),
.A2(n_151),
.A3(n_147),
.B(n_134),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_209),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

OAI21x1_ASAP7_75t_L g214 ( 
.A1(n_211),
.A2(n_206),
.B(n_134),
.Y(n_214)
);

NOR2xp67_ASAP7_75t_SL g216 ( 
.A(n_214),
.B(n_212),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_216),
.B(n_215),
.Y(n_217)
);


endmodule