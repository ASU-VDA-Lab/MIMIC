module fake_jpeg_22346_n_272 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_272);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_15),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_0),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_14),
.B(n_26),
.C(n_13),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_20),
.Y(n_50)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_41),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_30),
.Y(n_57)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_37),
.B1(n_32),
.B2(n_29),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_18),
.C(n_21),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_54),
.B(n_35),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_53),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_17),
.B1(n_27),
.B2(n_24),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_17),
.B1(n_37),
.B2(n_32),
.Y(n_69)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_60),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_68),
.B(n_48),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_64),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_35),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_66),
.C(n_67),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_35),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_72),
.B1(n_76),
.B2(n_48),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_25),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_25),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_38),
.Y(n_76)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_85),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_54),
.B1(n_32),
.B2(n_45),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_67),
.B1(n_63),
.B2(n_60),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_81),
.B(n_96),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_75),
.B(n_28),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_43),
.B1(n_17),
.B2(n_27),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_92),
.B1(n_58),
.B2(n_45),
.Y(n_101)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_56),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_28),
.C(n_44),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_28),
.C(n_70),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_44),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_59),
.Y(n_98)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_91),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_24),
.B1(n_33),
.B2(n_29),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_94),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_117),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_100),
.A2(n_102),
.B1(n_84),
.B2(n_77),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_111),
.B1(n_112),
.B2(n_114),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_57),
.B1(n_33),
.B2(n_29),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_95),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_106),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_73),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_80),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_94),
.B1(n_91),
.B2(n_87),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_88),
.B1(n_86),
.B2(n_93),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_93),
.A2(n_72),
.B1(n_73),
.B2(n_28),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_81),
.A2(n_28),
.B1(n_27),
.B2(n_40),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_74),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_71),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_40),
.B1(n_51),
.B2(n_53),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_87),
.B1(n_78),
.B2(n_80),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_127),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_84),
.B1(n_71),
.B2(n_89),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_126),
.B1(n_114),
.B2(n_112),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_118),
.B(n_16),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

AO22x1_ASAP7_75t_SL g126 ( 
.A1(n_110),
.A2(n_21),
.B1(n_13),
.B2(n_19),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_107),
.Y(n_127)
);

OAI21x1_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_21),
.B(n_19),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_128),
.A2(n_129),
.B(n_131),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_113),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_80),
.Y(n_136)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_108),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_31),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_100),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_76),
.Y(n_140)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_142),
.C(n_104),
.Y(n_155)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_62),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_147),
.B(n_149),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_111),
.C(n_105),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_150),
.C(n_160),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_139),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_98),
.B(n_115),
.Y(n_147)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_137),
.Y(n_170)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_31),
.B(n_51),
.C(n_19),
.D(n_26),
.Y(n_150)
);

OAI22x1_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_39),
.B1(n_116),
.B2(n_56),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_151),
.A2(n_14),
.B1(n_2),
.B2(n_3),
.Y(n_187)
);

AO21x1_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_14),
.B(n_26),
.Y(n_183)
);

AND2x4_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_39),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_14),
.B(n_2),
.Y(n_185)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_104),
.C(n_31),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_120),
.A2(n_138),
.B1(n_130),
.B2(n_123),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_163),
.B1(n_151),
.B2(n_122),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_120),
.A2(n_22),
.B1(n_15),
.B2(n_25),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_97),
.C(n_22),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_125),
.C(n_147),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_173),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_180),
.C(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_171),
.A2(n_176),
.B1(n_181),
.B2(n_187),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_121),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_174),
.A2(n_179),
.B(n_183),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_129),
.B1(n_124),
.B2(n_131),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_182),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_148),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_97),
.C(n_22),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_23),
.B1(n_26),
.B2(n_19),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_23),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_188),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_156),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_0),
.Y(n_186)
);

INVxp33_ASAP7_75t_SL g203 ( 
.A(n_186),
.Y(n_203)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_192),
.B(n_201),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_194),
.B(n_200),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_145),
.C(n_156),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_196),
.B(n_171),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_149),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_206),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_162),
.Y(n_199)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_169),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_158),
.C(n_165),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_175),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_204),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_156),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_198),
.A2(n_183),
.B1(n_150),
.B2(n_186),
.Y(n_211)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_189),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_213),
.B(n_220),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_R g214 ( 
.A1(n_203),
.A2(n_186),
.B1(n_167),
.B2(n_185),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_201),
.Y(n_227)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_217),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_180),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_187),
.Y(n_219)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_191),
.A2(n_181),
.B1(n_8),
.B2(n_9),
.Y(n_221)
);

OA21x2_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_194),
.B(n_12),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_206),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_8),
.B1(n_11),
.B2(n_10),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

NAND2xp33_ASAP7_75t_SL g247 ( 
.A(n_224),
.B(n_230),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_227),
.B(n_231),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_195),
.B1(n_192),
.B2(n_197),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_228),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_207),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_202),
.C(n_196),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_231),
.A2(n_234),
.B(n_222),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_209),
.B(n_221),
.Y(n_233)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_233),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_217),
.C(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_212),
.B(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_212),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_229),
.C(n_230),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_242),
.B(n_243),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_8),
.B(n_10),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_244),
.B(n_235),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_4),
.Y(n_246)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_250),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_256),
.B(n_240),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_232),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_224),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_255),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_246),
.B(n_224),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_4),
.C(n_5),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_251),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_258),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_254),
.A2(n_247),
.B1(n_5),
.B2(n_6),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_261),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_253),
.A2(n_247),
.B1(n_5),
.B2(n_6),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_262),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_260),
.A2(n_249),
.B(n_256),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_266),
.A2(n_259),
.B(n_5),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_268),
.B(n_263),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_4),
.C(n_7),
.Y(n_268)
);

BUFx24_ASAP7_75t_SL g270 ( 
.A(n_269),
.Y(n_270)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_264),
.B(n_7),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g272 ( 
.A(n_271),
.B(n_7),
.CI(n_235),
.CON(n_272),
.SN(n_272)
);


endmodule