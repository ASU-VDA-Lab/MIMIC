module fake_jpeg_24774_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g16 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_16),
.A2(n_23),
.B1(n_18),
.B2(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_21),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_10),
.A2(n_0),
.B(n_2),
.Y(n_20)
);

OAI21xp33_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_14),
.B(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_0),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_20),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g23 ( 
.A1(n_9),
.A2(n_4),
.B1(n_11),
.B2(n_6),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_23),
.A2(n_12),
.B1(n_11),
.B2(n_14),
.Y(n_24)
);

A2O1A1O1Ixp25_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_25),
.B(n_15),
.C(n_28),
.D(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_27),
.B(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_23),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_30),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_32),
.A2(n_34),
.B1(n_27),
.B2(n_30),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_33),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_29),
.B(n_28),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_32),
.C(n_34),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_39),
.B(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

AO221x1_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_41),
.B1(n_37),
.B2(n_30),
.C(n_35),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_24),
.B(n_26),
.Y(n_43)
);


endmodule