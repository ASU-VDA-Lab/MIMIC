module fake_jpeg_23631_n_135 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx6_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_11),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_17),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_20),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_22),
.A2(n_11),
.B1(n_17),
.B2(n_19),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_31),
.A2(n_38),
.B(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_20),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_11),
.B1(n_17),
.B2(n_12),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_21),
.B1(n_26),
.B2(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_23),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_24),
.A2(n_19),
.B1(n_21),
.B2(n_12),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_50),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_46),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_59)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_29),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_31),
.A2(n_36),
.B1(n_34),
.B2(n_39),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_33),
.A2(n_16),
.B1(n_20),
.B2(n_25),
.Y(n_53)
);

NOR3xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_35),
.C(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_63),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_49),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_65),
.Y(n_74)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_66),
.Y(n_67)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_32),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_73),
.Y(n_90)
);

AO21x2_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_52),
.B(n_39),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_70),
.A2(n_30),
.B1(n_25),
.B2(n_20),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_59),
.B1(n_55),
.B2(n_58),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_45),
.B1(n_61),
.B2(n_39),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_47),
.B(n_48),
.C(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_0),
.Y(n_83)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_80),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_61),
.C(n_30),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_39),
.B1(n_30),
.B2(n_29),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_82),
.A2(n_83),
.B(n_88),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_72),
.B(n_1),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_86),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_68),
.B(n_74),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_67),
.Y(n_89)
);

OA21x2_ASAP7_75t_SL g91 ( 
.A1(n_88),
.A2(n_78),
.B(n_71),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_2),
.B(n_3),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_70),
.B(n_74),
.C(n_85),
.D(n_79),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_95),
.C(n_84),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_87),
.B(n_70),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_2),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_104),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_87),
.C(n_75),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_4),
.C(n_5),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_97),
.A2(n_70),
.B1(n_82),
.B2(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_109),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_86),
.B1(n_83),
.B2(n_73),
.Y(n_106)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_107),
.A2(n_108),
.B(n_94),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_91),
.A2(n_92),
.B1(n_98),
.B2(n_93),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_98),
.B(n_96),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_101),
.B(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_114),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_3),
.C(n_4),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_4),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_110),
.B(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_117),
.B(n_120),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_122),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_6),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_127),
.C(n_7),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_116),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_8),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_120),
.B(n_8),
.Y(n_128)
);

AOI21x1_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_10),
.B(n_123),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_130),
.C(n_126),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_132),
.B(n_10),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_134),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);


endmodule