module real_jpeg_33431_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx2_ASAP7_75t_L g106 ( 
.A(n_0),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_0),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g200 ( 
.A(n_0),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_1),
.A2(n_14),
.B(n_393),
.Y(n_13)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_1),
.Y(n_395)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_2),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_2),
.B(n_177),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_2),
.A2(n_175),
.B1(n_374),
.B2(n_375),
.Y(n_373)
);

INVx3_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_3),
.A2(n_52),
.B1(n_97),
.B2(n_100),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_3),
.A2(n_52),
.B1(n_148),
.B2(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_3),
.B(n_25),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_3),
.B(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_3),
.B(n_323),
.C(n_326),
.Y(n_322)
);

NAND2xp67_ASAP7_75t_L g338 ( 
.A(n_3),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_3),
.B(n_188),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_5),
.Y(n_81)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_6),
.Y(n_99)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_6),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_6),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_6),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_7),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_8),
.Y(n_230)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_9),
.Y(n_129)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_9),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_9),
.Y(n_140)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_10),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_11),
.A2(n_110),
.B1(n_111),
.B2(n_115),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_11),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_11),
.A2(n_110),
.B1(n_181),
.B2(n_185),
.Y(n_180)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_12),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_364),
.Y(n_14)
);

AO21x1_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_237),
.B(n_362),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_204),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_20),
.B(n_204),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_158),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_21),
.B(n_159),
.C(n_390),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_93),
.B(n_154),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_22),
.A2(n_156),
.B(n_209),
.Y(n_208)
);

OAI21x1_ASAP7_75t_L g381 ( 
.A1(n_22),
.A2(n_154),
.B(n_197),
.Y(n_381)
);

NOR2x1p5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_60),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_23),
.B(n_123),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_23),
.Y(n_260)
);

AOI22x1_ASAP7_75t_L g386 ( 
.A1(n_23),
.A2(n_193),
.B1(n_387),
.B2(n_388),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_24),
.Y(n_157)
);

AO22x2_ASAP7_75t_L g195 ( 
.A1(n_24),
.A2(n_62),
.B1(n_157),
.B2(n_196),
.Y(n_195)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_38),
.B(n_51),
.Y(n_24)
);

OAI22x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_28),
.Y(n_218)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_32),
.Y(n_235)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2x1_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_45),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_49),
.Y(n_226)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B(n_56),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_87),
.B(n_91),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_52),
.B(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVxp33_ASAP7_75t_L g236 ( 
.A(n_56),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_61),
.B(n_123),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_61),
.B(n_371),
.Y(n_379)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_62),
.B(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_62),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_62),
.B(n_123),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_62),
.Y(n_265)
);

OA21x2_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_73),
.B(n_86),
.Y(n_62)
);

NOR2x1p5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_74),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_63),
.Y(n_313)
);

OAI22x1_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_66),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_66),
.Y(n_291)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_68),
.Y(n_184)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_72),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_72),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_78),
.B1(n_82),
.B2(n_83),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_85),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_90),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_91),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_94),
.B(n_195),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_123),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_95),
.A2(n_123),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_95),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_103),
.B1(n_109),
.B2(n_119),
.Y(n_95)
);

OR2x6_ASAP7_75t_L g211 ( 
.A(n_96),
.B(n_162),
.Y(n_211)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx4f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_103),
.A2(n_109),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_126),
.B1(n_130),
.B2(n_132),
.Y(n_125)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2x1p5_ASAP7_75t_L g197 ( 
.A(n_123),
.B(n_198),
.Y(n_197)
);

XOR2x2_ASAP7_75t_SL g207 ( 
.A(n_123),
.B(n_198),
.Y(n_207)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_123),
.Y(n_246)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_123),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_123),
.A2(n_210),
.B1(n_211),
.B2(n_246),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_123),
.A2(n_246),
.B1(n_317),
.B2(n_318),
.Y(n_346)
);

OA21x2_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_136),
.B(n_151),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_125),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_125),
.B(n_136),
.Y(n_192)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_129),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22x1_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_141),
.B1(n_145),
.B2(n_148),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_144),
.Y(n_282)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_149),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_151),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AND3x1_ASAP7_75t_L g249 ( 
.A(n_156),
.B(n_250),
.C(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_157),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_194),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_178),
.B1(n_179),
.B2(n_193),
.Y(n_159)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_160),
.A2(n_384),
.B(n_385),
.Y(n_383)
);

NAND2x1_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_169),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_168),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_167),
.Y(n_339)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

OAI21x1_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_175),
.B(n_176),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_188),
.B(n_190),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_180),
.A2(n_188),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_180),
.B(n_188),
.Y(n_385)
);

INVx3_ASAP7_75t_SL g181 ( 
.A(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_190),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_192),
.Y(n_372)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_193),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_194),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_197),
.B1(n_202),
.B2(n_203),
.Y(n_194)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_195),
.A2(n_202),
.B1(n_209),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.C(n_208),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_206),
.B(n_207),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_208),
.B(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_210),
.B(n_213),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_210),
.B(n_265),
.C(n_266),
.Y(n_264)
);

NAND2x1p5_ASAP7_75t_L g302 ( 
.A(n_210),
.B(n_275),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_210),
.A2(n_211),
.B1(n_266),
.B2(n_267),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_210),
.B(n_303),
.C(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_210),
.B(n_346),
.Y(n_345)
);

CKINVDCx11_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_211),
.B(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_211),
.B(n_337),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_211),
.B(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OA21x2_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_222),
.B(n_227),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx4f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_231),
.B(n_236),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx2_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AO21x1_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_268),
.B(n_356),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_254),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_241),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_252),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_242),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.C(n_248),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_245),
.A2(n_248),
.B1(n_249),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_246),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_250),
.Y(n_298)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_252),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

NOR2xp67_ASAP7_75t_L g361 ( 
.A(n_255),
.B(n_258),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.C(n_263),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_259),
.B(n_354),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_261),
.B(n_274),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_262),
.B(n_264),
.Y(n_354)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

O2A1O1Ixp33_ASAP7_75t_SL g271 ( 
.A1(n_265),
.A2(n_272),
.B(n_274),
.C(n_298),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_306),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_265),
.A2(n_370),
.B(n_378),
.Y(n_369)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21x1_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_351),
.B(n_355),
.Y(n_268)
);

AOI21x1_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_308),
.B(n_350),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_299),
.Y(n_270)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_271),
.B(n_299),
.Y(n_350)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_273),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_273),
.B(n_302),
.C(n_304),
.Y(n_352)
);

OAI21x1_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_279),
.B(n_287),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_292),
.B(n_296),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_295),
.Y(n_321)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_304),
.B1(n_305),
.B2(n_307),
.Y(n_299)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI21x1_ASAP7_75t_SL g308 ( 
.A1(n_309),
.A2(n_314),
.B(n_349),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_310),
.B(n_311),
.Y(n_349)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_312),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_315),
.A2(n_334),
.B(n_347),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_330),
.Y(n_315)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_316),
.Y(n_348)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_329),
.Y(n_342)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_331),
.B(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_345),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_343),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_340),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NOR2x1_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_352),
.B(n_353),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_360),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_365),
.B(n_391),
.Y(n_364)
);

INVxp33_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_389),
.Y(n_366)
);

NAND2x1p5_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_389),
.Y(n_392)
);

XNOR2x1_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_380),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx5_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

XNOR2x1_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

XOR2x1_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_386),
.Y(n_382)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_396),
.Y(n_393)
);

INVx5_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);


endmodule