module fake_aes_10869_n_671 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_671);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_671;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_466;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_24), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_17), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_68), .Y(n_81) );
BUFx10_ASAP7_75t_L g82 ( .A(n_63), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_78), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_15), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_43), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_69), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_58), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_65), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_67), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_70), .Y(n_90) );
HB1xp67_ASAP7_75t_L g91 ( .A(n_62), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_23), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_21), .Y(n_93) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_61), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_26), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_48), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_60), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_72), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_42), .Y(n_99) );
BUFx3_ASAP7_75t_L g100 ( .A(n_25), .Y(n_100) );
OR2x2_ASAP7_75t_L g101 ( .A(n_74), .B(n_59), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_52), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_19), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_16), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_13), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_45), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_6), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_47), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_7), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_28), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_75), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_30), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_32), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_5), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_73), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_53), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_50), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_1), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_34), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_41), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_57), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_38), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_88), .Y(n_123) );
BUFx8_ASAP7_75t_L g124 ( .A(n_115), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_112), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_115), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_109), .B(n_0), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_88), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_112), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_94), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_82), .B(n_0), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_90), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_90), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_109), .B(n_1), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_91), .B(n_2), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_79), .Y(n_136) );
AND3x2_ASAP7_75t_L g137 ( .A(n_107), .B(n_2), .C(n_3), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_82), .B(n_3), .Y(n_138) );
NOR2x1_ASAP7_75t_L g139 ( .A(n_114), .B(n_33), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_94), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_104), .B(n_4), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_80), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_94), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_89), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_81), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_83), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_84), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_89), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_118), .B(n_4), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_107), .B(n_5), .Y(n_150) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_105), .Y(n_151) );
AND2x2_ASAP7_75t_SL g152 ( .A(n_101), .B(n_36), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_100), .Y(n_153) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_86), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_85), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_82), .B(n_6), .Y(n_156) );
INVxp67_ASAP7_75t_L g157 ( .A(n_87), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_100), .B(n_7), .Y(n_158) );
BUFx10_ASAP7_75t_L g159 ( .A(n_86), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_154), .B(n_92), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_150), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_130), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_150), .Y(n_163) );
INVx4_ASAP7_75t_L g164 ( .A(n_158), .Y(n_164) );
NAND3x1_ASAP7_75t_L g165 ( .A(n_156), .B(n_119), .C(n_121), .Y(n_165) );
INVx4_ASAP7_75t_L g166 ( .A(n_158), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_150), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_127), .B(n_92), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_130), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_157), .B(n_122), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_153), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_150), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_126), .B(n_99), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_125), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_159), .B(n_99), .Y(n_175) );
INVxp67_ASAP7_75t_SL g176 ( .A(n_127), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_130), .Y(n_177) );
AND2x2_ASAP7_75t_SL g178 ( .A(n_152), .B(n_101), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_130), .Y(n_179) );
AND2x6_ASAP7_75t_L g180 ( .A(n_158), .B(n_120), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_130), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_159), .B(n_116), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_125), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_140), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_148), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_126), .B(n_106), .Y(n_186) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_151), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_159), .B(n_116), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_136), .B(n_106), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_129), .Y(n_190) );
AND2x6_ASAP7_75t_L g191 ( .A(n_156), .B(n_93), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_144), .Y(n_192) );
INVxp67_ASAP7_75t_SL g193 ( .A(n_134), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_124), .B(n_108), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_135), .B(n_96), .Y(n_195) );
INVx4_ASAP7_75t_L g196 ( .A(n_152), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_129), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_133), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_136), .B(n_110), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_133), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_140), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_140), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_140), .Y(n_203) );
INVxp67_ASAP7_75t_SL g204 ( .A(n_176), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_193), .B(n_135), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_189), .B(n_132), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_198), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_168), .B(n_132), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_168), .B(n_128), .Y(n_209) );
INVxp33_ASAP7_75t_L g210 ( .A(n_187), .Y(n_210) );
NOR2xp33_ASAP7_75t_SL g211 ( .A(n_196), .B(n_119), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_171), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_196), .A2(n_152), .B1(n_128), .B2(n_123), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_195), .B(n_123), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_195), .B(n_155), .Y(n_215) );
OR2x2_ASAP7_75t_L g216 ( .A(n_173), .B(n_144), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_171), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_182), .B(n_155), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_182), .B(n_124), .Y(n_219) );
INVx5_ASAP7_75t_L g220 ( .A(n_180), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_198), .Y(n_221) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_196), .A2(n_147), .B1(n_146), .B2(n_145), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_194), .B(n_131), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_196), .A2(n_145), .B1(n_147), .B2(n_146), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_188), .B(n_124), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_178), .A2(n_142), .B1(n_149), .B2(n_153), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_200), .Y(n_227) );
BUFx4f_ASAP7_75t_L g228 ( .A(n_191), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_171), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_188), .B(n_142), .Y(n_230) );
AOI22xp5_ASAP7_75t_SL g231 ( .A1(n_185), .A2(n_141), .B1(n_137), .B2(n_103), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_197), .Y(n_232) );
OR2x2_ASAP7_75t_L g233 ( .A(n_186), .B(n_138), .Y(n_233) );
NAND2x1p5_ASAP7_75t_L g234 ( .A(n_178), .B(n_139), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_170), .B(n_102), .Y(n_235) );
AND2x6_ASAP7_75t_L g236 ( .A(n_161), .B(n_111), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_164), .B(n_98), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_178), .A2(n_117), .B1(n_113), .B2(n_97), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_180), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_160), .B(n_95), .Y(n_240) );
NOR2x2_ASAP7_75t_L g241 ( .A(n_165), .B(n_8), .Y(n_241) );
OR2x6_ASAP7_75t_L g242 ( .A(n_165), .B(n_94), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_200), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_199), .B(n_8), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_175), .B(n_94), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_191), .B(n_143), .Y(n_246) );
INVxp67_ASAP7_75t_L g247 ( .A(n_191), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_174), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_164), .B(n_143), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_197), .Y(n_250) );
INVx2_ASAP7_75t_SL g251 ( .A(n_191), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_174), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_161), .B(n_143), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_197), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_183), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_191), .B(n_143), .Y(n_256) );
INVx4_ASAP7_75t_L g257 ( .A(n_164), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_213), .A2(n_180), .B1(n_191), .B2(n_172), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_208), .A2(n_167), .B(n_172), .C(n_163), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_204), .Y(n_260) );
NOR2x1_ASAP7_75t_L g261 ( .A(n_242), .B(n_197), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_204), .B(n_191), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_239), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_239), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_229), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_213), .A2(n_180), .B1(n_167), .B2(n_163), .Y(n_266) );
CKINVDCx6p67_ASAP7_75t_R g267 ( .A(n_242), .Y(n_267) );
CKINVDCx8_ASAP7_75t_R g268 ( .A(n_242), .Y(n_268) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_211), .A2(n_180), .B1(n_166), .B2(n_164), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_248), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_206), .A2(n_163), .B(n_183), .C(n_190), .Y(n_271) );
BUFx2_ASAP7_75t_L g272 ( .A(n_236), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_239), .Y(n_273) );
OAI21xp5_ASAP7_75t_L g274 ( .A1(n_253), .A2(n_163), .B(n_180), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_233), .B(n_166), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_205), .Y(n_276) );
INVx5_ASAP7_75t_L g277 ( .A(n_239), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_252), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_209), .Y(n_279) );
NOR3xp33_ASAP7_75t_L g280 ( .A(n_219), .B(n_192), .C(n_166), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_223), .B(n_166), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_218), .B(n_180), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_207), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_231), .Y(n_284) );
OAI22xp5_ASAP7_75t_L g285 ( .A1(n_238), .A2(n_190), .B1(n_140), .B2(n_143), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_229), .Y(n_286) );
INVx4_ASAP7_75t_L g287 ( .A(n_220), .Y(n_287) );
INVxp67_ASAP7_75t_L g288 ( .A(n_214), .Y(n_288) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_238), .A2(n_201), .B1(n_179), .B2(n_181), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_253), .A2(n_181), .B(n_202), .Y(n_290) );
BUFx12f_ASAP7_75t_L g291 ( .A(n_223), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_221), .Y(n_292) );
A2O1A1Ixp33_ASAP7_75t_L g293 ( .A1(n_215), .A2(n_201), .B(n_202), .C(n_179), .Y(n_293) );
INVx5_ASAP7_75t_L g294 ( .A(n_220), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_220), .Y(n_295) );
A2O1A1Ixp33_ASAP7_75t_SL g296 ( .A1(n_245), .A2(n_201), .B(n_177), .C(n_184), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_220), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_230), .B(n_9), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_229), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_225), .B(n_9), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_255), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_229), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_227), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_243), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_232), .Y(n_305) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_210), .A2(n_177), .B1(n_184), .B2(n_203), .C(n_169), .Y(n_306) );
NAND3xp33_ASAP7_75t_L g307 ( .A(n_271), .B(n_226), .C(n_245), .Y(n_307) );
INVx4_ASAP7_75t_L g308 ( .A(n_294), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_270), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_258), .A2(n_226), .B1(n_224), .B2(n_222), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_270), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_288), .B(n_224), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_278), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_288), .Y(n_314) );
CKINVDCx6p67_ASAP7_75t_R g315 ( .A(n_267), .Y(n_315) );
INVx4_ASAP7_75t_L g316 ( .A(n_294), .Y(n_316) );
OAI21x1_ASAP7_75t_L g317 ( .A1(n_261), .A2(n_256), .B(n_246), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_276), .B(n_222), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_277), .Y(n_319) );
INVxp67_ASAP7_75t_L g320 ( .A(n_279), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_291), .B(n_216), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_300), .A2(n_240), .B1(n_235), .B2(n_244), .C(n_234), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_263), .Y(n_323) );
AND2x6_ASAP7_75t_L g324 ( .A(n_264), .B(n_228), .Y(n_324) );
OAI21x1_ASAP7_75t_L g325 ( .A1(n_290), .A2(n_212), .B(n_217), .Y(n_325) );
OAI21x1_ASAP7_75t_L g326 ( .A1(n_274), .A2(n_234), .B(n_254), .Y(n_326) );
NOR2xp67_ASAP7_75t_L g327 ( .A(n_294), .B(n_277), .Y(n_327) );
BUFx12f_ASAP7_75t_L g328 ( .A(n_300), .Y(n_328) );
AOI22xp33_ASAP7_75t_SL g329 ( .A1(n_284), .A2(n_228), .B1(n_241), .B2(n_236), .Y(n_329) );
OAI21x1_ASAP7_75t_L g330 ( .A1(n_289), .A2(n_250), .B(n_237), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_278), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_301), .Y(n_332) );
AOI22xp33_ASAP7_75t_SL g333 ( .A1(n_272), .A2(n_236), .B1(n_251), .B2(n_247), .Y(n_333) );
OAI21xp5_ASAP7_75t_L g334 ( .A1(n_271), .A2(n_247), .B(n_236), .Y(n_334) );
OR2x6_ASAP7_75t_L g335 ( .A(n_281), .B(n_257), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_260), .B(n_257), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_281), .B(n_236), .Y(n_337) );
AO31x2_ASAP7_75t_L g338 ( .A1(n_293), .A2(n_249), .A3(n_11), .B(n_12), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_277), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_301), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_332), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_332), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_312), .B(n_283), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g344 ( .A1(n_320), .A2(n_275), .B1(n_280), .B2(n_298), .C(n_303), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_309), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_312), .B(n_292), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_309), .Y(n_347) );
OA21x2_ASAP7_75t_L g348 ( .A1(n_325), .A2(n_293), .B(n_266), .Y(n_348) );
O2A1O1Ixp33_ASAP7_75t_SL g349 ( .A1(n_311), .A2(n_296), .B(n_282), .C(n_262), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_328), .A2(n_322), .B1(n_314), .B2(n_329), .Y(n_350) );
AOI22xp33_ASAP7_75t_SL g351 ( .A1(n_328), .A2(n_275), .B1(n_268), .B2(n_304), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_311), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_314), .B(n_258), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_313), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_318), .A2(n_266), .B1(n_269), .B2(n_285), .Y(n_355) );
OA21x2_ASAP7_75t_L g356 ( .A1(n_325), .A2(n_306), .B(n_265), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_313), .Y(n_357) );
BUFx8_ASAP7_75t_L g358 ( .A(n_337), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_331), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_331), .Y(n_360) );
BUFx2_ASAP7_75t_L g361 ( .A(n_340), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_310), .A2(n_280), .B1(n_305), .B2(n_249), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_340), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_336), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_321), .A2(n_305), .B1(n_295), .B2(n_273), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_336), .Y(n_366) );
OAI21xp33_ASAP7_75t_L g367 ( .A1(n_307), .A2(n_334), .B(n_335), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_338), .Y(n_368) );
AO21x2_ASAP7_75t_L g369 ( .A1(n_368), .A2(n_307), .B(n_334), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_347), .B(n_338), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_341), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_341), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_358), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_342), .Y(n_374) );
INVx2_ASAP7_75t_SL g375 ( .A(n_361), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_342), .Y(n_376) );
OR2x2_ASAP7_75t_SL g377 ( .A(n_368), .B(n_315), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_347), .B(n_338), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_348), .A2(n_330), .B(n_326), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_345), .Y(n_380) );
AO21x2_ASAP7_75t_L g381 ( .A1(n_367), .A2(n_296), .B(n_330), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_343), .B(n_346), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_352), .Y(n_383) );
INVx3_ASAP7_75t_L g384 ( .A(n_345), .Y(n_384) );
INVxp67_ASAP7_75t_SL g385 ( .A(n_361), .Y(n_385) );
INVx5_ASAP7_75t_L g386 ( .A(n_359), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_350), .B(n_315), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_352), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_343), .B(n_338), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_354), .B(n_338), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_358), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_353), .A2(n_337), .B1(n_335), .B2(n_339), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_354), .B(n_326), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_359), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_363), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_346), .B(n_335), .Y(n_396) );
AO31x2_ASAP7_75t_L g397 ( .A1(n_355), .A2(n_357), .A3(n_360), .B(n_363), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_357), .B(n_339), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_360), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_370), .B(n_353), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_398), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_370), .B(n_366), .Y(n_402) );
NAND3xp33_ASAP7_75t_L g403 ( .A(n_386), .B(n_344), .C(n_362), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_370), .B(n_366), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_371), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_378), .B(n_364), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_380), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_378), .B(n_364), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_380), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_380), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_378), .B(n_327), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_395), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_395), .Y(n_413) );
NOR3xp33_ASAP7_75t_L g414 ( .A(n_387), .B(n_351), .C(n_308), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_390), .B(n_348), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_390), .B(n_348), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_371), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_372), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_372), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_390), .B(n_348), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_374), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_394), .B(n_356), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_382), .B(n_365), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_395), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_374), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_376), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_385), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_382), .B(n_358), .Y(n_428) );
NAND4xp25_ASAP7_75t_SL g429 ( .A(n_392), .B(n_333), .C(n_11), .D(n_12), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_376), .B(n_337), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_394), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_397), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_389), .B(n_356), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_383), .B(n_337), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_384), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_383), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_397), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_388), .B(n_335), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_389), .B(n_356), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_388), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_398), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_399), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_436), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_436), .Y(n_444) );
BUFx3_ASAP7_75t_L g445 ( .A(n_427), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_401), .B(n_385), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_441), .B(n_398), .Y(n_447) );
NAND2xp33_ASAP7_75t_R g448 ( .A(n_427), .B(n_384), .Y(n_448) );
BUFx2_ASAP7_75t_L g449 ( .A(n_431), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_402), .B(n_399), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_413), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_440), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_440), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_428), .B(n_396), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_400), .B(n_369), .Y(n_455) );
NAND2x1p5_ASAP7_75t_L g456 ( .A(n_431), .B(n_373), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_402), .B(n_375), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_442), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_400), .B(n_369), .Y(n_459) );
NOR2x1_ASAP7_75t_L g460 ( .A(n_403), .B(n_373), .Y(n_460) );
NOR3xp33_ASAP7_75t_L g461 ( .A(n_429), .B(n_391), .C(n_373), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_442), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_405), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_405), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_417), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_404), .B(n_375), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_404), .B(n_375), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_406), .B(n_396), .Y(n_468) );
NOR2xp33_ASAP7_75t_R g469 ( .A(n_438), .B(n_391), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_417), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_418), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_411), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_413), .Y(n_473) );
AND3x1_ASAP7_75t_L g474 ( .A(n_414), .B(n_392), .C(n_391), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_413), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_411), .B(n_393), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_423), .A2(n_396), .B1(n_386), .B2(n_393), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_408), .B(n_369), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_403), .A2(n_369), .B1(n_393), .B2(n_386), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_406), .B(n_384), .Y(n_480) );
BUFx3_ASAP7_75t_L g481 ( .A(n_407), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_408), .B(n_397), .Y(n_482) );
INVx3_ASAP7_75t_L g483 ( .A(n_411), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_424), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_418), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_408), .B(n_397), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_411), .Y(n_487) );
OAI21xp5_ASAP7_75t_SL g488 ( .A1(n_408), .A2(n_377), .B(n_384), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_415), .B(n_397), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_419), .B(n_386), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_419), .B(n_386), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_421), .B(n_386), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_415), .B(n_397), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_421), .B(n_377), .Y(n_494) );
NAND4xp75_ASAP7_75t_L g495 ( .A(n_434), .B(n_327), .C(n_356), .D(n_14), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_425), .B(n_386), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_416), .B(n_397), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_416), .B(n_379), .Y(n_498) );
INVx1_ASAP7_75t_SL g499 ( .A(n_422), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_451), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_443), .Y(n_501) );
NAND3xp33_ASAP7_75t_SL g502 ( .A(n_461), .B(n_469), .C(n_488), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_444), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_447), .B(n_425), .Y(n_504) );
OR2x6_ASAP7_75t_L g505 ( .A(n_460), .B(n_424), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_450), .B(n_426), .Y(n_506) );
OAI222xp33_ASAP7_75t_L g507 ( .A1(n_494), .A2(n_426), .B1(n_430), .B2(n_422), .C1(n_432), .C2(n_437), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_455), .B(n_420), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_455), .B(n_420), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_452), .Y(n_510) );
NOR2xp67_ASAP7_75t_L g511 ( .A(n_483), .B(n_437), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_454), .B(n_439), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_459), .B(n_439), .Y(n_513) );
INVxp33_ASAP7_75t_SL g514 ( .A(n_469), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_499), .B(n_424), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_453), .Y(n_516) );
INVx2_ASAP7_75t_SL g517 ( .A(n_456), .Y(n_517) );
NAND2x1p5_ASAP7_75t_L g518 ( .A(n_474), .B(n_308), .Y(n_518) );
AND2x2_ASAP7_75t_SL g519 ( .A(n_491), .B(n_433), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_458), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_459), .B(n_433), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_462), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_463), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_467), .B(n_437), .Y(n_524) );
NAND2x1_ASAP7_75t_L g525 ( .A(n_483), .B(n_409), .Y(n_525) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_479), .B(n_432), .C(n_435), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_451), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_473), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_464), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_465), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_470), .Y(n_531) );
AND2x4_ASAP7_75t_L g532 ( .A(n_483), .B(n_487), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_489), .B(n_432), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_476), .B(n_435), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_476), .B(n_412), .Y(n_535) );
INVxp67_ASAP7_75t_SL g536 ( .A(n_448), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_471), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_454), .B(n_10), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_489), .B(n_412), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_485), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_456), .A2(n_409), .B(n_407), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_468), .B(n_10), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_473), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_449), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_457), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_445), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_476), .B(n_410), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_482), .B(n_410), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_482), .B(n_379), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_486), .B(n_379), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_486), .B(n_381), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_466), .B(n_381), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_478), .B(n_472), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_493), .B(n_381), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_475), .Y(n_555) );
INVxp67_ASAP7_75t_SL g556 ( .A(n_448), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_493), .B(n_381), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_501), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_533), .B(n_446), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_544), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_514), .B(n_445), .Y(n_561) );
NOR2x1_ASAP7_75t_L g562 ( .A(n_502), .B(n_495), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_503), .Y(n_563) );
OAI22xp33_ASAP7_75t_SL g564 ( .A1(n_514), .A2(n_490), .B1(n_492), .B2(n_491), .Y(n_564) );
OA21x2_ASAP7_75t_L g565 ( .A1(n_536), .A2(n_479), .B(n_498), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_510), .Y(n_566) );
NOR4xp25_ASAP7_75t_SL g567 ( .A(n_536), .B(n_491), .C(n_496), .D(n_349), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_516), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_546), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_520), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_522), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_519), .B(n_478), .Y(n_572) );
NAND2x1_ASAP7_75t_L g573 ( .A(n_505), .B(n_496), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_544), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_539), .B(n_480), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_519), .A2(n_477), .B1(n_496), .B2(n_497), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_502), .A2(n_481), .B(n_484), .Y(n_577) );
AOI222xp33_ASAP7_75t_L g578 ( .A1(n_538), .A2(n_497), .B1(n_498), .B2(n_481), .C1(n_484), .C2(n_475), .Y(n_578) );
NAND3xp33_ASAP7_75t_SL g579 ( .A(n_518), .B(n_308), .C(n_316), .Y(n_579) );
NAND3xp33_ASAP7_75t_L g580 ( .A(n_538), .B(n_316), .C(n_319), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_523), .Y(n_581) );
AND2x4_ASAP7_75t_L g582 ( .A(n_556), .B(n_319), .Y(n_582) );
INVx1_ASAP7_75t_SL g583 ( .A(n_515), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_529), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_545), .A2(n_316), .B1(n_317), .B2(n_324), .Y(n_585) );
OAI21xp33_ASAP7_75t_L g586 ( .A1(n_556), .A2(n_317), .B(n_299), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_530), .Y(n_587) );
OAI211xp5_ASAP7_75t_L g588 ( .A1(n_542), .A2(n_259), .B(n_277), .C(n_294), .Y(n_588) );
INVxp33_ASAP7_75t_L g589 ( .A(n_542), .Y(n_589) );
OAI211xp5_ASAP7_75t_L g590 ( .A1(n_511), .A2(n_295), .B(n_14), .C(n_13), .Y(n_590) );
CKINVDCx14_ASAP7_75t_R g591 ( .A(n_504), .Y(n_591) );
OAI321xp33_ASAP7_75t_L g592 ( .A1(n_518), .A2(n_302), .A3(n_286), .B1(n_323), .B2(n_162), .C(n_203), .Y(n_592) );
O2A1O1Ixp33_ASAP7_75t_L g593 ( .A1(n_507), .A2(n_273), .B(n_264), .C(n_22), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_531), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_537), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_512), .B(n_18), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_512), .A2(n_323), .B1(n_287), .B2(n_263), .Y(n_597) );
OAI22xp33_ASAP7_75t_L g598 ( .A1(n_517), .A2(n_323), .B1(n_287), .B2(n_297), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_540), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_524), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_505), .A2(n_323), .B1(n_263), .B2(n_297), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_578), .B(n_521), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_589), .A2(n_507), .B1(n_506), .B2(n_513), .C(n_509), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_558), .Y(n_604) );
AOI21xp33_ASAP7_75t_SL g605 ( .A1(n_561), .A2(n_505), .B(n_532), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_563), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_591), .B(n_553), .Y(n_607) );
XNOR2xp5_ASAP7_75t_L g608 ( .A(n_569), .B(n_535), .Y(n_608) );
AOI322xp5_ASAP7_75t_L g609 ( .A1(n_562), .A2(n_508), .A3(n_549), .B1(n_550), .B2(n_551), .C1(n_557), .C2(n_554), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_566), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_568), .Y(n_611) );
XNOR2x2_ASAP7_75t_L g612 ( .A(n_580), .B(n_526), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_600), .B(n_548), .Y(n_613) );
A2O1A1Ixp33_ASAP7_75t_L g614 ( .A1(n_580), .A2(n_525), .B(n_532), .C(n_541), .Y(n_614) );
INVxp67_ASAP7_75t_SL g615 ( .A(n_560), .Y(n_615) );
AOI321xp33_ASAP7_75t_L g616 ( .A1(n_564), .A2(n_547), .A3(n_534), .B1(n_552), .B2(n_543), .C(n_555), .Y(n_616) );
AOI21xp33_ASAP7_75t_L g617 ( .A1(n_590), .A2(n_543), .B(n_528), .Y(n_617) );
AOI211xp5_ASAP7_75t_SL g618 ( .A1(n_579), .A2(n_555), .B(n_528), .C(n_527), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_574), .B(n_527), .Y(n_619) );
OAI21xp5_ASAP7_75t_SL g620 ( .A1(n_593), .A2(n_500), .B(n_323), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_570), .Y(n_621) );
XOR2xp5_ASAP7_75t_L g622 ( .A(n_576), .B(n_500), .Y(n_622) );
OAI22xp33_ASAP7_75t_SL g623 ( .A1(n_573), .A2(n_20), .B1(n_27), .B2(n_29), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_583), .B(n_31), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g625 ( .A1(n_577), .A2(n_203), .B1(n_184), .B2(n_169), .C(n_162), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_571), .B(n_35), .Y(n_626) );
XNOR2xp5_ASAP7_75t_L g627 ( .A(n_559), .B(n_37), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_581), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_614), .A2(n_592), .B(n_588), .Y(n_629) );
OAI22xp33_ASAP7_75t_L g630 ( .A1(n_618), .A2(n_565), .B1(n_572), .B2(n_575), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_607), .B(n_594), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_608), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_603), .A2(n_565), .B1(n_582), .B2(n_599), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_628), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_619), .B(n_613), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_622), .A2(n_582), .B1(n_567), .B2(n_596), .Y(n_636) );
NAND2x1_ASAP7_75t_L g637 ( .A(n_618), .B(n_584), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_605), .A2(n_567), .B1(n_585), .B2(n_595), .Y(n_638) );
XNOR2x1_ASAP7_75t_L g639 ( .A(n_627), .B(n_587), .Y(n_639) );
OAI21xp5_ASAP7_75t_L g640 ( .A1(n_617), .A2(n_586), .B(n_597), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_604), .Y(n_641) );
OAI211xp5_ASAP7_75t_L g642 ( .A1(n_609), .A2(n_601), .B(n_598), .C(n_297), .Y(n_642) );
AO21x1_ASAP7_75t_L g643 ( .A1(n_615), .A2(n_39), .B(n_40), .Y(n_643) );
OAI22xp33_ASAP7_75t_L g644 ( .A1(n_602), .A2(n_297), .B1(n_263), .B2(n_324), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_632), .A2(n_617), .B(n_623), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_632), .A2(n_636), .B1(n_630), .B2(n_633), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_629), .B(n_616), .Y(n_647) );
NAND3xp33_ASAP7_75t_SL g648 ( .A(n_643), .B(n_620), .C(n_612), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_642), .A2(n_621), .B1(n_611), .B2(n_610), .C(n_606), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g650 ( .A1(n_644), .A2(n_625), .B1(n_624), .B2(n_626), .C(n_203), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_637), .A2(n_626), .B(n_46), .C(n_49), .Y(n_651) );
AOI221xp5_ASAP7_75t_SL g652 ( .A1(n_638), .A2(n_203), .B1(n_184), .B2(n_169), .C(n_162), .Y(n_652) );
NOR4xp25_ASAP7_75t_L g653 ( .A(n_641), .B(n_44), .C(n_51), .D(n_54), .Y(n_653) );
OAI22xp33_ASAP7_75t_L g654 ( .A1(n_640), .A2(n_635), .B1(n_631), .B2(n_634), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_647), .A2(n_639), .B(n_203), .Y(n_655) );
NOR2xp67_ASAP7_75t_SL g656 ( .A(n_645), .B(n_324), .Y(n_656) );
NOR3xp33_ASAP7_75t_L g657 ( .A(n_648), .B(n_55), .C(n_56), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_646), .B(n_64), .Y(n_658) );
NAND3x1_ASAP7_75t_L g659 ( .A(n_649), .B(n_324), .C(n_71), .Y(n_659) );
NAND4xp75_ASAP7_75t_L g660 ( .A(n_652), .B(n_324), .C(n_76), .D(n_77), .Y(n_660) );
XNOR2xp5_ASAP7_75t_L g661 ( .A(n_655), .B(n_654), .Y(n_661) );
OR4x2_ASAP7_75t_L g662 ( .A(n_656), .B(n_651), .C(n_653), .D(n_650), .Y(n_662) );
OAI22x1_ASAP7_75t_L g663 ( .A1(n_658), .A2(n_324), .B1(n_66), .B2(n_169), .Y(n_663) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_661), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_662), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_664), .Y(n_666) );
AO22x1_ASAP7_75t_L g667 ( .A1(n_665), .A2(n_657), .B1(n_659), .B2(n_663), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_666), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_668), .A2(n_667), .B1(n_660), .B2(n_324), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_669), .A2(n_162), .B1(n_169), .B2(n_184), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_670), .A2(n_162), .B1(n_169), .B2(n_184), .C(n_664), .Y(n_671) );
endmodule