module fake_jpeg_15812_n_105 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_25),
.Y(n_39)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_23),
.B(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_2),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_26),
.B(n_16),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_18),
.Y(n_43)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_24),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_36),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_22),
.A2(n_14),
.B1(n_20),
.B2(n_18),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_32),
.A2(n_22),
.B1(n_28),
.B2(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_15),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_45),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_22),
.A2(n_17),
.B1(n_20),
.B2(n_14),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_27),
.B1(n_16),
.B2(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_30),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_58),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_37),
.B(n_41),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_59),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_36),
.Y(n_64)
);

BUFx24_ASAP7_75t_SL g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_44),
.B1(n_28),
.B2(n_38),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_68),
.B1(n_53),
.B2(n_59),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_38),
.B1(n_37),
.B2(n_34),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_57),
.B(n_50),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_70),
.B(n_39),
.Y(n_83)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_63),
.B1(n_67),
.B2(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_64),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_81),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_77),
.B(n_76),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_62),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_84),
.B(n_40),
.Y(n_87)
);

FAx1_ASAP7_75t_SL g92 ( 
.A(n_85),
.B(n_29),
.CI(n_35),
.CON(n_92),
.SN(n_92)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_79),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_3),
.B(n_4),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_94),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_35),
.C(n_55),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_3),
.B(n_4),
.Y(n_94)
);

OA21x2_ASAP7_75t_SL g97 ( 
.A1(n_93),
.A2(n_90),
.B(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_98),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_95),
.B(n_12),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_100),
.B(n_8),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_7),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_9),
.C(n_10),
.Y(n_104)
);

BUFx24_ASAP7_75t_SL g105 ( 
.A(n_104),
.Y(n_105)
);


endmodule