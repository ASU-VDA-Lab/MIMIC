module fake_jpeg_4353_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_31),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_29),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_29),
.Y(n_45)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx12_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_41),
.B(n_37),
.Y(n_60)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_45),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_23),
.B(n_27),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_46),
.A2(n_51),
.B1(n_26),
.B2(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_54),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_21),
.B1(n_23),
.B2(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_31),
.B(n_15),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_22),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_60),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_61),
.B(n_63),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_66),
.Y(n_83)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_32),
.B(n_38),
.C(n_19),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_68),
.B(n_72),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_21),
.B1(n_39),
.B2(n_36),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_69),
.A2(n_71),
.B1(n_21),
.B2(n_27),
.Y(n_82)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_57),
.B1(n_52),
.B2(n_48),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_88),
.B1(n_94),
.B2(n_66),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_86),
.B1(n_87),
.B2(n_93),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_82),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_70),
.B1(n_68),
.B2(n_64),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_45),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_19),
.B(n_28),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_55),
.B1(n_47),
.B2(n_40),
.Y(n_88)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_56),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_72),
.B(n_49),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_42),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_47),
.B1(n_42),
.B2(n_50),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_90),
.B1(n_92),
.B2(n_78),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_60),
.C(n_64),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_106),
.C(n_80),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_67),
.B(n_24),
.Y(n_128)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_101),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_107),
.B1(n_79),
.B2(n_73),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_105),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_104),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_28),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_47),
.C(n_36),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_77),
.A2(n_94),
.B1(n_90),
.B2(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_111),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_87),
.B(n_66),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_110),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_87),
.B(n_75),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_112),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_123),
.C(n_124),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_117),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_78),
.B(n_83),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_108),
.B(n_102),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_78),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_122),
.B(n_128),
.Y(n_139)
);

XNOR2x1_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_84),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_79),
.C(n_83),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_130),
.B1(n_98),
.B2(n_50),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_33),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_109),
.C(n_103),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_33),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_25),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_96),
.A2(n_73),
.B1(n_65),
.B2(n_56),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_132),
.A2(n_130),
.B1(n_116),
.B2(n_124),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_101),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_135),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_101),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_137),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_129),
.A2(n_111),
.B(n_99),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_25),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_144),
.C(n_113),
.Y(n_148)
);

NAND4xp25_ASAP7_75t_SL g141 ( 
.A(n_123),
.B(n_112),
.C(n_56),
.D(n_91),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_146),
.B1(n_127),
.B2(n_18),
.Y(n_153)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_117),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_18),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_158),
.C(n_140),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_155),
.B(n_132),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_128),
.C(n_126),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_152),
.B(n_145),
.Y(n_162)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_91),
.C(n_24),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_159),
.C(n_160),
.Y(n_163)
);

NAND2xp67_ASAP7_75t_SL g155 ( 
.A(n_141),
.B(n_25),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_25),
.C(n_18),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_25),
.C(n_18),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_164),
.C(n_166),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_162),
.B(n_167),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_154),
.C(n_159),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_165),
.A2(n_168),
.B(n_169),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_158),
.C(n_150),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_157),
.B(n_135),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_146),
.B(n_138),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_131),
.C(n_25),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_156),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_149),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_171),
.A2(n_17),
.B1(n_1),
.B2(n_3),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_177),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_17),
.B(n_1),
.C(n_2),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_176),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_171),
.A2(n_14),
.B1(n_3),
.B2(n_5),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_0),
.Y(n_177)
);

AO21x1_ASAP7_75t_L g180 ( 
.A1(n_163),
.A2(n_0),
.B(n_3),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_6),
.B(n_7),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_177),
.Y(n_183)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_186),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_174),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_185),
.A2(n_188),
.B(n_179),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_163),
.C(n_8),
.Y(n_188)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_181),
.B(n_180),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_190),
.A2(n_9),
.B(n_11),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_184),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_193),
.C(n_182),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_9),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_195),
.A2(n_191),
.B1(n_11),
.B2(n_12),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_194),
.A2(n_187),
.B(n_11),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_196),
.A2(n_197),
.B(n_12),
.Y(n_200)
);

OA21x2_ASAP7_75t_SL g201 ( 
.A1(n_199),
.A2(n_200),
.B(n_12),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_198),
.Y(n_202)
);


endmodule