module real_jpeg_601_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_1),
.A2(n_40),
.B1(n_41),
.B2(n_74),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_1),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_74),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_74),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_1),
.A2(n_62),
.B1(n_63),
.B2(n_74),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_51),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_51),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_2),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_3),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_120),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_120),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_120),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_4),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_5),
.B(n_52),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_5),
.B(n_25),
.C(n_27),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_5),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_5),
.B(n_24),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_5),
.B(n_59),
.C(n_62),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_209),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_5),
.B(n_110),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_5),
.B(n_64),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_209),
.Y(n_274)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_36),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_8),
.A2(n_36),
.B1(n_62),
.B2(n_63),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_8),
.A2(n_36),
.B1(n_40),
.B2(n_41),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_43),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_10),
.A2(n_43),
.B1(n_62),
.B2(n_63),
.Y(n_167)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_13),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_142),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_142),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_142),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_14),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_82),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_82),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_14),
.A2(n_62),
.B1(n_63),
.B2(n_82),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_15),
.A2(n_40),
.B1(n_41),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_15),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_174),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_174),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_15),
.A2(n_62),
.B1(n_63),
.B2(n_174),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_327),
.Y(n_17)
);

AOI21x1_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_87),
.B(n_326),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_75),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_20),
.B(n_75),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_55),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_37),
.B1(n_53),
.B2(n_54),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_22),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B(n_34),
.Y(n_22)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_23),
.B(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_30),
.Y(n_23)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_24),
.B(n_171),
.Y(n_275)
);

AO22x1_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_24)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_26),
.A2(n_27),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_27),
.B(n_248),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_32),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_31),
.B(n_199),
.Y(n_198)
);

NAND2xp33_ASAP7_75t_SL g223 ( 
.A(n_31),
.B(n_47),
.Y(n_223)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

AOI32xp33_ASAP7_75t_L g221 ( 
.A1(n_32),
.A2(n_41),
.A3(n_46),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_35),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_37),
.B(n_53),
.C(n_55),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_44),
.B1(n_50),
.B2(n_52),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_45),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_41),
.B1(n_46),
.B2(n_47),
.Y(n_49)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_41),
.A2(n_72),
.B(n_209),
.C(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_41),
.B(n_209),
.Y(n_210)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_44),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_44),
.A2(n_52),
.B1(n_141),
.B2(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_44),
.A2(n_50),
.B1(n_52),
.B2(n_330),
.Y(n_329)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_72),
.B1(n_73),
.B2(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_45),
.A2(n_81),
.B(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_45),
.B(n_119),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_45),
.A2(n_117),
.B(n_295),
.Y(n_294)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_67),
.C(n_71),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_67),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_80),
.C(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_56),
.A2(n_79),
.B1(n_84),
.B2(n_85),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_64),
.B(n_65),
.Y(n_56)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_57),
.A2(n_64),
.B1(n_115),
.B2(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_57),
.A2(n_64),
.B1(n_136),
.B2(n_165),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_57),
.A2(n_191),
.B(n_193),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_57),
.B(n_195),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_61),
.A2(n_66),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_61),
.A2(n_96),
.B1(n_97),
.B2(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_61),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_61),
.A2(n_216),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_61),
.A2(n_96),
.B1(n_192),
.B2(n_242),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_62),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_62),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_64),
.B(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_68),
.A2(n_69),
.B1(n_70),
.B2(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_68),
.A2(n_70),
.B1(n_86),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_68),
.A2(n_70),
.B1(n_94),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_68),
.A2(n_70),
.B1(n_182),
.B2(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_68),
.A2(n_274),
.B(n_275),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_68),
.A2(n_213),
.B(n_275),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_70),
.A2(n_138),
.B(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_70),
.A2(n_170),
.B(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_72),
.A2(n_140),
.B(n_143),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.C(n_83),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_76),
.A2(n_80),
.B1(n_99),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_76),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_80),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_83),
.B(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AO21x1_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_150),
.B(n_323),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_145),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_121),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_90),
.B(n_121),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_102),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_98),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_92),
.A2(n_93),
.B(n_95),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_92),
.B(n_98),
.C(n_102),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_96),
.A2(n_194),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_106),
.B(n_116),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_104),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_113),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_106),
.B1(n_116),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_105),
.A2(n_106),
.B1(n_113),
.B2(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_110),
.B(n_111),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_107),
.A2(n_110),
.B1(n_133),
.B2(n_167),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_107),
.A2(n_209),
.B(n_236),
.Y(n_256)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_108),
.A2(n_109),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_108),
.B(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_108),
.A2(n_109),
.B1(n_189),
.B2(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_108),
.A2(n_234),
.B(n_235),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_108),
.A2(n_109),
.B1(n_234),
.B2(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_109),
.A2(n_188),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_109),
.B(n_203),
.Y(n_236)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_110),
.A2(n_202),
.B(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_113),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_116),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_127),
.C(n_128),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_123),
.B1(n_127),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_137),
.C(n_139),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_130),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_131),
.A2(n_134),
.B1(n_135),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_131),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_137),
.B(n_139),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_144),
.B(n_208),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_145),
.A2(n_324),
.B(n_325),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_146),
.B(n_149),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_175),
.B(n_322),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_152),
.B(n_155),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_156),
.B(n_159),
.Y(n_320)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_161),
.B(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_168),
.C(n_172),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_162),
.A2(n_163),
.B1(n_310),
.B2(n_312),
.Y(n_309)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_164),
.B(n_166),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_165),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_167),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_168),
.A2(n_169),
.B1(n_172),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_172),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_173),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_317),
.B(n_321),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_286),
.B(n_314),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_228),
.B(n_285),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_204),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_179),
.B(n_204),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_190),
.C(n_196),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_180),
.B(n_282),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_181),
.B(n_184),
.C(n_187),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_190),
.B(n_196),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_200),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_218),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_205),
.B(n_219),
.C(n_227),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_211),
.B2(n_217),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_206),
.B(n_212),
.C(n_214),
.Y(n_299)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_210),
.Y(n_222)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_211),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_227),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_220),
.B(n_225),
.Y(n_290)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_280),
.B(n_284),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_269),
.B(n_279),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_251),
.B(n_268),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_245),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_245),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_237),
.B1(n_243),
.B2(n_244),
.Y(n_232)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_240),
.C(n_243),
.Y(n_270)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_246),
.A2(n_247),
.B1(n_249),
.B2(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_262),
.B(n_267),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_257),
.B(n_261),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_260),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_259),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_265),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_271),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_277),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_276),
.C(n_277),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_283),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_301),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_300),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_300),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_297),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_298),
.C(n_299),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_292),
.C(n_296),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_296),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_294),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_313),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_313),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_307),
.C(n_309),
.Y(n_318)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_310),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_319),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_332),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_329),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_331),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);


endmodule