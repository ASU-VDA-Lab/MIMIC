module fake_jpeg_19038_n_189 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_189);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_7),
.B(n_4),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_34),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_33),
.A2(n_20),
.B1(n_25),
.B2(n_21),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_20),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_33),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_48),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_52),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_38),
.B1(n_45),
.B2(n_62),
.Y(n_68)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_26),
.B1(n_16),
.B2(n_23),
.Y(n_88)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_41),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_81),
.C(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_67),
.B(n_71),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_27),
.B1(n_25),
.B2(n_38),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_69),
.A2(n_76),
.B1(n_63),
.B2(n_22),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_42),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_74),
.B(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_40),
.B1(n_31),
.B2(n_27),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_19),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_80),
.Y(n_103)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_78),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_19),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_32),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_36),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_85),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_44),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_29),
.C(n_18),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_24),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_90),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_44),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_43),
.B(n_53),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_9),
.B1(n_50),
.B2(n_4),
.Y(n_94)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

BUFx24_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_11),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_92),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_58),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_107),
.B1(n_108),
.B2(n_88),
.Y(n_132)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_93),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_67),
.A2(n_44),
.B1(n_55),
.B2(n_43),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_78),
.A2(n_63),
.B(n_3),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_68),
.B(n_87),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_9),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_1),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_65),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_120),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_77),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_121),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_99),
.B(n_65),
.CI(n_77),
.CON(n_122),
.SN(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_127),
.B(n_128),
.C(n_104),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_70),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_123),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_125),
.A2(n_131),
.B(n_102),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_110),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_66),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_80),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_130),
.A2(n_114),
.B(n_109),
.Y(n_135)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_115),
.B1(n_71),
.B2(n_92),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_109),
.C(n_103),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_122),
.C(n_116),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_142),
.B(n_134),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_138),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_125),
.A2(n_112),
.B(n_105),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_136),
.B(n_144),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_94),
.B1(n_107),
.B2(n_106),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_144),
.B1(n_145),
.B2(n_129),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_SL g142 ( 
.A1(n_132),
.A2(n_81),
.B(n_83),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_75),
.B1(n_90),
.B2(n_87),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_147),
.B(n_149),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_143),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_118),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_143),
.A2(n_131),
.B1(n_93),
.B2(n_96),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_152),
.A2(n_157),
.B1(n_101),
.B2(n_98),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_138),
.C(n_146),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_130),
.A3(n_122),
.B1(n_125),
.B2(n_121),
.C1(n_129),
.C2(n_96),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_154),
.A2(n_156),
.B(n_89),
.Y(n_163)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_96),
.C(n_4),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_139),
.C(n_89),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_101),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_163),
.C(n_153),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_167),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_95),
.B1(n_72),
.B2(n_124),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_170),
.B(n_173),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_161),
.A2(n_148),
.B(n_158),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_174),
.C(n_22),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_164),
.A2(n_149),
.B(n_124),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_124),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_167),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_177),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_166),
.B1(n_165),
.B2(n_162),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_124),
.B1(n_97),
.B2(n_6),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_178),
.A2(n_3),
.B(n_5),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_170),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_182),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_179),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_184),
.A2(n_3),
.B(n_5),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g185 ( 
.A(n_183),
.B(n_176),
.CI(n_175),
.CON(n_185),
.SN(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_186),
.C(n_6),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_6),
.C(n_8),
.Y(n_188)
);

BUFx24_ASAP7_75t_SL g189 ( 
.A(n_188),
.Y(n_189)
);


endmodule