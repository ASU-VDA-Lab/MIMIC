module fake_jpeg_2436_n_444 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_444);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_444;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_45),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_8),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_46),
.B(n_62),
.Y(n_100)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_50),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_31),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_51),
.B(n_78),
.Y(n_110)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_20),
.B(n_8),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_21),
.B(n_8),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_63),
.B(n_23),
.Y(n_121)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_22),
.B(n_34),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_80),
.Y(n_98)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_73),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_31),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_43),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_31),
.Y(n_82)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

BUFx24_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_85),
.Y(n_94)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_38),
.B(n_41),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_93),
.B(n_52),
.C(n_85),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_51),
.A2(n_36),
.B1(n_38),
.B2(n_43),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_95),
.A2(n_108),
.B1(n_112),
.B2(n_114),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_71),
.A2(n_32),
.B1(n_43),
.B2(n_41),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_107),
.A2(n_36),
.B1(n_74),
.B2(n_73),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_77),
.A2(n_36),
.B1(n_38),
.B2(n_43),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_29),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_109),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_45),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_55),
.A2(n_24),
.B1(n_22),
.B2(n_40),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_54),
.B(n_40),
.C(n_25),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_121),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_53),
.B(n_56),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_124),
.B(n_79),
.Y(n_159)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_137),
.Y(n_210)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_138),
.Y(n_216)
);

INVx4_ASAP7_75t_SL g139 ( 
.A(n_97),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_139),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_36),
.B1(n_19),
.B2(n_30),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_141),
.A2(n_142),
.B1(n_146),
.B2(n_179),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_86),
.B1(n_58),
.B2(n_59),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_93),
.A2(n_67),
.B1(n_60),
.B2(n_70),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_159),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

AO22x2_ASAP7_75t_L g151 ( 
.A1(n_109),
.A2(n_49),
.B1(n_50),
.B2(n_83),
.Y(n_151)
);

AO21x2_ASAP7_75t_L g192 ( 
.A1(n_151),
.A2(n_111),
.B(n_131),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_110),
.A2(n_19),
.B1(n_30),
.B2(n_23),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_153),
.Y(n_202)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_100),
.B(n_27),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_157),
.Y(n_186)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_27),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_94),
.B(n_75),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_158),
.Y(n_206)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_162),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_98),
.B(n_29),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_113),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_169),
.Y(n_199)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_117),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_76),
.B1(n_78),
.B2(n_65),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_167),
.A2(n_178),
.B1(n_136),
.B2(n_128),
.Y(n_209)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_171),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_120),
.B(n_29),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_89),
.B(n_29),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_176),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_91),
.B(n_29),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_99),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_101),
.A2(n_19),
.B1(n_28),
.B2(n_33),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_108),
.A2(n_28),
.B1(n_33),
.B2(n_2),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_95),
.A2(n_28),
.B1(n_33),
.B2(n_2),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_180),
.B(n_133),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_181),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_155),
.B(n_92),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_197),
.Y(n_225)
);

BUFx2_ASAP7_75t_SL g187 ( 
.A(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_187),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_151),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_192),
.A2(n_141),
.B1(n_142),
.B2(n_172),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_144),
.B(n_103),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_157),
.B(n_123),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_213),
.Y(n_239)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_209),
.A2(n_154),
.B1(n_156),
.B2(n_168),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_161),
.B(n_106),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_175),
.B(n_96),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_153),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_158),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_158),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_218),
.A2(n_222),
.B1(n_229),
.B2(n_234),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_165),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_221),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_166),
.B1(n_173),
.B2(n_149),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_224),
.A2(n_245),
.B(n_197),
.Y(n_261)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_203),
.A2(n_176),
.B1(n_167),
.B2(n_151),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_227),
.A2(n_215),
.B1(n_192),
.B2(n_213),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_182),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_243),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_190),
.A2(n_174),
.B1(n_151),
.B2(n_137),
.Y(n_229)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_231),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_232),
.B(n_198),
.Y(n_273)
);

AND2x2_ASAP7_75t_SL g233 ( 
.A(n_204),
.B(n_148),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_233),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_182),
.B(n_171),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_236),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_170),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_204),
.B(n_147),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_242),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_190),
.A2(n_119),
.B1(n_130),
.B2(n_177),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_240),
.A2(n_244),
.B1(n_192),
.B2(n_206),
.Y(n_265)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_241),
.Y(n_272)
);

AO22x1_ASAP7_75t_L g242 ( 
.A1(n_192),
.A2(n_130),
.B1(n_119),
.B2(n_128),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_199),
.B(n_126),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_185),
.A2(n_150),
.B1(n_99),
.B2(n_126),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_195),
.A2(n_115),
.B(n_153),
.Y(n_245)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_246),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_247),
.B(n_249),
.Y(n_267)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_189),
.Y(n_248)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_184),
.B(n_115),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_250),
.Y(n_279)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_188),
.Y(n_251)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_237),
.A2(n_191),
.B1(n_209),
.B2(n_205),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_254),
.A2(n_265),
.B1(n_266),
.B2(n_271),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_261),
.A2(n_270),
.B(n_280),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_235),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_263),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_186),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_225),
.C(n_233),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_228),
.B(n_196),
.Y(n_268)
);

OAI21x1_ASAP7_75t_L g297 ( 
.A1(n_268),
.A2(n_274),
.B(n_236),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_218),
.A2(n_192),
.B1(n_186),
.B2(n_193),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_269),
.A2(n_276),
.B1(n_265),
.B2(n_258),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_222),
.A2(n_193),
.B(n_181),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_237),
.A2(n_227),
.B1(n_246),
.B2(n_220),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_225),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_220),
.B(n_196),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_245),
.A2(n_192),
.B(n_207),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_219),
.A2(n_194),
.B1(n_216),
.B2(n_212),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_242),
.Y(n_302)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_283),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_232),
.B(n_249),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_284),
.A2(n_296),
.B(n_298),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_285),
.B(n_289),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_286),
.B(n_214),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_266),
.A2(n_229),
.B1(n_233),
.B2(n_239),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_287),
.A2(n_309),
.B1(n_272),
.B2(n_262),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_233),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_289),
.C(n_303),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_224),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_259),
.B(n_243),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_292),
.Y(n_320)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_255),
.Y(n_293)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_293),
.Y(n_334)
);

OAI32xp33_ASAP7_75t_L g294 ( 
.A1(n_276),
.A2(n_253),
.A3(n_256),
.B1(n_268),
.B2(n_274),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_279),
.Y(n_315)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_255),
.Y(n_295)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_267),
.A2(n_249),
.B(n_247),
.Y(n_296)
);

OAI21xp33_ASAP7_75t_L g322 ( 
.A1(n_297),
.A2(n_262),
.B(n_279),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_258),
.A2(n_242),
.B1(n_238),
.B2(n_240),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_256),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_300),
.B(n_311),
.Y(n_335)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_301),
.Y(n_323)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_302),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_270),
.C(n_263),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_305),
.A2(n_307),
.B1(n_308),
.B2(n_278),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_253),
.B(n_212),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_306),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_269),
.A2(n_244),
.B1(n_248),
.B2(n_250),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_280),
.A2(n_241),
.B1(n_231),
.B2(n_223),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_277),
.A2(n_226),
.B1(n_194),
.B2(n_230),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_267),
.B(n_188),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_310),
.B(n_252),
.C(n_210),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_260),
.B(n_211),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_283),
.Y(n_312)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_312),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_293),
.Y(n_313)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_313),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_315),
.A2(n_230),
.B1(n_257),
.B2(n_202),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_299),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_316),
.B(n_322),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_317),
.B(n_257),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_294),
.B(n_282),
.Y(n_319)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_319),
.Y(n_361)
);

OAI22x1_ASAP7_75t_L g324 ( 
.A1(n_298),
.A2(n_305),
.B1(n_308),
.B2(n_302),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_324),
.A2(n_325),
.B1(n_327),
.B2(n_257),
.Y(n_355)
);

OAI22x1_ASAP7_75t_SL g325 ( 
.A1(n_291),
.A2(n_282),
.B1(n_278),
.B2(n_272),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_328),
.A2(n_307),
.B1(n_301),
.B2(n_296),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_336),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_288),
.B(n_252),
.C(n_210),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_331),
.C(n_309),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_303),
.B(n_207),
.C(n_214),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_290),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_337),
.B(n_290),
.Y(n_342)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_295),
.Y(n_338)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_338),
.Y(n_351)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_339),
.Y(n_366)
);

AO22x1_ASAP7_75t_L g340 ( 
.A1(n_327),
.A2(n_304),
.B1(n_287),
.B2(n_291),
.Y(n_340)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_340),
.Y(n_368)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_342),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_343),
.B(n_357),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_315),
.A2(n_284),
.B(n_310),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_347),
.B(n_352),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_318),
.B(n_285),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_348),
.B(n_350),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_286),
.Y(n_349)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_349),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_318),
.B(n_115),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_214),
.C(n_200),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_353),
.B(n_356),
.C(n_329),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_354),
.B(n_331),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_355),
.A2(n_358),
.B1(n_328),
.B2(n_332),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_200),
.C(n_183),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_183),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_326),
.A2(n_164),
.B1(n_127),
.B2(n_122),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_313),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_360),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_333),
.A2(n_127),
.B(n_10),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_363),
.A2(n_378),
.B1(n_339),
.B2(n_345),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_369),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_317),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_370),
.B(n_323),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_346),
.B(n_333),
.C(n_325),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_371),
.B(n_376),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_346),
.B(n_324),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_377),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_344),
.B(n_335),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_375),
.B(n_356),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_349),
.B(n_320),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_312),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_361),
.A2(n_321),
.B1(n_323),
.B2(n_338),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_354),
.B(n_334),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_379),
.B(n_353),
.Y(n_384)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_383),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_384),
.B(n_390),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_374),
.A2(n_347),
.B(n_361),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_385),
.B(n_389),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_366),
.A2(n_340),
.B1(n_355),
.B2(n_357),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_386),
.A2(n_388),
.B1(n_377),
.B2(n_370),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_373),
.A2(n_360),
.B1(n_351),
.B2(n_341),
.Y(n_387)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_387),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_363),
.A2(n_340),
.B1(n_341),
.B2(n_343),
.Y(n_388)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_378),
.Y(n_391)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_391),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_365),
.B(n_314),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_393),
.B(n_365),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_380),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_394),
.B(n_371),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_362),
.A2(n_314),
.B(n_358),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_395),
.A2(n_364),
.B(n_369),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_367),
.B(n_28),
.C(n_0),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_396),
.B(n_379),
.C(n_364),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_399),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_383),
.B(n_368),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_403),
.B(n_408),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_404),
.B(n_406),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_392),
.B(n_372),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_407),
.A2(n_382),
.B1(n_386),
.B2(n_390),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_28),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_409),
.B(n_11),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_0),
.C(n_1),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_410),
.B(n_0),
.C(n_1),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_402),
.A2(n_381),
.B(n_384),
.Y(n_412)
);

OAI21x1_ASAP7_75t_L g426 ( 
.A1(n_412),
.A2(n_413),
.B(n_414),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_400),
.A2(n_396),
.B(n_395),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_398),
.A2(n_382),
.B1(n_9),
.B2(n_2),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_420),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_401),
.A2(n_33),
.B(n_9),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_418),
.A2(n_419),
.B(n_421),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_405),
.A2(n_33),
.B(n_10),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_R g421 ( 
.A(n_403),
.B(n_7),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_422),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_417),
.A2(n_399),
.B(n_398),
.Y(n_423)
);

OAI21xp33_ASAP7_75t_L g433 ( 
.A1(n_423),
.A2(n_424),
.B(n_425),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_415),
.A2(n_411),
.B(n_408),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_411),
.A2(n_407),
.B(n_405),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_421),
.B(n_410),
.C(n_397),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_428),
.B(n_420),
.Y(n_431)
);

NOR3xp33_ASAP7_75t_L g438 ( 
.A(n_431),
.B(n_434),
.C(n_435),
.Y(n_438)
);

A2O1A1O1Ixp25_ASAP7_75t_L g432 ( 
.A1(n_426),
.A2(n_11),
.B(n_3),
.C(n_4),
.D(n_5),
.Y(n_432)
);

NAND3xp33_ASAP7_75t_L g436 ( 
.A(n_432),
.B(n_430),
.C(n_3),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_429),
.B(n_6),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_427),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_436),
.A2(n_437),
.B(n_12),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_433),
.B(n_15),
.C(n_3),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_439),
.A2(n_440),
.B1(n_5),
.B2(n_13),
.Y(n_441)
);

A2O1A1O1Ixp25_ASAP7_75t_L g440 ( 
.A1(n_438),
.A2(n_12),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_441),
.A2(n_13),
.B(n_14),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_442),
.A2(n_14),
.B(n_15),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_443),
.A2(n_15),
.B(n_1),
.Y(n_444)
);


endmodule