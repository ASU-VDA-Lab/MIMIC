module fake_jpeg_23142_n_132 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_SL g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_13),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_9),
.B(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_35),
.Y(n_42)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_41),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_30),
.A2(n_24),
.B1(n_28),
.B2(n_23),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_17),
.B(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_29),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_27),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_57),
.B(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_31),
.B(n_22),
.Y(n_58)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_2),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_23),
.B(n_28),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_65),
.A2(n_67),
.B1(n_56),
.B2(n_59),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_39),
.B1(n_38),
.B2(n_40),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_74),
.B1(n_77),
.B2(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_50),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_49),
.B(n_21),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_59),
.C(n_47),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_21),
.B1(n_19),
.B2(n_16),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_2),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_45),
.B1(n_44),
.B2(n_61),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_62),
.B1(n_56),
.B2(n_47),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_77)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_81),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_6),
.Y(n_80)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_95),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_43),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_91),
.C(n_94),
.Y(n_98)
);

MAJx2_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_65),
.C(n_67),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_43),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_81),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_89),
.B(n_83),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_50),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_104),
.B(n_90),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_103),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_105),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_74),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_102),
.B(n_72),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_95),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_SL g104 ( 
.A1(n_93),
.A2(n_77),
.B(n_75),
.C(n_72),
.Y(n_104)
);

BUFx24_ASAP7_75t_SL g105 ( 
.A(n_84),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_82),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_108),
.C(n_109),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_94),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_64),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_104),
.A2(n_78),
.B1(n_90),
.B2(n_79),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_73),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_112),
.B(n_73),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_117),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_104),
.B(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_120),
.Y(n_121)
);

AOI322xp5_ASAP7_75t_SL g117 ( 
.A1(n_114),
.A2(n_78),
.A3(n_69),
.B1(n_86),
.B2(n_11),
.C1(n_10),
.C2(n_8),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_123),
.B(n_121),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_125),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_126),
.B(n_127),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_124),
.A2(n_107),
.B1(n_109),
.B2(n_69),
.Y(n_127)
);

MAJx2_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_11),
.C(n_54),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_130),
.C(n_128),
.Y(n_132)
);


endmodule