module fake_jpeg_17596_n_183 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_183);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

CKINVDCx12_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_37),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_18),
.B1(n_17),
.B2(n_27),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_18),
.B1(n_25),
.B2(n_26),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_15),
.C(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_55),
.B(n_36),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_18),
.B1(n_24),
.B2(n_17),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_56),
.A2(n_24),
.B1(n_19),
.B2(n_4),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_64),
.Y(n_81)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_71),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_62),
.A2(n_28),
.B1(n_47),
.B2(n_50),
.Y(n_78)
);

OR2x2_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_21),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_70),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_40),
.B(n_38),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_45),
.C(n_46),
.Y(n_87)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_49),
.Y(n_89)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_72),
.B1(n_24),
.B2(n_19),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_29),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_38),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_29),
.B1(n_27),
.B2(n_22),
.Y(n_72)
);

OR2x2_ASAP7_75t_SL g73 ( 
.A(n_44),
.B(n_22),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_75),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_44),
.B(n_21),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_15),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_80),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_86),
.B1(n_92),
.B2(n_65),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_15),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_28),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_45),
.B1(n_41),
.B2(n_46),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_61),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_0),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_96),
.Y(n_101)
);

INVx5_ASAP7_75t_SL g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_93),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_67),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_73),
.B(n_61),
.Y(n_112)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_95),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_57),
.C(n_56),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_77),
.C(n_79),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_103),
.Y(n_128)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_76),
.B(n_81),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_88),
.B(n_59),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_83),
.Y(n_108)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

CKINVDCx12_ASAP7_75t_R g111 ( 
.A(n_85),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_112),
.A2(n_94),
.B(n_79),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_3),
.Y(n_114)
);

AOI221xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_90),
.B1(n_62),
.B2(n_80),
.C(n_12),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_81),
.B1(n_95),
.B2(n_76),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_117),
.B1(n_126),
.B2(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_129),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_77),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_100),
.Y(n_132)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_102),
.A2(n_87),
.B1(n_86),
.B2(n_92),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_99),
.A2(n_86),
.B1(n_65),
.B2(n_69),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_101),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_130),
.B(n_103),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_114),
.C(n_13),
.Y(n_136)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_104),
.Y(n_134)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_118),
.B(n_80),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_110),
.Y(n_139)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_109),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_140),
.B(n_116),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_128),
.A2(n_113),
.B1(n_109),
.B2(n_97),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_142),
.B1(n_134),
.B2(n_132),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_113),
.B1(n_97),
.B2(n_112),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_144),
.B(n_86),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_142),
.A2(n_117),
.B(n_121),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_149),
.B(n_150),
.Y(n_159)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_118),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_148),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_86),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_151),
.B(n_156),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_129),
.C(n_115),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_133),
.C(n_127),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_154),
.A2(n_145),
.B1(n_135),
.B2(n_137),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_157),
.A2(n_150),
.B1(n_152),
.B2(n_155),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_146),
.A2(n_137),
.B(n_141),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_159),
.B(n_68),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_164),
.C(n_74),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_165),
.A2(n_167),
.B(n_168),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_153),
.B1(n_151),
.B2(n_74),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_170),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_162),
.B(n_8),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_169),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_68),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_163),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_160),
.A3(n_164),
.B1(n_9),
.B2(n_8),
.C1(n_10),
.C2(n_11),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_173),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_177),
.B(n_11),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_10),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_179),
.B(n_176),
.Y(n_181)
);

AOI221xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_180),
.B1(n_177),
.B2(n_5),
.C(n_7),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_3),
.Y(n_183)
);


endmodule