module fake_jpeg_5665_n_251 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_28),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_34),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_38),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_23),
.B1(n_15),
.B2(n_14),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_42),
.A2(n_57),
.B1(n_28),
.B2(n_18),
.Y(n_77)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_47),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_24),
.B1(n_15),
.B2(n_14),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_18),
.B1(n_22),
.B2(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_19),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_30),
.A2(n_15),
.B1(n_14),
.B2(n_24),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_18),
.B1(n_25),
.B2(n_26),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_58),
.Y(n_62)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_28),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_31),
.A2(n_24),
.B1(n_27),
.B2(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_16),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_55),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_59),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_75),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_69),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_33),
.B(n_20),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_20),
.B(n_39),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_40),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_72),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_41),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_74),
.A2(n_78),
.B1(n_42),
.B2(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_76),
.B(n_67),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_54),
.Y(n_103)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_100),
.B1(n_78),
.B2(n_68),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_94),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_97),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_42),
.B(n_54),
.C(n_48),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_91),
.B(n_61),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_42),
.C(n_46),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_90),
.C(n_94),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_46),
.Y(n_94)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_62),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_34),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_93),
.Y(n_124)
);

NAND2x1_ASAP7_75t_SL g102 ( 
.A(n_74),
.B(n_34),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_54),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_49),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_71),
.Y(n_105)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g106 ( 
.A1(n_102),
.A2(n_75),
.B1(n_61),
.B2(n_39),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_116),
.B(n_90),
.Y(n_140)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_110),
.B(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_59),
.Y(n_112)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_64),
.Y(n_113)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_72),
.Y(n_114)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_76),
.Y(n_115)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_65),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_117),
.B(n_122),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_78),
.B1(n_80),
.B2(n_62),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_102),
.A2(n_39),
.B1(n_32),
.B2(n_31),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_83),
.B1(n_103),
.B2(n_95),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_65),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_79),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_103),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_126),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_34),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_137),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_125),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_98),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_126),
.C(n_109),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_116),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_141),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_87),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_143),
.B(n_148),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_110),
.B1(n_120),
.B2(n_118),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_106),
.A2(n_91),
.B1(n_83),
.B2(n_31),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g155 ( 
.A1(n_146),
.A2(n_121),
.B(n_118),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_86),
.B1(n_96),
.B2(n_92),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_147),
.A2(n_88),
.B1(n_83),
.B2(n_89),
.Y(n_158)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_92),
.B(n_96),
.C(n_88),
.D(n_34),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_153),
.C(n_161),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_160),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_123),
.C(n_109),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_108),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_166),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_115),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_159),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_157),
.A2(n_158),
.B1(n_130),
.B2(n_129),
.Y(n_184)
);

NAND2xp33_ASAP7_75t_SL g159 ( 
.A(n_146),
.B(n_0),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_132),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_48),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_89),
.B1(n_79),
.B2(n_32),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_162),
.A2(n_167),
.B1(n_145),
.B2(n_134),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_53),
.Y(n_165)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_142),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_79),
.B1(n_32),
.B2(n_51),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_23),
.Y(n_168)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_177),
.B1(n_163),
.B2(n_21),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_149),
.A2(n_144),
.B1(n_147),
.B2(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_185),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_143),
.B1(n_144),
.B2(n_139),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_179),
.A2(n_184),
.B1(n_167),
.B2(n_164),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_143),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_181),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_140),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_135),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_186),
.C(n_171),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_163),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_53),
.C(n_48),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_20),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_172),
.A2(n_149),
.B1(n_159),
.B2(n_155),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_188),
.A2(n_191),
.B1(n_198),
.B2(n_23),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_183),
.A2(n_158),
.B(n_169),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_189),
.A2(n_193),
.B(n_0),
.Y(n_209)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_190),
.B(n_202),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_175),
.A2(n_155),
.B1(n_169),
.B2(n_162),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_200),
.C(n_196),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

O2A1O1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_182),
.B(n_173),
.C(n_21),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_176),
.B(n_21),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_200),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_51),
.C(n_23),
.Y(n_200)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_201),
.Y(n_210)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_180),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_206),
.C(n_213),
.Y(n_221)
);

AO21x1_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_176),
.B(n_181),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_204),
.A2(n_209),
.B(n_214),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_207),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_212),
.A2(n_188),
.B1(n_191),
.B2(n_8),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_7),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_7),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_215),
.Y(n_224)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_211),
.Y(n_217)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_217),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_205),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_219),
.B(n_222),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_204),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_225),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_210),
.B(n_206),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_212),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_213),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_228),
.A2(n_229),
.B(n_230),
.Y(n_237)
);

NOR2xp67_ASAP7_75t_SL g229 ( 
.A(n_221),
.B(n_203),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_6),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_231),
.B(n_8),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_0),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_238),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_227),
.A2(n_223),
.B1(n_6),
.B2(n_10),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_236),
.C(n_239),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_233),
.A2(n_6),
.B(n_12),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_10),
.B(n_12),
.Y(n_239)
);

AOI21xp33_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_226),
.B(n_11),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_243),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

AOI322xp5_ASAP7_75t_L g244 ( 
.A1(n_237),
.A2(n_5),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_2),
.C2(n_3),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_5),
.Y(n_246)
);

O2A1O1Ixp33_ASAP7_75t_SL g249 ( 
.A1(n_246),
.A2(n_1),
.B(n_13),
.C(n_245),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_11),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_240),
.C(n_2),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_249),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_1),
.Y(n_251)
);


endmodule