module fake_aes_2958_n_1382 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_241, n_95, n_238, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1382);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_241;
input n_95;
input n_238;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1382;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_1363;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g316 ( .A(n_264), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_239), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_259), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_56), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_83), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_16), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_14), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_223), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_291), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_193), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_55), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_115), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_58), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_148), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_31), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_248), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_133), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_190), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_165), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g335 ( .A(n_272), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_146), .Y(n_336) );
INVxp33_ASAP7_75t_SL g337 ( .A(n_246), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_124), .Y(n_338) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_89), .Y(n_339) );
CKINVDCx14_ASAP7_75t_R g340 ( .A(n_152), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_163), .Y(n_341) );
INVxp67_ASAP7_75t_L g342 ( .A(n_117), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_255), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_59), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_253), .Y(n_345) );
INVxp67_ASAP7_75t_SL g346 ( .A(n_195), .Y(n_346) );
INVxp33_ASAP7_75t_SL g347 ( .A(n_186), .Y(n_347) );
CKINVDCx14_ASAP7_75t_R g348 ( .A(n_249), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_69), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_228), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_285), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_221), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_45), .B(n_64), .Y(n_353) );
INVx4_ASAP7_75t_R g354 ( .A(n_103), .Y(n_354) );
CKINVDCx16_ASAP7_75t_R g355 ( .A(n_97), .Y(n_355) );
CKINVDCx20_ASAP7_75t_R g356 ( .A(n_260), .Y(n_356) );
BUFx2_ASAP7_75t_SL g357 ( .A(n_28), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_300), .Y(n_358) );
CKINVDCx14_ASAP7_75t_R g359 ( .A(n_2), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_20), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_44), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_313), .Y(n_362) );
CKINVDCx16_ASAP7_75t_R g363 ( .A(n_50), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_12), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_308), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_32), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_42), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_184), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_188), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_209), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_153), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_132), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_234), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_293), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_256), .Y(n_375) );
INVxp67_ASAP7_75t_L g376 ( .A(n_306), .Y(n_376) );
INVxp67_ASAP7_75t_L g377 ( .A(n_267), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_48), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_76), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_182), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_3), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_7), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_35), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_98), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_61), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_303), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_122), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_179), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_233), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_73), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_141), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_301), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_112), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_244), .Y(n_394) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_262), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_126), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_217), .Y(n_397) );
CKINVDCx16_ASAP7_75t_R g398 ( .A(n_198), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_63), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_40), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_55), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_160), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_104), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_86), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_298), .Y(n_405) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_79), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_22), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_92), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_150), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_206), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_238), .Y(n_411) );
BUFx3_ASAP7_75t_L g412 ( .A(n_136), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_13), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_108), .Y(n_414) );
BUFx3_ASAP7_75t_L g415 ( .A(n_174), .Y(n_415) );
CKINVDCx14_ASAP7_75t_R g416 ( .A(n_219), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_96), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_279), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_216), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_9), .Y(n_420) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_81), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_147), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_4), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_114), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_84), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_155), .Y(n_426) );
CKINVDCx16_ASAP7_75t_R g427 ( .A(n_203), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_18), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_247), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_314), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_72), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_56), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_68), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_47), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_315), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_289), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_109), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_30), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_286), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_296), .Y(n_440) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_243), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_106), .Y(n_442) );
CKINVDCx14_ASAP7_75t_R g443 ( .A(n_311), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_62), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_236), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_21), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_181), .Y(n_447) );
BUFx2_ASAP7_75t_L g448 ( .A(n_99), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_225), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_169), .Y(n_450) );
NOR2xp67_ASAP7_75t_L g451 ( .A(n_143), .B(n_197), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_35), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_120), .Y(n_453) );
CKINVDCx14_ASAP7_75t_R g454 ( .A(n_131), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_142), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_105), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_25), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_28), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_295), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_85), .Y(n_460) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_180), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_183), .Y(n_462) );
INVxp67_ASAP7_75t_SL g463 ( .A(n_222), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_139), .Y(n_464) );
CKINVDCx16_ASAP7_75t_R g465 ( .A(n_101), .Y(n_465) );
BUFx2_ASAP7_75t_L g466 ( .A(n_144), .Y(n_466) );
BUFx2_ASAP7_75t_L g467 ( .A(n_135), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_138), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_53), .Y(n_469) );
INVxp33_ASAP7_75t_SL g470 ( .A(n_23), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_66), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_382), .B(n_0), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_362), .B(n_0), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_362), .B(n_1), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_318), .Y(n_475) );
BUFx3_ASAP7_75t_L g476 ( .A(n_365), .Y(n_476) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_385), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_321), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_359), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_321), .B(n_1), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_383), .Y(n_481) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_385), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_359), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_318), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_382), .B(n_2), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_341), .B(n_3), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_349), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_363), .Y(n_488) );
INVx4_ASAP7_75t_L g489 ( .A(n_411), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_383), .Y(n_490) );
BUFx2_ASAP7_75t_L g491 ( .A(n_448), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_355), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_434), .Y(n_493) );
OAI22xp5_ASAP7_75t_SL g494 ( .A1(n_364), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_434), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_466), .B(n_8), .Y(n_496) );
OAI22xp5_ASAP7_75t_SL g497 ( .A1(n_364), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_497) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_385), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_316), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_398), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_349), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_317), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_467), .B(n_10), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_427), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_372), .Y(n_505) );
INVx6_ASAP7_75t_L g506 ( .A(n_385), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_320), .Y(n_507) );
AO22x2_ASAP7_75t_L g508 ( .A1(n_473), .A2(n_357), .B1(n_328), .B2(n_319), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_483), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_475), .Y(n_510) );
OAI22xp5_ASAP7_75t_SL g511 ( .A1(n_494), .A2(n_470), .B1(n_335), .B2(n_439), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_475), .Y(n_512) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_477), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_489), .B(n_461), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_489), .B(n_342), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_489), .B(n_491), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_477), .Y(n_517) );
AND2x2_ASAP7_75t_SL g518 ( .A(n_473), .B(n_465), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_477), .Y(n_519) );
INVx3_ASAP7_75t_L g520 ( .A(n_480), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_473), .B(n_360), .Y(n_521) );
INVxp67_ASAP7_75t_SL g522 ( .A(n_485), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_483), .B(n_376), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_491), .B(n_377), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_500), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_484), .Y(n_526) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_477), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_484), .Y(n_528) );
INVx3_ASAP7_75t_L g529 ( .A(n_480), .Y(n_529) );
INVx4_ASAP7_75t_L g530 ( .A(n_474), .Y(n_530) );
AND2x6_ASAP7_75t_L g531 ( .A(n_474), .B(n_353), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_487), .Y(n_532) );
INVx3_ASAP7_75t_L g533 ( .A(n_480), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_474), .B(n_324), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_496), .A2(n_339), .B1(n_439), .B2(n_335), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_477), .Y(n_536) );
INVxp67_ASAP7_75t_L g537 ( .A(n_500), .Y(n_537) );
AND2x4_ASAP7_75t_L g538 ( .A(n_496), .B(n_361), .Y(n_538) );
OAI22xp33_ASAP7_75t_SL g539 ( .A1(n_492), .A2(n_330), .B1(n_400), .B2(n_326), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_496), .B(n_366), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_487), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_482), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_476), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_501), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_501), .Y(n_545) );
BUFx3_ASAP7_75t_L g546 ( .A(n_476), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_505), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_505), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_482), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_482), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_482), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_546), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_520), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_520), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_520), .Y(n_555) );
INVx4_ASAP7_75t_L g556 ( .A(n_531), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_546), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_522), .B(n_503), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_534), .A2(n_503), .B(n_502), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_543), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_530), .B(n_486), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_530), .B(n_486), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_530), .B(n_503), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_518), .B(n_504), .Y(n_564) );
BUFx3_ASAP7_75t_L g565 ( .A(n_543), .Y(n_565) );
NAND2x1p5_ASAP7_75t_L g566 ( .A(n_518), .B(n_472), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_529), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_508), .A2(n_472), .B1(n_504), .B2(n_479), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_510), .Y(n_569) );
INVx5_ASAP7_75t_L g570 ( .A(n_531), .Y(n_570) );
O2A1O1Ixp5_ASAP7_75t_L g571 ( .A1(n_529), .A2(n_502), .B(n_507), .C(n_499), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_538), .B(n_337), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_538), .B(n_347), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_529), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_538), .B(n_485), .Y(n_575) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_531), .Y(n_576) );
INVx3_ASAP7_75t_L g577 ( .A(n_533), .Y(n_577) );
AND2x4_ASAP7_75t_L g578 ( .A(n_540), .B(n_499), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_521), .B(n_507), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_508), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_533), .Y(n_581) );
AOI21xp33_ASAP7_75t_L g582 ( .A1(n_516), .A2(n_348), .B(n_340), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_521), .B(n_340), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_533), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_510), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_514), .B(n_488), .Y(n_586) );
NOR2x1p5_ASAP7_75t_L g587 ( .A(n_525), .B(n_407), .Y(n_587) );
INVx3_ASAP7_75t_L g588 ( .A(n_512), .Y(n_588) );
NOR2xp33_ASAP7_75t_SL g589 ( .A(n_509), .B(n_339), .Y(n_589) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_531), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_512), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_525), .Y(n_592) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_535), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_521), .B(n_348), .Y(n_594) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_508), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_540), .B(n_327), .Y(n_596) );
INVxp67_ASAP7_75t_L g597 ( .A(n_531), .Y(n_597) );
BUFx2_ASAP7_75t_L g598 ( .A(n_508), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_531), .A2(n_443), .B1(n_454), .B2(n_416), .Y(n_599) );
A2O1A1Ixp33_ASAP7_75t_L g600 ( .A1(n_526), .A2(n_481), .B(n_490), .C(n_478), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_526), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_528), .Y(n_602) );
INVx4_ASAP7_75t_L g603 ( .A(n_540), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_515), .B(n_333), .Y(n_604) );
INVx6_ASAP7_75t_L g605 ( .A(n_513), .Y(n_605) );
BUFx3_ASAP7_75t_L g606 ( .A(n_528), .Y(n_606) );
INVxp67_ASAP7_75t_L g607 ( .A(n_532), .Y(n_607) );
AND2x4_ASAP7_75t_L g608 ( .A(n_523), .B(n_459), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_532), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_524), .B(n_416), .Y(n_610) );
BUFx3_ASAP7_75t_L g611 ( .A(n_541), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_541), .Y(n_612) );
NAND2x1p5_ASAP7_75t_L g613 ( .A(n_544), .B(n_367), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_539), .A2(n_459), .B1(n_497), .B2(n_356), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_544), .A2(n_374), .B(n_372), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_545), .B(n_443), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_545), .B(n_454), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_547), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_547), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_548), .B(n_346), .Y(n_620) );
CKINVDCx5p33_ASAP7_75t_R g621 ( .A(n_537), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_548), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g623 ( .A(n_511), .Y(n_623) );
OR2x6_ASAP7_75t_L g624 ( .A(n_517), .B(n_378), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_517), .A2(n_399), .B1(n_429), .B2(n_332), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_519), .B(n_395), .Y(n_626) );
INVx3_ASAP7_75t_L g627 ( .A(n_513), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_519), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_536), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_536), .Y(n_630) );
INVx2_ASAP7_75t_SL g631 ( .A(n_613), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_606), .Y(n_632) );
INVx4_ASAP7_75t_L g633 ( .A(n_570), .Y(n_633) );
AO21x1_ASAP7_75t_L g634 ( .A1(n_615), .A2(n_325), .B(n_323), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_611), .Y(n_635) );
OR2x6_ASAP7_75t_L g636 ( .A(n_566), .B(n_381), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_577), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_612), .B(n_445), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_577), .Y(n_639) );
A2O1A1Ixp33_ASAP7_75t_SL g640 ( .A1(n_599), .A2(n_495), .B(n_481), .C(n_490), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_553), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_588), .Y(n_642) );
INVx2_ASAP7_75t_SL g643 ( .A(n_613), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_607), .B(n_413), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_SL g645 ( .A1(n_582), .A2(n_495), .B(n_493), .C(n_478), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_576), .B(n_344), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_586), .B(n_432), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_607), .B(n_578), .Y(n_648) );
BUFx3_ASAP7_75t_L g649 ( .A(n_621), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_598), .A2(n_420), .B1(n_423), .B2(n_401), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_580), .A2(n_493), .B(n_438), .C(n_446), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_554), .Y(n_652) );
O2A1O1Ixp33_ASAP7_75t_L g653 ( .A1(n_580), .A2(n_452), .B(n_457), .C(n_428), .Y(n_653) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_592), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_588), .Y(n_655) );
OAI21x1_ASAP7_75t_L g656 ( .A1(n_571), .A2(n_384), .B(n_374), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_564), .B(n_458), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_563), .A2(n_463), .B(n_331), .Y(n_658) );
BUFx12f_ASAP7_75t_L g659 ( .A(n_587), .Y(n_659) );
INVx4_ASAP7_75t_L g660 ( .A(n_570), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_568), .A2(n_595), .B1(n_566), .B2(n_575), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_572), .B(n_469), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_563), .A2(n_334), .B(n_329), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_555), .Y(n_664) );
BUFx10_ASAP7_75t_L g665 ( .A(n_558), .Y(n_665) );
INVx4_ASAP7_75t_L g666 ( .A(n_570), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_569), .Y(n_667) );
A2O1A1Ixp33_ASAP7_75t_L g668 ( .A1(n_571), .A2(n_336), .B(n_343), .C(n_338), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_567), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_561), .A2(n_351), .B(n_345), .Y(n_670) );
BUFx8_ASAP7_75t_L g671 ( .A(n_608), .Y(n_671) );
INVx3_ASAP7_75t_L g672 ( .A(n_556), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_561), .A2(n_358), .B(n_352), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_585), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_591), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_574), .Y(n_676) );
INVx4_ASAP7_75t_L g677 ( .A(n_570), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_576), .B(n_350), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_558), .A2(n_322), .B1(n_495), .B2(n_369), .Y(n_679) );
INVx3_ASAP7_75t_L g680 ( .A(n_556), .Y(n_680) );
OAI221xp5_ASAP7_75t_L g681 ( .A1(n_579), .A2(n_442), .B1(n_368), .B2(n_370), .C(n_371), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_601), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_581), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_562), .A2(n_375), .B(n_373), .Y(n_684) );
BUFx3_ASAP7_75t_L g685 ( .A(n_552), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_578), .A2(n_322), .B1(n_380), .B2(n_379), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_562), .B(n_387), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_576), .B(n_388), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_589), .B(n_322), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_584), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_609), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_590), .B(n_418), .Y(n_692) );
INVx1_ASAP7_75t_SL g693 ( .A(n_590), .Y(n_693) );
O2A1O1Ixp33_ASAP7_75t_L g694 ( .A1(n_600), .A2(n_579), .B(n_610), .C(n_616), .Y(n_694) );
NOR2xp67_ASAP7_75t_L g695 ( .A(n_614), .B(n_11), .Y(n_695) );
AND2x4_ASAP7_75t_SL g696 ( .A(n_603), .B(n_322), .Y(n_696) );
AOI21x1_ASAP7_75t_L g697 ( .A1(n_615), .A2(n_549), .B(n_542), .Y(n_697) );
INVx2_ASAP7_75t_SL g698 ( .A(n_603), .Y(n_698) );
INVx3_ASAP7_75t_L g699 ( .A(n_590), .Y(n_699) );
A2O1A1Ixp33_ASAP7_75t_SL g700 ( .A1(n_610), .A2(n_549), .B(n_550), .C(n_542), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_619), .Y(n_701) );
CKINVDCx16_ASAP7_75t_R g702 ( .A(n_625), .Y(n_702) );
INVx4_ASAP7_75t_L g703 ( .A(n_624), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_602), .B(n_389), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_618), .Y(n_705) );
A2O1A1Ixp33_ASAP7_75t_L g706 ( .A1(n_559), .A2(n_391), .B(n_392), .C(n_390), .Y(n_706) );
BUFx2_ASAP7_75t_L g707 ( .A(n_608), .Y(n_707) );
AND2x4_ASAP7_75t_L g708 ( .A(n_596), .B(n_393), .Y(n_708) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_622), .Y(n_709) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_624), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_559), .B(n_620), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_616), .A2(n_397), .B(n_394), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_617), .A2(n_403), .B(n_402), .Y(n_713) );
BUFx3_ASAP7_75t_L g714 ( .A(n_557), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_620), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_560), .Y(n_716) );
BUFx2_ASAP7_75t_L g717 ( .A(n_597), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_617), .B(n_404), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_624), .Y(n_719) );
AND2x4_ASAP7_75t_L g720 ( .A(n_573), .B(n_405), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_583), .B(n_409), .Y(n_721) );
INVxp67_ASAP7_75t_L g722 ( .A(n_583), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_597), .A2(n_414), .B1(n_417), .B2(n_410), .Y(n_723) );
INVx3_ASAP7_75t_L g724 ( .A(n_565), .Y(n_724) );
INVx4_ASAP7_75t_L g725 ( .A(n_605), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_594), .B(n_419), .Y(n_726) );
INVx1_ASAP7_75t_SL g727 ( .A(n_594), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_626), .Y(n_728) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_593), .Y(n_729) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_623), .Y(n_730) );
CKINVDCx5p33_ASAP7_75t_R g731 ( .A(n_604), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_626), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_629), .A2(n_426), .B1(n_430), .B2(n_424), .Y(n_733) );
INVx2_ASAP7_75t_SL g734 ( .A(n_605), .Y(n_734) );
NOR3xp33_ASAP7_75t_L g735 ( .A(n_630), .B(n_456), .C(n_433), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_628), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_627), .B(n_11), .Y(n_737) );
INVx2_ASAP7_75t_SL g738 ( .A(n_605), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_627), .B(n_422), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_577), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_606), .Y(n_741) );
INVx3_ASAP7_75t_L g742 ( .A(n_710), .Y(n_742) );
OAI21x1_ASAP7_75t_L g743 ( .A1(n_697), .A2(n_386), .B(n_384), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_705), .Y(n_744) );
AOI21xp33_ASAP7_75t_L g745 ( .A1(n_645), .A2(n_436), .B(n_431), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_654), .B(n_12), .Y(n_746) );
NAND2x1p5_ASAP7_75t_L g747 ( .A(n_703), .B(n_365), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_681), .A2(n_447), .B1(n_450), .B2(n_437), .Y(n_748) );
OAI21x1_ASAP7_75t_L g749 ( .A1(n_656), .A2(n_711), .B(n_712), .Y(n_749) );
OAI221xp5_ASAP7_75t_L g750 ( .A1(n_722), .A2(n_468), .B1(n_455), .B2(n_453), .C(n_471), .Y(n_750) );
AO32x2_ASAP7_75t_L g751 ( .A1(n_631), .A2(n_506), .A3(n_498), .B1(n_482), .B2(n_451), .Y(n_751) );
BUFx4f_ASAP7_75t_SL g752 ( .A(n_659), .Y(n_752) );
OAI21x1_ASAP7_75t_L g753 ( .A1(n_711), .A2(n_396), .B(n_386), .Y(n_753) );
OAI21x1_ASAP7_75t_L g754 ( .A1(n_712), .A2(n_408), .B(n_396), .Y(n_754) );
OA21x2_ASAP7_75t_L g755 ( .A1(n_668), .A2(n_425), .B(n_408), .Y(n_755) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_710), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_709), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_713), .A2(n_464), .B(n_425), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g759 ( .A1(n_681), .A2(n_464), .B1(n_415), .B2(n_412), .Y(n_759) );
OAI21x1_ASAP7_75t_L g760 ( .A1(n_713), .A2(n_551), .B(n_550), .Y(n_760) );
AO21x2_ASAP7_75t_L g761 ( .A1(n_700), .A2(n_551), .B(n_498), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_715), .Y(n_762) );
AOI21xp5_ASAP7_75t_L g763 ( .A1(n_694), .A2(n_527), .B(n_513), .Y(n_763) );
OAI21x1_ASAP7_75t_L g764 ( .A1(n_663), .A2(n_421), .B(n_406), .Y(n_764) );
AOI21x1_ASAP7_75t_L g765 ( .A1(n_634), .A2(n_354), .B(n_406), .Y(n_765) );
INVx4_ASAP7_75t_L g766 ( .A(n_710), .Y(n_766) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_703), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_704), .Y(n_768) );
INVxp67_ASAP7_75t_SL g769 ( .A(n_648), .Y(n_769) );
A2O1A1Ixp33_ASAP7_75t_L g770 ( .A1(n_694), .A2(n_412), .B(n_415), .C(n_406), .Y(n_770) );
BUFx2_ASAP7_75t_L g771 ( .A(n_649), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_667), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_674), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_704), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_648), .A2(n_406), .B1(n_421), .B2(n_441), .Y(n_775) );
INVx5_ASAP7_75t_L g776 ( .A(n_665), .Y(n_776) );
CKINVDCx5p33_ASAP7_75t_R g777 ( .A(n_671), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_641), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_652), .Y(n_779) );
OAI21x1_ASAP7_75t_L g780 ( .A1(n_663), .A2(n_441), .B(n_421), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_675), .Y(n_781) );
OAI21x1_ASAP7_75t_L g782 ( .A1(n_670), .A2(n_441), .B(n_421), .Y(n_782) );
NAND2xp5_ASAP7_75t_SL g783 ( .A(n_643), .B(n_441), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_664), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_669), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_671), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_676), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_683), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_690), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_636), .B(n_13), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_716), .Y(n_791) );
INVx4_ASAP7_75t_L g792 ( .A(n_665), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_687), .A2(n_506), .B1(n_435), .B2(n_460), .Y(n_793) );
OR2x6_ASAP7_75t_L g794 ( .A(n_636), .B(n_506), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_732), .Y(n_795) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_658), .A2(n_444), .B(n_440), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_682), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_636), .B(n_14), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_691), .Y(n_799) );
AND2x4_ASAP7_75t_L g800 ( .A(n_724), .B(n_15), .Y(n_800) );
OAI21x1_ASAP7_75t_L g801 ( .A1(n_670), .A2(n_65), .B(n_60), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_661), .B(n_15), .Y(n_802) );
BUFx6f_ASAP7_75t_L g803 ( .A(n_633), .Y(n_803) );
O2A1O1Ixp33_ASAP7_75t_SL g804 ( .A1(n_640), .A2(n_170), .B(n_254), .C(n_252), .Y(n_804) );
OAI21x1_ASAP7_75t_L g805 ( .A1(n_673), .A2(n_70), .B(n_67), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_707), .B(n_16), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_701), .Y(n_807) );
O2A1O1Ixp33_ASAP7_75t_SL g808 ( .A1(n_706), .A2(n_171), .B(n_257), .C(n_251), .Y(n_808) );
AOI22xp33_ASAP7_75t_SL g809 ( .A1(n_702), .A2(n_449), .B1(n_462), .B2(n_506), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_728), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_638), .B(n_17), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_687), .Y(n_812) );
O2A1O1Ixp33_ASAP7_75t_L g813 ( .A1(n_651), .A2(n_17), .B(n_18), .C(n_19), .Y(n_813) );
INVx2_ASAP7_75t_L g814 ( .A(n_737), .Y(n_814) );
OAI21x1_ASAP7_75t_L g815 ( .A1(n_673), .A2(n_74), .B(n_71), .Y(n_815) );
BUFx3_ASAP7_75t_L g816 ( .A(n_696), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_736), .Y(n_817) );
OAI21x1_ASAP7_75t_L g818 ( .A1(n_684), .A2(n_77), .B(n_75), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_638), .A2(n_498), .B1(n_513), .B2(n_527), .Y(n_819) );
AOI221xp5_ASAP7_75t_L g820 ( .A1(n_662), .A2(n_498), .B1(n_527), .B2(n_513), .C(n_22), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_689), .Y(n_821) );
NOR2x1_ASAP7_75t_R g822 ( .A(n_731), .B(n_19), .Y(n_822) );
INVx2_ASAP7_75t_L g823 ( .A(n_642), .Y(n_823) );
INVx2_ASAP7_75t_SL g824 ( .A(n_724), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_655), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_718), .Y(n_826) );
OAI21x1_ASAP7_75t_L g827 ( .A1(n_684), .A2(n_80), .B(n_78), .Y(n_827) );
BUFx8_ASAP7_75t_L g828 ( .A(n_708), .Y(n_828) );
AND2x4_ASAP7_75t_L g829 ( .A(n_722), .B(n_20), .Y(n_829) );
OAI21xp5_ASAP7_75t_L g830 ( .A1(n_658), .A2(n_498), .B(n_527), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_727), .B(n_21), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_718), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_721), .Y(n_833) );
INVx2_ASAP7_75t_L g834 ( .A(n_639), .Y(n_834) );
INVx2_ASAP7_75t_SL g835 ( .A(n_708), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_637), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_721), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_727), .A2(n_527), .B1(n_24), .B2(n_25), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_650), .B(n_23), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_644), .Y(n_840) );
OAI21x1_ASAP7_75t_SL g841 ( .A1(n_651), .A2(n_24), .B(n_26), .Y(n_841) );
AOI21x1_ASAP7_75t_L g842 ( .A1(n_726), .A2(n_87), .B(n_82), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_644), .Y(n_843) );
BUFx3_ASAP7_75t_L g844 ( .A(n_685), .Y(n_844) );
INVx3_ASAP7_75t_L g845 ( .A(n_633), .Y(n_845) );
OAI21x1_ASAP7_75t_L g846 ( .A1(n_740), .A2(n_90), .B(n_88), .Y(n_846) );
BUFx3_ASAP7_75t_L g847 ( .A(n_714), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_720), .Y(n_848) );
OAI21x1_ASAP7_75t_L g849 ( .A1(n_719), .A2(n_93), .B(n_91), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_695), .A2(n_26), .B1(n_27), .B2(n_29), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_720), .Y(n_851) );
AOI21xp5_ASAP7_75t_L g852 ( .A1(n_653), .A2(n_95), .B(n_94), .Y(n_852) );
A2O1A1Ixp33_ASAP7_75t_L g853 ( .A1(n_653), .A2(n_27), .B(n_29), .C(n_30), .Y(n_853) );
INVx2_ASAP7_75t_SL g854 ( .A(n_729), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_647), .B(n_31), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_657), .A2(n_32), .B1(n_33), .B2(n_34), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_730), .B(n_33), .Y(n_857) );
OAI22xp33_ASAP7_75t_L g858 ( .A1(n_723), .A2(n_34), .B1(n_36), .B2(n_37), .Y(n_858) );
OAI21xp5_ASAP7_75t_L g859 ( .A1(n_679), .A2(n_36), .B(n_37), .Y(n_859) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_693), .Y(n_860) );
INVx2_ASAP7_75t_L g861 ( .A(n_632), .Y(n_861) );
OAI21x1_ASAP7_75t_L g862 ( .A1(n_672), .A2(n_102), .B(n_100), .Y(n_862) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_693), .Y(n_863) );
OAI21x1_ASAP7_75t_L g864 ( .A1(n_672), .A2(n_199), .B(n_310), .Y(n_864) );
AOI21xp5_ASAP7_75t_L g865 ( .A1(n_646), .A2(n_196), .B(n_309), .Y(n_865) );
BUFx2_ASAP7_75t_L g866 ( .A(n_828), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_802), .A2(n_735), .B1(n_635), .B2(n_741), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_802), .A2(n_686), .B1(n_717), .B2(n_733), .Y(n_868) );
BUFx8_ASAP7_75t_L g869 ( .A(n_771), .Y(n_869) );
AOI22xp33_ASAP7_75t_SL g870 ( .A1(n_790), .A2(n_680), .B1(n_666), .B2(n_677), .Y(n_870) );
OR2x6_ASAP7_75t_L g871 ( .A(n_794), .B(n_698), .Y(n_871) );
NAND2x1_ASAP7_75t_L g872 ( .A(n_803), .B(n_660), .Y(n_872) );
AOI22xp33_ASAP7_75t_SL g873 ( .A1(n_798), .A2(n_680), .B1(n_666), .B2(n_677), .Y(n_873) );
BUFx6f_ASAP7_75t_L g874 ( .A(n_803), .Y(n_874) );
AOI221xp5_ASAP7_75t_L g875 ( .A1(n_840), .A2(n_678), .B1(n_688), .B2(n_692), .C(n_739), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_769), .A2(n_699), .B1(n_660), .B2(n_725), .Y(n_876) );
INVx2_ASAP7_75t_SL g877 ( .A(n_776), .Y(n_877) );
INVx2_ASAP7_75t_SL g878 ( .A(n_776), .Y(n_878) );
AOI22xp33_ASAP7_75t_SL g879 ( .A1(n_829), .A2(n_699), .B1(n_725), .B2(n_734), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_812), .B(n_738), .Y(n_880) );
AND2x4_ASAP7_75t_L g881 ( .A(n_769), .B(n_38), .Y(n_881) );
AOI22xp33_ASAP7_75t_SL g882 ( .A1(n_829), .A2(n_38), .B1(n_39), .B2(n_40), .Y(n_882) );
AOI21xp5_ASAP7_75t_L g883 ( .A1(n_763), .A2(n_200), .B(n_307), .Y(n_883) );
OAI221xp5_ASAP7_75t_L g884 ( .A1(n_835), .A2(n_39), .B1(n_41), .B2(n_42), .C(n_43), .Y(n_884) );
HB1xp67_ASAP7_75t_L g885 ( .A(n_828), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_826), .B(n_41), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_832), .A2(n_43), .B1(n_44), .B2(n_45), .Y(n_887) );
INVx2_ASAP7_75t_L g888 ( .A(n_762), .Y(n_888) );
CKINVDCx5p33_ASAP7_75t_R g889 ( .A(n_786), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_768), .A2(n_46), .B1(n_47), .B2(n_48), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_833), .A2(n_46), .B1(n_49), .B2(n_50), .Y(n_891) );
OAI22xp33_ASAP7_75t_L g892 ( .A1(n_750), .A2(n_49), .B1(n_51), .B2(n_52), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_795), .B(n_51), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_810), .Y(n_894) );
AOI21xp5_ASAP7_75t_L g895 ( .A1(n_763), .A2(n_208), .B(n_305), .Y(n_895) );
OR2x2_ASAP7_75t_L g896 ( .A(n_854), .B(n_52), .Y(n_896) );
AOI21xp5_ASAP7_75t_L g897 ( .A1(n_830), .A2(n_210), .B(n_304), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_837), .A2(n_53), .B1(n_54), .B2(n_57), .Y(n_898) );
OAI221xp5_ASAP7_75t_L g899 ( .A1(n_843), .A2(n_54), .B1(n_57), .B2(n_58), .C(n_107), .Y(n_899) );
OAI221xp5_ASAP7_75t_L g900 ( .A1(n_809), .A2(n_110), .B1(n_111), .B2(n_113), .C(n_116), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_774), .A2(n_118), .B1(n_119), .B2(n_121), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_748), .A2(n_123), .B1(n_125), .B2(n_127), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_848), .B(n_312), .Y(n_903) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_748), .A2(n_128), .B1(n_129), .B2(n_130), .Y(n_904) );
OAI33xp33_ASAP7_75t_L g905 ( .A1(n_858), .A2(n_134), .A3(n_137), .B1(n_140), .B2(n_145), .B3(n_149), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_757), .B(n_151), .Y(n_906) );
AOI221xp5_ASAP7_75t_L g907 ( .A1(n_750), .A2(n_154), .B1(n_156), .B2(n_157), .C(n_158), .Y(n_907) );
AND2x2_ASAP7_75t_L g908 ( .A(n_746), .B(n_159), .Y(n_908) );
OAI221xp5_ASAP7_75t_L g909 ( .A1(n_809), .A2(n_161), .B1(n_162), .B2(n_164), .C(n_166), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_744), .Y(n_910) );
AND2x2_ASAP7_75t_L g911 ( .A(n_851), .B(n_167), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_759), .A2(n_168), .B1(n_172), .B2(n_173), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_811), .A2(n_175), .B1(n_176), .B2(n_177), .Y(n_913) );
OA21x2_ASAP7_75t_L g914 ( .A1(n_743), .A2(n_753), .B(n_749), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_855), .A2(n_178), .B1(n_185), .B2(n_187), .Y(n_915) );
AOI22xp33_ASAP7_75t_SL g916 ( .A1(n_800), .A2(n_189), .B1(n_191), .B2(n_192), .Y(n_916) );
AND2x4_ASAP7_75t_L g917 ( .A(n_776), .B(n_194), .Y(n_917) );
OAI21x1_ASAP7_75t_L g918 ( .A1(n_760), .A2(n_201), .B(n_202), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_806), .B(n_204), .Y(n_919) );
OA21x2_ASAP7_75t_L g920 ( .A1(n_770), .A2(n_782), .B(n_780), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_778), .Y(n_921) );
OAI21x1_ASAP7_75t_L g922 ( .A1(n_764), .A2(n_205), .B(n_207), .Y(n_922) );
HB1xp67_ASAP7_75t_L g923 ( .A(n_794), .Y(n_923) );
INVx2_ASAP7_75t_L g924 ( .A(n_772), .Y(n_924) );
HB1xp67_ASAP7_75t_L g925 ( .A(n_794), .Y(n_925) );
AND2x2_ASAP7_75t_L g926 ( .A(n_792), .B(n_211), .Y(n_926) );
AOI21xp5_ASAP7_75t_L g927 ( .A1(n_830), .A2(n_212), .B(n_213), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_792), .B(n_214), .Y(n_928) );
AOI22xp33_ASAP7_75t_SL g929 ( .A1(n_800), .A2(n_215), .B1(n_218), .B2(n_220), .Y(n_929) );
AOI21xp5_ASAP7_75t_SL g930 ( .A1(n_759), .A2(n_775), .B(n_783), .Y(n_930) );
OA21x2_ASAP7_75t_L g931 ( .A1(n_754), .A2(n_224), .B(n_226), .Y(n_931) );
OR2x2_ASAP7_75t_L g932 ( .A(n_844), .B(n_227), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_779), .Y(n_933) );
AOI221xp5_ASAP7_75t_L g934 ( .A1(n_858), .A2(n_229), .B1(n_230), .B2(n_231), .C(n_232), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_784), .B(n_235), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_821), .A2(n_237), .B1(n_240), .B2(n_241), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_831), .A2(n_242), .B1(n_245), .B2(n_250), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_847), .B(n_258), .Y(n_938) );
AOI22xp33_ASAP7_75t_SL g939 ( .A1(n_841), .A2(n_261), .B1(n_263), .B2(n_265), .Y(n_939) );
NOR2xp33_ASAP7_75t_L g940 ( .A(n_785), .B(n_266), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_839), .A2(n_814), .B1(n_857), .B2(n_831), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_839), .A2(n_268), .B1(n_269), .B2(n_270), .Y(n_942) );
AOI221xp5_ASAP7_75t_L g943 ( .A1(n_813), .A2(n_271), .B1(n_273), .B2(n_274), .C(n_275), .Y(n_943) );
AOI221xp5_ASAP7_75t_L g944 ( .A1(n_813), .A2(n_276), .B1(n_277), .B2(n_278), .C(n_280), .Y(n_944) );
INVx2_ASAP7_75t_L g945 ( .A(n_773), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_850), .A2(n_281), .B1(n_282), .B2(n_283), .Y(n_946) );
A2O1A1Ixp33_ASAP7_75t_L g947 ( .A1(n_852), .A2(n_284), .B(n_287), .C(n_288), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_787), .Y(n_948) );
CKINVDCx11_ASAP7_75t_R g949 ( .A(n_752), .Y(n_949) );
INVxp67_ASAP7_75t_SL g950 ( .A(n_816), .Y(n_950) );
BUFx2_ASAP7_75t_L g951 ( .A(n_777), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_850), .A2(n_290), .B1(n_292), .B2(n_294), .Y(n_952) );
AOI22xp5_ASAP7_75t_L g953 ( .A1(n_793), .A2(n_776), .B1(n_788), .B2(n_789), .Y(n_953) );
OR2x6_ASAP7_75t_L g954 ( .A(n_747), .B(n_297), .Y(n_954) );
INVxp67_ASAP7_75t_L g955 ( .A(n_822), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_838), .A2(n_299), .B1(n_302), .B2(n_775), .Y(n_956) );
OAI21xp5_ASAP7_75t_L g957 ( .A1(n_758), .A2(n_852), .B(n_755), .Y(n_957) );
INVx4_ASAP7_75t_L g958 ( .A(n_752), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_791), .B(n_799), .Y(n_959) );
INVx2_ASAP7_75t_L g960 ( .A(n_781), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_859), .A2(n_796), .B1(n_861), .B2(n_797), .Y(n_961) );
AO21x1_ASAP7_75t_L g962 ( .A1(n_783), .A2(n_859), .B(n_765), .Y(n_962) );
BUFx2_ASAP7_75t_L g963 ( .A(n_756), .Y(n_963) );
INVx2_ASAP7_75t_L g964 ( .A(n_807), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_817), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_796), .A2(n_856), .B1(n_793), .B2(n_756), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_856), .A2(n_767), .B1(n_766), .B2(n_820), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_767), .A2(n_766), .B1(n_820), .B2(n_742), .Y(n_968) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_767), .Y(n_969) );
CKINVDCx6p67_ASAP7_75t_R g970 ( .A(n_803), .Y(n_970) );
AOI221xp5_ASAP7_75t_L g971 ( .A1(n_745), .A2(n_853), .B1(n_758), .B2(n_838), .C(n_824), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_836), .Y(n_972) );
OAI221xp5_ASAP7_75t_L g973 ( .A1(n_745), .A2(n_747), .B1(n_819), .B2(n_755), .C(n_834), .Y(n_973) );
OA21x2_ASAP7_75t_L g974 ( .A1(n_849), .A2(n_827), .B(n_818), .Y(n_974) );
INVx3_ASAP7_75t_L g975 ( .A(n_845), .Y(n_975) );
INVx2_ASAP7_75t_L g976 ( .A(n_823), .Y(n_976) );
OR2x2_ASAP7_75t_L g977 ( .A(n_742), .B(n_825), .Y(n_977) );
OAI22xp33_ASAP7_75t_L g978 ( .A1(n_845), .A2(n_863), .B1(n_860), .B2(n_865), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g979 ( .A1(n_860), .A2(n_863), .B1(n_865), .B2(n_842), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_751), .Y(n_980) );
OA21x2_ASAP7_75t_L g981 ( .A1(n_801), .A2(n_805), .B(n_815), .Y(n_981) );
OR2x2_ASAP7_75t_L g982 ( .A(n_864), .B(n_862), .Y(n_982) );
OAI22xp33_ASAP7_75t_L g983 ( .A1(n_808), .A2(n_804), .B1(n_846), .B2(n_751), .Y(n_983) );
OAI21xp5_ASAP7_75t_SL g984 ( .A1(n_808), .A2(n_804), .B(n_751), .Y(n_984) );
OAI221xp5_ASAP7_75t_L g985 ( .A1(n_751), .A2(n_568), .B1(n_695), .B2(n_566), .C(n_589), .Y(n_985) );
INVx2_ASAP7_75t_L g986 ( .A(n_761), .Y(n_986) );
CKINVDCx5p33_ASAP7_75t_R g987 ( .A(n_761), .Y(n_987) );
INVx2_ASAP7_75t_SL g988 ( .A(n_970), .Y(n_988) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_881), .Y(n_989) );
NOR2x1_ASAP7_75t_SL g990 ( .A(n_954), .B(n_912), .Y(n_990) );
INVx2_ASAP7_75t_L g991 ( .A(n_914), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_921), .Y(n_992) );
NOR2xp33_ASAP7_75t_L g993 ( .A(n_955), .B(n_958), .Y(n_993) );
HB1xp67_ASAP7_75t_L g994 ( .A(n_881), .Y(n_994) );
AND2x4_ASAP7_75t_L g995 ( .A(n_954), .B(n_874), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_933), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_948), .Y(n_997) );
INVx2_ASAP7_75t_L g998 ( .A(n_914), .Y(n_998) );
INVx2_ASAP7_75t_L g999 ( .A(n_986), .Y(n_999) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_894), .B(n_910), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_924), .B(n_945), .Y(n_1001) );
HB1xp67_ASAP7_75t_L g1002 ( .A(n_869), .Y(n_1002) );
BUFx2_ASAP7_75t_L g1003 ( .A(n_963), .Y(n_1003) );
INVx2_ASAP7_75t_L g1004 ( .A(n_888), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_959), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_965), .Y(n_1006) );
HB1xp67_ASAP7_75t_L g1007 ( .A(n_869), .Y(n_1007) );
BUFx2_ASAP7_75t_L g1008 ( .A(n_871), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_960), .Y(n_1009) );
INVx2_ASAP7_75t_L g1010 ( .A(n_920), .Y(n_1010) );
BUFx3_ASAP7_75t_L g1011 ( .A(n_874), .Y(n_1011) );
INVxp67_ASAP7_75t_SL g1012 ( .A(n_874), .Y(n_1012) );
BUFx2_ASAP7_75t_L g1013 ( .A(n_871), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_964), .B(n_972), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_980), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_886), .Y(n_1016) );
OR2x2_ASAP7_75t_L g1017 ( .A(n_886), .B(n_941), .Y(n_1017) );
AND2x4_ASAP7_75t_L g1018 ( .A(n_954), .B(n_975), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_935), .Y(n_1019) );
INVx2_ASAP7_75t_L g1020 ( .A(n_931), .Y(n_1020) );
BUFx2_ASAP7_75t_L g1021 ( .A(n_871), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_867), .B(n_893), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_976), .B(n_890), .Y(n_1023) );
HB1xp67_ASAP7_75t_L g1024 ( .A(n_969), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_935), .Y(n_1025) );
INVx2_ASAP7_75t_SL g1026 ( .A(n_877), .Y(n_1026) );
INVx2_ASAP7_75t_L g1027 ( .A(n_931), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_890), .B(n_961), .Y(n_1028) );
BUFx6f_ASAP7_75t_L g1029 ( .A(n_922), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_880), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_880), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_953), .B(n_975), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_982), .Y(n_1033) );
INVx2_ASAP7_75t_L g1034 ( .A(n_918), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_977), .B(n_906), .Y(n_1035) );
INVx2_ASAP7_75t_L g1036 ( .A(n_974), .Y(n_1036) );
NOR2x1_ASAP7_75t_L g1037 ( .A(n_958), .B(n_866), .Y(n_1037) );
BUFx2_ASAP7_75t_L g1038 ( .A(n_876), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_882), .B(n_919), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_985), .A2(n_868), .B1(n_892), .B2(n_967), .Y(n_1040) );
BUFx6f_ASAP7_75t_L g1041 ( .A(n_917), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_908), .B(n_966), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_896), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_911), .B(n_917), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_962), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_923), .B(n_925), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_940), .B(n_926), .Y(n_1047) );
INVx3_ASAP7_75t_L g1048 ( .A(n_872), .Y(n_1048) );
INVx2_ASAP7_75t_L g1049 ( .A(n_981), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_950), .B(n_878), .Y(n_1050) );
INVxp67_ASAP7_75t_SL g1051 ( .A(n_912), .Y(n_1051) );
INVxp67_ASAP7_75t_SL g1052 ( .A(n_876), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_928), .B(n_898), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_887), .B(n_891), .Y(n_1054) );
OAI22xp33_ASAP7_75t_L g1055 ( .A1(n_884), .A2(n_885), .B1(n_899), .B2(n_956), .Y(n_1055) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_932), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_938), .Y(n_1057) );
INVx2_ASAP7_75t_L g1058 ( .A(n_981), .Y(n_1058) );
INVx2_ASAP7_75t_L g1059 ( .A(n_987), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_903), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_879), .B(n_870), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_873), .B(n_957), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_957), .B(n_939), .Y(n_1063) );
INVx2_ASAP7_75t_L g1064 ( .A(n_973), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_968), .B(n_971), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_978), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_937), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_930), .B(n_929), .Y(n_1068) );
AO21x2_ASAP7_75t_L g1069 ( .A1(n_983), .A2(n_984), .B(n_979), .Y(n_1069) );
INVx2_ASAP7_75t_L g1070 ( .A(n_979), .Y(n_1070) );
NAND2x1p5_ASAP7_75t_L g1071 ( .A(n_904), .B(n_927), .Y(n_1071) );
INVx2_ASAP7_75t_L g1072 ( .A(n_937), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_934), .A2(n_956), .B1(n_943), .B2(n_944), .Y(n_1073) );
INVx2_ASAP7_75t_L g1074 ( .A(n_900), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_951), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_875), .B(n_907), .Y(n_1076) );
BUFx2_ASAP7_75t_L g1077 ( .A(n_947), .Y(n_1077) );
OAI22xp5_ASAP7_75t_L g1078 ( .A1(n_916), .A2(n_909), .B1(n_952), .B2(n_946), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_984), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_942), .B(n_902), .Y(n_1080) );
NAND3xp33_ASAP7_75t_SL g1081 ( .A(n_889), .B(n_915), .C(n_913), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_883), .Y(n_1082) );
OAI221xp5_ASAP7_75t_L g1083 ( .A1(n_936), .A2(n_901), .B1(n_895), .B2(n_897), .C(n_905), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_949), .Y(n_1084) );
INVx2_ASAP7_75t_L g1085 ( .A(n_914), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_894), .B(n_910), .Y(n_1086) );
NOR2xp33_ASAP7_75t_L g1087 ( .A(n_955), .B(n_702), .Y(n_1087) );
AND2x4_ASAP7_75t_L g1088 ( .A(n_954), .B(n_874), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_894), .B(n_910), .Y(n_1089) );
INVx2_ASAP7_75t_L g1090 ( .A(n_914), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_921), .Y(n_1091) );
AND2x4_ASAP7_75t_L g1092 ( .A(n_954), .B(n_874), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_921), .B(n_762), .Y(n_1093) );
OR2x2_ASAP7_75t_L g1094 ( .A(n_963), .B(n_769), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_992), .Y(n_1095) );
AO21x2_ASAP7_75t_L g1096 ( .A1(n_1020), .A2(n_1027), .B(n_1034), .Y(n_1096) );
HB1xp67_ASAP7_75t_L g1097 ( .A(n_1033), .Y(n_1097) );
NAND3xp33_ASAP7_75t_L g1098 ( .A(n_1059), .B(n_989), .C(n_994), .Y(n_1098) );
OAI22xp5_ASAP7_75t_SL g1099 ( .A1(n_1002), .A2(n_1007), .B1(n_1037), .B2(n_1084), .Y(n_1099) );
AOI21xp5_ASAP7_75t_L g1100 ( .A1(n_990), .A2(n_1072), .B(n_1067), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1014), .B(n_1000), .Y(n_1101) );
AND2x4_ASAP7_75t_L g1102 ( .A(n_1032), .B(n_1033), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_992), .Y(n_1103) );
BUFx2_ASAP7_75t_L g1104 ( .A(n_988), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1014), .B(n_1000), .Y(n_1105) );
OR2x2_ASAP7_75t_L g1106 ( .A(n_1003), .B(n_1094), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_1005), .B(n_1030), .Y(n_1107) );
INVx4_ASAP7_75t_L g1108 ( .A(n_1041), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1086), .B(n_1089), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1086), .B(n_1089), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_996), .Y(n_1111) );
BUFx2_ASAP7_75t_L g1112 ( .A(n_988), .Y(n_1112) );
NOR2xp33_ASAP7_75t_R g1113 ( .A(n_1041), .B(n_1081), .Y(n_1113) );
INVx2_ASAP7_75t_L g1114 ( .A(n_1036), .Y(n_1114) );
BUFx2_ASAP7_75t_L g1115 ( .A(n_1003), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1046), .B(n_1001), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_1046), .B(n_1001), .Y(n_1117) );
OR2x2_ASAP7_75t_L g1118 ( .A(n_1094), .B(n_1004), .Y(n_1118) );
NAND3xp33_ASAP7_75t_L g1119 ( .A(n_1059), .B(n_1045), .C(n_1056), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_996), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_997), .Y(n_1121) );
INVx2_ASAP7_75t_SL g1122 ( .A(n_995), .Y(n_1122) );
AND2x4_ASAP7_75t_L g1123 ( .A(n_1032), .B(n_1062), .Y(n_1123) );
OR2x2_ASAP7_75t_L g1124 ( .A(n_1004), .B(n_1024), .Y(n_1124) );
OAI221xp5_ASAP7_75t_SL g1125 ( .A1(n_1040), .A2(n_1055), .B1(n_1017), .B2(n_1022), .C(n_1039), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1043), .B(n_1035), .Y(n_1126) );
BUFx3_ASAP7_75t_L g1127 ( .A(n_1011), .Y(n_1127) );
OR2x2_ASAP7_75t_L g1128 ( .A(n_1005), .B(n_1030), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1031), .B(n_997), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1035), .B(n_1026), .Y(n_1130) );
OR2x2_ASAP7_75t_L g1131 ( .A(n_1031), .B(n_1006), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1091), .Y(n_1132) );
OR2x2_ASAP7_75t_L g1133 ( .A(n_1006), .B(n_1091), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1093), .Y(n_1134) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1009), .Y(n_1135) );
OR2x2_ASAP7_75t_L g1136 ( .A(n_1009), .B(n_1017), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_1016), .B(n_1039), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1026), .Y(n_1138) );
NAND3xp33_ASAP7_75t_L g1139 ( .A(n_1045), .B(n_1075), .C(n_1065), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1050), .B(n_1044), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1015), .Y(n_1141) );
HB1xp67_ASAP7_75t_L g1142 ( .A(n_999), .Y(n_1142) );
INVxp67_ASAP7_75t_L g1143 ( .A(n_990), .Y(n_1143) );
OAI22xp33_ASAP7_75t_L g1144 ( .A1(n_1051), .A2(n_1038), .B1(n_1041), .B2(n_1072), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_1028), .A2(n_1054), .B1(n_1042), .B2(n_1076), .Y(n_1145) );
OAI21xp5_ASAP7_75t_L g1146 ( .A1(n_1054), .A2(n_1074), .B(n_1016), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1015), .Y(n_1147) );
NOR2x1_ASAP7_75t_L g1148 ( .A(n_1018), .B(n_995), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1023), .Y(n_1149) );
HB1xp67_ASAP7_75t_L g1150 ( .A(n_991), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1044), .B(n_1057), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1023), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_1028), .A2(n_1042), .B1(n_1067), .B2(n_1053), .Y(n_1153) );
INVxp67_ASAP7_75t_SL g1154 ( .A(n_1041), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1008), .B(n_1013), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1008), .B(n_1013), .Y(n_1156) );
BUFx3_ASAP7_75t_L g1157 ( .A(n_1011), .Y(n_1157) );
OAI22xp5_ASAP7_75t_L g1158 ( .A1(n_1038), .A2(n_1041), .B1(n_1047), .B2(n_1073), .Y(n_1158) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1049), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1021), .Y(n_1160) );
INVx3_ASAP7_75t_L g1161 ( .A(n_1018), .Y(n_1161) );
AOI21x1_ASAP7_75t_L g1162 ( .A1(n_1020), .A2(n_1027), .B(n_1077), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1021), .B(n_1061), .Y(n_1163) );
INVxp67_ASAP7_75t_SL g1164 ( .A(n_991), .Y(n_1164) );
AOI221xp5_ASAP7_75t_L g1165 ( .A1(n_1079), .A2(n_1087), .B1(n_1066), .B2(n_1061), .C(n_1053), .Y(n_1165) );
NAND2xp5_ASAP7_75t_L g1166 ( .A(n_1047), .B(n_1018), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1079), .Y(n_1167) );
AOI22xp5_ASAP7_75t_L g1168 ( .A1(n_1080), .A2(n_1060), .B1(n_993), .B2(n_1074), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1084), .B(n_995), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1088), .B(n_1092), .Y(n_1170) );
HB1xp67_ASAP7_75t_L g1171 ( .A(n_998), .Y(n_1171) );
INVxp67_ASAP7_75t_SL g1172 ( .A(n_998), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1088), .Y(n_1173) );
OR2x2_ASAP7_75t_L g1174 ( .A(n_1088), .B(n_1092), .Y(n_1174) );
HB1xp67_ASAP7_75t_L g1175 ( .A(n_1085), .Y(n_1175) );
AND2x4_ASAP7_75t_L g1176 ( .A(n_1062), .B(n_1092), .Y(n_1176) );
HB1xp67_ASAP7_75t_L g1177 ( .A(n_1085), .Y(n_1177) );
BUFx2_ASAP7_75t_L g1178 ( .A(n_1012), .Y(n_1178) );
OAI221xp5_ASAP7_75t_L g1179 ( .A1(n_1077), .A2(n_1078), .B1(n_1019), .B2(n_1025), .C(n_1068), .Y(n_1179) );
INVx5_ASAP7_75t_L g1180 ( .A(n_1048), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1181 ( .A(n_1019), .B(n_1025), .Y(n_1181) );
INVx1_ASAP7_75t_SL g1182 ( .A(n_1048), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1149), .B(n_1066), .Y(n_1183) );
INVx2_ASAP7_75t_L g1184 ( .A(n_1114), .Y(n_1184) );
OR2x2_ASAP7_75t_L g1185 ( .A(n_1152), .B(n_1052), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1123), .B(n_1069), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1187 ( .A(n_1101), .B(n_1068), .Y(n_1187) );
HB1xp67_ASAP7_75t_L g1188 ( .A(n_1115), .Y(n_1188) );
HB1xp67_ASAP7_75t_L g1189 ( .A(n_1124), .Y(n_1189) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_1105), .B(n_1063), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1109), .B(n_1063), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1141), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1123), .B(n_1069), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1110), .B(n_1064), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1147), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_1126), .B(n_1064), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1145), .B(n_1080), .Y(n_1197) );
OR2x2_ASAP7_75t_L g1198 ( .A(n_1123), .B(n_1069), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1102), .B(n_1070), .Y(n_1199) );
AND2x2_ASAP7_75t_SL g1200 ( .A(n_1176), .B(n_1070), .Y(n_1200) );
HB1xp67_ASAP7_75t_L g1201 ( .A(n_1178), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1102), .B(n_1010), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1095), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1102), .B(n_1010), .Y(n_1204) );
AOI222xp33_ASAP7_75t_L g1205 ( .A1(n_1165), .A2(n_1145), .B1(n_1146), .B2(n_1153), .C1(n_1179), .C2(n_1099), .Y(n_1205) );
AOI221x1_ASAP7_75t_L g1206 ( .A1(n_1139), .A2(n_1119), .B1(n_1098), .B2(n_1138), .C(n_1100), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1103), .Y(n_1207) );
OR2x2_ASAP7_75t_L g1208 ( .A(n_1097), .B(n_1058), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1111), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1120), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1116), .B(n_1048), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1142), .B(n_1167), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1121), .Y(n_1213) );
NOR2x1_ASAP7_75t_L g1214 ( .A(n_1127), .B(n_1082), .Y(n_1214) );
AND2x4_ASAP7_75t_L g1215 ( .A(n_1143), .B(n_1090), .Y(n_1215) );
INVx3_ASAP7_75t_L g1216 ( .A(n_1180), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1176), .B(n_1082), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1132), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1176), .B(n_1034), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1117), .B(n_1071), .Y(n_1220) );
OR2x2_ASAP7_75t_L g1221 ( .A(n_1097), .B(n_1071), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1134), .B(n_1071), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1151), .B(n_1029), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1163), .B(n_1029), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1150), .B(n_1029), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_1137), .B(n_1029), .Y(n_1226) );
NAND4xp25_ASAP7_75t_L g1227 ( .A(n_1125), .B(n_1029), .C(n_1083), .D(n_1153), .Y(n_1227) );
HB1xp67_ASAP7_75t_L g1228 ( .A(n_1106), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1150), .B(n_1171), .Y(n_1229) );
HB1xp67_ASAP7_75t_L g1230 ( .A(n_1130), .Y(n_1230) );
NAND5xp2_ASAP7_75t_L g1231 ( .A(n_1168), .B(n_1143), .C(n_1169), .D(n_1170), .E(n_1166), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1171), .B(n_1175), .Y(n_1232) );
OR2x2_ASAP7_75t_L g1233 ( .A(n_1136), .B(n_1118), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1175), .B(n_1177), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1133), .B(n_1131), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1177), .B(n_1159), .Y(n_1236) );
OAI211xp5_ASAP7_75t_L g1237 ( .A1(n_1113), .A2(n_1104), .B(n_1112), .C(n_1148), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1135), .Y(n_1238) );
OR2x2_ASAP7_75t_L g1239 ( .A(n_1128), .B(n_1181), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1107), .B(n_1140), .Y(n_1240) );
NOR2xp33_ASAP7_75t_L g1241 ( .A(n_1161), .B(n_1129), .Y(n_1241) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_1189), .B(n_1160), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1192), .Y(n_1243) );
AOI21xp33_ASAP7_75t_SL g1244 ( .A1(n_1205), .A2(n_1158), .B(n_1144), .Y(n_1244) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1192), .Y(n_1245) );
INVx2_ASAP7_75t_L g1246 ( .A(n_1236), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1195), .Y(n_1247) );
CKINVDCx20_ASAP7_75t_R g1248 ( .A(n_1230), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1186), .B(n_1164), .Y(n_1249) );
NOR2x1_ASAP7_75t_L g1250 ( .A(n_1237), .B(n_1157), .Y(n_1250) );
OR2x2_ASAP7_75t_L g1251 ( .A(n_1228), .B(n_1172), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1195), .Y(n_1252) );
OR2x2_ASAP7_75t_L g1253 ( .A(n_1233), .B(n_1172), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1203), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1186), .B(n_1164), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1203), .Y(n_1256) );
OR2x2_ASAP7_75t_L g1257 ( .A(n_1233), .B(n_1235), .Y(n_1257) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1207), .Y(n_1258) );
INVxp67_ASAP7_75t_L g1259 ( .A(n_1201), .Y(n_1259) );
NOR3xp33_ASAP7_75t_L g1260 ( .A(n_1227), .B(n_1161), .C(n_1182), .Y(n_1260) );
OAI21xp33_ASAP7_75t_L g1261 ( .A1(n_1193), .A2(n_1113), .B(n_1173), .Y(n_1261) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1207), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1209), .Y(n_1263) );
AO21x2_ASAP7_75t_L g1264 ( .A1(n_1222), .A2(n_1162), .B(n_1144), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1197), .B(n_1155), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1193), .B(n_1154), .Y(n_1266) );
INVxp67_ASAP7_75t_L g1267 ( .A(n_1188), .Y(n_1267) );
OR2x2_ASAP7_75t_L g1268 ( .A(n_1235), .B(n_1174), .Y(n_1268) );
INVx2_ASAP7_75t_L g1269 ( .A(n_1236), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1199), .B(n_1217), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1194), .B(n_1156), .Y(n_1271) );
NAND2xp5_ASAP7_75t_L g1272 ( .A(n_1183), .B(n_1122), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1199), .B(n_1154), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1217), .B(n_1096), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1223), .B(n_1096), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1223), .B(n_1122), .Y(n_1276) );
INVx2_ASAP7_75t_L g1277 ( .A(n_1184), .Y(n_1277) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_1231), .A2(n_1127), .B1(n_1157), .B2(n_1108), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1202), .B(n_1108), .Y(n_1279) );
BUFx2_ASAP7_75t_L g1280 ( .A(n_1229), .Y(n_1280) );
NOR2xp33_ASAP7_75t_L g1281 ( .A(n_1240), .B(n_1180), .Y(n_1281) );
NAND2xp5_ASAP7_75t_L g1282 ( .A(n_1183), .B(n_1180), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1202), .B(n_1108), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1204), .B(n_1180), .Y(n_1284) );
BUFx2_ASAP7_75t_SL g1285 ( .A(n_1216), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1196), .B(n_1190), .Y(n_1286) );
INVx2_ASAP7_75t_SL g1287 ( .A(n_1229), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1204), .B(n_1224), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1224), .B(n_1219), .Y(n_1289) );
INVx2_ASAP7_75t_L g1290 ( .A(n_1251), .Y(n_1290) );
OAI21xp33_ASAP7_75t_SL g1291 ( .A1(n_1250), .A2(n_1200), .B(n_1216), .Y(n_1291) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_1286), .B(n_1191), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1257), .Y(n_1293) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1257), .Y(n_1294) );
AOI22xp5_ASAP7_75t_L g1295 ( .A1(n_1248), .A2(n_1220), .B1(n_1241), .B2(n_1200), .Y(n_1295) );
HB1xp67_ASAP7_75t_L g1296 ( .A(n_1280), .Y(n_1296) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1245), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1245), .Y(n_1298) );
BUFx3_ASAP7_75t_L g1299 ( .A(n_1248), .Y(n_1299) );
AOI31xp33_ASAP7_75t_L g1300 ( .A1(n_1244), .A2(n_1239), .A3(n_1211), .B(n_1198), .Y(n_1300) );
AOI221xp5_ASAP7_75t_L g1301 ( .A1(n_1259), .A2(n_1187), .B1(n_1218), .B2(n_1210), .C(n_1213), .Y(n_1301) );
O2A1O1Ixp5_ASAP7_75t_L g1302 ( .A1(n_1281), .A2(n_1216), .B(n_1238), .C(n_1218), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1247), .Y(n_1303) );
INVx1_ASAP7_75t_SL g1304 ( .A(n_1253), .Y(n_1304) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1247), .Y(n_1305) );
OR2x2_ASAP7_75t_L g1306 ( .A(n_1253), .B(n_1239), .Y(n_1306) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_1265), .B(n_1212), .Y(n_1307) );
AOI22xp5_ASAP7_75t_L g1308 ( .A1(n_1260), .A2(n_1220), .B1(n_1200), .B2(n_1219), .Y(n_1308) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1254), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1280), .B(n_1212), .Y(n_1310) );
INVxp67_ASAP7_75t_L g1311 ( .A(n_1251), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1312 ( .A(n_1267), .B(n_1185), .Y(n_1312) );
AOI322xp5_ASAP7_75t_L g1313 ( .A1(n_1270), .A2(n_1209), .A3(n_1210), .B1(n_1213), .B2(n_1238), .C1(n_1232), .C2(n_1234), .Y(n_1313) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1254), .Y(n_1314) );
NAND2xp5_ASAP7_75t_SL g1315 ( .A(n_1278), .B(n_1215), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1268), .Y(n_1316) );
AOI221xp5_ASAP7_75t_L g1317 ( .A1(n_1271), .A2(n_1198), .B1(n_1185), .B2(n_1232), .C(n_1234), .Y(n_1317) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1268), .Y(n_1318) );
INVxp67_ASAP7_75t_L g1319 ( .A(n_1285), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1242), .Y(n_1320) );
INVx2_ASAP7_75t_L g1321 ( .A(n_1296), .Y(n_1321) );
A2O1A1Ixp33_ASAP7_75t_L g1322 ( .A1(n_1291), .A2(n_1261), .B(n_1285), .C(n_1287), .Y(n_1322) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1306), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g1324 ( .A(n_1313), .B(n_1274), .Y(n_1324) );
NAND2x1_ASAP7_75t_L g1325 ( .A(n_1300), .B(n_1214), .Y(n_1325) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1311), .Y(n_1326) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_1317), .B(n_1274), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1297), .Y(n_1328) );
A2O1A1Ixp33_ASAP7_75t_L g1329 ( .A1(n_1302), .A2(n_1287), .B(n_1270), .C(n_1282), .Y(n_1329) );
AOI222xp33_ASAP7_75t_L g1330 ( .A1(n_1299), .A2(n_1243), .B1(n_1252), .B2(n_1256), .C1(n_1258), .C2(n_1262), .Y(n_1330) );
OAI32xp33_ASAP7_75t_L g1331 ( .A1(n_1296), .A2(n_1242), .A3(n_1221), .B1(n_1272), .B2(n_1246), .Y(n_1331) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1298), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1301), .B(n_1275), .Y(n_1333) );
OAI21xp33_ASAP7_75t_L g1334 ( .A1(n_1308), .A2(n_1289), .B(n_1288), .Y(n_1334) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1293), .B(n_1263), .Y(n_1335) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1303), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1337 ( .A(n_1294), .B(n_1275), .Y(n_1337) );
XNOR2xp5_ASAP7_75t_L g1338 ( .A(n_1295), .B(n_1288), .Y(n_1338) );
OR2x2_ASAP7_75t_L g1339 ( .A(n_1304), .B(n_1246), .Y(n_1339) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1305), .Y(n_1340) );
OAI21xp33_ASAP7_75t_L g1341 ( .A1(n_1334), .A2(n_1312), .B(n_1310), .Y(n_1341) );
NAND2xp5_ASAP7_75t_SL g1342 ( .A(n_1322), .B(n_1302), .Y(n_1342) );
OAI21xp33_ASAP7_75t_L g1343 ( .A1(n_1324), .A2(n_1320), .B(n_1292), .Y(n_1343) );
OAI221xp5_ASAP7_75t_SL g1344 ( .A1(n_1329), .A2(n_1319), .B1(n_1318), .B2(n_1316), .C(n_1307), .Y(n_1344) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1335), .Y(n_1345) );
INVx2_ASAP7_75t_L g1346 ( .A(n_1321), .Y(n_1346) );
OAI322xp33_ASAP7_75t_L g1347 ( .A1(n_1327), .A2(n_1319), .A3(n_1315), .B1(n_1290), .B2(n_1309), .C1(n_1314), .C2(n_1221), .Y(n_1347) );
BUFx6f_ASAP7_75t_L g1348 ( .A(n_1325), .Y(n_1348) );
AOI21xp5_ASAP7_75t_L g1349 ( .A1(n_1331), .A2(n_1206), .B(n_1283), .Y(n_1349) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1335), .Y(n_1350) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1326), .Y(n_1351) );
AOI21xp33_ASAP7_75t_SL g1352 ( .A1(n_1330), .A2(n_1284), .B(n_1264), .Y(n_1352) );
OAI21xp33_ASAP7_75t_L g1353 ( .A1(n_1333), .A2(n_1276), .B(n_1266), .Y(n_1353) );
INVx1_ASAP7_75t_SL g1354 ( .A(n_1348), .Y(n_1354) );
NAND2xp5_ASAP7_75t_L g1355 ( .A(n_1345), .B(n_1330), .Y(n_1355) );
OAI211xp5_ASAP7_75t_SL g1356 ( .A1(n_1342), .A2(n_1323), .B(n_1337), .C(n_1328), .Y(n_1356) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1350), .Y(n_1357) );
A2O1A1Ixp33_ASAP7_75t_L g1358 ( .A1(n_1344), .A2(n_1284), .B(n_1339), .C(n_1279), .Y(n_1358) );
OAI321xp33_ASAP7_75t_L g1359 ( .A1(n_1343), .A2(n_1336), .A3(n_1332), .B1(n_1340), .B2(n_1283), .C(n_1279), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1341), .B(n_1338), .Y(n_1360) );
NAND3xp33_ASAP7_75t_SL g1361 ( .A(n_1352), .B(n_1249), .C(n_1255), .Y(n_1361) );
OAI22xp5_ASAP7_75t_L g1362 ( .A1(n_1360), .A2(n_1348), .B1(n_1353), .B2(n_1349), .Y(n_1362) );
AND2x4_ASAP7_75t_L g1363 ( .A(n_1354), .B(n_1351), .Y(n_1363) );
NOR4xp75_ASAP7_75t_L g1364 ( .A(n_1361), .B(n_1347), .C(n_1348), .D(n_1276), .Y(n_1364) );
NAND4xp25_ASAP7_75t_L g1365 ( .A(n_1358), .B(n_1206), .C(n_1214), .D(n_1346), .Y(n_1365) );
NAND2xp5_ASAP7_75t_L g1366 ( .A(n_1355), .B(n_1289), .Y(n_1366) );
OAI22xp5_ASAP7_75t_L g1367 ( .A1(n_1358), .A2(n_1269), .B1(n_1266), .B2(n_1249), .Y(n_1367) );
NOR3xp33_ASAP7_75t_L g1368 ( .A(n_1362), .B(n_1356), .C(n_1359), .Y(n_1368) );
INVxp67_ASAP7_75t_L g1369 ( .A(n_1363), .Y(n_1369) );
OR4x2_ASAP7_75t_L g1370 ( .A(n_1364), .B(n_1357), .C(n_1255), .D(n_1273), .Y(n_1370) );
NOR3xp33_ASAP7_75t_L g1371 ( .A(n_1365), .B(n_1226), .C(n_1277), .Y(n_1371) );
XOR2x2_ASAP7_75t_L g1372 ( .A(n_1368), .B(n_1366), .Y(n_1372) );
NOR2xp67_ASAP7_75t_L g1373 ( .A(n_1369), .B(n_1367), .Y(n_1373) );
INVx1_ASAP7_75t_SL g1374 ( .A(n_1370), .Y(n_1374) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1373), .Y(n_1375) );
NAND2xp5_ASAP7_75t_L g1376 ( .A(n_1372), .B(n_1371), .Y(n_1376) );
OAI21xp5_ASAP7_75t_L g1377 ( .A1(n_1375), .A2(n_1374), .B(n_1273), .Y(n_1377) );
OAI22xp5_ASAP7_75t_SL g1378 ( .A1(n_1376), .A2(n_1269), .B1(n_1215), .B2(n_1208), .Y(n_1378) );
OR2x2_ASAP7_75t_L g1379 ( .A(n_1377), .B(n_1264), .Y(n_1379) );
AOI21xp33_ASAP7_75t_SL g1380 ( .A1(n_1378), .A2(n_1264), .B(n_1208), .Y(n_1380) );
HB1xp67_ASAP7_75t_L g1381 ( .A(n_1379), .Y(n_1381) );
AOI21xp33_ASAP7_75t_L g1382 ( .A1(n_1381), .A2(n_1380), .B(n_1225), .Y(n_1382) );
endmodule