module fake_jpeg_18780_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_5),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_29),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_23),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_21),
.B(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_68),
.Y(n_74)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_60),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_62),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_79),
.Y(n_95)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_60),
.B1(n_48),
.B2(n_56),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_61),
.B1(n_49),
.B2(n_43),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_54),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_80),
.A2(n_57),
.B1(n_58),
.B2(n_52),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_91),
.B1(n_93),
.B2(n_74),
.Y(n_98)
);

OA21x2_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_51),
.B(n_59),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_104)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_92),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_9),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_63),
.B1(n_44),
.B2(n_45),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_65),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_103),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_55),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_102),
.C(n_107),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_64),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_0),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_105),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_22),
.B1(n_38),
.B2(n_37),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_2),
.Y(n_106)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

AND2x4_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_3),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g110 ( 
.A(n_108),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_117),
.Y(n_118)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_121),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_112),
.A2(n_104),
.B1(n_107),
.B2(n_13),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_113),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_11),
.C(n_12),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_122),
.B(n_111),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_124),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_118),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_110),
.A3(n_118),
.B1(n_123),
.B2(n_114),
.C1(n_32),
.C2(n_34),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_110),
.C(n_24),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_14),
.C(n_28),
.Y(n_130)
);

AO21x1_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_30),
.B(n_35),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_36),
.Y(n_132)
);


endmodule