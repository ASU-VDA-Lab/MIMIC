module fake_jpeg_18729_n_109 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_109);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_109;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_23),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_25),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx4f_ASAP7_75t_SL g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_54),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_0),
.Y(n_60)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_49),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_51),
.A2(n_48),
.B1(n_47),
.B2(n_45),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_39),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_1),
.B(n_2),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_36),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_80),
.B1(n_82),
.B2(n_66),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_44),
.B1(n_42),
.B2(n_38),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_74),
.B1(n_78),
.B2(n_81),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_37),
.B1(n_19),
.B2(n_21),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_18),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_2),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_77),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_6),
.B1(n_12),
.B2(n_13),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_27),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_91),
.C(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_86),
.Y(n_97)
);

AOI221xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_99),
.B1(n_94),
.B2(n_93),
.C(n_85),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_95),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

AOI221xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_86),
.B1(n_87),
.B2(n_84),
.C(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_101),
.C(n_96),
.Y(n_106)
);

NOR4xp25_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_70),
.C(n_29),
.D(n_30),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_SL g108 ( 
.A1(n_107),
.A2(n_28),
.B(n_31),
.C(n_32),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_34),
.Y(n_109)
);


endmodule