module fake_jpeg_4069_n_141 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_30),
.Y(n_43)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_35),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_23),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_34),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_37),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_49),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_28),
.B1(n_22),
.B2(n_25),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_50),
.B1(n_20),
.B2(n_18),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_28),
.B(n_15),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_21),
.C(n_15),
.Y(n_64)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_25),
.B1(n_20),
.B2(n_21),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_53),
.B(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_24),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_13),
.Y(n_59)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_13),
.Y(n_60)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_18),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_66),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_71),
.B1(n_72),
.B2(n_27),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_32),
.B1(n_17),
.B2(n_14),
.Y(n_81)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_68),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_70),
.Y(n_85)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_38),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_32),
.C(n_31),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_52),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_76),
.B(n_63),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_71),
.B1(n_57),
.B2(n_51),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_30),
.B1(n_17),
.B2(n_14),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_70),
.B1(n_66),
.B2(n_6),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_95),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_86),
.B(n_1),
.Y(n_93)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_78),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_74),
.A2(n_1),
.B(n_5),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_101),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_100),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_79),
.B(n_6),
.Y(n_102)
);

XOR2x2_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_80),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_82),
.Y(n_117)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_82),
.B(n_97),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_118),
.C(n_120),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_83),
.B(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_104),
.A2(n_81),
.B1(n_95),
.B2(n_84),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_119),
.A2(n_103),
.B1(n_109),
.B2(n_111),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_111),
.B(n_91),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_119),
.B1(n_101),
.B2(n_99),
.Y(n_130)
);

NOR2xp67_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_120),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_127),
.A2(n_130),
.B(n_106),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_107),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_129),
.C(n_131),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_121),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_73),
.C(n_75),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_127),
.A2(n_125),
.B1(n_122),
.B2(n_108),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_133),
.C(n_134),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_77),
.B(n_106),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_135),
.B(n_77),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_137),
.B(n_87),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_136),
.B(n_11),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_8),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_12),
.Y(n_141)
);


endmodule