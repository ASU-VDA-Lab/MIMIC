module fake_netlist_5_512_n_5399 (n_924, n_1263, n_977, n_611, n_1126, n_1166, n_469, n_82, n_785, n_549, n_532, n_1161, n_1150, n_226, n_667, n_790, n_1055, n_111, n_880, n_544, n_1007, n_155, n_552, n_1198, n_1099, n_956, n_564, n_423, n_21, n_105, n_1021, n_4, n_551, n_688, n_800, n_671, n_819, n_1022, n_915, n_864, n_173, n_859, n_951, n_1264, n_447, n_247, n_292, n_625, n_854, n_674, n_417, n_516, n_933, n_1152, n_497, n_606, n_275, n_26, n_877, n_2, n_755, n_1118, n_6, n_947, n_1285, n_373, n_307, n_530, n_87, n_150, n_1107, n_556, n_1230, n_668, n_375, n_301, n_929, n_1124, n_902, n_191, n_1104, n_659, n_51, n_1257, n_171, n_1182, n_579, n_1261, n_938, n_1098, n_320, n_1154, n_1242, n_1135, n_24, n_406, n_519, n_1016, n_1243, n_546, n_101, n_1280, n_281, n_240, n_291, n_231, n_257, n_731, n_371, n_709, n_317, n_1236, n_569, n_227, n_920, n_1289, n_94, n_335, n_370, n_976, n_343, n_308, n_297, n_156, n_1078, n_775, n_219, n_157, n_600, n_223, n_264, n_955, n_163, n_339, n_1146, n_882, n_183, n_243, n_1036, n_1097, n_347, n_59, n_550, n_696, n_897, n_215, n_350, n_196, n_798, n_646, n_436, n_1216, n_290, n_580, n_1040, n_578, n_926, n_344, n_1218, n_422, n_475, n_777, n_1070, n_1030, n_72, n_415, n_1071, n_485, n_1165, n_1267, n_496, n_958, n_1034, n_670, n_48, n_521, n_663, n_845, n_673, n_837, n_1239, n_528, n_680, n_395, n_164, n_553, n_901, n_813, n_1284, n_214, n_675, n_888, n_1167, n_637, n_184, n_446, n_1064, n_144, n_858, n_114, n_96, n_923, n_691, n_1151, n_881, n_468, n_213, n_129, n_342, n_464, n_363, n_197, n_1069, n_1075, n_460, n_889, n_973, n_477, n_571, n_461, n_1211, n_1197, n_907, n_190, n_989, n_1039, n_34, n_228, n_283, n_488, n_736, n_892, n_1000, n_1202, n_1278, n_1002, n_49, n_310, n_54, n_593, n_12, n_748, n_586, n_1058, n_838, n_332, n_1053, n_1224, n_349, n_1248, n_230, n_953, n_279, n_1014, n_1241, n_70, n_289, n_963, n_1052, n_954, n_627, n_440, n_793, n_478, n_476, n_534, n_884, n_345, n_944, n_91, n_182, n_143, n_647, n_237, n_407, n_1072, n_832, n_857, n_207, n_561, n_18, n_1027, n_971, n_1156, n_117, n_326, n_794, n_404, n_686, n_847, n_596, n_558, n_702, n_1276, n_822, n_728, n_266, n_1162, n_272, n_1199, n_352, n_53, n_1038, n_520, n_409, n_887, n_154, n_71, n_300, n_809, n_870, n_931, n_599, n_434, n_868, n_639, n_914, n_411, n_414, n_965, n_935, n_121, n_1175, n_817, n_360, n_36, n_64, n_759, n_28, n_806, n_324, n_187, n_1189, n_103, n_97, n_11, n_7, n_1259, n_706, n_746, n_747, n_52, n_784, n_110, n_1244, n_431, n_1194, n_615, n_851, n_843, n_523, n_913, n_705, n_865, n_61, n_678, n_697, n_127, n_1222, n_75, n_776, n_367, n_452, n_525, n_1260, n_649, n_547, n_43, n_1191, n_116, n_284, n_1128, n_139, n_744, n_590, n_629, n_254, n_1233, n_23, n_526, n_293, n_372, n_677, n_244, n_47, n_1121, n_314, n_368, n_433, n_604, n_8, n_949, n_100, n_1008, n_946, n_1001, n_498, n_689, n_738, n_640, n_252, n_624, n_295, n_133, n_1010, n_1231, n_739, n_1279, n_1195, n_610, n_936, n_568, n_39, n_1090, n_757, n_633, n_439, n_106, n_259, n_448, n_758, n_999, n_93, n_1158, n_563, n_1145, n_878, n_524, n_204, n_394, n_1049, n_1153, n_741, n_1068, n_122, n_331, n_10, n_906, n_1163, n_1207, n_919, n_908, n_90, n_724, n_658, n_456, n_959, n_535, n_152, n_940, n_9, n_592, n_1169, n_45, n_1017, n_123, n_978, n_1054, n_1269, n_1095, n_267, n_514, n_457, n_1079, n_1045, n_1208, n_603, n_484, n_1033, n_442, n_131, n_636, n_660, n_1009, n_1148, n_109, n_742, n_750, n_995, n_454, n_374, n_185, n_396, n_1073, n_255, n_662, n_459, n_218, n_962, n_1215, n_1171, n_723, n_1065, n_473, n_1043, n_355, n_486, n_614, n_337, n_88, n_1286, n_1177, n_168, n_974, n_727, n_1159, n_957, n_773, n_208, n_142, n_743, n_299, n_303, n_296, n_613, n_1119, n_1240, n_65, n_829, n_361, n_700, n_1237, n_573, n_69, n_1132, n_388, n_1127, n_761, n_1006, n_329, n_274, n_1270, n_582, n_73, n_19, n_309, n_30, n_512, n_84, n_130, n_322, n_1249, n_652, n_1111, n_25, n_1093, n_288, n_1031, n_263, n_609, n_1041, n_1265, n_44, n_224, n_383, n_834, n_112, n_765, n_893, n_1015, n_1140, n_891, n_239, n_630, n_55, n_504, n_511, n_874, n_358, n_1101, n_77, n_102, n_1106, n_987, n_261, n_174, n_767, n_993, n_545, n_441, n_860, n_450, n_429, n_948, n_1217, n_628, n_365, n_729, n_1131, n_1084, n_970, n_911, n_83, n_513, n_1094, n_560, n_340, n_1044, n_1205, n_346, n_1209, n_495, n_602, n_574, n_879, n_16, n_58, n_623, n_405, n_824, n_359, n_490, n_996, n_921, n_233, n_572, n_366, n_815, n_128, n_120, n_327, n_135, n_1037, n_1080, n_1274, n_426, n_1082, n_589, n_716, n_562, n_62, n_952, n_1229, n_391, n_701, n_1023, n_645, n_539, n_803, n_1092, n_238, n_531, n_890, n_764, n_1056, n_162, n_960, n_222, n_1290, n_1123, n_1047, n_634, n_199, n_32, n_1252, n_348, n_1029, n_925, n_1206, n_424, n_256, n_950, n_380, n_419, n_444, n_1060, n_1141, n_316, n_389, n_418, n_248, n_136, n_86, n_146, n_912, n_315, n_968, n_451, n_619, n_408, n_376, n_967, n_74, n_1139, n_515, n_57, n_351, n_885, n_397, n_483, n_683, n_1057, n_1051, n_1085, n_1066, n_721, n_1157, n_841, n_1050, n_22, n_802, n_46, n_983, n_38, n_280, n_873, n_378, n_1112, n_762, n_1283, n_17, n_690, n_33, n_583, n_302, n_1203, n_821, n_321, n_1179, n_621, n_753, n_455, n_1048, n_1288, n_212, n_385, n_507, n_330, n_1228, n_972, n_692, n_820, n_1200, n_1185, n_991, n_828, n_779, n_576, n_1143, n_804, n_537, n_945, n_492, n_153, n_943, n_341, n_250, n_992, n_543, n_260, n_842, n_650, n_984, n_694, n_286, n_883, n_470, n_325, n_449, n_132, n_1214, n_900, n_856, n_918, n_942, n_189, n_1147, n_13, n_1077, n_540, n_618, n_896, n_323, n_195, n_356, n_894, n_831, n_964, n_1096, n_234, n_833, n_5, n_225, n_988, n_814, n_192, n_1201, n_1114, n_655, n_669, n_472, n_1176, n_387, n_1149, n_398, n_635, n_763, n_1020, n_1062, n_211, n_1219, n_3, n_1204, n_178, n_1035, n_287, n_555, n_783, n_1188, n_661, n_41, n_849, n_15, n_336, n_584, n_681, n_50, n_430, n_510, n_216, n_311, n_830, n_801, n_241, n_875, n_357, n_1110, n_445, n_749, n_1134, n_717, n_165, n_939, n_482, n_1088, n_588, n_1173, n_789, n_1232, n_734, n_638, n_866, n_107, n_969, n_1019, n_1105, n_249, n_304, n_577, n_338, n_149, n_693, n_14, n_836, n_990, n_975, n_1256, n_567, n_778, n_1122, n_151, n_306, n_458, n_770, n_1102, n_711, n_85, n_1187, n_1164, n_489, n_1174, n_617, n_876, n_1190, n_118, n_601, n_917, n_966, n_253, n_1116, n_1212, n_172, n_206, n_217, n_726, n_982, n_818, n_861, n_1183, n_899, n_1253, n_210, n_774, n_1059, n_176, n_1133, n_557, n_1005, n_607, n_1003, n_679, n_710, n_527, n_1168, n_707, n_937, n_393, n_108, n_487, n_665, n_66, n_177, n_421, n_910, n_768, n_205, n_1136, n_754, n_179, n_1125, n_125, n_410, n_708, n_529, n_735, n_232, n_1109, n_126, n_895, n_202, n_427, n_791, n_732, n_193, n_808, n_797, n_1025, n_500, n_1067, n_148, n_435, n_159, n_766, n_541, n_538, n_1117, n_799, n_687, n_715, n_1213, n_1266, n_536, n_872, n_594, n_200, n_1291, n_1155, n_89, n_115, n_1011, n_1184, n_985, n_869, n_810, n_416, n_827, n_401, n_626, n_1144, n_1137, n_1170, n_305, n_137, n_676, n_294, n_318, n_653, n_642, n_194, n_855, n_1178, n_850, n_684, n_124, n_268, n_664, n_503, n_235, n_605, n_1273, n_353, n_620, n_643, n_916, n_1081, n_493, n_1235, n_703, n_698, n_980, n_1115, n_1282, n_780, n_998, n_467, n_1227, n_840, n_501, n_823, n_245, n_725, n_672, n_581, n_382, n_554, n_898, n_1013, n_718, n_265, n_1120, n_719, n_443, n_198, n_714, n_909, n_997, n_932, n_612, n_788, n_119, n_1268, n_559, n_825, n_508, n_506, n_737, n_986, n_509, n_147, n_1281, n_67, n_1192, n_1024, n_1063, n_209, n_733, n_941, n_981, n_68, n_867, n_186, n_134, n_587, n_63, n_792, n_756, n_399, n_1238, n_548, n_812, n_298, n_518, n_505, n_282, n_752, n_905, n_1108, n_782, n_1100, n_862, n_760, n_381, n_220, n_390, n_31, n_481, n_769, n_42, n_1046, n_271, n_934, n_826, n_886, n_1221, n_654, n_1172, n_167, n_379, n_428, n_570, n_853, n_377, n_751, n_786, n_1083, n_1142, n_1129, n_392, n_158, n_704, n_787, n_138, n_961, n_771, n_276, n_95, n_1225, n_169, n_522, n_1287, n_1262, n_400, n_930, n_181, n_221, n_622, n_1087, n_386, n_994, n_848, n_1223, n_1272, n_104, n_682, n_56, n_141, n_1247, n_922, n_816, n_591, n_145, n_313, n_631, n_479, n_1246, n_432, n_839, n_1210, n_328, n_140, n_1250, n_369, n_871, n_598, n_685, n_928, n_608, n_78, n_772, n_499, n_517, n_98, n_402, n_413, n_1086, n_796, n_236, n_1012, n_1, n_903, n_740, n_203, n_384, n_80, n_35, n_277, n_1061, n_92, n_333, n_462, n_1193, n_1255, n_258, n_1113, n_29, n_79, n_1226, n_722, n_1277, n_188, n_844, n_201, n_471, n_852, n_40, n_1028, n_781, n_474, n_542, n_463, n_595, n_502, n_466, n_420, n_632, n_699, n_979, n_1245, n_846, n_465, n_76, n_362, n_170, n_27, n_161, n_273, n_585, n_270, n_616, n_81, n_745, n_1103, n_648, n_312, n_1076, n_1091, n_494, n_641, n_730, n_354, n_575, n_480, n_425, n_795, n_695, n_180, n_656, n_1220, n_37, n_229, n_437, n_60, n_403, n_453, n_1130, n_720, n_0, n_863, n_805, n_1275, n_113, n_712, n_246, n_1042, n_269, n_285, n_412, n_657, n_644, n_1160, n_491, n_1258, n_1074, n_251, n_160, n_566, n_565, n_597, n_1181, n_1196, n_651, n_334, n_811, n_807, n_835, n_175, n_666, n_262, n_99, n_1254, n_1026, n_1234, n_319, n_364, n_1138, n_927, n_20, n_1089, n_1004, n_1186, n_1032, n_242, n_1018, n_438, n_713, n_904, n_166, n_1180, n_1271, n_533, n_1251, n_278, n_5399);

input n_924;
input n_1263;
input n_977;
input n_611;
input n_1126;
input n_1166;
input n_469;
input n_82;
input n_785;
input n_549;
input n_532;
input n_1161;
input n_1150;
input n_226;
input n_667;
input n_790;
input n_1055;
input n_111;
input n_880;
input n_544;
input n_1007;
input n_155;
input n_552;
input n_1198;
input n_1099;
input n_956;
input n_564;
input n_423;
input n_21;
input n_105;
input n_1021;
input n_4;
input n_551;
input n_688;
input n_800;
input n_671;
input n_819;
input n_1022;
input n_915;
input n_864;
input n_173;
input n_859;
input n_951;
input n_1264;
input n_447;
input n_247;
input n_292;
input n_625;
input n_854;
input n_674;
input n_417;
input n_516;
input n_933;
input n_1152;
input n_497;
input n_606;
input n_275;
input n_26;
input n_877;
input n_2;
input n_755;
input n_1118;
input n_6;
input n_947;
input n_1285;
input n_373;
input n_307;
input n_530;
input n_87;
input n_150;
input n_1107;
input n_556;
input n_1230;
input n_668;
input n_375;
input n_301;
input n_929;
input n_1124;
input n_902;
input n_191;
input n_1104;
input n_659;
input n_51;
input n_1257;
input n_171;
input n_1182;
input n_579;
input n_1261;
input n_938;
input n_1098;
input n_320;
input n_1154;
input n_1242;
input n_1135;
input n_24;
input n_406;
input n_519;
input n_1016;
input n_1243;
input n_546;
input n_101;
input n_1280;
input n_281;
input n_240;
input n_291;
input n_231;
input n_257;
input n_731;
input n_371;
input n_709;
input n_317;
input n_1236;
input n_569;
input n_227;
input n_920;
input n_1289;
input n_94;
input n_335;
input n_370;
input n_976;
input n_343;
input n_308;
input n_297;
input n_156;
input n_1078;
input n_775;
input n_219;
input n_157;
input n_600;
input n_223;
input n_264;
input n_955;
input n_163;
input n_339;
input n_1146;
input n_882;
input n_183;
input n_243;
input n_1036;
input n_1097;
input n_347;
input n_59;
input n_550;
input n_696;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_646;
input n_436;
input n_1216;
input n_290;
input n_580;
input n_1040;
input n_578;
input n_926;
input n_344;
input n_1218;
input n_422;
input n_475;
input n_777;
input n_1070;
input n_1030;
input n_72;
input n_415;
input n_1071;
input n_485;
input n_1165;
input n_1267;
input n_496;
input n_958;
input n_1034;
input n_670;
input n_48;
input n_521;
input n_663;
input n_845;
input n_673;
input n_837;
input n_1239;
input n_528;
input n_680;
input n_395;
input n_164;
input n_553;
input n_901;
input n_813;
input n_1284;
input n_214;
input n_675;
input n_888;
input n_1167;
input n_637;
input n_184;
input n_446;
input n_1064;
input n_144;
input n_858;
input n_114;
input n_96;
input n_923;
input n_691;
input n_1151;
input n_881;
input n_468;
input n_213;
input n_129;
input n_342;
input n_464;
input n_363;
input n_197;
input n_1069;
input n_1075;
input n_460;
input n_889;
input n_973;
input n_477;
input n_571;
input n_461;
input n_1211;
input n_1197;
input n_907;
input n_190;
input n_989;
input n_1039;
input n_34;
input n_228;
input n_283;
input n_488;
input n_736;
input n_892;
input n_1000;
input n_1202;
input n_1278;
input n_1002;
input n_49;
input n_310;
input n_54;
input n_593;
input n_12;
input n_748;
input n_586;
input n_1058;
input n_838;
input n_332;
input n_1053;
input n_1224;
input n_349;
input n_1248;
input n_230;
input n_953;
input n_279;
input n_1014;
input n_1241;
input n_70;
input n_289;
input n_963;
input n_1052;
input n_954;
input n_627;
input n_440;
input n_793;
input n_478;
input n_476;
input n_534;
input n_884;
input n_345;
input n_944;
input n_91;
input n_182;
input n_143;
input n_647;
input n_237;
input n_407;
input n_1072;
input n_832;
input n_857;
input n_207;
input n_561;
input n_18;
input n_1027;
input n_971;
input n_1156;
input n_117;
input n_326;
input n_794;
input n_404;
input n_686;
input n_847;
input n_596;
input n_558;
input n_702;
input n_1276;
input n_822;
input n_728;
input n_266;
input n_1162;
input n_272;
input n_1199;
input n_352;
input n_53;
input n_1038;
input n_520;
input n_409;
input n_887;
input n_154;
input n_71;
input n_300;
input n_809;
input n_870;
input n_931;
input n_599;
input n_434;
input n_868;
input n_639;
input n_914;
input n_411;
input n_414;
input n_965;
input n_935;
input n_121;
input n_1175;
input n_817;
input n_360;
input n_36;
input n_64;
input n_759;
input n_28;
input n_806;
input n_324;
input n_187;
input n_1189;
input n_103;
input n_97;
input n_11;
input n_7;
input n_1259;
input n_706;
input n_746;
input n_747;
input n_52;
input n_784;
input n_110;
input n_1244;
input n_431;
input n_1194;
input n_615;
input n_851;
input n_843;
input n_523;
input n_913;
input n_705;
input n_865;
input n_61;
input n_678;
input n_697;
input n_127;
input n_1222;
input n_75;
input n_776;
input n_367;
input n_452;
input n_525;
input n_1260;
input n_649;
input n_547;
input n_43;
input n_1191;
input n_116;
input n_284;
input n_1128;
input n_139;
input n_744;
input n_590;
input n_629;
input n_254;
input n_1233;
input n_23;
input n_526;
input n_293;
input n_372;
input n_677;
input n_244;
input n_47;
input n_1121;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_949;
input n_100;
input n_1008;
input n_946;
input n_1001;
input n_498;
input n_689;
input n_738;
input n_640;
input n_252;
input n_624;
input n_295;
input n_133;
input n_1010;
input n_1231;
input n_739;
input n_1279;
input n_1195;
input n_610;
input n_936;
input n_568;
input n_39;
input n_1090;
input n_757;
input n_633;
input n_439;
input n_106;
input n_259;
input n_448;
input n_758;
input n_999;
input n_93;
input n_1158;
input n_563;
input n_1145;
input n_878;
input n_524;
input n_204;
input n_394;
input n_1049;
input n_1153;
input n_741;
input n_1068;
input n_122;
input n_331;
input n_10;
input n_906;
input n_1163;
input n_1207;
input n_919;
input n_908;
input n_90;
input n_724;
input n_658;
input n_456;
input n_959;
input n_535;
input n_152;
input n_940;
input n_9;
input n_592;
input n_1169;
input n_45;
input n_1017;
input n_123;
input n_978;
input n_1054;
input n_1269;
input n_1095;
input n_267;
input n_514;
input n_457;
input n_1079;
input n_1045;
input n_1208;
input n_603;
input n_484;
input n_1033;
input n_442;
input n_131;
input n_636;
input n_660;
input n_1009;
input n_1148;
input n_109;
input n_742;
input n_750;
input n_995;
input n_454;
input n_374;
input n_185;
input n_396;
input n_1073;
input n_255;
input n_662;
input n_459;
input n_218;
input n_962;
input n_1215;
input n_1171;
input n_723;
input n_1065;
input n_473;
input n_1043;
input n_355;
input n_486;
input n_614;
input n_337;
input n_88;
input n_1286;
input n_1177;
input n_168;
input n_974;
input n_727;
input n_1159;
input n_957;
input n_773;
input n_208;
input n_142;
input n_743;
input n_299;
input n_303;
input n_296;
input n_613;
input n_1119;
input n_1240;
input n_65;
input n_829;
input n_361;
input n_700;
input n_1237;
input n_573;
input n_69;
input n_1132;
input n_388;
input n_1127;
input n_761;
input n_1006;
input n_329;
input n_274;
input n_1270;
input n_582;
input n_73;
input n_19;
input n_309;
input n_30;
input n_512;
input n_84;
input n_130;
input n_322;
input n_1249;
input n_652;
input n_1111;
input n_25;
input n_1093;
input n_288;
input n_1031;
input n_263;
input n_609;
input n_1041;
input n_1265;
input n_44;
input n_224;
input n_383;
input n_834;
input n_112;
input n_765;
input n_893;
input n_1015;
input n_1140;
input n_891;
input n_239;
input n_630;
input n_55;
input n_504;
input n_511;
input n_874;
input n_358;
input n_1101;
input n_77;
input n_102;
input n_1106;
input n_987;
input n_261;
input n_174;
input n_767;
input n_993;
input n_545;
input n_441;
input n_860;
input n_450;
input n_429;
input n_948;
input n_1217;
input n_628;
input n_365;
input n_729;
input n_1131;
input n_1084;
input n_970;
input n_911;
input n_83;
input n_513;
input n_1094;
input n_560;
input n_340;
input n_1044;
input n_1205;
input n_346;
input n_1209;
input n_495;
input n_602;
input n_574;
input n_879;
input n_16;
input n_58;
input n_623;
input n_405;
input n_824;
input n_359;
input n_490;
input n_996;
input n_921;
input n_233;
input n_572;
input n_366;
input n_815;
input n_128;
input n_120;
input n_327;
input n_135;
input n_1037;
input n_1080;
input n_1274;
input n_426;
input n_1082;
input n_589;
input n_716;
input n_562;
input n_62;
input n_952;
input n_1229;
input n_391;
input n_701;
input n_1023;
input n_645;
input n_539;
input n_803;
input n_1092;
input n_238;
input n_531;
input n_890;
input n_764;
input n_1056;
input n_162;
input n_960;
input n_222;
input n_1290;
input n_1123;
input n_1047;
input n_634;
input n_199;
input n_32;
input n_1252;
input n_348;
input n_1029;
input n_925;
input n_1206;
input n_424;
input n_256;
input n_950;
input n_380;
input n_419;
input n_444;
input n_1060;
input n_1141;
input n_316;
input n_389;
input n_418;
input n_248;
input n_136;
input n_86;
input n_146;
input n_912;
input n_315;
input n_968;
input n_451;
input n_619;
input n_408;
input n_376;
input n_967;
input n_74;
input n_1139;
input n_515;
input n_57;
input n_351;
input n_885;
input n_397;
input n_483;
input n_683;
input n_1057;
input n_1051;
input n_1085;
input n_1066;
input n_721;
input n_1157;
input n_841;
input n_1050;
input n_22;
input n_802;
input n_46;
input n_983;
input n_38;
input n_280;
input n_873;
input n_378;
input n_1112;
input n_762;
input n_1283;
input n_17;
input n_690;
input n_33;
input n_583;
input n_302;
input n_1203;
input n_821;
input n_321;
input n_1179;
input n_621;
input n_753;
input n_455;
input n_1048;
input n_1288;
input n_212;
input n_385;
input n_507;
input n_330;
input n_1228;
input n_972;
input n_692;
input n_820;
input n_1200;
input n_1185;
input n_991;
input n_828;
input n_779;
input n_576;
input n_1143;
input n_804;
input n_537;
input n_945;
input n_492;
input n_153;
input n_943;
input n_341;
input n_250;
input n_992;
input n_543;
input n_260;
input n_842;
input n_650;
input n_984;
input n_694;
input n_286;
input n_883;
input n_470;
input n_325;
input n_449;
input n_132;
input n_1214;
input n_900;
input n_856;
input n_918;
input n_942;
input n_189;
input n_1147;
input n_13;
input n_1077;
input n_540;
input n_618;
input n_896;
input n_323;
input n_195;
input n_356;
input n_894;
input n_831;
input n_964;
input n_1096;
input n_234;
input n_833;
input n_5;
input n_225;
input n_988;
input n_814;
input n_192;
input n_1201;
input n_1114;
input n_655;
input n_669;
input n_472;
input n_1176;
input n_387;
input n_1149;
input n_398;
input n_635;
input n_763;
input n_1020;
input n_1062;
input n_211;
input n_1219;
input n_3;
input n_1204;
input n_178;
input n_1035;
input n_287;
input n_555;
input n_783;
input n_1188;
input n_661;
input n_41;
input n_849;
input n_15;
input n_336;
input n_584;
input n_681;
input n_50;
input n_430;
input n_510;
input n_216;
input n_311;
input n_830;
input n_801;
input n_241;
input n_875;
input n_357;
input n_1110;
input n_445;
input n_749;
input n_1134;
input n_717;
input n_165;
input n_939;
input n_482;
input n_1088;
input n_588;
input n_1173;
input n_789;
input n_1232;
input n_734;
input n_638;
input n_866;
input n_107;
input n_969;
input n_1019;
input n_1105;
input n_249;
input n_304;
input n_577;
input n_338;
input n_149;
input n_693;
input n_14;
input n_836;
input n_990;
input n_975;
input n_1256;
input n_567;
input n_778;
input n_1122;
input n_151;
input n_306;
input n_458;
input n_770;
input n_1102;
input n_711;
input n_85;
input n_1187;
input n_1164;
input n_489;
input n_1174;
input n_617;
input n_876;
input n_1190;
input n_118;
input n_601;
input n_917;
input n_966;
input n_253;
input n_1116;
input n_1212;
input n_172;
input n_206;
input n_217;
input n_726;
input n_982;
input n_818;
input n_861;
input n_1183;
input n_899;
input n_1253;
input n_210;
input n_774;
input n_1059;
input n_176;
input n_1133;
input n_557;
input n_1005;
input n_607;
input n_1003;
input n_679;
input n_710;
input n_527;
input n_1168;
input n_707;
input n_937;
input n_393;
input n_108;
input n_487;
input n_665;
input n_66;
input n_177;
input n_421;
input n_910;
input n_768;
input n_205;
input n_1136;
input n_754;
input n_179;
input n_1125;
input n_125;
input n_410;
input n_708;
input n_529;
input n_735;
input n_232;
input n_1109;
input n_126;
input n_895;
input n_202;
input n_427;
input n_791;
input n_732;
input n_193;
input n_808;
input n_797;
input n_1025;
input n_500;
input n_1067;
input n_148;
input n_435;
input n_159;
input n_766;
input n_541;
input n_538;
input n_1117;
input n_799;
input n_687;
input n_715;
input n_1213;
input n_1266;
input n_536;
input n_872;
input n_594;
input n_200;
input n_1291;
input n_1155;
input n_89;
input n_115;
input n_1011;
input n_1184;
input n_985;
input n_869;
input n_810;
input n_416;
input n_827;
input n_401;
input n_626;
input n_1144;
input n_1137;
input n_1170;
input n_305;
input n_137;
input n_676;
input n_294;
input n_318;
input n_653;
input n_642;
input n_194;
input n_855;
input n_1178;
input n_850;
input n_684;
input n_124;
input n_268;
input n_664;
input n_503;
input n_235;
input n_605;
input n_1273;
input n_353;
input n_620;
input n_643;
input n_916;
input n_1081;
input n_493;
input n_1235;
input n_703;
input n_698;
input n_980;
input n_1115;
input n_1282;
input n_780;
input n_998;
input n_467;
input n_1227;
input n_840;
input n_501;
input n_823;
input n_245;
input n_725;
input n_672;
input n_581;
input n_382;
input n_554;
input n_898;
input n_1013;
input n_718;
input n_265;
input n_1120;
input n_719;
input n_443;
input n_198;
input n_714;
input n_909;
input n_997;
input n_932;
input n_612;
input n_788;
input n_119;
input n_1268;
input n_559;
input n_825;
input n_508;
input n_506;
input n_737;
input n_986;
input n_509;
input n_147;
input n_1281;
input n_67;
input n_1192;
input n_1024;
input n_1063;
input n_209;
input n_733;
input n_941;
input n_981;
input n_68;
input n_867;
input n_186;
input n_134;
input n_587;
input n_63;
input n_792;
input n_756;
input n_399;
input n_1238;
input n_548;
input n_812;
input n_298;
input n_518;
input n_505;
input n_282;
input n_752;
input n_905;
input n_1108;
input n_782;
input n_1100;
input n_862;
input n_760;
input n_381;
input n_220;
input n_390;
input n_31;
input n_481;
input n_769;
input n_42;
input n_1046;
input n_271;
input n_934;
input n_826;
input n_886;
input n_1221;
input n_654;
input n_1172;
input n_167;
input n_379;
input n_428;
input n_570;
input n_853;
input n_377;
input n_751;
input n_786;
input n_1083;
input n_1142;
input n_1129;
input n_392;
input n_158;
input n_704;
input n_787;
input n_138;
input n_961;
input n_771;
input n_276;
input n_95;
input n_1225;
input n_169;
input n_522;
input n_1287;
input n_1262;
input n_400;
input n_930;
input n_181;
input n_221;
input n_622;
input n_1087;
input n_386;
input n_994;
input n_848;
input n_1223;
input n_1272;
input n_104;
input n_682;
input n_56;
input n_141;
input n_1247;
input n_922;
input n_816;
input n_591;
input n_145;
input n_313;
input n_631;
input n_479;
input n_1246;
input n_432;
input n_839;
input n_1210;
input n_328;
input n_140;
input n_1250;
input n_369;
input n_871;
input n_598;
input n_685;
input n_928;
input n_608;
input n_78;
input n_772;
input n_499;
input n_517;
input n_98;
input n_402;
input n_413;
input n_1086;
input n_796;
input n_236;
input n_1012;
input n_1;
input n_903;
input n_740;
input n_203;
input n_384;
input n_80;
input n_35;
input n_277;
input n_1061;
input n_92;
input n_333;
input n_462;
input n_1193;
input n_1255;
input n_258;
input n_1113;
input n_29;
input n_79;
input n_1226;
input n_722;
input n_1277;
input n_188;
input n_844;
input n_201;
input n_471;
input n_852;
input n_40;
input n_1028;
input n_781;
input n_474;
input n_542;
input n_463;
input n_595;
input n_502;
input n_466;
input n_420;
input n_632;
input n_699;
input n_979;
input n_1245;
input n_846;
input n_465;
input n_76;
input n_362;
input n_170;
input n_27;
input n_161;
input n_273;
input n_585;
input n_270;
input n_616;
input n_81;
input n_745;
input n_1103;
input n_648;
input n_312;
input n_1076;
input n_1091;
input n_494;
input n_641;
input n_730;
input n_354;
input n_575;
input n_480;
input n_425;
input n_795;
input n_695;
input n_180;
input n_656;
input n_1220;
input n_37;
input n_229;
input n_437;
input n_60;
input n_403;
input n_453;
input n_1130;
input n_720;
input n_0;
input n_863;
input n_805;
input n_1275;
input n_113;
input n_712;
input n_246;
input n_1042;
input n_269;
input n_285;
input n_412;
input n_657;
input n_644;
input n_1160;
input n_491;
input n_1258;
input n_1074;
input n_251;
input n_160;
input n_566;
input n_565;
input n_597;
input n_1181;
input n_1196;
input n_651;
input n_334;
input n_811;
input n_807;
input n_835;
input n_175;
input n_666;
input n_262;
input n_99;
input n_1254;
input n_1026;
input n_1234;
input n_319;
input n_364;
input n_1138;
input n_927;
input n_20;
input n_1089;
input n_1004;
input n_1186;
input n_1032;
input n_242;
input n_1018;
input n_438;
input n_713;
input n_904;
input n_166;
input n_1180;
input n_1271;
input n_533;
input n_1251;
input n_278;

output n_5399;

wire n_2253;
wire n_2417;
wire n_2756;
wire n_4706;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_5287;
wire n_2327;
wire n_1488;
wire n_2899;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_2395;
wire n_5161;
wire n_5207;
wire n_2347;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_2021;
wire n_2391;
wire n_5035;
wire n_5282;
wire n_1960;
wire n_2843;
wire n_3615;
wire n_2059;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_3202;
wire n_4977;
wire n_3813;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_5033;
wire n_1462;
wire n_4211;
wire n_3448;
wire n_3019;
wire n_2096;
wire n_3776;
wire n_2530;
wire n_4517;
wire n_2483;
wire n_1696;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1860;
wire n_4615;
wire n_1728;
wire n_2076;
wire n_2147;
wire n_3010;
wire n_2770;
wire n_4131;
wire n_2584;
wire n_3188;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_3283;
wire n_2323;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_5202;
wire n_1314;
wire n_1512;
wire n_1490;
wire n_3214;
wire n_2091;
wire n_1517;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_1449;
wire n_4678;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_3947;
wire n_3490;
wire n_1948;
wire n_3868;
wire n_3183;
wire n_3437;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_5241;
wire n_2384;
wire n_3156;
wire n_3376;
wire n_5037;
wire n_4468;
wire n_3653;
wire n_3702;
wire n_4976;
wire n_2202;
wire n_2648;
wire n_5008;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_2439;
wire n_4811;
wire n_5398;
wire n_2276;
wire n_2089;
wire n_3420;
wire n_1561;
wire n_5144;
wire n_3361;
wire n_4758;
wire n_1600;
wire n_4255;
wire n_1796;
wire n_4484;
wire n_3668;
wire n_4237;
wire n_2934;
wire n_1672;
wire n_1880;
wire n_3550;
wire n_1626;
wire n_2079;
wire n_2238;
wire n_1405;
wire n_1706;
wire n_3418;
wire n_4901;
wire n_2859;
wire n_3395;
wire n_4917;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_2968;
wire n_1585;
wire n_2684;
wire n_3593;
wire n_5343;
wire n_1599;
wire n_4421;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_1377;
wire n_4469;
wire n_4414;
wire n_5184;
wire n_4532;
wire n_3339;
wire n_3735;
wire n_3349;
wire n_2248;
wire n_3007;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_2100;
wire n_5236;
wire n_3310;
wire n_3487;
wire n_2258;
wire n_1667;
wire n_3983;
wire n_4405;
wire n_1926;
wire n_1331;
wire n_4195;
wire n_4969;
wire n_4504;
wire n_1385;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_4531;
wire n_2987;
wire n_1527;
wire n_4567;
wire n_4164;
wire n_5315;
wire n_4234;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_5348;
wire n_2175;
wire n_5055;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_5397;
wire n_4471;
wire n_5031;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_3208;
wire n_3331;
wire n_2379;
wire n_4983;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_3649;
wire n_4302;
wire n_2514;
wire n_5189;
wire n_5381;
wire n_4786;
wire n_3257;
wire n_4160;
wire n_2293;
wire n_4051;
wire n_2028;
wire n_3009;
wire n_1412;
wire n_3981;
wire n_1841;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_1711;
wire n_1891;
wire n_5254;
wire n_3526;
wire n_2546;
wire n_3790;
wire n_3491;
wire n_4613;
wire n_4649;
wire n_1888;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_4028;
wire n_1690;
wire n_3819;
wire n_2449;
wire n_5083;
wire n_2297;
wire n_4186;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_3747;
wire n_2227;
wire n_4618;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_2876;
wire n_4099;
wire n_3484;
wire n_3620;
wire n_1746;
wire n_2479;
wire n_1464;
wire n_4295;
wire n_5303;
wire n_1444;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_4697;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_4810;
wire n_3317;
wire n_4391;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_1503;
wire n_4638;
wire n_1468;
wire n_3455;
wire n_5047;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_5346;
wire n_1994;
wire n_4707;
wire n_2577;
wire n_4527;
wire n_5109;
wire n_2796;
wire n_2342;
wire n_4156;
wire n_1851;
wire n_4848;
wire n_2937;
wire n_3095;
wire n_2805;
wire n_4918;
wire n_3856;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_5010;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_2857;
wire n_5358;
wire n_4528;
wire n_3932;
wire n_4619;
wire n_4673;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1596;
wire n_2947;
wire n_4299;
wire n_4801;
wire n_1474;
wire n_1665;
wire n_3515;
wire n_2886;
wire n_2093;
wire n_2473;
wire n_3287;
wire n_3378;
wire n_1431;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_5373;
wire n_4294;
wire n_1732;
wire n_5279;
wire n_4125;
wire n_4232;
wire n_4949;
wire n_2941;
wire n_2457;
wire n_4790;
wire n_2536;
wire n_1336;
wire n_1758;
wire n_2952;
wire n_4847;
wire n_5321;
wire n_3058;
wire n_5096;
wire n_4365;
wire n_1878;
wire n_3505;
wire n_4610;
wire n_3730;
wire n_4489;
wire n_5210;
wire n_4967;
wire n_4992;
wire n_3001;
wire n_3945;
wire n_4542;
wire n_2261;
wire n_2729;
wire n_3597;
wire n_1612;
wire n_2897;
wire n_2077;
wire n_4198;
wire n_2909;
wire n_4534;
wire n_4500;
wire n_5014;
wire n_3185;
wire n_1300;
wire n_3523;
wire n_1785;
wire n_2829;
wire n_4597;
wire n_4329;
wire n_4087;
wire n_3811;
wire n_1664;
wire n_3200;
wire n_2231;
wire n_2017;
wire n_2604;
wire n_4257;
wire n_3453;
wire n_2390;
wire n_3213;
wire n_3077;
wire n_1562;
wire n_3474;
wire n_3984;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_1913;
wire n_1823;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_4189;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_3707;
wire n_1846;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_4687;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_4037;
wire n_2922;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2727;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_1552;
wire n_3618;
wire n_2593;
wire n_5262;
wire n_3683;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_1327;
wire n_4763;
wire n_1684;
wire n_3590;
wire n_5310;
wire n_4594;
wire n_3424;
wire n_1381;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_2419;
wire n_3215;
wire n_5146;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_2786;
wire n_3171;
wire n_1437;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_3468;
wire n_2910;
wire n_1893;
wire n_1467;
wire n_2163;
wire n_2254;
wire n_1382;
wire n_3546;
wire n_2647;
wire n_1311;
wire n_1519;
wire n_4443;
wire n_4507;
wire n_2443;
wire n_1811;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_3244;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_4452;
wire n_4348;
wire n_5362;
wire n_4355;
wire n_3494;
wire n_5050;
wire n_5063;
wire n_5229;
wire n_2125;
wire n_3771;
wire n_5199;
wire n_3110;
wire n_3073;
wire n_4572;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_1608;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_1305;
wire n_5266;
wire n_3178;
wire n_5355;
wire n_2334;
wire n_4521;
wire n_4488;
wire n_2289;
wire n_3051;
wire n_1343;
wire n_2783;
wire n_2263;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_4519;
wire n_3715;
wire n_3040;
wire n_1938;
wire n_2499;
wire n_3568;
wire n_3737;
wire n_1967;
wire n_1329;
wire n_3255;
wire n_4856;
wire n_2997;
wire n_4400;
wire n_5168;
wire n_3326;
wire n_3734;
wire n_4778;
wire n_2429;
wire n_5322;
wire n_1793;
wire n_4352;
wire n_4441;
wire n_4761;
wire n_1804;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_2533;
wire n_2364;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_5371;
wire n_2291;
wire n_4043;
wire n_1636;
wire n_3601;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_2094;
wire n_1575;
wire n_2393;
wire n_1697;
wire n_5316;
wire n_3831;
wire n_3801;
wire n_2043;
wire n_2751;
wire n_4893;
wire n_5032;
wire n_1549;
wire n_1934;
wire n_4948;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_1446;
wire n_4406;
wire n_2758;
wire n_1458;
wire n_1807;
wire n_2618;
wire n_5112;
wire n_5386;
wire n_2559;
wire n_4748;
wire n_2295;
wire n_3931;
wire n_4010;
wire n_2840;
wire n_5017;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_4607;
wire n_5123;
wire n_4117;
wire n_3636;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_2795;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_3380;
wire n_2098;
wire n_1296;
wire n_3460;
wire n_3409;
wire n_3538;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_4728;
wire n_4247;
wire n_4933;
wire n_4018;
wire n_3900;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_3872;
wire n_4336;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_3877;
wire n_2995;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_4052;
wire n_3459;
wire n_1499;
wire n_4398;
wire n_3155;
wire n_2633;
wire n_4954;
wire n_2435;
wire n_1392;
wire n_2097;
wire n_4304;
wire n_3911;
wire n_5333;
wire n_1303;
wire n_4431;
wire n_4192;
wire n_3736;
wire n_4805;
wire n_4885;
wire n_1661;
wire n_3565;
wire n_4701;
wire n_2575;
wire n_5040;
wire n_1658;
wire n_1904;
wire n_1345;
wire n_1899;
wire n_2067;
wire n_2219;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_1726;
wire n_4631;
wire n_3035;
wire n_5194;
wire n_1657;
wire n_1475;
wire n_1725;
wire n_1313;
wire n_1491;
wire n_3639;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_1915;
wire n_5239;
wire n_1310;
wire n_2605;
wire n_4747;
wire n_5197;
wire n_1399;
wire n_1979;
wire n_2924;
wire n_4111;
wire n_2484;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_5305;
wire n_4538;
wire n_2754;
wire n_1742;
wire n_5376;
wire n_2489;
wire n_5204;
wire n_2012;
wire n_4094;
wire n_3503;
wire n_2866;
wire n_3561;
wire n_1418;
wire n_2917;
wire n_2425;
wire n_3536;
wire n_3661;
wire n_4150;
wire n_4878;
wire n_1703;
wire n_1650;
wire n_3934;
wire n_4985;
wire n_3922;
wire n_3846;
wire n_2103;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_3074;
wire n_1999;
wire n_2372;
wire n_3673;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_2430;
wire n_2433;
wire n_3293;
wire n_4022;
wire n_1531;
wire n_1334;
wire n_4852;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_3415;
wire n_2284;
wire n_2817;
wire n_3139;
wire n_5292;
wire n_2598;
wire n_4601;
wire n_2687;
wire n_1890;
wire n_4220;
wire n_1944;
wire n_1497;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_4515;
wire n_4351;
wire n_5264;
wire n_3126;
wire n_4403;
wire n_1981;
wire n_1663;
wire n_1718;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_1518;
wire n_4223;
wire n_1889;
wire n_1489;
wire n_5025;
wire n_2966;
wire n_1376;
wire n_2326;
wire n_1569;
wire n_2188;
wire n_1429;
wire n_4644;
wire n_4456;
wire n_5060;
wire n_5334;
wire n_2448;
wire n_4346;
wire n_3170;
wire n_2748;
wire n_3311;
wire n_3272;
wire n_2898;
wire n_2717;
wire n_1861;
wire n_3628;
wire n_3691;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_2573;
wire n_4435;
wire n_2939;
wire n_3807;
wire n_2447;
wire n_4764;
wire n_5394;
wire n_2774;
wire n_1707;
wire n_4655;
wire n_3161;
wire n_4581;
wire n_4827;
wire n_2488;
wire n_3477;
wire n_2476;
wire n_4399;
wire n_2781;
wire n_5309;
wire n_2778;
wire n_4782;
wire n_1520;
wire n_4363;
wire n_2887;
wire n_4864;
wire n_2691;
wire n_1411;
wire n_3054;
wire n_4335;
wire n_2526;
wire n_2703;
wire n_2167;
wire n_3391;
wire n_4259;
wire n_2709;
wire n_1536;
wire n_4865;
wire n_4056;
wire n_1344;
wire n_4564;
wire n_3840;
wire n_1339;
wire n_5085;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_2173;
wire n_1842;
wire n_3738;
wire n_5116;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_1555;
wire n_3245;
wire n_4417;
wire n_4899;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_2453;
wire n_4798;
wire n_1525;
wire n_3509;
wire n_3352;
wire n_3076;
wire n_3535;
wire n_2182;
wire n_3251;
wire n_2931;
wire n_5185;
wire n_3118;
wire n_3511;
wire n_3443;
wire n_2146;
wire n_1487;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_3521;
wire n_5379;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_1515;
wire n_2918;
wire n_3232;
wire n_1673;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_4981;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_4430;
wire n_4081;
wire n_3132;
wire n_4407;
wire n_3951;
wire n_4894;
wire n_3238;
wire n_3210;
wire n_2036;
wire n_3267;
wire n_4995;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_3884;
wire n_3726;
wire n_2525;
wire n_2892;
wire n_2907;
wire n_3577;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1741;
wire n_4057;
wire n_4332;
wire n_4314;
wire n_3347;
wire n_3216;
wire n_1621;
wire n_3809;
wire n_2113;
wire n_1448;
wire n_4288;
wire n_3567;
wire n_5066;
wire n_1634;
wire n_3939;
wire n_4241;
wire n_3321;
wire n_3212;
wire n_1433;
wire n_2256;
wire n_3152;
wire n_5106;
wire n_2920;
wire n_4265;
wire n_5319;
wire n_2247;
wire n_1622;
wire n_3705;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_2268;
wire n_3778;
wire n_5337;
wire n_3304;
wire n_1378;
wire n_3912;
wire n_1729;
wire n_2739;
wire n_2771;
wire n_4604;
wire n_5223;
wire n_3795;
wire n_5020;
wire n_4419;
wire n_4477;
wire n_3179;
wire n_3256;
wire n_2386;
wire n_1501;
wire n_3086;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_5074;
wire n_2568;
wire n_5364;
wire n_1738;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_4639;
wire n_3713;
wire n_3663;
wire n_5046;
wire n_5166;
wire n_3246;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_5088;
wire n_2302;
wire n_1494;
wire n_2069;
wire n_3434;
wire n_1806;
wire n_1563;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_4243;
wire n_4982;
wire n_3695;
wire n_4330;
wire n_2482;
wire n_2677;
wire n_3832;
wire n_3987;
wire n_5352;
wire n_4991;
wire n_1698;
wire n_2329;
wire n_2142;
wire n_3332;
wire n_3048;
wire n_3937;
wire n_2203;
wire n_4525;
wire n_3782;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_3786;
wire n_2888;
wire n_3638;
wire n_1633;
wire n_4177;
wire n_3763;
wire n_2669;
wire n_1778;
wire n_2306;
wire n_3022;
wire n_4264;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_5129;
wire n_2149;
wire n_3060;
wire n_4276;
wire n_5219;
wire n_3013;
wire n_1984;
wire n_5170;
wire n_2408;
wire n_5320;
wire n_1877;
wire n_3049;
wire n_1723;
wire n_5107;
wire n_4485;
wire n_4626;
wire n_2659;
wire n_1414;
wire n_4975;
wire n_1852;
wire n_3089;
wire n_2470;
wire n_3985;
wire n_5253;
wire n_1391;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_2551;
wire n_1587;
wire n_2682;
wire n_3440;
wire n_1748;
wire n_4569;
wire n_2699;
wire n_4897;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_2615;
wire n_3940;
wire n_2985;
wire n_5065;
wire n_2753;
wire n_1582;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_3141;
wire n_5084;
wire n_3164;
wire n_3570;
wire n_5260;
wire n_4919;
wire n_4025;
wire n_2712;
wire n_5328;
wire n_3936;
wire n_4503;
wire n_3507;
wire n_3821;
wire n_2700;
wire n_3367;
wire n_4464;
wire n_3096;
wire n_3496;
wire n_4114;
wire n_2544;
wire n_2356;
wire n_4556;
wire n_2620;
wire n_1581;
wire n_4089;
wire n_2919;
wire n_4327;
wire n_4218;
wire n_2150;
wire n_3146;
wire n_5165;
wire n_2241;
wire n_2757;
wire n_4353;
wire n_2042;
wire n_1754;
wire n_1623;
wire n_2921;
wire n_2720;
wire n_1854;
wire n_4990;
wire n_1856;
wire n_4959;
wire n_4161;
wire n_1319;
wire n_3992;
wire n_2616;
wire n_1906;
wire n_4103;
wire n_1387;
wire n_4466;
wire n_2262;
wire n_2462;
wire n_1532;
wire n_3625;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2837;
wire n_4844;
wire n_2979;
wire n_5257;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_2548;
wire n_5180;
wire n_2108;
wire n_3640;
wire n_4388;
wire n_4206;
wire n_1538;
wire n_1779;
wire n_4738;
wire n_1369;
wire n_3909;
wire n_3207;
wire n_3944;
wire n_4434;
wire n_4837;
wire n_3042;
wire n_1942;
wire n_2510;
wire n_4219;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_5012;
wire n_1293;
wire n_1876;
wire n_4620;
wire n_1810;
wire n_2813;
wire n_4438;
wire n_2009;
wire n_2222;
wire n_3510;
wire n_3218;
wire n_2667;
wire n_3150;
wire n_4325;
wire n_1733;
wire n_2413;
wire n_3775;
wire n_4133;
wire n_4184;
wire n_5203;
wire n_2518;
wire n_2629;
wire n_4481;
wire n_3416;
wire n_4379;
wire n_2181;
wire n_1829;
wire n_4030;
wire n_4490;
wire n_3138;
wire n_4397;
wire n_1710;
wire n_2928;
wire n_1734;
wire n_4820;
wire n_3770;
wire n_1308;
wire n_5094;
wire n_4938;
wire n_4179;
wire n_3469;
wire n_5336;
wire n_2723;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_3855;
wire n_2054;
wire n_5339;
wire n_1559;
wire n_4931;
wire n_1765;
wire n_3158;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_3113;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_2856;
wire n_1832;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_3828;
wire n_3288;
wire n_4404;
wire n_5091;
wire n_1509;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_3667;
wire n_1306;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_4356;
wire n_2061;
wire n_4432;
wire n_5251;
wire n_2378;
wire n_1740;
wire n_1586;
wire n_4291;
wire n_4386;
wire n_4149;
wire n_1492;
wire n_1692;
wire n_2982;
wire n_2481;
wire n_3545;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_1614;
wire n_2339;
wire n_4637;
wire n_4935;
wire n_4785;
wire n_3426;
wire n_3454;
wire n_3820;
wire n_3741;
wire n_3410;
wire n_2029;
wire n_1609;
wire n_5298;
wire n_1887;
wire n_4413;
wire n_2346;
wire n_3990;
wire n_4493;
wire n_3475;
wire n_1592;
wire n_2882;
wire n_1721;
wire n_2338;
wire n_3672;
wire n_5290;
wire n_3197;
wire n_3109;
wire n_2721;
wire n_5095;
wire n_3002;
wire n_5324;
wire n_3897;
wire n_3845;
wire n_2081;
wire n_4570;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_1820;
wire n_5019;
wire n_2418;
wire n_2179;
wire n_1416;
wire n_2521;
wire n_1724;
wire n_3458;
wire n_1420;
wire n_3330;
wire n_4606;
wire n_4774;
wire n_2477;
wire n_3887;
wire n_4093;
wire n_1486;
wire n_4672;
wire n_3519;
wire n_4174;
wire n_3374;
wire n_3045;
wire n_2367;
wire n_1870;
wire n_4766;
wire n_2896;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_1927;
wire n_1349;
wire n_4460;
wire n_3645;
wire n_3223;
wire n_3929;
wire n_2255;
wire n_2272;
wire n_1965;
wire n_1902;
wire n_1941;
wire n_3938;
wire n_5377;
wire n_2878;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_3189;
wire n_2066;
wire n_3154;
wire n_1551;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_2220;
wire n_4349;
wire n_3788;
wire n_2410;
wire n_4313;
wire n_1935;
wire n_3366;
wire n_1534;
wire n_1351;
wire n_2696;
wire n_4863;
wire n_3242;
wire n_3525;
wire n_3486;
wire n_2405;
wire n_3995;
wire n_2953;
wire n_2088;
wire n_4036;
wire n_5100;
wire n_1795;
wire n_2578;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_5367;
wire n_2656;
wire n_3524;
wire n_5034;
wire n_1708;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_2092;
wire n_2075;
wire n_3658;
wire n_1776;
wire n_4807;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_1757;
wire n_1919;
wire n_4230;
wire n_3419;
wire n_2053;
wire n_1958;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_1553;
wire n_3678;
wire n_2664;
wire n_3456;
wire n_1808;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_5003;
wire n_5252;
wire n_2731;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_1357;
wire n_3979;
wire n_4582;
wire n_2998;
wire n_4684;
wire n_4840;
wire n_3162;
wire n_2760;
wire n_3377;
wire n_3749;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_5325;
wire n_2637;
wire n_5375;
wire n_4384;
wire n_4423;
wire n_4096;
wire n_2881;
wire n_3282;
wire n_1763;
wire n_3231;
wire n_1966;
wire n_4996;
wire n_2475;
wire n_4598;
wire n_5064;
wire n_4478;
wire n_2646;
wire n_1605;
wire n_5173;
wire n_3920;
wire n_4890;
wire n_5027;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_4106;
wire n_3717;
wire n_2743;
wire n_2675;
wire n_1439;
wire n_3052;
wire n_5215;
wire n_3743;
wire n_1932;
wire n_4721;
wire n_1983;
wire n_4029;
wire n_1594;
wire n_3870;
wire n_4496;
wire n_3529;
wire n_1977;
wire n_2153;
wire n_4338;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_1470;
wire n_2318;
wire n_1735;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_3442;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_5121;
wire n_1824;
wire n_3386;
wire n_1917;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_2446;
wire n_3488;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_4668;
wire n_4953;
wire n_3898;
wire n_1786;
wire n_5284;
wire n_4997;
wire n_5308;
wire n_4274;
wire n_2627;
wire n_4759;
wire n_1413;
wire n_4467;
wire n_2377;
wire n_2080;
wire n_2340;
wire n_3552;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_2361;
wire n_1603;
wire n_1401;
wire n_4113;
wire n_1998;
wire n_4686;
wire n_3759;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_3933;
wire n_3206;
wire n_3966;
wire n_5243;
wire n_1702;
wire n_5221;
wire n_4183;
wire n_4068;
wire n_4872;
wire n_4233;
wire n_3192;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_2649;
wire n_1929;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_3324;
wire n_3914;
wire n_4625;
wire n_2558;
wire n_2063;
wire n_3803;
wire n_3742;
wire n_2252;
wire n_4819;
wire n_1685;
wire n_1714;
wire n_1541;
wire n_2576;
wire n_4900;
wire n_3390;
wire n_1573;
wire n_3746;
wire n_2373;
wire n_1713;
wire n_3817;
wire n_2745;
wire n_1737;
wire n_2493;
wire n_4930;
wire n_5276;
wire n_5078;
wire n_4537;
wire n_2885;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_4282;
wire n_3485;
wire n_4180;
wire n_3839;
wire n_1440;
wire n_5205;
wire n_3333;
wire n_2845;
wire n_4143;
wire n_4659;
wire n_2602;
wire n_4579;
wire n_4616;
wire n_1496;
wire n_3014;
wire n_2547;
wire n_5023;
wire n_1812;
wire n_4105;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_5351;
wire n_3905;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_2401;
wire n_3135;
wire n_2003;
wire n_1457;
wire n_4895;
wire n_3573;
wire n_3148;
wire n_2264;
wire n_3534;
wire n_1482;
wire n_4275;
wire n_3970;
wire n_3438;
wire n_4098;
wire n_1297;
wire n_4789;
wire n_1972;
wire n_2806;
wire n_2184;
wire n_5312;
wire n_3217;
wire n_3425;
wire n_3404;
wire n_5111;
wire n_4055;
wire n_2926;
wire n_3540;
wire n_3670;
wire n_3973;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_5113;
wire n_4442;
wire n_4698;
wire n_1602;
wire n_4779;
wire n_2286;
wire n_4966;
wire n_2065;
wire n_4017;
wire n_3397;
wire n_3740;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1318;
wire n_2977;
wire n_1454;
wire n_3723;
wire n_3600;
wire n_4134;
wire n_1388;
wire n_2836;
wire n_1625;
wire n_2130;
wire n_5167;
wire n_3239;
wire n_5117;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_1452;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_4251;
wire n_1817;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_1326;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_4740;
wire n_5301;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_2221;
wire n_3576;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_4049;
wire n_3862;
wire n_5214;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_4724;
wire n_1772;
wire n_1476;
wire n_2818;
wire n_3646;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_4546;
wire n_3584;
wire n_3756;
wire n_2889;
wire n_5021;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_4382;
wire n_1554;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_5211;
wire n_5230;
wire n_2260;
wire n_5389;
wire n_1813;
wire n_4833;
wire n_3056;
wire n_2345;
wire n_5110;
wire n_1341;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_3289;
wire n_1973;
wire n_2579;
wire n_1770;
wire n_4228;
wire n_4401;
wire n_1756;
wire n_1716;
wire n_2788;
wire n_2984;
wire n_3364;
wire n_1873;
wire n_3201;
wire n_3472;
wire n_2874;
wire n_5179;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_4968;
wire n_5030;
wire n_3949;
wire n_3543;
wire n_3050;
wire n_1478;
wire n_3903;
wire n_4834;
wire n_1364;
wire n_5272;
wire n_2183;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_5361;
wire n_4171;
wire n_4045;
wire n_1367;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_1460;
wire n_2834;
wire n_2531;
wire n_5015;
wire n_2702;
wire n_2030;
wire n_3115;
wire n_4749;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_1404;
wire n_1794;
wire n_2234;
wire n_4804;
wire n_2209;
wire n_4270;
wire n_2797;
wire n_5152;
wire n_2321;
wire n_3680;
wire n_3497;
wire n_1601;
wire n_2940;
wire n_2612;
wire n_1495;
wire n_5128;
wire n_4566;
wire n_2841;
wire n_3322;
wire n_4576;
wire n_2427;
wire n_2505;
wire n_4061;
wire n_3250;
wire n_2070;
wire n_2594;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_5307;
wire n_4767;
wire n_4328;
wire n_3004;
wire n_3112;
wire n_2349;
wire n_1379;
wire n_3874;
wire n_4676;
wire n_4544;
wire n_2170;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_4591;
wire n_3266;
wire n_4646;
wire n_4563;
wire n_4725;
wire n_2210;
wire n_4169;
wire n_5331;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_2426;
wire n_4320;
wire n_5341;
wire n_4881;
wire n_5271;
wire n_5089;
wire n_5263;
wire n_3613;
wire n_3444;
wire n_1505;
wire n_4012;
wire n_4636;
wire n_4584;
wire n_3910;
wire n_4711;
wire n_3319;
wire n_5240;
wire n_3335;
wire n_3413;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_2689;
wire n_3259;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_2010;
wire n_3688;
wire n_3016;
wire n_1693;
wire n_5393;
wire n_2599;
wire n_3338;
wire n_3414;
wire n_1827;
wire n_4671;
wire n_4209;
wire n_1542;
wire n_5041;
wire n_1423;
wire n_1751;
wire n_1508;
wire n_2200;
wire n_3261;
wire n_5026;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_5059;
wire n_3127;
wire n_1780;
wire n_3732;
wire n_4250;
wire n_5329;
wire n_3596;
wire n_4699;
wire n_3906;
wire n_4127;
wire n_3297;
wire n_2683;
wire n_1370;
wire n_1360;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_4202;
wire n_5212;
wire n_5000;
wire n_2853;
wire n_1323;
wire n_3766;
wire n_1353;
wire n_2880;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_4412;
wire n_3407;
wire n_3599;
wire n_3621;
wire n_1580;
wire n_5234;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_1607;
wire n_2538;
wire n_2105;
wire n_5259;
wire n_3163;
wire n_1686;
wire n_3710;
wire n_4155;
wire n_1359;
wire n_2031;
wire n_3891;
wire n_4144;
wire n_2165;
wire n_3379;
wire n_4374;
wire n_3532;
wire n_5131;
wire n_2127;
wire n_1818;
wire n_1576;
wire n_1294;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_4548;
wire n_3258;
wire n_4989;
wire n_4622;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_1845;
wire n_2193;
wire n_2478;
wire n_5140;
wire n_4816;
wire n_1483;
wire n_2983;
wire n_3810;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_5306;
wire n_4483;
wire n_5342;
wire n_2782;
wire n_2672;
wire n_1670;
wire n_2651;
wire n_4358;
wire n_5147;
wire n_3656;
wire n_2071;
wire n_2561;
wire n_2643;
wire n_1374;
wire n_4793;
wire n_4168;
wire n_3446;
wire n_3028;
wire n_4806;
wire n_4350;
wire n_5280;
wire n_1428;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1931;
wire n_4187;
wire n_4166;
wire n_5206;
wire n_3222;
wire n_1801;
wire n_1513;
wire n_2970;
wire n_2235;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_1473;
wire n_3755;
wire n_4258;
wire n_4498;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_5285;
wire n_3563;
wire n_2506;
wire n_4064;
wire n_4936;
wire n_5387;
wire n_1556;
wire n_1863;
wire n_3841;
wire n_2118;
wire n_4770;
wire n_2944;
wire n_2407;
wire n_4907;
wire n_5058;
wire n_3262;
wire n_1450;
wire n_5018;
wire n_4006;
wire n_4861;
wire n_1322;
wire n_3690;
wire n_2358;
wire n_5192;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_2370;
wire n_5159;
wire n_3954;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_5097;
wire n_2750;
wire n_3899;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_4069;
wire n_2784;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_2557;
wire n_5300;
wire n_4850;
wire n_3781;
wire n_4813;
wire n_4912;
wire n_2590;
wire n_2330;
wire n_2942;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_3889;
wire n_4256;
wire n_4224;
wire n_3508;
wire n_4024;
wire n_2218;
wire n_2267;
wire n_2636;
wire n_1951;
wire n_1825;
wire n_1883;
wire n_2759;
wire n_4415;
wire n_4702;
wire n_4252;
wire n_4457;
wire n_5139;
wire n_1393;
wire n_2319;
wire n_3481;
wire n_2808;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_4491;
wire n_2930;
wire n_1838;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_2611;
wire n_4261;
wire n_1660;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_2698;
wire n_5043;
wire n_1662;
wire n_1481;
wire n_4001;
wire n_3047;
wire n_2454;
wire n_4371;
wire n_5281;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_4268;
wire n_5048;
wire n_5028;
wire n_1479;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_4194;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_2990;
wire n_1766;
wire n_1571;
wire n_3119;
wire n_4142;
wire n_4082;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_4260;
wire n_1649;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_3279;
wire n_2621;
wire n_5073;
wire n_5024;
wire n_1537;
wire n_4262;
wire n_2671;
wire n_1798;
wire n_1790;
wire n_4720;
wire n_1647;
wire n_4685;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_1674;
wire n_1830;
wire n_2073;
wire n_4511;
wire n_4014;
wire n_5250;
wire n_3144;
wire n_4757;
wire n_2913;
wire n_2336;
wire n_1615;
wire n_4175;
wire n_2005;
wire n_1916;
wire n_4648;
wire n_1333;
wire n_5006;
wire n_1443;
wire n_1539;
wire n_4892;
wire n_3823;
wire n_1866;
wire n_4173;
wire n_1624;
wire n_4970;
wire n_3816;
wire n_4108;
wire n_4486;
wire n_2960;
wire n_4627;
wire n_2290;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_2145;
wire n_1639;
wire n_3030;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_5163;
wire n_2039;
wire n_4961;
wire n_3753;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_5190;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_1362;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_3396;
wire n_1445;
wire n_4023;
wire n_4420;
wire n_1923;
wire n_5138;
wire n_5374;
wire n_2116;
wire n_1434;
wire n_1828;
wire n_2320;
wire n_5349;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_4640;
wire n_2583;
wire n_4396;
wire n_5127;
wire n_4367;
wire n_2087;
wire n_5216;
wire n_1989;
wire n_3818;
wire n_2523;
wire n_4387;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_1578;
wire n_3719;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_4308;
wire n_2812;
wire n_2355;
wire n_2133;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_2725;
wire n_5175;
wire n_3883;
wire n_1355;
wire n_2565;
wire n_4152;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_3466;
wire n_4962;
wire n_2595;
wire n_3411;
wire n_4958;
wire n_4271;
wire n_5171;
wire n_3586;
wire n_1390;
wire n_4071;
wire n_4921;
wire n_1980;
wire n_3065;
wire n_4361;
wire n_4614;
wire n_2681;
wire n_3103;
wire n_4945;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_1651;
wire n_2775;
wire n_4693;
wire n_4326;
wire n_3557;
wire n_2230;
wire n_5383;
wire n_4744;
wire n_2851;
wire n_4305;
wire n_1455;
wire n_2490;
wire n_1407;
wire n_4213;
wire n_2849;
wire n_3692;
wire n_2204;
wire n_4929;
wire n_1961;
wire n_4964;
wire n_1430;
wire n_4802;
wire n_1354;
wire n_4139;
wire n_3029;
wire n_2508;
wire n_4031;
wire n_2416;
wire n_3881;
wire n_2461;
wire n_2243;
wire n_4583;
wire n_4210;
wire n_5245;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_1611;
wire n_2368;
wire n_2890;
wire n_2554;
wire n_3698;
wire n_3927;
wire n_1840;
wire n_4540;
wire n_3961;
wire n_1630;
wire n_4891;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_3993;
wire n_4940;
wire n_5208;
wire n_3588;
wire n_2308;
wire n_4590;
wire n_4830;
wire n_5231;
wire n_5237;
wire n_4664;
wire n_3860;
wire n_3160;
wire n_2191;
wire n_5093;
wire n_2428;
wire n_3847;
wire n_4946;
wire n_1346;
wire n_4906;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_5390;
wire n_5347;
wire n_2824;
wire n_3033;
wire n_3298;
wire n_2440;
wire n_4883;
wire n_1386;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_2333;
wire n_2916;
wire n_4297;
wire n_1632;
wire n_3800;
wire n_2403;
wire n_4608;
wire n_5232;
wire n_2792;
wire n_2870;
wire n_3991;
wire n_3134;
wire n_4172;
wire n_4791;
wire n_4536;
wire n_5149;
wire n_2463;
wire n_5151;
wire n_4773;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_2472;
wire n_4611;
wire n_4755;
wire n_1768;
wire n_2294;
wire n_4960;
wire n_2993;
wire n_1719;
wire n_3864;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2309;
wire n_2948;
wire n_1560;
wire n_4362;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_4422;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_3482;
wire n_2233;
wire n_1312;
wire n_4555;
wire n_2827;
wire n_5136;
wire n_5228;
wire n_1504;
wire n_3956;
wire n_5323;
wire n_3572;
wire n_4215;
wire n_4280;
wire n_3375;
wire n_4047;
wire n_2082;
wire n_1643;
wire n_3167;
wire n_5350;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_5338;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3854;
wire n_2468;
wire n_1610;
wire n_1422;
wire n_3078;
wire n_3253;
wire n_4027;
wire n_2280;
wire n_4599;
wire n_3363;
wire n_4812;
wire n_1511;
wire n_3689;
wire n_2020;
wire n_4628;
wire n_1881;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_3950;
wire n_4458;
wire n_4121;
wire n_1616;
wire n_5090;
wire n_4476;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_2303;
wire n_2810;
wire n_2747;
wire n_1848;
wire n_2126;
wire n_4573;
wire n_5289;
wire n_4118;
wire n_4803;
wire n_4079;
wire n_4091;
wire n_1638;
wire n_2002;
wire n_5145;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_5132;
wire n_5191;
wire n_3085;
wire n_1655;
wire n_5359;
wire n_2574;
wire n_5293;
wire n_1358;
wire n_4316;
wire n_3697;
wire n_2638;
wire n_4044;
wire n_4062;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_2711;
wire n_5363;
wire n_5200;
wire n_1653;
wire n_1506;
wire n_2867;
wire n_1894;
wire n_2794;
wire n_3145;
wire n_3124;
wire n_4253;
wire n_5356;
wire n_5369;
wire n_2608;
wire n_5258;
wire n_2657;
wire n_5255;
wire n_2852;
wire n_2392;
wire n_3517;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_1834;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_5080;
wire n_1516;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_2409;
wire n_3402;
wire n_5295;
wire n_4679;
wire n_4115;
wire n_4998;
wire n_2988;
wire n_1731;
wire n_1970;
wire n_2766;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_2205;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_1912;
wire n_3401;
wire n_3226;
wire n_1410;
wire n_3902;
wire n_4730;
wire n_2779;
wire n_1584;
wire n_3654;
wire n_2164;
wire n_2115;
wire n_2232;
wire n_5327;
wire n_1302;
wire n_1774;
wire n_4713;
wire n_5137;
wire n_2811;
wire n_3348;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_4204;
wire n_5098;
wire n_1543;
wire n_2224;
wire n_1991;
wire n_4743;
wire n_3805;
wire n_3825;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_2692;
wire n_2008;
wire n_4654;
wire n_4733;
wire n_3792;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_1753;
wire n_2283;
wire n_3278;
wire n_1689;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_3312;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_5069;
wire n_3285;
wire n_3968;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_2480;
wire n_2363;
wire n_4072;
wire n_4781;
wire n_3606;
wire n_5004;
wire n_2550;
wire n_4424;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_3878;
wire n_4450;
wire n_3553;
wire n_4746;
wire n_1683;
wire n_1530;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_1409;
wire n_3850;
wire n_4459;
wire n_2996;
wire n_1320;
wire n_4050;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_2102;
wire n_4853;
wire n_2422;
wire n_2239;
wire n_5256;
wire n_2950;
wire n_5220;
wire n_3852;
wire n_5178;
wire n_4520;
wire n_2057;
wire n_4008;
wire n_5077;
wire n_3858;
wire n_1901;
wire n_4502;
wire n_3032;
wire n_4851;
wire n_1330;
wire n_3072;
wire n_3081;
wire n_3313;
wire n_2710;
wire n_1745;
wire n_3924;
wire n_4571;
wire n_2006;
wire n_5314;
wire n_1618;
wire n_2343;
wire n_3439;
wire n_5049;
wire n_2535;
wire n_4205;
wire n_2726;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_2799;
wire n_4454;
wire n_4229;
wire n_4739;
wire n_2376;
wire n_3017;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_4879;
wire n_5051;
wire n_3926;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2854;
wire n_1701;
wire n_4181;
wire n_1550;
wire n_2764;
wire n_1498;
wire n_4225;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_1648;
wire n_4153;
wire n_5156;
wire n_3627;
wire n_4300;
wire n_3551;
wire n_1769;
wire n_4783;
wire n_2964;
wire n_3769;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_2442;
wire n_1943;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_3351;
wire n_3527;
wire n_1396;
wire n_1348;
wire n_2883;
wire n_1752;
wire n_4182;
wire n_2912;
wire n_1315;
wire n_4825;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_5120;
wire n_4565;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_4839;
wire n_5222;
wire n_4016;
wire n_3435;
wire n_3575;
wire n_1546;
wire n_4231;
wire n_3165;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_4083;
wire n_1937;
wire n_4461;
wire n_3234;
wire n_5392;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3916;
wire n_2569;
wire n_3556;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3024;
wire n_3512;
wire n_4939;
wire n_5169;
wire n_4389;
wire n_3930;
wire n_4448;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_2503;
wire n_1540;
wire n_1936;
wire n_2027;
wire n_2642;
wire n_2500;
wire n_1918;
wire n_4831;
wire n_2513;
wire n_2695;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_2414;
wire n_1402;
wire n_3662;
wire n_4319;
wire n_2229;
wire n_1397;
wire n_4596;
wire n_2004;
wire n_3694;
wire n_2586;
wire n_4726;
wire n_1398;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_4119;
wire n_3799;
wire n_4298;
wire n_5201;
wire n_4474;
wire n_5217;
wire n_2511;
wire n_1681;
wire n_3383;
wire n_3585;
wire n_2975;
wire n_5029;
wire n_2704;
wire n_4214;
wire n_5158;
wire n_4884;
wire n_4366;
wire n_4009;
wire n_4580;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_1859;
wire n_1677;
wire n_2955;
wire n_4112;
wire n_4337;
wire n_4138;
wire n_5396;
wire n_1528;
wire n_5335;
wire n_1292;
wire n_2520;
wire n_2134;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_1347;
wire n_5143;
wire n_4238;
wire n_1451;
wire n_2374;
wire n_1545;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_2396;
wire n_1799;
wire n_4734;
wire n_1939;
wire n_2486;
wire n_4635;
wire n_3501;
wire n_1869;
wire n_4013;
wire n_3039;
wire n_2011;
wire n_4242;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_3036;
wire n_1896;
wire n_3180;
wire n_5283;
wire n_5268;
wire n_1705;
wire n_4561;
wire n_2639;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_5122;
wire n_3186;
wire n_4955;
wire n_4501;
wire n_3696;
wire n_3650;
wire n_2761;
wire n_3157;
wire n_2537;
wire n_2144;
wire n_2515;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_1949;
wire n_2936;
wire n_1946;
wire n_1484;
wire n_1328;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_4369;
wire n_5378;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_1831;
wire n_1598;
wire n_4394;
wire n_1850;
wire n_1749;
wire n_3101;
wire n_3669;
wire n_5278;
wire n_2663;
wire n_1394;
wire n_2693;
wire n_3798;
wire n_4065;
wire n_5187;
wire n_4944;
wire n_2180;
wire n_2249;
wire n_4135;
wire n_2632;
wire n_1547;
wire n_1755;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_2915;
wire n_2300;
wire n_3291;
wire n_4716;
wire n_4942;
wire n_2432;
wire n_1521;
wire n_3405;
wire n_4745;
wire n_2337;
wire n_1384;
wire n_3907;
wire n_5344;
wire n_4629;
wire n_2932;
wire n_2980;
wire n_5225;
wire n_3306;
wire n_1784;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1986;
wire n_1471;
wire n_4752;
wire n_5265;
wire n_1750;
wire n_1459;
wire n_3986;
wire n_4376;
wire n_4753;
wire n_4552;
wire n_3885;
wire n_2713;
wire n_5196;
wire n_5181;
wire n_2644;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_5126;
wire n_2214;
wire n_3427;
wire n_2055;
wire n_4067;
wire n_1403;
wire n_4042;
wire n_4176;
wire n_4385;
wire n_3320;
wire n_5009;
wire n_2688;
wire n_5368;
wire n_1463;
wire n_3651;
wire n_4333;
wire n_3359;
wire n_2865;
wire n_2706;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_4815;
wire n_4246;
wire n_3580;
wire n_2139;
wire n_4609;
wire n_5291;
wire n_5114;
wire n_2674;
wire n_1565;
wire n_4088;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_4462;
wire n_4472;
wire n_3433;
wire n_5288;
wire n_2305;
wire n_2450;
wire n_3447;
wire n_3305;
wire n_4151;
wire n_4148;
wire n_1712;
wire n_3528;
wire n_4373;
wire n_4934;
wire n_5218;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_4630;
wire n_4643;
wire n_4331;
wire n_3989;
wire n_4475;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_1775;
wire n_3296;
wire n_1368;
wire n_2762;
wire n_4683;
wire n_5366;
wire n_1847;
wire n_2767;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_3602;
wire n_2967;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_3923;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_1544;
wire n_5086;
wire n_1629;
wire n_2801;
wire n_4011;
wire n_4905;
wire n_2763;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_1997;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_4278;
wire n_1635;
wire n_4623;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_2215;
wire n_5053;
wire n_4553;
wire n_3978;
wire n_4809;
wire n_5226;
wire n_1925;
wire n_3660;
wire n_1815;
wire n_2491;
wire n_1788;
wire n_5079;
wire n_3833;
wire n_1679;
wire n_4841;
wire n_2022;
wire n_3814;
wire n_1415;
wire n_2592;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_3513;
wire n_3133;
wire n_4645;
wire n_2992;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_2517;
wire n_3128;
wire n_2631;
wire n_2178;
wire n_1767;
wire n_1529;
wire n_2469;
wire n_3355;
wire n_2007;
wire n_3917;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_3000;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_1839;
wire n_1837;
wire n_4557;
wire n_5248;
wire n_4451;
wire n_2875;
wire n_1500;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_3471;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_1656;
wire n_3564;
wire n_3988;
wire n_3457;
wire n_1678;
wire n_4324;
wire n_4821;
wire n_1871;
wire n_3630;
wire n_3271;
wire n_4771;
wire n_4086;
wire n_2412;
wire n_4814;
wire n_1781;
wire n_2084;
wire n_3648;
wire n_3075;
wire n_3173;
wire n_5332;
wire n_5108;
wire n_4692;
wire n_3031;
wire n_3701;
wire n_1773;
wire n_3243;
wire n_2666;
wire n_3385;
wire n_2171;
wire n_4708;
wire n_2768;
wire n_2314;
wire n_4826;
wire n_2420;
wire n_3343;
wire n_1593;
wire n_3767;
wire n_2299;
wire n_2873;
wire n_2540;
wire n_4589;
wire n_5057;
wire n_4578;
wire n_1640;
wire n_2162;
wire n_2847;
wire n_2051;
wire n_3221;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_2359;
wire n_3674;
wire n_5286;
wire n_3502;
wire n_3098;
wire n_1383;
wire n_5013;
wire n_2312;
wire n_3015;
wire n_1920;
wire n_4147;
wire n_2048;
wire n_3607;
wire n_4925;
wire n_1921;
wire n_1309;
wire n_4974;
wire n_1800;
wire n_1548;
wire n_4932;
wire n_1421;
wire n_4510;
wire n_2571;
wire n_3276;
wire n_3787;
wire n_5119;
wire n_2124;
wire n_3827;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_4447;
wire n_4285;
wire n_4651;
wire n_4818;
wire n_4514;
wire n_1366;
wire n_4800;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_1568;
wire n_2110;
wire n_1332;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_1591;
wire n_2033;
wire n_4341;
wire n_1682;
wire n_4312;
wire n_2628;
wire n_3399;
wire n_2132;
wire n_2400;
wire n_4633;
wire n_3838;
wire n_1909;
wire n_4277;
wire n_4140;
wire n_3675;
wire n_5092;
wire n_3387;
wire n_5186;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_2831;
wire n_1456;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_4832;
wire n_4207;
wire n_4545;
wire n_3037;
wire n_4868;
wire n_1885;
wire n_2452;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_5238;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_1849;
wire n_5054;
wire n_2467;
wire n_2288;
wire n_4063;
wire n_3592;
wire n_4650;
wire n_4888;
wire n_5326;
wire n_1435;
wire n_3394;
wire n_4874;
wire n_3793;
wire n_4669;
wire n_4339;
wire n_1645;
wire n_4041;
wire n_2858;
wire n_4060;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_2128;
wire n_3097;
wire n_5391;
wire n_4541;
wire n_3824;
wire n_3388;
wire n_5267;
wire n_4494;
wire n_3059;
wire n_3465;
wire n_1316;
wire n_4796;
wire n_1438;
wire n_3589;
wire n_2534;
wire n_4799;
wire n_5153;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_2789;
wire n_4775;
wire n_2216;
wire n_5044;
wire n_1897;
wire n_1424;
wire n_5365;
wire n_2933;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_5354;
wire n_4455;
wire n_2328;
wire n_4248;
wire n_4754;
wire n_4554;
wire n_4845;
wire n_3053;
wire n_1299;
wire n_3893;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_1699;
wire n_3334;
wire n_2541;
wire n_4383;
wire n_1432;
wire n_3875;
wire n_5370;
wire n_4003;
wire n_5372;
wire n_5299;
wire n_2402;
wire n_4301;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_1844;
wire n_3777;
wire n_4784;
wire n_2999;
wire n_1644;
wire n_5082;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_5209;
wire n_3080;
wire n_4199;
wire n_2701;
wire n_3362;
wire n_1631;
wire n_3105;
wire n_4286;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_4470;
wire n_2236;
wire n_2816;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3664;
wire n_4188;
wire n_1668;
wire n_3913;
wire n_3417;
wire n_1579;
wire n_4034;
wire n_1688;
wire n_3327;
wire n_5275;
wire n_4689;
wire n_5071;
wire n_3067;
wire n_2755;
wire n_3237;
wire n_1992;
wire n_4402;
wire n_4239;
wire n_3400;
wire n_4550;
wire n_1400;
wire n_1342;
wire n_3382;
wire n_3574;
wire n_5227;
wire n_2169;
wire n_1557;
wire n_4201;
wire n_3316;
wire n_5242;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_1730;
wire n_3603;
wire n_4123;
wire n_2192;
wire n_3633;
wire n_4479;
wire n_1373;
wire n_2670;
wire n_1646;
wire n_1307;
wire n_4416;
wire n_3372;
wire n_4539;
wire n_2707;
wire n_2471;
wire n_1472;
wire n_1671;
wire n_3230;
wire n_3342;
wire n_4682;
wire n_5353;
wire n_3708;
wire n_5294;
wire n_3729;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_3861;
wire n_4736;
wire n_3780;
wire n_1928;
wire n_5244;
wire n_5382;
wire n_3957;
wire n_5274;
wire n_3848;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_5384;
wire n_3608;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_2352;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_2619;
wire n_2444;
wire n_3123;
wire n_5056;
wire n_5249;
wire n_3393;
wire n_5198;
wire n_5360;
wire n_5233;
wire n_4887;
wire n_4617;
wire n_5269;
wire n_3520;
wire n_2492;
wire n_4005;
wire n_1687;
wire n_1637;
wire n_4904;
wire n_1419;
wire n_4792;
wire n_3578;
wire n_3812;
wire n_1886;
wire n_1389;
wire n_4980;
wire n_1465;
wire n_4290;
wire n_5247;
wire n_1375;
wire n_3727;
wire n_5317;
wire n_3774;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_1597;
wire n_1659;
wire n_2431;
wire n_1371;
wire n_4956;
wire n_5380;
wire n_2206;
wire n_3182;
wire n_2564;
wire n_4947;
wire n_4656;
wire n_3896;
wire n_3958;
wire n_3450;
wire n_4729;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_2000;
wire n_2074;
wire n_3174;
wire n_1453;
wire n_2217;
wire n_3398;
wire n_2307;
wire n_3408;
wire n_2722;
wire n_5388;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_1628;
wire n_3432;
wire n_1514;
wire n_1771;
wire n_3090;
wire n_2437;
wire n_3762;
wire n_2445;
wire n_1427;
wire n_1835;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_4529;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_3972;
wire n_3308;
wire n_1533;
wire n_5036;
wire n_4772;
wire n_3467;
wire n_4322;
wire n_1720;
wire n_2830;
wire n_4354;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_5273;
wire n_4677;
wire n_3901;
wire n_1480;
wire n_5261;
wire n_3757;
wire n_3381;
wire n_5193;
wire n_2245;
wire n_1782;
wire n_4909;
wire n_1524;
wire n_1485;
wire n_2965;
wire n_3635;
wire n_5022;
wire n_5005;
wire n_2814;
wire n_1570;
wire n_3882;
wire n_3046;
wire n_2213;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_4634;
wire n_3337;
wire n_2527;
wire n_1461;
wire n_3204;
wire n_2136;
wire n_5174;
wire n_1822;
wire n_4952;
wire n_5157;
wire n_3005;
wire n_4380;
wire n_3129;
wire n_4126;
wire n_1783;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_4880;
wire n_1907;
wire n_2686;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_1417;
wire n_1295;
wire n_5061;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_2187;
wire n_1762;
wire n_3023;
wire n_4193;
wire n_4075;
wire n_3104;
wire n_4737;
wire n_3647;
wire n_2819;
wire n_5195;
wire n_3609;
wire n_4136;
wire n_1715;
wire n_1952;
wire n_4393;
wire n_3720;
wire n_4535;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_4794;
wire n_3959;
wire n_3140;
wire n_5246;
wire n_3724;
wire n_2104;
wire n_3011;
wire n_5164;
wire n_4196;
wire n_1425;
wire n_4592;
wire n_4675;
wire n_5340;
wire n_3069;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_5183;
wire n_3084;
wire n_1727;
wire n_2735;
wire n_2497;
wire n_3412;
wire n_1995;
wire n_2411;
wire n_3761;
wire n_4889;
wire n_2014;
wire n_2986;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_4828;
wire n_5385;
wire n_4558;
wire n_2172;
wire n_4722;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_2250;
wire n_4092;
wire n_3908;
wire n_2423;
wire n_3671;
wire n_3344;
wire n_2194;
wire n_4465;
wire n_3302;
wire n_5304;
wire n_2680;
wire n_5130;
wire n_1567;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_3842;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_1797;
wire n_2957;
wire n_2357;
wire n_3309;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_1589;
wire n_4116;
wire n_2570;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_3754;
wire n_4612;
wire n_1469;
wire n_2744;
wire n_4287;
wire n_2397;
wire n_2208;
wire n_3063;
wire n_5177;
wire n_3617;
wire n_1298;
wire n_1652;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_1676;
wire n_2591;
wire n_3384;
wire n_4602;
wire n_5172;
wire n_4449;
wire n_1864;
wire n_5070;
wire n_1337;
wire n_4445;
wire n_1627;
wire n_4870;
wire n_2438;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_3181;
wire n_2278;
wire n_4915;
wire n_5296;
wire n_2135;
wire n_3493;
wire n_5313;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_2823;
wire n_1408;
wire n_1761;
wire n_5270;
wire n_4345;
wire n_5188;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_1694;
wire n_4318;
wire n_2485;
wire n_2655;
wire n_4185;
wire n_4797;
wire n_2366;
wire n_1526;
wire n_3997;
wire n_1604;
wire n_4032;
wire n_1764;
wire n_3582;
wire n_1583;
wire n_2826;
wire n_3539;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_4124;
wire n_4492;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_4245;
wire n_4364;
wire n_4928;
wire n_2225;
wire n_1507;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3853;
wire n_4216;
wire n_2019;
wire n_1340;
wire n_1558;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_1704;
wire n_3721;
wire n_2026;
wire n_2109;
wire n_2013;
wire n_1990;
wire n_2614;
wire n_2991;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_3473;
wire n_4560;
wire n_5318;
wire n_2839;
wire n_1588;
wire n_5395;
wire n_2237;
wire n_3463;
wire n_3699;
wire n_5067;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_2728;
wire n_3857;

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_154),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1134),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1061),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_25),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1266),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1261),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1271),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_92),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_1187),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_547),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_132),
.Y(n_1302)
);

CKINVDCx16_ASAP7_75t_R g1303 ( 
.A(n_115),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_613),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_561),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_459),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_901),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1265),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_136),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1181),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_143),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_629),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1252),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_75),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_86),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_868),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_314),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_618),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_464),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_533),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_32),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_30),
.Y(n_1322)
);

CKINVDCx20_ASAP7_75t_R g1323 ( 
.A(n_575),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_159),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_9),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_341),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1188),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1280),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_81),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1075),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_761),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_701),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_54),
.Y(n_1333)
);

BUFx6f_ASAP7_75t_L g1334 ( 
.A(n_1167),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_997),
.Y(n_1335)
);

INVxp67_ASAP7_75t_L g1336 ( 
.A(n_1277),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1173),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1151),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1208),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_53),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_431),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_485),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1286),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1288),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_916),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1228),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_486),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_54),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1198),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_119),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_336),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1098),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_508),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1170),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_427),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_1064),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_795),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_517),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1206),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_746),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1149),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_291),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_989),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1060),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_715),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1140),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_854),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_758),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_318),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_320),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_770),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1178),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_265),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_907),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_361),
.Y(n_1375)
);

INVx1_ASAP7_75t_SL g1376 ( 
.A(n_1087),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_251),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1027),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1229),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_2),
.Y(n_1380)
);

BUFx10_ASAP7_75t_L g1381 ( 
.A(n_157),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_367),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_479),
.Y(n_1383)
);

BUFx5_ASAP7_75t_L g1384 ( 
.A(n_1204),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1090),
.Y(n_1385)
);

BUFx10_ASAP7_75t_L g1386 ( 
.A(n_99),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1033),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_469),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_818),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1041),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_852),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1285),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_1150),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1182),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1289),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1012),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_729),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1256),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_294),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_769),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_156),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_452),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_884),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_311),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_742),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_896),
.Y(n_1406)
);

CKINVDCx20_ASAP7_75t_R g1407 ( 
.A(n_496),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1011),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1185),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_1146),
.Y(n_1410)
);

BUFx2_ASAP7_75t_L g1411 ( 
.A(n_375),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_124),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1032),
.Y(n_1413)
);

INVx2_ASAP7_75t_SL g1414 ( 
.A(n_832),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_191),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_899),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1046),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_368),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1023),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_808),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_308),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_304),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_97),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1093),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_907),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_982),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_647),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_543),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1239),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1209),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1074),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1177),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_822),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_284),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_576),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_757),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_157),
.Y(n_1437)
);

CKINVDCx16_ASAP7_75t_R g1438 ( 
.A(n_563),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_644),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_28),
.Y(n_1440)
);

CKINVDCx14_ASAP7_75t_R g1441 ( 
.A(n_27),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_631),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_867),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1153),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_966),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_707),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1222),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1245),
.Y(n_1448)
);

BUFx10_ASAP7_75t_L g1449 ( 
.A(n_541),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_703),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_198),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1136),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1219),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_109),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_626),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_1238),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_561),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_244),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1031),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_120),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_1038),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_361),
.Y(n_1462)
);

INVx1_ASAP7_75t_SL g1463 ( 
.A(n_1127),
.Y(n_1463)
);

CKINVDCx20_ASAP7_75t_R g1464 ( 
.A(n_263),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_483),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1179),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_420),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_792),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_694),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_94),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_474),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_581),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_697),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_198),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1133),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_476),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1069),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_1210),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_521),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1013),
.Y(n_1480)
);

CKINVDCx20_ASAP7_75t_R g1481 ( 
.A(n_851),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_674),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1251),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_287),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_38),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_15),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_976),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1202),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_736),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_26),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_564),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_591),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1043),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_759),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_634),
.Y(n_1495)
);

CKINVDCx20_ASAP7_75t_R g1496 ( 
.A(n_1040),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_630),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_490),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1207),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_60),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_472),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_114),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1094),
.Y(n_1503)
);

INVxp67_ASAP7_75t_L g1504 ( 
.A(n_123),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1247),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_1165),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_248),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_816),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_865),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1290),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_115),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1272),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1104),
.Y(n_1513)
);

CKINVDCx12_ASAP7_75t_R g1514 ( 
.A(n_981),
.Y(n_1514)
);

CKINVDCx16_ASAP7_75t_R g1515 ( 
.A(n_1131),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_422),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_134),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1034),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_274),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_825),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1049),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_702),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_882),
.Y(n_1523)
);

CKINVDCx20_ASAP7_75t_R g1524 ( 
.A(n_1291),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1257),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1066),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_792),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_670),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_558),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_476),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_730),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_312),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_58),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_279),
.Y(n_1534)
);

BUFx10_ASAP7_75t_L g1535 ( 
.A(n_105),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1108),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1020),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_788),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_247),
.Y(n_1539)
);

CKINVDCx20_ASAP7_75t_R g1540 ( 
.A(n_41),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_326),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_337),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_797),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_734),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_371),
.Y(n_1545)
);

BUFx10_ASAP7_75t_L g1546 ( 
.A(n_971),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_97),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1112),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_821),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_100),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_170),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1044),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1139),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_959),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_832),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_296),
.Y(n_1556)
);

CKINVDCx20_ASAP7_75t_R g1557 ( 
.A(n_1194),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_175),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_866),
.Y(n_1559)
);

CKINVDCx20_ASAP7_75t_R g1560 ( 
.A(n_8),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_885),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1154),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_744),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_804),
.Y(n_1564)
);

CKINVDCx20_ASAP7_75t_R g1565 ( 
.A(n_1255),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_99),
.Y(n_1566)
);

INVx4_ASAP7_75t_R g1567 ( 
.A(n_1218),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1160),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_270),
.Y(n_1569)
);

CKINVDCx20_ASAP7_75t_R g1570 ( 
.A(n_1054),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1235),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_335),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_337),
.Y(n_1573)
);

CKINVDCx20_ASAP7_75t_R g1574 ( 
.A(n_1230),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_861),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_868),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_631),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_16),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_1262),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_571),
.Y(n_1580)
);

CKINVDCx20_ASAP7_75t_R g1581 ( 
.A(n_860),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_100),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_479),
.Y(n_1583)
);

BUFx10_ASAP7_75t_L g1584 ( 
.A(n_1138),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_233),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_766),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_415),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_646),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_758),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1225),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1163),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_843),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_893),
.Y(n_1593)
);

CKINVDCx20_ASAP7_75t_R g1594 ( 
.A(n_931),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_10),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_784),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1282),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_863),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1115),
.Y(n_1599)
);

CKINVDCx20_ASAP7_75t_R g1600 ( 
.A(n_1172),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1215),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_203),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_429),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_623),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1279),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_638),
.Y(n_1606)
);

BUFx5_ASAP7_75t_L g1607 ( 
.A(n_641),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_924),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_78),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_123),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_1162),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_710),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_710),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_946),
.Y(n_1614)
);

CKINVDCx14_ASAP7_75t_R g1615 ( 
.A(n_624),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1236),
.Y(n_1616)
);

BUFx6f_ASAP7_75t_L g1617 ( 
.A(n_1007),
.Y(n_1617)
);

BUFx3_ASAP7_75t_L g1618 ( 
.A(n_518),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1056),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1055),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_195),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1158),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1070),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_86),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_114),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_78),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_833),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_209),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_315),
.Y(n_1629)
);

CKINVDCx20_ASAP7_75t_R g1630 ( 
.A(n_926),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1086),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1145),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_1258),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_766),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_108),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1111),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1184),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_176),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1101),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_987),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1242),
.Y(n_1641)
);

CKINVDCx20_ASAP7_75t_R g1642 ( 
.A(n_599),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1095),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_449),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_397),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_1237),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_828),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1176),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_1232),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_24),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_632),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_893),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_268),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_460),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_328),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1244),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1144),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_151),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1067),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1049),
.Y(n_1660)
);

CKINVDCx20_ASAP7_75t_R g1661 ( 
.A(n_1114),
.Y(n_1661)
);

INVx1_ASAP7_75t_SL g1662 ( 
.A(n_1032),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_186),
.Y(n_1663)
);

CKINVDCx20_ASAP7_75t_R g1664 ( 
.A(n_1201),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_113),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1224),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_134),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_878),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1231),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_289),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1100),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_518),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1039),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_548),
.Y(n_1674)
);

BUFx10_ASAP7_75t_L g1675 ( 
.A(n_1017),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1260),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1141),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_843),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_418),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_357),
.Y(n_1680)
);

CKINVDCx20_ASAP7_75t_R g1681 ( 
.A(n_1122),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_1096),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1099),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_1227),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_194),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_128),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_188),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_587),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_1267),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1259),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_52),
.Y(n_1691)
);

BUFx10_ASAP7_75t_L g1692 ( 
.A(n_151),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1156),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1082),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_987),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_806),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_906),
.Y(n_1697)
);

CKINVDCx20_ASAP7_75t_R g1698 ( 
.A(n_800),
.Y(n_1698)
);

CKINVDCx20_ASAP7_75t_R g1699 ( 
.A(n_1166),
.Y(n_1699)
);

INVx2_ASAP7_75t_SL g1700 ( 
.A(n_1246),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1161),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_31),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_109),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_636),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_1221),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_1155),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_37),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_213),
.Y(n_1708)
);

CKINVDCx20_ASAP7_75t_R g1709 ( 
.A(n_1169),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_1103),
.Y(n_1710)
);

CKINVDCx20_ASAP7_75t_R g1711 ( 
.A(n_202),
.Y(n_1711)
);

CKINVDCx20_ASAP7_75t_R g1712 ( 
.A(n_1022),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_236),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_434),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_1053),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_84),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1211),
.Y(n_1717)
);

CKINVDCx20_ASAP7_75t_R g1718 ( 
.A(n_324),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1043),
.Y(n_1719)
);

INVx2_ASAP7_75t_SL g1720 ( 
.A(n_1287),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_464),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_511),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_231),
.Y(n_1724)
);

BUFx6f_ASAP7_75t_L g1725 ( 
.A(n_976),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_281),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_89),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_789),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1041),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_807),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_395),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_47),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_142),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_818),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1026),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_887),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_849),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1183),
.Y(n_1738)
);

BUFx10_ASAP7_75t_L g1739 ( 
.A(n_615),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1046),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_470),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_686),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_236),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1106),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_636),
.Y(n_1745)
);

CKINVDCx20_ASAP7_75t_R g1746 ( 
.A(n_1234),
.Y(n_1746)
);

CKINVDCx20_ASAP7_75t_R g1747 ( 
.A(n_994),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_1189),
.Y(n_1748)
);

INVx1_ASAP7_75t_SL g1749 ( 
.A(n_848),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_199),
.Y(n_1750)
);

BUFx6f_ASAP7_75t_L g1751 ( 
.A(n_1152),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_716),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_483),
.Y(n_1753)
);

BUFx2_ASAP7_75t_L g1754 ( 
.A(n_486),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_471),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1058),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1056),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_174),
.Y(n_1758)
);

CKINVDCx16_ASAP7_75t_R g1759 ( 
.A(n_1030),
.Y(n_1759)
);

INVx2_ASAP7_75t_SL g1760 ( 
.A(n_1269),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_77),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1196),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_747),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_89),
.Y(n_1764)
);

CKINVDCx20_ASAP7_75t_R g1765 ( 
.A(n_1171),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1199),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1175),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_993),
.Y(n_1768)
);

CKINVDCx20_ASAP7_75t_R g1769 ( 
.A(n_1159),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1024),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1016),
.Y(n_1771)
);

INVx2_ASAP7_75t_SL g1772 ( 
.A(n_1195),
.Y(n_1772)
);

INVxp33_ASAP7_75t_SL g1773 ( 
.A(n_64),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1135),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1214),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1012),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_1121),
.Y(n_1777)
);

CKINVDCx20_ASAP7_75t_R g1778 ( 
.A(n_630),
.Y(n_1778)
);

BUFx6f_ASAP7_75t_L g1779 ( 
.A(n_16),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_1281),
.Y(n_1780)
);

INVx1_ASAP7_75t_SL g1781 ( 
.A(n_355),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1035),
.Y(n_1782)
);

INVx2_ASAP7_75t_SL g1783 ( 
.A(n_428),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_632),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1097),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1042),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_1142),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_390),
.Y(n_1788)
);

CKINVDCx16_ASAP7_75t_R g1789 ( 
.A(n_102),
.Y(n_1789)
);

INVx2_ASAP7_75t_SL g1790 ( 
.A(n_540),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_1072),
.Y(n_1791)
);

CKINVDCx20_ASAP7_75t_R g1792 ( 
.A(n_365),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1096),
.Y(n_1793)
);

BUFx2_ASAP7_75t_SL g1794 ( 
.A(n_682),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_110),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_516),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_939),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1050),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1029),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_246),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_431),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_437),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1078),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1197),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1061),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_311),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_498),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1190),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_814),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1168),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_412),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1028),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_90),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1212),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_234),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1091),
.Y(n_1816)
);

INVxp67_ASAP7_75t_L g1817 ( 
.A(n_773),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_957),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_684),
.Y(n_1819)
);

INVx1_ASAP7_75t_SL g1820 ( 
.A(n_831),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_506),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_58),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1193),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_700),
.Y(n_1824)
);

INVx1_ASAP7_75t_SL g1825 ( 
.A(n_427),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_7),
.Y(n_1826)
);

CKINVDCx16_ASAP7_75t_R g1827 ( 
.A(n_23),
.Y(n_1827)
);

INVx1_ASAP7_75t_SL g1828 ( 
.A(n_396),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1248),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1243),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_75),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_839),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_576),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_936),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1233),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_968),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1015),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1270),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_456),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_654),
.Y(n_1840)
);

BUFx8_ASAP7_75t_SL g1841 ( 
.A(n_120),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_611),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_1223),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_793),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_514),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1217),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1253),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1078),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_1079),
.Y(n_1849)
);

BUFx2_ASAP7_75t_L g1850 ( 
.A(n_1057),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_1068),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_1110),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1284),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_321),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_1254),
.Y(n_1855)
);

INVx2_ASAP7_75t_SL g1856 ( 
.A(n_1113),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_988),
.Y(n_1857)
);

BUFx3_ASAP7_75t_L g1858 ( 
.A(n_88),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_637),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_153),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_713),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_673),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1164),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_451),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_743),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1278),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1105),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_1025),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_666),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_571),
.Y(n_1870)
);

CKINVDCx20_ASAP7_75t_R g1871 ( 
.A(n_175),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_709),
.Y(n_1872)
);

INVx1_ASAP7_75t_SL g1873 ( 
.A(n_1018),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_380),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_819),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_344),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1105),
.Y(n_1877)
);

BUFx3_ASAP7_75t_L g1878 ( 
.A(n_340),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_1077),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1240),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_755),
.Y(n_1881)
);

CKINVDCx20_ASAP7_75t_R g1882 ( 
.A(n_610),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_92),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_257),
.Y(n_1884)
);

CKINVDCx20_ASAP7_75t_R g1885 ( 
.A(n_953),
.Y(n_1885)
);

BUFx2_ASAP7_75t_L g1886 ( 
.A(n_652),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_775),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_894),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_865),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_730),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_161),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_936),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_497),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_669),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_798),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_795),
.Y(n_1896)
);

INVx1_ASAP7_75t_SL g1897 ( 
.A(n_998),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_6),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_1109),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1080),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_1051),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_254),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_1034),
.Y(n_1903)
);

INVx1_ASAP7_75t_SL g1904 ( 
.A(n_142),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1249),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_968),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_210),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_273),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_329),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_1080),
.Y(n_1910)
);

CKINVDCx20_ASAP7_75t_R g1911 ( 
.A(n_1113),
.Y(n_1911)
);

INVx2_ASAP7_75t_SL g1912 ( 
.A(n_273),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_423),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_301),
.Y(n_1914)
);

CKINVDCx20_ASAP7_75t_R g1915 ( 
.A(n_217),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_546),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_214),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_219),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_870),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_399),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1147),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_253),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_447),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_1126),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_117),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1024),
.Y(n_1926)
);

BUFx5_ASAP7_75t_L g1927 ( 
.A(n_1088),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_1059),
.Y(n_1928)
);

CKINVDCx16_ASAP7_75t_R g1929 ( 
.A(n_1037),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_17),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_840),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1059),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_524),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_1275),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_649),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1250),
.Y(n_1936)
);

CKINVDCx20_ASAP7_75t_R g1937 ( 
.A(n_1092),
.Y(n_1937)
);

BUFx3_ASAP7_75t_L g1938 ( 
.A(n_721),
.Y(n_1938)
);

CKINVDCx5p33_ASAP7_75t_R g1939 ( 
.A(n_245),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1276),
.Y(n_1940)
);

CKINVDCx5p33_ASAP7_75t_R g1941 ( 
.A(n_1273),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_127),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_842),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_641),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1021),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_240),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_269),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1203),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_974),
.Y(n_1949)
);

INVxp67_ASAP7_75t_L g1950 ( 
.A(n_1081),
.Y(n_1950)
);

HB1xp67_ASAP7_75t_L g1951 ( 
.A(n_1016),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_650),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_139),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1226),
.Y(n_1954)
);

CKINVDCx20_ASAP7_75t_R g1955 ( 
.A(n_1031),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1086),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_887),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_74),
.Y(n_1958)
);

BUFx2_ASAP7_75t_L g1959 ( 
.A(n_415),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_910),
.Y(n_1960)
);

BUFx2_ASAP7_75t_L g1961 ( 
.A(n_1083),
.Y(n_1961)
);

BUFx2_ASAP7_75t_L g1962 ( 
.A(n_532),
.Y(n_1962)
);

CKINVDCx5p33_ASAP7_75t_R g1963 ( 
.A(n_362),
.Y(n_1963)
);

BUFx2_ASAP7_75t_SL g1964 ( 
.A(n_883),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_172),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_824),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1107),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_388),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_689),
.Y(n_1969)
);

CKINVDCx20_ASAP7_75t_R g1970 ( 
.A(n_1205),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_517),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_64),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1072),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1264),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_1014),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_1084),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1063),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_360),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1263),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1192),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_1090),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1137),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_429),
.Y(n_1983)
);

BUFx3_ASAP7_75t_L g1984 ( 
.A(n_757),
.Y(n_1984)
);

CKINVDCx20_ASAP7_75t_R g1985 ( 
.A(n_931),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_801),
.Y(n_1986)
);

CKINVDCx20_ASAP7_75t_R g1987 ( 
.A(n_647),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1089),
.Y(n_1988)
);

CKINVDCx5p33_ASAP7_75t_R g1989 ( 
.A(n_161),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_1186),
.Y(n_1990)
);

CKINVDCx5p33_ASAP7_75t_R g1991 ( 
.A(n_386),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1057),
.Y(n_1992)
);

INVx1_ASAP7_75t_SL g1993 ( 
.A(n_543),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_597),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1047),
.Y(n_1995)
);

CKINVDCx11_ASAP7_75t_R g1996 ( 
.A(n_681),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_492),
.Y(n_1997)
);

CKINVDCx20_ASAP7_75t_R g1998 ( 
.A(n_919),
.Y(n_1998)
);

CKINVDCx5p33_ASAP7_75t_R g1999 ( 
.A(n_1036),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1017),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_682),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_388),
.Y(n_2002)
);

INVxp67_ASAP7_75t_SL g2003 ( 
.A(n_938),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_330),
.Y(n_2004)
);

BUFx8_ASAP7_75t_SL g2005 ( 
.A(n_1070),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_49),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1191),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_727),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_40),
.Y(n_2009)
);

CKINVDCx5p33_ASAP7_75t_R g2010 ( 
.A(n_720),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_1274),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_316),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_167),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_496),
.Y(n_2014)
);

CKINVDCx16_ASAP7_75t_R g2015 ( 
.A(n_1076),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_812),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_232),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_65),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_1085),
.Y(n_2019)
);

CKINVDCx5p33_ASAP7_75t_R g2020 ( 
.A(n_138),
.Y(n_2020)
);

CKINVDCx16_ASAP7_75t_R g2021 ( 
.A(n_139),
.Y(n_2021)
);

CKINVDCx20_ASAP7_75t_R g2022 ( 
.A(n_424),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_60),
.Y(n_2023)
);

CKINVDCx20_ASAP7_75t_R g2024 ( 
.A(n_15),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_1220),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_520),
.Y(n_2026)
);

HB1xp67_ASAP7_75t_L g2027 ( 
.A(n_1213),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_66),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1065),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_913),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_1048),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_776),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_413),
.Y(n_2033)
);

INVx2_ASAP7_75t_SL g2034 ( 
.A(n_869),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_502),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_896),
.Y(n_2036)
);

INVxp67_ASAP7_75t_L g2037 ( 
.A(n_184),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_610),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_801),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_1019),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_281),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_332),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_1062),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_67),
.Y(n_2044)
);

CKINVDCx20_ASAP7_75t_R g2045 ( 
.A(n_583),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_79),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_920),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1129),
.Y(n_2048)
);

BUFx10_ASAP7_75t_L g2049 ( 
.A(n_268),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_869),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_1102),
.Y(n_2051)
);

BUFx10_ASAP7_75t_L g2052 ( 
.A(n_840),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_398),
.Y(n_2053)
);

CKINVDCx20_ASAP7_75t_R g2054 ( 
.A(n_172),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_1143),
.Y(n_2055)
);

BUFx3_ASAP7_75t_L g2056 ( 
.A(n_852),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_1025),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_722),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_330),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_352),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_44),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_960),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1241),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_524),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_307),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_504),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_1099),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1268),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_320),
.Y(n_2069)
);

CKINVDCx5p33_ASAP7_75t_R g2070 ( 
.A(n_845),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_747),
.Y(n_2071)
);

BUFx10_ASAP7_75t_L g2072 ( 
.A(n_392),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_19),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_912),
.Y(n_2074)
);

CKINVDCx5p33_ASAP7_75t_R g2075 ( 
.A(n_445),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1085),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1174),
.Y(n_2077)
);

CKINVDCx5p33_ASAP7_75t_R g2078 ( 
.A(n_344),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1073),
.Y(n_2079)
);

CKINVDCx5p33_ASAP7_75t_R g2080 ( 
.A(n_845),
.Y(n_2080)
);

CKINVDCx5p33_ASAP7_75t_R g2081 ( 
.A(n_910),
.Y(n_2081)
);

BUFx6f_ASAP7_75t_L g2082 ( 
.A(n_1052),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_81),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_321),
.Y(n_2084)
);

CKINVDCx5p33_ASAP7_75t_R g2085 ( 
.A(n_1065),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_377),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_883),
.Y(n_2087)
);

CKINVDCx5p33_ASAP7_75t_R g2088 ( 
.A(n_2),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_13),
.Y(n_2089)
);

CKINVDCx5p33_ASAP7_75t_R g2090 ( 
.A(n_84),
.Y(n_2090)
);

CKINVDCx20_ASAP7_75t_R g2091 ( 
.A(n_652),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1148),
.Y(n_2092)
);

CKINVDCx20_ASAP7_75t_R g2093 ( 
.A(n_788),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_455),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1045),
.Y(n_2095)
);

CKINVDCx5p33_ASAP7_75t_R g2096 ( 
.A(n_1071),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1283),
.Y(n_2097)
);

CKINVDCx5p33_ASAP7_75t_R g2098 ( 
.A(n_1200),
.Y(n_2098)
);

BUFx2_ASAP7_75t_L g2099 ( 
.A(n_468),
.Y(n_2099)
);

CKINVDCx5p33_ASAP7_75t_R g2100 ( 
.A(n_1216),
.Y(n_2100)
);

CKINVDCx5p33_ASAP7_75t_R g2101 ( 
.A(n_338),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_1180),
.Y(n_2102)
);

CKINVDCx5p33_ASAP7_75t_R g2103 ( 
.A(n_1157),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_276),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_191),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1607),
.Y(n_2106)
);

INVxp67_ASAP7_75t_SL g2107 ( 
.A(n_2027),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1607),
.Y(n_2108)
);

INVxp33_ASAP7_75t_SL g2109 ( 
.A(n_1663),
.Y(n_2109)
);

BUFx3_ASAP7_75t_L g2110 ( 
.A(n_1584),
.Y(n_2110)
);

INVxp67_ASAP7_75t_SL g2111 ( 
.A(n_1393),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1607),
.Y(n_2112)
);

CKINVDCx20_ASAP7_75t_R g2113 ( 
.A(n_1410),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1607),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1607),
.Y(n_2115)
);

HB1xp67_ASAP7_75t_L g2116 ( 
.A(n_1514),
.Y(n_2116)
);

BUFx5_ASAP7_75t_L g2117 ( 
.A(n_1293),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1927),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1927),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1927),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1927),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1927),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1302),
.Y(n_2123)
);

INVxp67_ASAP7_75t_SL g2124 ( 
.A(n_1553),
.Y(n_2124)
);

INVxp67_ASAP7_75t_SL g2125 ( 
.A(n_1336),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1302),
.Y(n_2126)
);

INVxp33_ASAP7_75t_SL g2127 ( 
.A(n_1436),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1302),
.Y(n_2128)
);

CKINVDCx16_ASAP7_75t_R g2129 ( 
.A(n_1303),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1306),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1306),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1306),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1311),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1311),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1311),
.Y(n_2135)
);

CKINVDCx20_ASAP7_75t_R g2136 ( 
.A(n_1524),
.Y(n_2136)
);

BUFx6f_ASAP7_75t_L g2137 ( 
.A(n_1364),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1364),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1364),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1365),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1365),
.Y(n_2141)
);

INVxp67_ASAP7_75t_SL g2142 ( 
.A(n_1466),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1365),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1370),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1370),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1370),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1383),
.Y(n_2147)
);

INVxp67_ASAP7_75t_L g2148 ( 
.A(n_1411),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1383),
.Y(n_2149)
);

INVxp67_ASAP7_75t_L g2150 ( 
.A(n_1564),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1383),
.Y(n_2151)
);

CKINVDCx20_ASAP7_75t_R g2152 ( 
.A(n_1557),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1406),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1406),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1406),
.Y(n_2155)
);

INVxp67_ASAP7_75t_SL g2156 ( 
.A(n_1680),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1437),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1437),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1437),
.Y(n_2159)
);

CKINVDCx5p33_ASAP7_75t_R g2160 ( 
.A(n_1996),
.Y(n_2160)
);

BUFx6f_ASAP7_75t_L g2161 ( 
.A(n_1473),
.Y(n_2161)
);

INVxp67_ASAP7_75t_L g2162 ( 
.A(n_1754),
.Y(n_2162)
);

INVxp67_ASAP7_75t_SL g2163 ( 
.A(n_1695),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1473),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1473),
.Y(n_2165)
);

CKINVDCx20_ASAP7_75t_R g2166 ( 
.A(n_1565),
.Y(n_2166)
);

INVxp67_ASAP7_75t_SL g2167 ( 
.A(n_1951),
.Y(n_2167)
);

CKINVDCx5p33_ASAP7_75t_R g2168 ( 
.A(n_1841),
.Y(n_2168)
);

BUFx3_ASAP7_75t_L g2169 ( 
.A(n_1584),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_2005),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1479),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1479),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1479),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1484),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1484),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1484),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1516),
.Y(n_2177)
);

INVxp33_ASAP7_75t_SL g2178 ( 
.A(n_1986),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1516),
.Y(n_2179)
);

INVxp33_ASAP7_75t_L g2180 ( 
.A(n_1776),
.Y(n_2180)
);

CKINVDCx16_ASAP7_75t_R g2181 ( 
.A(n_1438),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_1296),
.Y(n_2182)
);

BUFx2_ASAP7_75t_L g2183 ( 
.A(n_1793),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_1297),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1516),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1519),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1519),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_1298),
.Y(n_2188)
);

CKINVDCx5p33_ASAP7_75t_R g2189 ( 
.A(n_1310),
.Y(n_2189)
);

INVxp33_ASAP7_75t_SL g2190 ( 
.A(n_1850),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1519),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_1617),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1617),
.Y(n_2193)
);

CKINVDCx20_ASAP7_75t_R g2194 ( 
.A(n_1574),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1617),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1725),
.Y(n_2196)
);

INVxp67_ASAP7_75t_L g2197 ( 
.A(n_1886),
.Y(n_2197)
);

INVxp33_ASAP7_75t_SL g2198 ( 
.A(n_1959),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1725),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1725),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1779),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1779),
.Y(n_2202)
);

INVxp33_ASAP7_75t_SL g2203 ( 
.A(n_1961),
.Y(n_2203)
);

CKINVDCx20_ASAP7_75t_R g2204 ( 
.A(n_1579),
.Y(n_2204)
);

INVxp67_ASAP7_75t_L g2205 ( 
.A(n_1962),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1779),
.Y(n_2206)
);

CKINVDCx20_ASAP7_75t_R g2207 ( 
.A(n_1600),
.Y(n_2207)
);

INVxp33_ASAP7_75t_SL g2208 ( 
.A(n_2099),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1887),
.Y(n_2209)
);

INVxp67_ASAP7_75t_SL g2210 ( 
.A(n_1887),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1887),
.Y(n_2211)
);

INVxp67_ASAP7_75t_SL g2212 ( 
.A(n_1969),
.Y(n_2212)
);

INVxp33_ASAP7_75t_SL g2213 ( 
.A(n_1292),
.Y(n_2213)
);

CKINVDCx16_ASAP7_75t_R g2214 ( 
.A(n_1759),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1969),
.Y(n_2215)
);

CKINVDCx16_ASAP7_75t_R g2216 ( 
.A(n_1789),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1969),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2082),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2082),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2082),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1312),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1417),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1618),
.Y(n_2223)
);

CKINVDCx20_ASAP7_75t_R g2224 ( 
.A(n_1664),
.Y(n_2224)
);

INVxp33_ASAP7_75t_SL g2225 ( 
.A(n_1294),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_1384),
.Y(n_2226)
);

CKINVDCx16_ASAP7_75t_R g2227 ( 
.A(n_1827),
.Y(n_2227)
);

BUFx2_ASAP7_75t_L g2228 ( 
.A(n_1441),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1729),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1858),
.Y(n_2230)
);

CKINVDCx20_ASAP7_75t_R g2231 ( 
.A(n_1681),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1878),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1938),
.Y(n_2233)
);

INVx3_ASAP7_75t_L g2234 ( 
.A(n_1984),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2056),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2094),
.Y(n_2236)
);

INVxp33_ASAP7_75t_L g2237 ( 
.A(n_1307),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2105),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1314),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1320),
.Y(n_2240)
);

CKINVDCx5p33_ASAP7_75t_R g2241 ( 
.A(n_1327),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1322),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1331),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1332),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1345),
.Y(n_2245)
);

INVxp33_ASAP7_75t_L g2246 ( 
.A(n_1352),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1355),
.Y(n_2247)
);

CKINVDCx20_ASAP7_75t_R g2248 ( 
.A(n_1699),
.Y(n_2248)
);

CKINVDCx20_ASAP7_75t_R g2249 ( 
.A(n_1709),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1357),
.Y(n_2250)
);

CKINVDCx20_ASAP7_75t_R g2251 ( 
.A(n_1746),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_1384),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2089),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1373),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1374),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1375),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1390),
.Y(n_2257)
);

INVxp67_ASAP7_75t_SL g2258 ( 
.A(n_1308),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1391),
.Y(n_2259)
);

CKINVDCx5p33_ASAP7_75t_R g2260 ( 
.A(n_1328),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1399),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_1400),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_1334),
.Y(n_2263)
);

CKINVDCx16_ASAP7_75t_R g2264 ( 
.A(n_1929),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1402),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1412),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1413),
.Y(n_2267)
);

BUFx2_ASAP7_75t_SL g2268 ( 
.A(n_1765),
.Y(n_2268)
);

INVxp67_ASAP7_75t_SL g2269 ( 
.A(n_1313),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1418),
.Y(n_2270)
);

INVxp67_ASAP7_75t_SL g2271 ( 
.A(n_1339),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2126),
.Y(n_2272)
);

AND2x4_ASAP7_75t_L g2273 ( 
.A(n_2228),
.B(n_1300),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2263),
.Y(n_2274)
);

BUFx2_ASAP7_75t_L g2275 ( 
.A(n_2160),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2182),
.B(n_1525),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2263),
.Y(n_2277)
);

CKINVDCx11_ASAP7_75t_R g2278 ( 
.A(n_2113),
.Y(n_2278)
);

INVxp67_ASAP7_75t_L g2279 ( 
.A(n_2110),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2111),
.B(n_1615),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2210),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2184),
.B(n_1700),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2188),
.B(n_1701),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2145),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2212),
.Y(n_2285)
);

OAI22x1_ASAP7_75t_R g2286 ( 
.A1(n_2136),
.A2(n_1321),
.B1(n_1323),
.B2(n_1317),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2137),
.Y(n_2287)
);

BUFx6f_ASAP7_75t_L g2288 ( 
.A(n_2137),
.Y(n_2288)
);

INVxp67_ASAP7_75t_L g2289 ( 
.A(n_2169),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2155),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2186),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2161),
.Y(n_2292)
);

CKINVDCx11_ASAP7_75t_R g2293 ( 
.A(n_2152),
.Y(n_2293)
);

BUFx2_ASAP7_75t_L g2294 ( 
.A(n_2189),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2161),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2191),
.Y(n_2296)
);

BUFx2_ASAP7_75t_L g2297 ( 
.A(n_2241),
.Y(n_2297)
);

BUFx6f_ASAP7_75t_L g2298 ( 
.A(n_2192),
.Y(n_2298)
);

CKINVDCx5p33_ASAP7_75t_R g2299 ( 
.A(n_2260),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2124),
.B(n_1720),
.Y(n_2300)
);

BUFx12f_ASAP7_75t_L g2301 ( 
.A(n_2168),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2125),
.B(n_2015),
.Y(n_2302)
);

INVxp67_ASAP7_75t_L g2303 ( 
.A(n_2183),
.Y(n_2303)
);

INVx5_ASAP7_75t_L g2304 ( 
.A(n_2234),
.Y(n_2304)
);

BUFx3_ASAP7_75t_L g2305 ( 
.A(n_2221),
.Y(n_2305)
);

AND2x4_ASAP7_75t_L g2306 ( 
.A(n_2156),
.B(n_1463),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2193),
.Y(n_2307)
);

INVx3_ASAP7_75t_L g2308 ( 
.A(n_2123),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2128),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2130),
.Y(n_2310)
);

AND2x4_ASAP7_75t_L g2311 ( 
.A(n_2163),
.B(n_1760),
.Y(n_2311)
);

BUFx6f_ASAP7_75t_L g2312 ( 
.A(n_2131),
.Y(n_2312)
);

INVx5_ASAP7_75t_L g2313 ( 
.A(n_2129),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2132),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2133),
.Y(n_2315)
);

BUFx6f_ASAP7_75t_L g2316 ( 
.A(n_2134),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2135),
.Y(n_2317)
);

INVxp67_ASAP7_75t_L g2318 ( 
.A(n_2116),
.Y(n_2318)
);

BUFx12f_ASAP7_75t_L g2319 ( 
.A(n_2170),
.Y(n_2319)
);

HB1xp67_ASAP7_75t_L g2320 ( 
.A(n_2181),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2138),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2139),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2140),
.Y(n_2323)
);

CKINVDCx5p33_ASAP7_75t_R g2324 ( 
.A(n_2268),
.Y(n_2324)
);

AOI22xp5_ASAP7_75t_L g2325 ( 
.A1(n_2190),
.A2(n_1773),
.B1(n_1515),
.B2(n_2021),
.Y(n_2325)
);

OAI21x1_ASAP7_75t_L g2326 ( 
.A1(n_2108),
.A2(n_1366),
.B(n_1337),
.Y(n_2326)
);

BUFx6f_ASAP7_75t_L g2327 ( 
.A(n_2141),
.Y(n_2327)
);

OA21x2_ASAP7_75t_L g2328 ( 
.A1(n_2106),
.A2(n_1379),
.B(n_1346),
.Y(n_2328)
);

NOR2x1_ASAP7_75t_L g2329 ( 
.A(n_2112),
.B(n_1398),
.Y(n_2329)
);

INVx2_ASAP7_75t_SL g2330 ( 
.A(n_2222),
.Y(n_2330)
);

AND2x2_ASAP7_75t_SL g2331 ( 
.A(n_2214),
.B(n_1420),
.Y(n_2331)
);

AND2x4_ASAP7_75t_L g2332 ( 
.A(n_2167),
.B(n_1772),
.Y(n_2332)
);

CKINVDCx20_ASAP7_75t_R g2333 ( 
.A(n_2166),
.Y(n_2333)
);

OA21x2_ASAP7_75t_L g2334 ( 
.A1(n_2114),
.A2(n_1448),
.B(n_1409),
.Y(n_2334)
);

BUFx2_ASAP7_75t_L g2335 ( 
.A(n_2216),
.Y(n_2335)
);

INVx3_ASAP7_75t_L g2336 ( 
.A(n_2143),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2144),
.Y(n_2337)
);

BUFx6f_ASAP7_75t_L g2338 ( 
.A(n_2146),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2147),
.Y(n_2339)
);

OA21x2_ASAP7_75t_L g2340 ( 
.A1(n_2119),
.A2(n_1562),
.B(n_1453),
.Y(n_2340)
);

AND2x4_ASAP7_75t_L g2341 ( 
.A(n_2107),
.B(n_1590),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2149),
.Y(n_2342)
);

BUFx8_ASAP7_75t_SL g2343 ( 
.A(n_2194),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2151),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2153),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2142),
.B(n_1429),
.Y(n_2346)
);

NOR2x1_ASAP7_75t_L g2347 ( 
.A(n_2120),
.B(n_1601),
.Y(n_2347)
);

OAI22xp5_ASAP7_75t_L g2348 ( 
.A1(n_2198),
.A2(n_1451),
.B1(n_1504),
.B2(n_1450),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2154),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2157),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2158),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2159),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2180),
.B(n_2003),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2164),
.Y(n_2354)
);

OAI21x1_ASAP7_75t_L g2355 ( 
.A1(n_2115),
.A2(n_1512),
.B(n_1499),
.Y(n_2355)
);

INVx4_ASAP7_75t_L g2356 ( 
.A(n_2117),
.Y(n_2356)
);

OA21x2_ASAP7_75t_L g2357 ( 
.A1(n_2121),
.A2(n_1762),
.B(n_1738),
.Y(n_2357)
);

AND2x4_ASAP7_75t_L g2358 ( 
.A(n_2148),
.B(n_1767),
.Y(n_2358)
);

BUFx3_ASAP7_75t_L g2359 ( 
.A(n_2223),
.Y(n_2359)
);

INVx4_ASAP7_75t_L g2360 ( 
.A(n_2117),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2258),
.B(n_1622),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2165),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2171),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2172),
.Y(n_2364)
);

HB1xp67_ASAP7_75t_L g2365 ( 
.A(n_2227),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2173),
.Y(n_2366)
);

INVx3_ASAP7_75t_L g2367 ( 
.A(n_2174),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2175),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_2204),
.Y(n_2369)
);

BUFx2_ASAP7_75t_L g2370 ( 
.A(n_2264),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2176),
.Y(n_2371)
);

AND2x4_ASAP7_75t_L g2372 ( 
.A(n_2150),
.B(n_1775),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2177),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2179),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2185),
.Y(n_2375)
);

NOR2xp33_ASAP7_75t_L g2376 ( 
.A(n_2213),
.B(n_1804),
.Y(n_2376)
);

INVx3_ASAP7_75t_L g2377 ( 
.A(n_2187),
.Y(n_2377)
);

BUFx12f_ASAP7_75t_L g2378 ( 
.A(n_2225),
.Y(n_2378)
);

BUFx3_ASAP7_75t_L g2379 ( 
.A(n_2229),
.Y(n_2379)
);

AOI22xp5_ASAP7_75t_L g2380 ( 
.A1(n_2203),
.A2(n_2208),
.B1(n_2127),
.B2(n_2178),
.Y(n_2380)
);

BUFx8_ASAP7_75t_L g2381 ( 
.A(n_2230),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2195),
.Y(n_2382)
);

BUFx6f_ASAP7_75t_L g2383 ( 
.A(n_2196),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2269),
.B(n_1676),
.Y(n_2384)
);

BUFx6f_ASAP7_75t_L g2385 ( 
.A(n_2199),
.Y(n_2385)
);

HB1xp67_ASAP7_75t_L g2386 ( 
.A(n_2162),
.Y(n_2386)
);

OAI22xp5_ASAP7_75t_L g2387 ( 
.A1(n_2109),
.A2(n_2205),
.B1(n_2197),
.B2(n_2271),
.Y(n_2387)
);

INVx5_ASAP7_75t_L g2388 ( 
.A(n_2118),
.Y(n_2388)
);

AND2x6_ASAP7_75t_L g2389 ( 
.A(n_2232),
.B(n_1304),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_2237),
.B(n_1295),
.Y(n_2390)
);

INVx3_ASAP7_75t_L g2391 ( 
.A(n_2200),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2117),
.B(n_1835),
.Y(n_2392)
);

HB1xp67_ASAP7_75t_L g2393 ( 
.A(n_2233),
.Y(n_2393)
);

NAND2xp33_ASAP7_75t_L g2394 ( 
.A(n_2117),
.B(n_1299),
.Y(n_2394)
);

INVx5_ASAP7_75t_L g2395 ( 
.A(n_2226),
.Y(n_2395)
);

AND2x4_ASAP7_75t_L g2396 ( 
.A(n_2235),
.B(n_1810),
.Y(n_2396)
);

INVx6_ASAP7_75t_L g2397 ( 
.A(n_2246),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2201),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2202),
.B(n_1414),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2206),
.Y(n_2400)
);

CKINVDCx6p67_ASAP7_75t_R g2401 ( 
.A(n_2207),
.Y(n_2401)
);

BUFx3_ASAP7_75t_L g2402 ( 
.A(n_2209),
.Y(n_2402)
);

INVxp67_ASAP7_75t_L g2403 ( 
.A(n_2236),
.Y(n_2403)
);

BUFx6f_ASAP7_75t_L g2404 ( 
.A(n_2211),
.Y(n_2404)
);

BUFx6f_ASAP7_75t_L g2405 ( 
.A(n_2215),
.Y(n_2405)
);

OAI21x1_ASAP7_75t_L g2406 ( 
.A1(n_2252),
.A2(n_2068),
.B(n_1921),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2217),
.Y(n_2407)
);

BUFx12f_ASAP7_75t_L g2408 ( 
.A(n_2224),
.Y(n_2408)
);

BUFx3_ASAP7_75t_L g2409 ( 
.A(n_2218),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2219),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_2220),
.Y(n_2411)
);

INVx6_ASAP7_75t_L g2412 ( 
.A(n_2238),
.Y(n_2412)
);

INVx5_ASAP7_75t_L g2413 ( 
.A(n_2239),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2122),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2240),
.Y(n_2415)
);

BUFx3_ASAP7_75t_L g2416 ( 
.A(n_2242),
.Y(n_2416)
);

OAI22xp5_ASAP7_75t_L g2417 ( 
.A1(n_2231),
.A2(n_1602),
.B1(n_1608),
.B2(n_1550),
.Y(n_2417)
);

CKINVDCx20_ASAP7_75t_R g2418 ( 
.A(n_2248),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2243),
.Y(n_2419)
);

CKINVDCx5p33_ASAP7_75t_R g2420 ( 
.A(n_2249),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2244),
.Y(n_2421)
);

BUFx3_ASAP7_75t_L g2422 ( 
.A(n_2245),
.Y(n_2422)
);

AND2x4_ASAP7_75t_L g2423 ( 
.A(n_2247),
.B(n_1823),
.Y(n_2423)
);

AND2x4_ASAP7_75t_L g2424 ( 
.A(n_2250),
.B(n_1830),
.Y(n_2424)
);

BUFx6f_ASAP7_75t_L g2425 ( 
.A(n_2253),
.Y(n_2425)
);

BUFx12f_ASAP7_75t_L g2426 ( 
.A(n_2251),
.Y(n_2426)
);

BUFx6f_ASAP7_75t_L g2427 ( 
.A(n_2254),
.Y(n_2427)
);

NOR2x1_ASAP7_75t_L g2428 ( 
.A(n_2255),
.B(n_1838),
.Y(n_2428)
);

BUFx2_ASAP7_75t_L g2429 ( 
.A(n_2256),
.Y(n_2429)
);

OAI22xp5_ASAP7_75t_L g2430 ( 
.A1(n_2257),
.A2(n_1877),
.B1(n_1950),
.B2(n_1817),
.Y(n_2430)
);

INVx6_ASAP7_75t_L g2431 ( 
.A(n_2259),
.Y(n_2431)
);

CKINVDCx11_ASAP7_75t_R g2432 ( 
.A(n_2261),
.Y(n_2432)
);

OAI22xp5_ASAP7_75t_L g2433 ( 
.A1(n_2262),
.A2(n_2037),
.B1(n_1305),
.B2(n_1309),
.Y(n_2433)
);

BUFx6f_ASAP7_75t_L g2434 ( 
.A(n_2265),
.Y(n_2434)
);

OAI22xp5_ASAP7_75t_SL g2435 ( 
.A1(n_2266),
.A2(n_1350),
.B1(n_1407),
.B2(n_1405),
.Y(n_2435)
);

BUFx3_ASAP7_75t_L g2436 ( 
.A(n_2267),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2270),
.Y(n_2437)
);

INVx6_ASAP7_75t_L g2438 ( 
.A(n_2137),
.Y(n_2438)
);

HB1xp67_ASAP7_75t_L g2439 ( 
.A(n_2129),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2126),
.Y(n_2440)
);

AND2x4_ASAP7_75t_L g2441 ( 
.A(n_2228),
.B(n_1846),
.Y(n_2441)
);

AOI22xp5_ASAP7_75t_L g2442 ( 
.A1(n_2190),
.A2(n_1970),
.B1(n_1769),
.B2(n_1315),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2126),
.Y(n_2443)
);

BUFx6f_ASAP7_75t_L g2444 ( 
.A(n_2137),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_2182),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2228),
.B(n_1443),
.Y(n_2446)
);

INVx6_ASAP7_75t_L g2447 ( 
.A(n_2137),
.Y(n_2447)
);

AND2x4_ASAP7_75t_L g2448 ( 
.A(n_2228),
.B(n_1847),
.Y(n_2448)
);

HB1xp67_ASAP7_75t_L g2449 ( 
.A(n_2129),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2126),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2182),
.B(n_2077),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2263),
.Y(n_2452)
);

HB1xp67_ASAP7_75t_L g2453 ( 
.A(n_2129),
.Y(n_2453)
);

HB1xp67_ASAP7_75t_L g2454 ( 
.A(n_2129),
.Y(n_2454)
);

INVx5_ASAP7_75t_L g2455 ( 
.A(n_2137),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2263),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2126),
.Y(n_2457)
);

BUFx6f_ASAP7_75t_L g2458 ( 
.A(n_2137),
.Y(n_2458)
);

BUFx2_ASAP7_75t_L g2459 ( 
.A(n_2160),
.Y(n_2459)
);

AOI22xp5_ASAP7_75t_L g2460 ( 
.A1(n_2190),
.A2(n_1316),
.B1(n_1318),
.B2(n_1301),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2263),
.Y(n_2461)
);

BUFx6f_ASAP7_75t_L g2462 ( 
.A(n_2137),
.Y(n_2462)
);

AOI22xp5_ASAP7_75t_L g2463 ( 
.A1(n_2190),
.A2(n_1324),
.B1(n_1325),
.B2(n_1319),
.Y(n_2463)
);

BUFx6f_ASAP7_75t_L g2464 ( 
.A(n_2137),
.Y(n_2464)
);

BUFx6f_ASAP7_75t_L g2465 ( 
.A(n_2137),
.Y(n_2465)
);

BUFx3_ASAP7_75t_L g2466 ( 
.A(n_2234),
.Y(n_2466)
);

AND2x4_ASAP7_75t_L g2467 ( 
.A(n_2228),
.B(n_1866),
.Y(n_2467)
);

INVx3_ASAP7_75t_L g2468 ( 
.A(n_2137),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2182),
.B(n_1880),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2126),
.Y(n_2470)
);

INVx3_ASAP7_75t_L g2471 ( 
.A(n_2137),
.Y(n_2471)
);

BUFx2_ASAP7_75t_L g2472 ( 
.A(n_2160),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2263),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2263),
.Y(n_2474)
);

CKINVDCx6p67_ASAP7_75t_R g2475 ( 
.A(n_2129),
.Y(n_2475)
);

BUFx6f_ASAP7_75t_L g2476 ( 
.A(n_2137),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2126),
.Y(n_2477)
);

AND2x4_ASAP7_75t_L g2478 ( 
.A(n_2228),
.B(n_1974),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2263),
.Y(n_2479)
);

BUFx12f_ASAP7_75t_L g2480 ( 
.A(n_2168),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2126),
.Y(n_2481)
);

AOI22x1_ASAP7_75t_SL g2482 ( 
.A1(n_2113),
.A2(n_1454),
.B1(n_1461),
.B2(n_1419),
.Y(n_2482)
);

BUFx6f_ASAP7_75t_L g2483 ( 
.A(n_2137),
.Y(n_2483)
);

INVx3_ASAP7_75t_L g2484 ( 
.A(n_2137),
.Y(n_2484)
);

INVx3_ASAP7_75t_L g2485 ( 
.A(n_2137),
.Y(n_2485)
);

HB1xp67_ASAP7_75t_L g2486 ( 
.A(n_2129),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2126),
.Y(n_2487)
);

OAI22x1_ASAP7_75t_L g2488 ( 
.A1(n_2183),
.A2(n_1356),
.B1(n_1376),
.B2(n_1333),
.Y(n_2488)
);

OA21x2_ASAP7_75t_L g2489 ( 
.A1(n_2106),
.A2(n_1982),
.B(n_1979),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2126),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2182),
.B(n_2007),
.Y(n_2491)
);

BUFx6f_ASAP7_75t_L g2492 ( 
.A(n_2137),
.Y(n_2492)
);

AOI22xp5_ASAP7_75t_L g2493 ( 
.A1(n_2190),
.A2(n_1329),
.B1(n_1330),
.B2(n_1326),
.Y(n_2493)
);

INVx2_ASAP7_75t_SL g2494 ( 
.A(n_2110),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2263),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2228),
.B(n_1764),
.Y(n_2496)
);

AND2x4_ASAP7_75t_L g2497 ( 
.A(n_2228),
.B(n_2048),
.Y(n_2497)
);

OAI21x1_ASAP7_75t_L g2498 ( 
.A1(n_2108),
.A2(n_2092),
.B(n_2063),
.Y(n_2498)
);

AND2x4_ASAP7_75t_L g2499 ( 
.A(n_2228),
.B(n_2097),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2228),
.B(n_1783),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2126),
.Y(n_2501)
);

AND2x2_ASAP7_75t_SL g2502 ( 
.A(n_2129),
.B(n_1421),
.Y(n_2502)
);

NOR2x1_ASAP7_75t_L g2503 ( 
.A(n_2110),
.B(n_1334),
.Y(n_2503)
);

AND2x4_ASAP7_75t_L g2504 ( 
.A(n_2228),
.B(n_1790),
.Y(n_2504)
);

INVx3_ASAP7_75t_L g2505 ( 
.A(n_2137),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2263),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2263),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2182),
.B(n_1338),
.Y(n_2508)
);

BUFx2_ASAP7_75t_L g2509 ( 
.A(n_2160),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_2182),
.B(n_1343),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2263),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2126),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2126),
.Y(n_2513)
);

OAI21x1_ASAP7_75t_L g2514 ( 
.A1(n_2108),
.A2(n_1442),
.B(n_1424),
.Y(n_2514)
);

BUFx6f_ASAP7_75t_L g2515 ( 
.A(n_2137),
.Y(n_2515)
);

OA21x2_ASAP7_75t_L g2516 ( 
.A1(n_2106),
.A2(n_1349),
.B(n_1344),
.Y(n_2516)
);

AOI22xp5_ASAP7_75t_L g2517 ( 
.A1(n_2190),
.A2(n_1335),
.B1(n_1341),
.B2(n_1340),
.Y(n_2517)
);

OAI22x1_ASAP7_75t_R g2518 ( 
.A1(n_2113),
.A2(n_1481),
.B1(n_1495),
.B2(n_1464),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2263),
.Y(n_2519)
);

NOR2x1_ASAP7_75t_L g2520 ( 
.A(n_2110),
.B(n_1334),
.Y(n_2520)
);

INVx6_ASAP7_75t_L g2521 ( 
.A(n_2137),
.Y(n_2521)
);

INVx3_ASAP7_75t_L g2522 ( 
.A(n_2137),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2263),
.Y(n_2523)
);

OAI22xp5_ASAP7_75t_L g2524 ( 
.A1(n_2190),
.A2(n_1347),
.B1(n_1348),
.B2(n_1342),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2228),
.B(n_1856),
.Y(n_2525)
);

BUFx12f_ASAP7_75t_L g2526 ( 
.A(n_2168),
.Y(n_2526)
);

BUFx6f_ASAP7_75t_L g2527 ( 
.A(n_2137),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2126),
.Y(n_2528)
);

CKINVDCx5p33_ASAP7_75t_R g2529 ( 
.A(n_2182),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2263),
.Y(n_2530)
);

INVx3_ASAP7_75t_L g2531 ( 
.A(n_2137),
.Y(n_2531)
);

HB1xp67_ASAP7_75t_L g2532 ( 
.A(n_2129),
.Y(n_2532)
);

BUFx3_ASAP7_75t_L g2533 ( 
.A(n_2234),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2263),
.Y(n_2534)
);

HB1xp67_ASAP7_75t_L g2535 ( 
.A(n_2129),
.Y(n_2535)
);

INVx3_ASAP7_75t_L g2536 ( 
.A(n_2137),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2263),
.Y(n_2537)
);

AOI22xp5_ASAP7_75t_L g2538 ( 
.A1(n_2190),
.A2(n_1353),
.B1(n_1358),
.B2(n_1351),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2263),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2263),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2126),
.Y(n_2541)
);

INVx2_ASAP7_75t_SL g2542 ( 
.A(n_2110),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2263),
.Y(n_2543)
);

AND2x4_ASAP7_75t_L g2544 ( 
.A(n_2228),
.B(n_1912),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_2182),
.B(n_1359),
.Y(n_2545)
);

OAI22xp5_ASAP7_75t_SL g2546 ( 
.A1(n_2190),
.A2(n_1529),
.B1(n_1540),
.B2(n_1496),
.Y(n_2546)
);

BUFx8_ASAP7_75t_L g2547 ( 
.A(n_2228),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2263),
.Y(n_2548)
);

BUFx2_ASAP7_75t_L g2549 ( 
.A(n_2160),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2182),
.B(n_1361),
.Y(n_2550)
);

NAND2xp33_ASAP7_75t_L g2551 ( 
.A(n_2182),
.B(n_1360),
.Y(n_2551)
);

INVxp67_ASAP7_75t_L g2552 ( 
.A(n_2110),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2126),
.Y(n_2553)
);

BUFx3_ASAP7_75t_L g2554 ( 
.A(n_2234),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2263),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_2126),
.Y(n_2556)
);

INVx3_ASAP7_75t_L g2557 ( 
.A(n_2137),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2263),
.Y(n_2558)
);

BUFx6f_ASAP7_75t_L g2559 ( 
.A(n_2137),
.Y(n_2559)
);

AND2x4_ASAP7_75t_L g2560 ( 
.A(n_2228),
.B(n_2034),
.Y(n_2560)
);

BUFx6f_ASAP7_75t_L g2561 ( 
.A(n_2137),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2228),
.B(n_1381),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2263),
.Y(n_2563)
);

INVx4_ASAP7_75t_L g2564 ( 
.A(n_2182),
.Y(n_2564)
);

BUFx3_ASAP7_75t_L g2565 ( 
.A(n_2234),
.Y(n_2565)
);

NOR2xp33_ASAP7_75t_L g2566 ( 
.A(n_2213),
.B(n_1372),
.Y(n_2566)
);

HB1xp67_ASAP7_75t_L g2567 ( 
.A(n_2129),
.Y(n_2567)
);

BUFx3_ASAP7_75t_L g2568 ( 
.A(n_2234),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2126),
.Y(n_2569)
);

BUFx6f_ASAP7_75t_L g2570 ( 
.A(n_2137),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2126),
.Y(n_2571)
);

BUFx2_ASAP7_75t_L g2572 ( 
.A(n_2160),
.Y(n_2572)
);

BUFx12f_ASAP7_75t_L g2573 ( 
.A(n_2168),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2182),
.B(n_1392),
.Y(n_2574)
);

BUFx6f_ASAP7_75t_L g2575 ( 
.A(n_2137),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2263),
.Y(n_2576)
);

HB1xp67_ASAP7_75t_L g2577 ( 
.A(n_2129),
.Y(n_2577)
);

INVx4_ASAP7_75t_L g2578 ( 
.A(n_2182),
.Y(n_2578)
);

HB1xp67_ASAP7_75t_L g2579 ( 
.A(n_2129),
.Y(n_2579)
);

BUFx6f_ASAP7_75t_L g2580 ( 
.A(n_2137),
.Y(n_2580)
);

AND2x2_ASAP7_75t_SL g2581 ( 
.A(n_2129),
.B(n_1493),
.Y(n_2581)
);

BUFx6f_ASAP7_75t_L g2582 ( 
.A(n_2137),
.Y(n_2582)
);

BUFx6f_ASAP7_75t_L g2583 ( 
.A(n_2137),
.Y(n_2583)
);

INVx2_ASAP7_75t_L g2584 ( 
.A(n_2126),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2263),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2263),
.Y(n_2586)
);

INVx2_ASAP7_75t_SL g2587 ( 
.A(n_2110),
.Y(n_2587)
);

HB1xp67_ASAP7_75t_L g2588 ( 
.A(n_2129),
.Y(n_2588)
);

HB1xp67_ASAP7_75t_L g2589 ( 
.A(n_2129),
.Y(n_2589)
);

BUFx8_ASAP7_75t_L g2590 ( 
.A(n_2228),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2126),
.Y(n_2591)
);

OAI21x1_ASAP7_75t_L g2592 ( 
.A1(n_2108),
.A2(n_1522),
.B(n_1520),
.Y(n_2592)
);

INVx4_ASAP7_75t_L g2593 ( 
.A(n_2182),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2263),
.Y(n_2594)
);

AND2x2_ASAP7_75t_SL g2595 ( 
.A(n_2129),
.B(n_1527),
.Y(n_2595)
);

BUFx6f_ASAP7_75t_L g2596 ( 
.A(n_2137),
.Y(n_2596)
);

AND2x6_ASAP7_75t_L g2597 ( 
.A(n_2110),
.B(n_1422),
.Y(n_2597)
);

OA21x2_ASAP7_75t_L g2598 ( 
.A1(n_2106),
.A2(n_1395),
.B(n_1394),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2228),
.B(n_1381),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2415),
.Y(n_2600)
);

BUFx6f_ASAP7_75t_L g2601 ( 
.A(n_2288),
.Y(n_2601)
);

BUFx6f_ASAP7_75t_L g2602 ( 
.A(n_2444),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2419),
.Y(n_2603)
);

AND2x4_ASAP7_75t_L g2604 ( 
.A(n_2466),
.B(n_1427),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2298),
.Y(n_2605)
);

BUFx3_ASAP7_75t_L g2606 ( 
.A(n_2533),
.Y(n_2606)
);

AND2x4_ASAP7_75t_L g2607 ( 
.A(n_2554),
.B(n_1440),
.Y(n_2607)
);

AND2x4_ASAP7_75t_L g2608 ( 
.A(n_2565),
.B(n_1455),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2421),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2437),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2416),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2422),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2436),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2425),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2272),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2427),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2284),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2290),
.Y(n_2618)
);

INVx3_ASAP7_75t_L g2619 ( 
.A(n_2397),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2291),
.Y(n_2620)
);

INVx3_ASAP7_75t_L g2621 ( 
.A(n_2458),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2434),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2414),
.Y(n_2623)
);

XOR2xp5_ASAP7_75t_L g2624 ( 
.A(n_2333),
.B(n_1430),
.Y(n_2624)
);

BUFx3_ASAP7_75t_L g2625 ( 
.A(n_2568),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2305),
.Y(n_2626)
);

BUFx6f_ASAP7_75t_L g2627 ( 
.A(n_2462),
.Y(n_2627)
);

AND2x4_ASAP7_75t_L g2628 ( 
.A(n_2494),
.B(n_1458),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2440),
.Y(n_2629)
);

HB1xp67_ASAP7_75t_L g2630 ( 
.A(n_2320),
.Y(n_2630)
);

BUFx2_ASAP7_75t_L g2631 ( 
.A(n_2335),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2359),
.Y(n_2632)
);

AND2x4_ASAP7_75t_L g2633 ( 
.A(n_2542),
.B(n_1462),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2379),
.Y(n_2634)
);

BUFx6f_ASAP7_75t_L g2635 ( 
.A(n_2464),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2412),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2280),
.B(n_1432),
.Y(n_2637)
);

NOR2xp33_ASAP7_75t_SL g2638 ( 
.A(n_2378),
.B(n_1560),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2443),
.Y(n_2639)
);

BUFx6f_ASAP7_75t_L g2640 ( 
.A(n_2465),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2450),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2431),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2451),
.B(n_1444),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2457),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2402),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2409),
.Y(n_2646)
);

BUFx6f_ASAP7_75t_L g2647 ( 
.A(n_2476),
.Y(n_2647)
);

BUFx6f_ASAP7_75t_L g2648 ( 
.A(n_2483),
.Y(n_2648)
);

INVx3_ASAP7_75t_L g2649 ( 
.A(n_2492),
.Y(n_2649)
);

HB1xp67_ASAP7_75t_L g2650 ( 
.A(n_2365),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2281),
.Y(n_2651)
);

BUFx8_ASAP7_75t_L g2652 ( 
.A(n_2370),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2285),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2393),
.Y(n_2654)
);

INVx2_ASAP7_75t_L g2655 ( 
.A(n_2470),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2274),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2277),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2452),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2469),
.B(n_1447),
.Y(n_2659)
);

INVx3_ASAP7_75t_L g2660 ( 
.A(n_2515),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2477),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2456),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2461),
.Y(n_2663)
);

AND2x4_ASAP7_75t_L g2664 ( 
.A(n_2587),
.B(n_1465),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2473),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2481),
.Y(n_2666)
);

INVx3_ASAP7_75t_L g2667 ( 
.A(n_2527),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_SL g2668 ( 
.A(n_2273),
.B(n_1452),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2474),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2491),
.B(n_1456),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2479),
.Y(n_2671)
);

NOR2xp33_ASAP7_75t_L g2672 ( 
.A(n_2276),
.B(n_1362),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2376),
.B(n_1475),
.Y(n_2673)
);

NOR2xp33_ASAP7_75t_L g2674 ( 
.A(n_2282),
.B(n_1363),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2495),
.Y(n_2675)
);

AND2x4_ASAP7_75t_L g2676 ( 
.A(n_2441),
.B(n_2448),
.Y(n_2676)
);

BUFx2_ASAP7_75t_L g2677 ( 
.A(n_2439),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2390),
.B(n_2302),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2487),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2506),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2507),
.Y(n_2681)
);

BUFx6f_ASAP7_75t_L g2682 ( 
.A(n_2559),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2511),
.Y(n_2683)
);

INVx3_ASAP7_75t_L g2684 ( 
.A(n_2561),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2519),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2523),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2508),
.B(n_1478),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2490),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2501),
.Y(n_2689)
);

HB1xp67_ASAP7_75t_L g2690 ( 
.A(n_2449),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2530),
.Y(n_2691)
);

OAI22xp5_ASAP7_75t_SL g2692 ( 
.A1(n_2546),
.A2(n_1576),
.B1(n_1581),
.B2(n_1570),
.Y(n_2692)
);

NOR2xp33_ASAP7_75t_L g2693 ( 
.A(n_2283),
.B(n_1367),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2534),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2537),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2539),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2540),
.Y(n_2697)
);

AND2x4_ASAP7_75t_L g2698 ( 
.A(n_2467),
.B(n_1476),
.Y(n_2698)
);

CKINVDCx5p33_ASAP7_75t_R g2699 ( 
.A(n_2343),
.Y(n_2699)
);

HB1xp67_ASAP7_75t_L g2700 ( 
.A(n_2453),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2512),
.Y(n_2701)
);

INVx3_ASAP7_75t_L g2702 ( 
.A(n_2570),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2543),
.Y(n_2703)
);

INVx3_ASAP7_75t_L g2704 ( 
.A(n_2575),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2510),
.B(n_1483),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2548),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2513),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2545),
.B(n_1488),
.Y(n_2708)
);

BUFx3_ASAP7_75t_L g2709 ( 
.A(n_2408),
.Y(n_2709)
);

HB1xp67_ASAP7_75t_L g2710 ( 
.A(n_2454),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2555),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2528),
.Y(n_2712)
);

AND2x6_ASAP7_75t_L g2713 ( 
.A(n_2329),
.B(n_1354),
.Y(n_2713)
);

AND2x6_ASAP7_75t_L g2714 ( 
.A(n_2347),
.B(n_1354),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2541),
.Y(n_2715)
);

CKINVDCx8_ASAP7_75t_R g2716 ( 
.A(n_2313),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2558),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_SL g2718 ( 
.A(n_2306),
.B(n_1505),
.Y(n_2718)
);

INVx3_ASAP7_75t_L g2719 ( 
.A(n_2580),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2563),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2576),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2585),
.Y(n_2722)
);

BUFx6f_ASAP7_75t_L g2723 ( 
.A(n_2582),
.Y(n_2723)
);

INVxp67_ASAP7_75t_L g2724 ( 
.A(n_2386),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2586),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2594),
.Y(n_2726)
);

CKINVDCx8_ASAP7_75t_R g2727 ( 
.A(n_2313),
.Y(n_2727)
);

AND2x4_ASAP7_75t_L g2728 ( 
.A(n_2478),
.B(n_1486),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_2553),
.Y(n_2729)
);

INVxp67_ASAP7_75t_L g2730 ( 
.A(n_2599),
.Y(n_2730)
);

INVx3_ASAP7_75t_L g2731 ( 
.A(n_2583),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2315),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2321),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2556),
.Y(n_2734)
);

INVx3_ASAP7_75t_L g2735 ( 
.A(n_2596),
.Y(n_2735)
);

BUFx6f_ASAP7_75t_L g2736 ( 
.A(n_2312),
.Y(n_2736)
);

OA21x2_ASAP7_75t_L g2737 ( 
.A1(n_2326),
.A2(n_1510),
.B(n_1506),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2339),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2569),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2344),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2571),
.Y(n_2741)
);

BUFx6f_ASAP7_75t_L g2742 ( 
.A(n_2316),
.Y(n_2742)
);

BUFx2_ASAP7_75t_L g2743 ( 
.A(n_2486),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2584),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2591),
.Y(n_2745)
);

AND2x4_ASAP7_75t_L g2746 ( 
.A(n_2497),
.B(n_1489),
.Y(n_2746)
);

INVx3_ASAP7_75t_L g2747 ( 
.A(n_2438),
.Y(n_2747)
);

BUFx2_ASAP7_75t_L g2748 ( 
.A(n_2532),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2349),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2309),
.Y(n_2750)
);

CKINVDCx8_ASAP7_75t_R g2751 ( 
.A(n_2597),
.Y(n_2751)
);

HB1xp67_ASAP7_75t_L g2752 ( 
.A(n_2535),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2350),
.Y(n_2753)
);

AND2x2_ASAP7_75t_L g2754 ( 
.A(n_2353),
.B(n_1386),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2351),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2310),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2352),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2562),
.B(n_1386),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2314),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2354),
.Y(n_2760)
);

AND2x4_ASAP7_75t_L g2761 ( 
.A(n_2499),
.B(n_1498),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2363),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2368),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2371),
.Y(n_2764)
);

AND2x4_ASAP7_75t_L g2765 ( 
.A(n_2429),
.B(n_1502),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_SL g2766 ( 
.A(n_2331),
.B(n_1568),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2374),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2550),
.B(n_1571),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2574),
.B(n_1591),
.Y(n_2769)
);

HB1xp67_ASAP7_75t_L g2770 ( 
.A(n_2567),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2566),
.B(n_1597),
.Y(n_2771)
);

BUFx6f_ASAP7_75t_L g2772 ( 
.A(n_2327),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2300),
.B(n_1599),
.Y(n_2773)
);

INVxp67_ASAP7_75t_L g2774 ( 
.A(n_2446),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2375),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2317),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2398),
.Y(n_2777)
);

NAND3xp33_ASAP7_75t_L g2778 ( 
.A(n_2348),
.B(n_1369),
.C(n_1368),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2400),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2410),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2287),
.Y(n_2781)
);

BUFx2_ASAP7_75t_L g2782 ( 
.A(n_2577),
.Y(n_2782)
);

BUFx3_ASAP7_75t_L g2783 ( 
.A(n_2426),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2322),
.Y(n_2784)
);

INVx5_ASAP7_75t_L g2785 ( 
.A(n_2597),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2292),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2295),
.Y(n_2787)
);

INVx2_ASAP7_75t_SL g2788 ( 
.A(n_2579),
.Y(n_2788)
);

INVx3_ASAP7_75t_L g2789 ( 
.A(n_2447),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2496),
.B(n_1449),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2330),
.Y(n_2791)
);

AND2x2_ASAP7_75t_L g2792 ( 
.A(n_2500),
.B(n_1449),
.Y(n_2792)
);

HB1xp67_ASAP7_75t_L g2793 ( 
.A(n_2588),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2323),
.Y(n_2794)
);

INVx1_ASAP7_75t_SL g2795 ( 
.A(n_2418),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2514),
.Y(n_2796)
);

BUFx6f_ASAP7_75t_L g2797 ( 
.A(n_2338),
.Y(n_2797)
);

HB1xp67_ASAP7_75t_L g2798 ( 
.A(n_2589),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2337),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2342),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2592),
.Y(n_2801)
);

INVx1_ASAP7_75t_SL g2802 ( 
.A(n_2278),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2308),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2336),
.Y(n_2804)
);

BUFx6f_ASAP7_75t_L g2805 ( 
.A(n_2383),
.Y(n_2805)
);

OA21x2_ASAP7_75t_L g2806 ( 
.A1(n_2355),
.A2(n_1611),
.B(n_1605),
.Y(n_2806)
);

BUFx6f_ASAP7_75t_L g2807 ( 
.A(n_2385),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2367),
.Y(n_2808)
);

INVx3_ASAP7_75t_L g2809 ( 
.A(n_2521),
.Y(n_2809)
);

AOI22xp5_ASAP7_75t_L g2810 ( 
.A1(n_2502),
.A2(n_1547),
.B1(n_1640),
.B2(n_1431),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2377),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2361),
.B(n_1616),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2391),
.Y(n_2813)
);

OAI22xp5_ASAP7_75t_L g2814 ( 
.A1(n_2325),
.A2(n_1371),
.B1(n_1378),
.B2(n_1377),
.Y(n_2814)
);

OA21x2_ASAP7_75t_L g2815 ( 
.A1(n_2406),
.A2(n_2498),
.B(n_2392),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2345),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2362),
.Y(n_2817)
);

INVx3_ASAP7_75t_L g2818 ( 
.A(n_2468),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2364),
.Y(n_2819)
);

NOR2xp33_ASAP7_75t_L g2820 ( 
.A(n_2564),
.B(n_1380),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2525),
.B(n_1535),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2366),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2373),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2384),
.B(n_1632),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2311),
.B(n_1633),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2382),
.Y(n_2826)
);

INVx3_ASAP7_75t_L g2827 ( 
.A(n_2471),
.Y(n_2827)
);

INVx3_ASAP7_75t_L g2828 ( 
.A(n_2484),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2407),
.Y(n_2829)
);

OA21x2_ASAP7_75t_L g2830 ( 
.A1(n_2346),
.A2(n_1641),
.B(n_1637),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2411),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2485),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2505),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2522),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2531),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2404),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2405),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2296),
.Y(n_2838)
);

BUFx6f_ASAP7_75t_L g2839 ( 
.A(n_2536),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2307),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2557),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2388),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2403),
.Y(n_2843)
);

HB1xp67_ASAP7_75t_L g2844 ( 
.A(n_2303),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2328),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2334),
.Y(n_2846)
);

BUFx2_ASAP7_75t_L g2847 ( 
.A(n_2279),
.Y(n_2847)
);

AND2x2_ASAP7_75t_L g2848 ( 
.A(n_2504),
.B(n_1535),
.Y(n_2848)
);

BUFx6f_ASAP7_75t_L g2849 ( 
.A(n_2455),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2340),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2357),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2489),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2423),
.Y(n_2853)
);

INVx3_ASAP7_75t_L g2854 ( 
.A(n_2455),
.Y(n_2854)
);

AND2x2_ASAP7_75t_L g2855 ( 
.A(n_2544),
.B(n_1546),
.Y(n_2855)
);

NOR2xp33_ASAP7_75t_L g2856 ( 
.A(n_2578),
.B(n_1382),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2424),
.Y(n_2857)
);

AND2x6_ASAP7_75t_L g2858 ( 
.A(n_2396),
.B(n_1354),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2428),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2332),
.B(n_1646),
.Y(n_2860)
);

AND2x2_ASAP7_75t_L g2861 ( 
.A(n_2560),
.B(n_2581),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2388),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2399),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2395),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2395),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2413),
.Y(n_2866)
);

BUFx2_ASAP7_75t_L g2867 ( 
.A(n_2289),
.Y(n_2867)
);

AND2x4_ASAP7_75t_L g2868 ( 
.A(n_2552),
.B(n_1503),
.Y(n_2868)
);

OAI21x1_ASAP7_75t_L g2869 ( 
.A1(n_2516),
.A2(n_1629),
.B(n_1612),
.Y(n_2869)
);

CKINVDCx5p33_ASAP7_75t_R g2870 ( 
.A(n_2299),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2341),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_SL g2872 ( 
.A(n_2595),
.B(n_1648),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2413),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2503),
.Y(n_2874)
);

INVxp67_ASAP7_75t_L g2875 ( 
.A(n_2389),
.Y(n_2875)
);

HB1xp67_ASAP7_75t_L g2876 ( 
.A(n_2318),
.Y(n_2876)
);

OA21x2_ASAP7_75t_L g2877 ( 
.A1(n_2358),
.A2(n_1656),
.B(n_1649),
.Y(n_2877)
);

INVx3_ASAP7_75t_L g2878 ( 
.A(n_2304),
.Y(n_2878)
);

AND2x6_ASAP7_75t_L g2879 ( 
.A(n_2520),
.B(n_1657),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2394),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2372),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2356),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2360),
.Y(n_2883)
);

AND2x2_ASAP7_75t_L g2884 ( 
.A(n_2294),
.B(n_1546),
.Y(n_2884)
);

BUFx2_ASAP7_75t_L g2885 ( 
.A(n_2389),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2598),
.Y(n_2886)
);

AND2x2_ASAP7_75t_L g2887 ( 
.A(n_2297),
.B(n_1675),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2304),
.Y(n_2888)
);

INVx1_ASAP7_75t_SL g2889 ( 
.A(n_2293),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2551),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2433),
.Y(n_2891)
);

INVx3_ASAP7_75t_L g2892 ( 
.A(n_2432),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2430),
.Y(n_2893)
);

BUFx6f_ASAP7_75t_L g2894 ( 
.A(n_2475),
.Y(n_2894)
);

INVxp67_ASAP7_75t_L g2895 ( 
.A(n_2380),
.Y(n_2895)
);

HB1xp67_ASAP7_75t_L g2896 ( 
.A(n_2488),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2417),
.Y(n_2897)
);

BUFx6f_ASAP7_75t_L g2898 ( 
.A(n_2275),
.Y(n_2898)
);

NAND2xp33_ASAP7_75t_SL g2899 ( 
.A(n_2435),
.B(n_1594),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2387),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2524),
.Y(n_2901)
);

OAI22xp5_ASAP7_75t_L g2902 ( 
.A1(n_2460),
.A2(n_1385),
.B1(n_1388),
.B2(n_1387),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2463),
.Y(n_2903)
);

AND2x2_ASAP7_75t_L g2904 ( 
.A(n_2324),
.B(n_1675),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2593),
.Y(n_2905)
);

OA21x2_ASAP7_75t_L g2906 ( 
.A1(n_2493),
.A2(n_1669),
.B(n_1666),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2517),
.B(n_1677),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2445),
.B(n_1692),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2538),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2529),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2381),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2442),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2890),
.B(n_1684),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_2615),
.Y(n_2914)
);

AOI22xp5_ASAP7_75t_L g2915 ( 
.A1(n_2903),
.A2(n_1689),
.B1(n_1693),
.B2(n_1690),
.Y(n_2915)
);

INVx4_ASAP7_75t_L g2916 ( 
.A(n_2619),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2672),
.B(n_1705),
.Y(n_2917)
);

BUFx8_ASAP7_75t_SL g2918 ( 
.A(n_2699),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_SL g2919 ( 
.A(n_2678),
.B(n_1706),
.Y(n_2919)
);

INVx5_ASAP7_75t_L g2920 ( 
.A(n_2894),
.Y(n_2920)
);

AOI22xp5_ASAP7_75t_L g2921 ( 
.A1(n_2909),
.A2(n_1717),
.B1(n_1766),
.B2(n_1748),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2617),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_SL g2923 ( 
.A(n_2785),
.B(n_1774),
.Y(n_2923)
);

AND2x6_ASAP7_75t_L g2924 ( 
.A(n_2886),
.B(n_1657),
.Y(n_2924)
);

BUFx6f_ASAP7_75t_L g2925 ( 
.A(n_2601),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_SL g2926 ( 
.A(n_2785),
.B(n_1777),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2674),
.B(n_1780),
.Y(n_2927)
);

NOR2xp33_ASAP7_75t_SL g2928 ( 
.A(n_2870),
.B(n_2301),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2754),
.B(n_2459),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2600),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_L g2931 ( 
.A(n_2673),
.B(n_2472),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2618),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2693),
.B(n_1787),
.Y(n_2933)
);

CKINVDCx5p33_ASAP7_75t_R g2934 ( 
.A(n_2795),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_SL g2935 ( 
.A(n_2774),
.B(n_2730),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2603),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_SL g2937 ( 
.A(n_2861),
.B(n_1808),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2812),
.B(n_1814),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2609),
.Y(n_2939)
);

AND3x1_ASAP7_75t_L g2940 ( 
.A(n_2810),
.B(n_1528),
.C(n_1513),
.Y(n_2940)
);

BUFx4f_ASAP7_75t_L g2941 ( 
.A(n_2894),
.Y(n_2941)
);

NOR2xp33_ASAP7_75t_SL g2942 ( 
.A(n_2751),
.B(n_2319),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2620),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2629),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2639),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2610),
.Y(n_2946)
);

OAI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2901),
.A2(n_1843),
.B1(n_1853),
.B2(n_1829),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2824),
.B(n_1855),
.Y(n_2948)
);

INVx6_ASAP7_75t_L g2949 ( 
.A(n_2652),
.Y(n_2949)
);

AOI22xp33_ASAP7_75t_L g2950 ( 
.A1(n_2845),
.A2(n_1794),
.B1(n_1964),
.B2(n_1384),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2771),
.B(n_1863),
.Y(n_2951)
);

OR2x6_ASAP7_75t_L g2952 ( 
.A(n_2898),
.B(n_2480),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2732),
.Y(n_2953)
);

INVx2_ASAP7_75t_L g2954 ( 
.A(n_2641),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2644),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_SL g2956 ( 
.A(n_2820),
.B(n_1905),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2733),
.Y(n_2957)
);

INVx4_ASAP7_75t_L g2958 ( 
.A(n_2736),
.Y(n_2958)
);

AOI22xp5_ASAP7_75t_L g2959 ( 
.A1(n_2912),
.A2(n_1924),
.B1(n_1936),
.B2(n_1934),
.Y(n_2959)
);

OR2x6_ASAP7_75t_L g2960 ( 
.A(n_2898),
.B(n_2788),
.Y(n_2960)
);

BUFx10_ASAP7_75t_L g2961 ( 
.A(n_2910),
.Y(n_2961)
);

NOR2xp33_ASAP7_75t_L g2962 ( 
.A(n_2724),
.B(n_2659),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2687),
.B(n_2705),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2708),
.B(n_1940),
.Y(n_2964)
);

INVx4_ASAP7_75t_L g2965 ( 
.A(n_2736),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_SL g2966 ( 
.A(n_2856),
.B(n_1941),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2738),
.Y(n_2967)
);

BUFx2_ASAP7_75t_L g2968 ( 
.A(n_2631),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2740),
.Y(n_2969)
);

INVx4_ASAP7_75t_L g2970 ( 
.A(n_2742),
.Y(n_2970)
);

OAI22xp5_ASAP7_75t_L g2971 ( 
.A1(n_2880),
.A2(n_1954),
.B1(n_1980),
.B2(n_1948),
.Y(n_2971)
);

AO22x2_ASAP7_75t_L g2972 ( 
.A1(n_2897),
.A2(n_2482),
.B1(n_2518),
.B2(n_2286),
.Y(n_2972)
);

NOR2xp33_ASAP7_75t_L g2973 ( 
.A(n_2670),
.B(n_2509),
.Y(n_2973)
);

AND2x4_ASAP7_75t_L g2974 ( 
.A(n_2606),
.B(n_2549),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2749),
.Y(n_2975)
);

AND2x4_ASAP7_75t_L g2976 ( 
.A(n_2625),
.B(n_2572),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_SL g2977 ( 
.A(n_2758),
.B(n_1990),
.Y(n_2977)
);

INVx5_ASAP7_75t_L g2978 ( 
.A(n_2849),
.Y(n_2978)
);

INVx1_ASAP7_75t_SL g2979 ( 
.A(n_2677),
.Y(n_2979)
);

NOR2xp33_ASAP7_75t_L g2980 ( 
.A(n_2643),
.B(n_2369),
.Y(n_2980)
);

AND2x4_ASAP7_75t_L g2981 ( 
.A(n_2747),
.B(n_2420),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2753),
.Y(n_2982)
);

NOR2xp33_ASAP7_75t_L g2983 ( 
.A(n_2844),
.B(n_2401),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2755),
.Y(n_2984)
);

INVx4_ASAP7_75t_SL g2985 ( 
.A(n_2709),
.Y(n_2985)
);

OR2x2_ASAP7_75t_L g2986 ( 
.A(n_2900),
.B(n_1662),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2768),
.B(n_2011),
.Y(n_2987)
);

AND2x4_ASAP7_75t_L g2988 ( 
.A(n_2789),
.B(n_1530),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2769),
.B(n_2025),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_SL g2990 ( 
.A(n_2637),
.B(n_2055),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2757),
.Y(n_2991)
);

OR2x2_ASAP7_75t_L g2992 ( 
.A(n_2743),
.B(n_1679),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2623),
.B(n_2098),
.Y(n_2993)
);

AND2x6_ASAP7_75t_L g2994 ( 
.A(n_2846),
.B(n_1657),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2655),
.Y(n_2995)
);

NOR3xp33_ASAP7_75t_L g2996 ( 
.A(n_2692),
.B(n_1749),
.C(n_1685),
.Y(n_2996)
);

AND2x2_ASAP7_75t_L g2997 ( 
.A(n_2790),
.B(n_1692),
.Y(n_2997)
);

INVx3_ASAP7_75t_L g2998 ( 
.A(n_2601),
.Y(n_2998)
);

BUFx3_ASAP7_75t_L g2999 ( 
.A(n_2602),
.Y(n_2999)
);

AND2x2_ASAP7_75t_L g3000 ( 
.A(n_2792),
.B(n_2821),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2661),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2760),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2773),
.B(n_2100),
.Y(n_3003)
);

HB1xp67_ASAP7_75t_L g3004 ( 
.A(n_2630),
.Y(n_3004)
);

BUFx6f_ASAP7_75t_L g3005 ( 
.A(n_2602),
.Y(n_3005)
);

OR2x2_ASAP7_75t_L g3006 ( 
.A(n_2748),
.B(n_1781),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2762),
.Y(n_3007)
);

AOI22xp5_ASAP7_75t_L g3008 ( 
.A1(n_2891),
.A2(n_2906),
.B1(n_2907),
.B2(n_2877),
.Y(n_3008)
);

INVx2_ASAP7_75t_SL g3009 ( 
.A(n_2628),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_SL g3010 ( 
.A(n_2884),
.B(n_2887),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2651),
.B(n_2102),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_SL g3012 ( 
.A(n_2843),
.B(n_2103),
.Y(n_3012)
);

NOR2xp33_ASAP7_75t_L g3013 ( 
.A(n_2875),
.B(n_2526),
.Y(n_3013)
);

INVx1_ASAP7_75t_SL g3014 ( 
.A(n_2782),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2763),
.Y(n_3015)
);

NOR2xp33_ASAP7_75t_L g3016 ( 
.A(n_2766),
.B(n_2872),
.Y(n_3016)
);

NOR2xp33_ASAP7_75t_L g3017 ( 
.A(n_2876),
.B(n_2573),
.Y(n_3017)
);

INVx2_ASAP7_75t_L g3018 ( 
.A(n_2666),
.Y(n_3018)
);

AND2x6_ASAP7_75t_L g3019 ( 
.A(n_2850),
.B(n_1751),
.Y(n_3019)
);

CKINVDCx16_ASAP7_75t_R g3020 ( 
.A(n_2638),
.Y(n_3020)
);

BUFx3_ASAP7_75t_L g3021 ( 
.A(n_2627),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2679),
.Y(n_3022)
);

AND2x6_ASAP7_75t_L g3023 ( 
.A(n_2851),
.B(n_1751),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2764),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2688),
.Y(n_3025)
);

BUFx3_ASAP7_75t_L g3026 ( 
.A(n_2627),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_SL g3027 ( 
.A(n_2885),
.B(n_2547),
.Y(n_3027)
);

AOI22xp33_ASAP7_75t_L g3028 ( 
.A1(n_2852),
.A2(n_1384),
.B1(n_1691),
.B2(n_1674),
.Y(n_3028)
);

AOI22xp33_ASAP7_75t_L g3029 ( 
.A1(n_2893),
.A2(n_1384),
.B1(n_1741),
.B2(n_1702),
.Y(n_3029)
);

AOI22xp5_ASAP7_75t_L g3030 ( 
.A1(n_2653),
.A2(n_1642),
.B1(n_1661),
.B2(n_1630),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_SL g3031 ( 
.A(n_2676),
.B(n_2590),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2859),
.B(n_1751),
.Y(n_3032)
);

OR2x2_ASAP7_75t_L g3033 ( 
.A(n_2650),
.B(n_1820),
.Y(n_3033)
);

OR2x6_ASAP7_75t_L g3034 ( 
.A(n_2783),
.B(n_1744),
.Y(n_3034)
);

AND2x2_ASAP7_75t_SL g3035 ( 
.A(n_2847),
.B(n_1831),
.Y(n_3035)
);

AND2x2_ASAP7_75t_L g3036 ( 
.A(n_2867),
.B(n_1739),
.Y(n_3036)
);

INVx6_ASAP7_75t_L g3037 ( 
.A(n_2635),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_2689),
.Y(n_3038)
);

INVx5_ASAP7_75t_L g3039 ( 
.A(n_2849),
.Y(n_3039)
);

AND2x2_ASAP7_75t_L g3040 ( 
.A(n_2904),
.B(n_1739),
.Y(n_3040)
);

INVx4_ASAP7_75t_L g3041 ( 
.A(n_2742),
.Y(n_3041)
);

NOR2xp33_ASAP7_75t_SL g3042 ( 
.A(n_2716),
.B(n_1698),
.Y(n_3042)
);

INVx3_ASAP7_75t_L g3043 ( 
.A(n_2635),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_SL g3044 ( 
.A(n_2905),
.B(n_1389),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_SL g3045 ( 
.A(n_2825),
.B(n_1396),
.Y(n_3045)
);

BUFx6f_ASAP7_75t_L g3046 ( 
.A(n_2640),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2767),
.Y(n_3047)
);

NAND3xp33_ASAP7_75t_L g3048 ( 
.A(n_2778),
.B(n_1401),
.C(n_1397),
.Y(n_3048)
);

AND2x2_ASAP7_75t_L g3049 ( 
.A(n_2848),
.B(n_2049),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_SL g3050 ( 
.A(n_2860),
.B(n_1403),
.Y(n_3050)
);

AOI22xp33_ASAP7_75t_L g3051 ( 
.A1(n_2830),
.A2(n_1860),
.B1(n_1890),
.B2(n_1848),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_L g3052 ( 
.A(n_2882),
.B(n_1404),
.Y(n_3052)
);

BUFx10_ASAP7_75t_L g3053 ( 
.A(n_2698),
.Y(n_3053)
);

AND2x2_ASAP7_75t_SL g3054 ( 
.A(n_2908),
.B(n_1913),
.Y(n_3054)
);

NOR2xp33_ASAP7_75t_L g3055 ( 
.A(n_2895),
.B(n_1825),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_SL g3056 ( 
.A(n_2871),
.B(n_1408),
.Y(n_3056)
);

NAND2xp33_ASAP7_75t_SL g3057 ( 
.A(n_2855),
.B(n_1711),
.Y(n_3057)
);

AND2x2_ASAP7_75t_SL g3058 ( 
.A(n_2690),
.B(n_1926),
.Y(n_3058)
);

AOI22xp33_ASAP7_75t_L g3059 ( 
.A1(n_2796),
.A2(n_2801),
.B1(n_2765),
.B2(n_2863),
.Y(n_3059)
);

INVxp67_ASAP7_75t_SL g3060 ( 
.A(n_2883),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2775),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_SL g3062 ( 
.A(n_2611),
.B(n_1415),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_2777),
.B(n_1416),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2779),
.Y(n_3064)
);

NOR2xp33_ASAP7_75t_L g3065 ( 
.A(n_2654),
.B(n_1828),
.Y(n_3065)
);

OR2x2_ASAP7_75t_L g3066 ( 
.A(n_2700),
.B(n_1873),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_2701),
.Y(n_3067)
);

INVx3_ASAP7_75t_L g3068 ( 
.A(n_2640),
.Y(n_3068)
);

OR2x2_ASAP7_75t_L g3069 ( 
.A(n_2710),
.B(n_1897),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_SL g3070 ( 
.A(n_2612),
.B(n_1423),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_SL g3071 ( 
.A(n_2613),
.B(n_1425),
.Y(n_3071)
);

BUFx6f_ASAP7_75t_L g3072 ( 
.A(n_2647),
.Y(n_3072)
);

AND2x4_ASAP7_75t_L g3073 ( 
.A(n_2809),
.B(n_1537),
.Y(n_3073)
);

BUFx2_ASAP7_75t_L g3074 ( 
.A(n_2752),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2780),
.Y(n_3075)
);

BUFx6f_ASAP7_75t_L g3076 ( 
.A(n_2647),
.Y(n_3076)
);

INVxp67_ASAP7_75t_SL g3077 ( 
.A(n_2772),
.Y(n_3077)
);

AOI22xp33_ASAP7_75t_L g3078 ( 
.A1(n_2728),
.A2(n_1933),
.B1(n_1965),
.B2(n_1930),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_2707),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2712),
.B(n_1426),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2715),
.B(n_1428),
.Y(n_3081)
);

BUFx6f_ASAP7_75t_L g3082 ( 
.A(n_2648),
.Y(n_3082)
);

INVx3_ASAP7_75t_L g3083 ( 
.A(n_2648),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_SL g3084 ( 
.A(n_2626),
.B(n_1433),
.Y(n_3084)
);

BUFx3_ASAP7_75t_L g3085 ( 
.A(n_2682),
.Y(n_3085)
);

NAND3xp33_ASAP7_75t_L g3086 ( 
.A(n_2902),
.B(n_1435),
.C(n_1434),
.Y(n_3086)
);

AND2x4_ASAP7_75t_L g3087 ( 
.A(n_2818),
.B(n_1538),
.Y(n_3087)
);

INVx5_ASAP7_75t_L g3088 ( 
.A(n_2682),
.Y(n_3088)
);

BUFx10_ASAP7_75t_L g3089 ( 
.A(n_2746),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2729),
.B(n_1439),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2734),
.B(n_1445),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_SL g3092 ( 
.A(n_2632),
.B(n_1446),
.Y(n_3092)
);

OR2x6_ASAP7_75t_L g3093 ( 
.A(n_2911),
.B(n_1966),
.Y(n_3093)
);

AND2x6_ASAP7_75t_L g3094 ( 
.A(n_2853),
.B(n_1542),
.Y(n_3094)
);

AOI22xp5_ASAP7_75t_L g3095 ( 
.A1(n_2718),
.A2(n_1718),
.B1(n_1747),
.B2(n_1712),
.Y(n_3095)
);

AOI22xp33_ASAP7_75t_L g3096 ( 
.A1(n_2761),
.A2(n_1988),
.B1(n_2071),
.B2(n_1967),
.Y(n_3096)
);

BUFx3_ASAP7_75t_L g3097 ( 
.A(n_2723),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2739),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2741),
.Y(n_3099)
);

INVx2_ASAP7_75t_L g3100 ( 
.A(n_2744),
.Y(n_3100)
);

INVx4_ASAP7_75t_SL g3101 ( 
.A(n_2879),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2745),
.Y(n_3102)
);

NAND2xp33_ASAP7_75t_SL g3103 ( 
.A(n_2668),
.B(n_2896),
.Y(n_3103)
);

AOI22xp33_ASAP7_75t_L g3104 ( 
.A1(n_2869),
.A2(n_2095),
.B1(n_2086),
.B2(n_1554),
.Y(n_3104)
);

INVxp67_ASAP7_75t_SL g3105 ( 
.A(n_2772),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2750),
.B(n_1457),
.Y(n_3106)
);

AND2x2_ASAP7_75t_SL g3107 ( 
.A(n_2770),
.B(n_1545),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_SL g3108 ( 
.A(n_2634),
.B(n_1459),
.Y(n_3108)
);

INVx5_ASAP7_75t_L g3109 ( 
.A(n_2723),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_SL g3110 ( 
.A(n_2791),
.B(n_1460),
.Y(n_3110)
);

INVx4_ASAP7_75t_L g3111 ( 
.A(n_2797),
.Y(n_3111)
);

AOI22xp5_ASAP7_75t_L g3112 ( 
.A1(n_2881),
.A2(n_1792),
.B1(n_1871),
.B2(n_1778),
.Y(n_3112)
);

INVx4_ASAP7_75t_L g3113 ( 
.A(n_2797),
.Y(n_3113)
);

INVx4_ASAP7_75t_L g3114 ( 
.A(n_2805),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2838),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2756),
.Y(n_3116)
);

INVx5_ASAP7_75t_L g3117 ( 
.A(n_2879),
.Y(n_3117)
);

INVx3_ASAP7_75t_L g3118 ( 
.A(n_2839),
.Y(n_3118)
);

INVx2_ASAP7_75t_L g3119 ( 
.A(n_2759),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2776),
.B(n_1467),
.Y(n_3120)
);

BUFx2_ASAP7_75t_L g3121 ( 
.A(n_2793),
.Y(n_3121)
);

AND2x4_ASAP7_75t_L g3122 ( 
.A(n_2827),
.B(n_1561),
.Y(n_3122)
);

BUFx3_ASAP7_75t_L g3123 ( 
.A(n_2805),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2784),
.B(n_1468),
.Y(n_3124)
);

AND2x4_ASAP7_75t_L g3125 ( 
.A(n_2828),
.B(n_1563),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2840),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2794),
.B(n_2799),
.Y(n_3127)
);

INVx1_ASAP7_75t_SL g3128 ( 
.A(n_2798),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2800),
.B(n_1469),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2816),
.Y(n_3130)
);

BUFx6f_ASAP7_75t_L g3131 ( 
.A(n_2839),
.Y(n_3131)
);

NAND2xp33_ASAP7_75t_L g3132 ( 
.A(n_2713),
.B(n_1470),
.Y(n_3132)
);

NAND2xp33_ASAP7_75t_SL g3133 ( 
.A(n_2814),
.B(n_1882),
.Y(n_3133)
);

AOI22xp5_ASAP7_75t_L g3134 ( 
.A1(n_2857),
.A2(n_1911),
.B1(n_1915),
.B2(n_1885),
.Y(n_3134)
);

INVx4_ASAP7_75t_L g3135 ( 
.A(n_2807),
.Y(n_3135)
);

NOR2xp33_ASAP7_75t_L g3136 ( 
.A(n_2645),
.B(n_1904),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2829),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_2817),
.B(n_1471),
.Y(n_3138)
);

AND2x6_ASAP7_75t_L g3139 ( 
.A(n_2646),
.B(n_1575),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2819),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2822),
.Y(n_3141)
);

NAND2xp33_ASAP7_75t_R g3142 ( 
.A(n_2868),
.B(n_1472),
.Y(n_3142)
);

CKINVDCx5p33_ASAP7_75t_R g3143 ( 
.A(n_2727),
.Y(n_3143)
);

INVx4_ASAP7_75t_L g3144 ( 
.A(n_2807),
.Y(n_3144)
);

AND2x2_ASAP7_75t_L g3145 ( 
.A(n_2633),
.B(n_2049),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_2823),
.Y(n_3146)
);

INVx1_ASAP7_75t_SL g3147 ( 
.A(n_2624),
.Y(n_3147)
);

AOI22xp33_ASAP7_75t_L g3148 ( 
.A1(n_2664),
.A2(n_1582),
.B1(n_1589),
.B2(n_1580),
.Y(n_3148)
);

OR2x2_ASAP7_75t_L g3149 ( 
.A(n_2604),
.B(n_1993),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2826),
.Y(n_3150)
);

NOR2xp33_ASAP7_75t_L g3151 ( 
.A(n_2874),
.B(n_2656),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2831),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_2607),
.B(n_2608),
.Y(n_3153)
);

AND2x6_ASAP7_75t_L g3154 ( 
.A(n_2888),
.B(n_1595),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_SL g3155 ( 
.A(n_3000),
.B(n_2803),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_SL g3156 ( 
.A(n_2962),
.B(n_2804),
.Y(n_3156)
);

O2A1O1Ixp5_ASAP7_75t_L g3157 ( 
.A1(n_3016),
.A2(n_2811),
.B(n_2813),
.C(n_2808),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2914),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2963),
.B(n_2713),
.Y(n_3159)
);

NOR2xp67_ASAP7_75t_L g3160 ( 
.A(n_2920),
.B(n_2636),
.Y(n_3160)
);

OR2x6_ASAP7_75t_L g3161 ( 
.A(n_2960),
.B(n_2892),
.Y(n_3161)
);

AOI21xp5_ASAP7_75t_L g3162 ( 
.A1(n_3060),
.A2(n_2806),
.B(n_2737),
.Y(n_3162)
);

INVx2_ASAP7_75t_SL g3163 ( 
.A(n_2968),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_L g3164 ( 
.A(n_2917),
.B(n_2927),
.Y(n_3164)
);

AND2x4_ASAP7_75t_L g3165 ( 
.A(n_2920),
.B(n_2642),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2933),
.B(n_2713),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_SL g3167 ( 
.A(n_3035),
.B(n_2899),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2930),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_SL g3169 ( 
.A(n_3054),
.B(n_2614),
.Y(n_3169)
);

BUFx5_ASAP7_75t_L g3170 ( 
.A(n_2936),
.Y(n_3170)
);

O2A1O1Ixp33_ASAP7_75t_L g3171 ( 
.A1(n_3010),
.A2(n_2939),
.B(n_2953),
.C(n_2946),
.Y(n_3171)
);

BUFx6f_ASAP7_75t_SL g3172 ( 
.A(n_2952),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_SL g3173 ( 
.A(n_2929),
.B(n_2616),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2951),
.B(n_2714),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_2922),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2957),
.Y(n_3176)
);

INVx3_ASAP7_75t_L g3177 ( 
.A(n_2925),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_SL g3178 ( 
.A(n_3058),
.B(n_2622),
.Y(n_3178)
);

AND2x2_ASAP7_75t_L g3179 ( 
.A(n_3055),
.B(n_2997),
.Y(n_3179)
);

OAI22xp33_ASAP7_75t_L g3180 ( 
.A1(n_3008),
.A2(n_2658),
.B1(n_2662),
.B2(n_2657),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2931),
.B(n_2980),
.Y(n_3181)
);

INVx2_ASAP7_75t_SL g3182 ( 
.A(n_3037),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_2967),
.Y(n_3183)
);

NOR2xp33_ASAP7_75t_L g3184 ( 
.A(n_2973),
.B(n_3128),
.Y(n_3184)
);

A2O1A1Ixp33_ASAP7_75t_L g3185 ( 
.A1(n_3065),
.A2(n_2665),
.B(n_2669),
.C(n_2663),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2969),
.Y(n_3186)
);

OR2x6_ASAP7_75t_L g3187 ( 
.A(n_2949),
.B(n_2605),
.Y(n_3187)
);

A2O1A1Ixp33_ASAP7_75t_L g3188 ( 
.A1(n_3059),
.A2(n_2675),
.B(n_2680),
.C(n_2671),
.Y(n_3188)
);

INVx2_ASAP7_75t_SL g3189 ( 
.A(n_3074),
.Y(n_3189)
);

NOR2xp33_ASAP7_75t_L g3190 ( 
.A(n_2934),
.B(n_2802),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2975),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_2964),
.B(n_2714),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2982),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_2987),
.B(n_2714),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2932),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_2989),
.B(n_3003),
.Y(n_3196)
);

INVxp67_ASAP7_75t_SL g3197 ( 
.A(n_2925),
.Y(n_3197)
);

INVx2_ASAP7_75t_SL g3198 ( 
.A(n_3121),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_SL g3199 ( 
.A(n_3107),
.B(n_2681),
.Y(n_3199)
);

OR2x2_ASAP7_75t_SL g3200 ( 
.A(n_3020),
.B(n_2836),
.Y(n_3200)
);

NOR2xp33_ASAP7_75t_L g3201 ( 
.A(n_2979),
.B(n_2889),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_2943),
.Y(n_3202)
);

CKINVDCx5p33_ASAP7_75t_R g3203 ( 
.A(n_2918),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2938),
.B(n_2858),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_SL g3205 ( 
.A(n_3117),
.B(n_2683),
.Y(n_3205)
);

OAI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_2913),
.A2(n_1955),
.B1(n_1985),
.B2(n_1937),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2948),
.B(n_2858),
.Y(n_3207)
);

NAND2xp33_ASAP7_75t_L g3208 ( 
.A(n_3117),
.B(n_2879),
.Y(n_3208)
);

NOR2xp33_ASAP7_75t_L g3209 ( 
.A(n_3014),
.B(n_2685),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2984),
.Y(n_3210)
);

NOR2xp33_ASAP7_75t_L g3211 ( 
.A(n_2992),
.B(n_2686),
.Y(n_3211)
);

INVx2_ASAP7_75t_SL g3212 ( 
.A(n_3088),
.Y(n_3212)
);

AOI22xp5_ASAP7_75t_L g3213 ( 
.A1(n_3133),
.A2(n_2694),
.B1(n_2695),
.B2(n_2691),
.Y(n_3213)
);

AND2x4_ASAP7_75t_L g3214 ( 
.A(n_2985),
.B(n_2837),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_SL g3215 ( 
.A(n_2961),
.B(n_2696),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2991),
.Y(n_3216)
);

NOR2xp67_ASAP7_75t_L g3217 ( 
.A(n_2916),
.B(n_2978),
.Y(n_3217)
);

INVx2_ASAP7_75t_L g3218 ( 
.A(n_2944),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_3002),
.B(n_2858),
.Y(n_3219)
);

NOR2xp33_ASAP7_75t_L g3220 ( 
.A(n_3006),
.B(n_2697),
.Y(n_3220)
);

AND2x2_ASAP7_75t_L g3221 ( 
.A(n_3040),
.B(n_2703),
.Y(n_3221)
);

NOR2x1p5_ASAP7_75t_L g3222 ( 
.A(n_3143),
.B(n_2621),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_3007),
.B(n_2706),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_SL g3224 ( 
.A(n_3009),
.B(n_2711),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_2945),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_3015),
.B(n_2717),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3024),
.Y(n_3227)
);

AOI21xp5_ASAP7_75t_L g3228 ( 
.A1(n_3127),
.A2(n_2815),
.B(n_2721),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_2954),
.Y(n_3229)
);

OR2x6_ASAP7_75t_L g3230 ( 
.A(n_2981),
.B(n_2649),
.Y(n_3230)
);

NOR2xp33_ASAP7_75t_L g3231 ( 
.A(n_3004),
.B(n_2720),
.Y(n_3231)
);

BUFx6f_ASAP7_75t_L g3232 ( 
.A(n_3005),
.Y(n_3232)
);

OAI22xp33_ASAP7_75t_L g3233 ( 
.A1(n_3095),
.A2(n_2986),
.B1(n_3042),
.B2(n_3047),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3061),
.Y(n_3234)
);

HB1xp67_ASAP7_75t_L g3235 ( 
.A(n_3005),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_SL g3236 ( 
.A(n_2915),
.B(n_2722),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_3064),
.B(n_2725),
.Y(n_3237)
);

NAND2x1_ASAP7_75t_L g3238 ( 
.A(n_2924),
.B(n_2726),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_3075),
.B(n_2781),
.Y(n_3239)
);

NAND2xp33_ASAP7_75t_L g3240 ( 
.A(n_3094),
.B(n_2786),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_3136),
.B(n_2787),
.Y(n_3241)
);

BUFx4_ASAP7_75t_L g3242 ( 
.A(n_2941),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_SL g3243 ( 
.A(n_2921),
.B(n_2959),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_2955),
.B(n_2842),
.Y(n_3244)
);

NOR2xp33_ASAP7_75t_L g3245 ( 
.A(n_3033),
.B(n_3066),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_2995),
.B(n_2862),
.Y(n_3246)
);

INVxp33_ASAP7_75t_L g3247 ( 
.A(n_3069),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_3001),
.B(n_2865),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_3018),
.B(n_2864),
.Y(n_3249)
);

INVx4_ASAP7_75t_L g3250 ( 
.A(n_2978),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_3098),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_3099),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3102),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_3022),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_SL g3255 ( 
.A(n_3011),
.B(n_2878),
.Y(n_3255)
);

INVx2_ASAP7_75t_L g3256 ( 
.A(n_3025),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_3038),
.B(n_2832),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_3067),
.B(n_2833),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_SL g3259 ( 
.A(n_3052),
.B(n_2866),
.Y(n_3259)
);

AND2x4_ASAP7_75t_L g3260 ( 
.A(n_3088),
.B(n_2660),
.Y(n_3260)
);

AND2x4_ASAP7_75t_L g3261 ( 
.A(n_3109),
.B(n_2667),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_3079),
.B(n_2834),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_3140),
.Y(n_3263)
);

INVx5_ASAP7_75t_L g3264 ( 
.A(n_3139),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_SL g3265 ( 
.A(n_2993),
.B(n_2873),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3141),
.Y(n_3266)
);

NOR2xp33_ASAP7_75t_L g3267 ( 
.A(n_2935),
.B(n_1987),
.Y(n_3267)
);

INVxp33_ASAP7_75t_L g3268 ( 
.A(n_3036),
.Y(n_3268)
);

NOR2xp33_ASAP7_75t_L g3269 ( 
.A(n_3030),
.B(n_3134),
.Y(n_3269)
);

INVx2_ASAP7_75t_SL g3270 ( 
.A(n_3109),
.Y(n_3270)
);

AOI22xp5_ASAP7_75t_L g3271 ( 
.A1(n_3146),
.A2(n_2841),
.B1(n_2835),
.B2(n_2022),
.Y(n_3271)
);

INVxp67_ASAP7_75t_L g3272 ( 
.A(n_3049),
.Y(n_3272)
);

NOR2xp33_ASAP7_75t_L g3273 ( 
.A(n_3112),
.B(n_1998),
.Y(n_3273)
);

AND2x2_ASAP7_75t_L g3274 ( 
.A(n_3145),
.B(n_2684),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_3100),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3150),
.Y(n_3276)
);

OAI22xp5_ASAP7_75t_L g3277 ( 
.A1(n_2950),
.A2(n_2045),
.B1(n_2054),
.B2(n_2024),
.Y(n_3277)
);

INVx2_ASAP7_75t_SL g3278 ( 
.A(n_3046),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_3116),
.B(n_1474),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_3119),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_SL g3281 ( 
.A(n_3048),
.B(n_2854),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_SL g3282 ( 
.A(n_3151),
.B(n_2091),
.Y(n_3282)
);

AND2x2_ASAP7_75t_L g3283 ( 
.A(n_3149),
.B(n_3153),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_SL g3284 ( 
.A(n_3063),
.B(n_2093),
.Y(n_3284)
);

NOR2xp67_ASAP7_75t_L g3285 ( 
.A(n_3039),
.B(n_2702),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3152),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3137),
.B(n_3130),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3115),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_L g3289 ( 
.A(n_2956),
.B(n_1477),
.Y(n_3289)
);

NOR2xp67_ASAP7_75t_L g3290 ( 
.A(n_3039),
.B(n_2704),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_2966),
.B(n_1480),
.Y(n_3291)
);

NOR2xp67_ASAP7_75t_L g3292 ( 
.A(n_3017),
.B(n_2719),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_3126),
.B(n_1482),
.Y(n_3293)
);

NOR2xp33_ASAP7_75t_L g3294 ( 
.A(n_2947),
.B(n_2731),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3028),
.B(n_1485),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_2990),
.B(n_1487),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_3029),
.B(n_1490),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_3032),
.B(n_1491),
.Y(n_3298)
);

HB1xp67_ASAP7_75t_L g3299 ( 
.A(n_3046),
.Y(n_3299)
);

NAND3xp33_ASAP7_75t_L g3300 ( 
.A(n_2996),
.B(n_1494),
.C(n_1492),
.Y(n_3300)
);

CKINVDCx5p33_ASAP7_75t_R g3301 ( 
.A(n_3147),
.Y(n_3301)
);

INVxp67_ASAP7_75t_SL g3302 ( 
.A(n_3072),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_3080),
.B(n_1497),
.Y(n_3303)
);

OAI22xp5_ASAP7_75t_L g3304 ( 
.A1(n_3104),
.A2(n_1501),
.B1(n_1507),
.B2(n_1500),
.Y(n_3304)
);

BUFx2_ASAP7_75t_L g3305 ( 
.A(n_3072),
.Y(n_3305)
);

BUFx8_ASAP7_75t_L g3306 ( 
.A(n_2974),
.Y(n_3306)
);

AND2x6_ASAP7_75t_L g3307 ( 
.A(n_3013),
.B(n_1596),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_3081),
.B(n_1508),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3087),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_3090),
.B(n_3091),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3122),
.Y(n_3311)
);

OAI22xp33_ASAP7_75t_L g3312 ( 
.A1(n_3138),
.A2(n_1511),
.B1(n_1517),
.B2(n_1509),
.Y(n_3312)
);

INVx2_ASAP7_75t_L g3313 ( 
.A(n_3125),
.Y(n_3313)
);

NOR2xp33_ASAP7_75t_L g3314 ( 
.A(n_2919),
.B(n_2735),
.Y(n_3314)
);

INVx4_ASAP7_75t_L g3315 ( 
.A(n_3076),
.Y(n_3315)
);

BUFx6f_ASAP7_75t_L g3316 ( 
.A(n_3232),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_SL g3317 ( 
.A(n_3181),
.B(n_2928),
.Y(n_3317)
);

INVxp67_ASAP7_75t_SL g3318 ( 
.A(n_3170),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_3179),
.B(n_3094),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3168),
.Y(n_3320)
);

NOR2xp33_ASAP7_75t_L g3321 ( 
.A(n_3184),
.B(n_2983),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3158),
.Y(n_3322)
);

INVx2_ASAP7_75t_L g3323 ( 
.A(n_3175),
.Y(n_3323)
);

AOI22xp5_ASAP7_75t_L g3324 ( 
.A1(n_3269),
.A2(n_3103),
.B1(n_3094),
.B2(n_3057),
.Y(n_3324)
);

OAI22xp5_ASAP7_75t_SL g3325 ( 
.A1(n_3273),
.A2(n_3301),
.B1(n_3267),
.B2(n_2940),
.Y(n_3325)
);

INVxp67_ASAP7_75t_SL g3326 ( 
.A(n_3170),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3176),
.Y(n_3327)
);

AND2x2_ASAP7_75t_L g3328 ( 
.A(n_3245),
.B(n_2976),
.Y(n_3328)
);

NOR2xp33_ASAP7_75t_L g3329 ( 
.A(n_3247),
.B(n_2977),
.Y(n_3329)
);

HB1xp67_ASAP7_75t_L g3330 ( 
.A(n_3189),
.Y(n_3330)
);

AOI22xp33_ASAP7_75t_L g3331 ( 
.A1(n_3243),
.A2(n_3086),
.B1(n_3139),
.B2(n_3051),
.Y(n_3331)
);

INVx2_ASAP7_75t_L g3332 ( 
.A(n_3195),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_SL g3333 ( 
.A(n_3233),
.B(n_2942),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_SL g3334 ( 
.A(n_3241),
.B(n_3106),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3183),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_3164),
.B(n_3139),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_3196),
.B(n_3120),
.Y(n_3337)
);

AOI22xp5_ASAP7_75t_L g3338 ( 
.A1(n_3167),
.A2(n_2937),
.B1(n_3050),
.B2(n_3045),
.Y(n_3338)
);

BUFx6f_ASAP7_75t_L g3339 ( 
.A(n_3232),
.Y(n_3339)
);

BUFx6f_ASAP7_75t_L g3340 ( 
.A(n_3305),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_3310),
.B(n_3186),
.Y(n_3341)
);

INVx2_ASAP7_75t_L g3342 ( 
.A(n_3202),
.Y(n_3342)
);

AOI22xp5_ASAP7_75t_L g3343 ( 
.A1(n_3272),
.A2(n_3012),
.B1(n_3044),
.B2(n_3062),
.Y(n_3343)
);

INVx2_ASAP7_75t_L g3344 ( 
.A(n_3218),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_3191),
.B(n_3124),
.Y(n_3345)
);

NOR2xp33_ASAP7_75t_L g3346 ( 
.A(n_3282),
.B(n_3056),
.Y(n_3346)
);

NOR2xp33_ASAP7_75t_L g3347 ( 
.A(n_3206),
.B(n_3129),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_3193),
.B(n_3148),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3210),
.Y(n_3349)
);

BUFx6f_ASAP7_75t_L g3350 ( 
.A(n_3315),
.Y(n_3350)
);

AOI22xp5_ASAP7_75t_L g3351 ( 
.A1(n_3284),
.A2(n_3071),
.B1(n_3084),
.B2(n_3070),
.Y(n_3351)
);

AOI22xp5_ASAP7_75t_L g3352 ( 
.A1(n_3221),
.A2(n_3108),
.B1(n_3092),
.B2(n_2972),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_SL g3353 ( 
.A(n_3170),
.B(n_3101),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3216),
.Y(n_3354)
);

BUFx8_ASAP7_75t_L g3355 ( 
.A(n_3172),
.Y(n_3355)
);

BUFx3_ASAP7_75t_L g3356 ( 
.A(n_3306),
.Y(n_3356)
);

AOI22xp33_ASAP7_75t_L g3357 ( 
.A1(n_3227),
.A2(n_3110),
.B1(n_3154),
.B2(n_3132),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3234),
.Y(n_3358)
);

CKINVDCx5p33_ASAP7_75t_R g3359 ( 
.A(n_3203),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_SL g3360 ( 
.A(n_3170),
.B(n_3053),
.Y(n_3360)
);

INVx3_ASAP7_75t_L g3361 ( 
.A(n_3250),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_SL g3362 ( 
.A(n_3264),
.B(n_3089),
.Y(n_3362)
);

BUFx6f_ASAP7_75t_L g3363 ( 
.A(n_3260),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_SL g3364 ( 
.A(n_3264),
.B(n_2971),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3263),
.Y(n_3365)
);

OR2x2_ASAP7_75t_L g3366 ( 
.A(n_3198),
.B(n_3118),
.Y(n_3366)
);

AND2x4_ASAP7_75t_L g3367 ( 
.A(n_3165),
.B(n_3123),
.Y(n_3367)
);

HB1xp67_ASAP7_75t_L g3368 ( 
.A(n_3163),
.Y(n_3368)
);

INVx2_ASAP7_75t_SL g3369 ( 
.A(n_3235),
.Y(n_3369)
);

BUFx4f_ASAP7_75t_L g3370 ( 
.A(n_3161),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_3225),
.Y(n_3371)
);

BUFx3_ASAP7_75t_L g3372 ( 
.A(n_3261),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3159),
.B(n_3077),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3211),
.B(n_3105),
.Y(n_3374)
);

NOR2xp33_ASAP7_75t_L g3375 ( 
.A(n_3277),
.B(n_2958),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_3220),
.B(n_3154),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_3266),
.B(n_3154),
.Y(n_3377)
);

OR2x4_ASAP7_75t_L g3378 ( 
.A(n_3190),
.B(n_3076),
.Y(n_3378)
);

INVx4_ASAP7_75t_L g3379 ( 
.A(n_3187),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_3229),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3276),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_3254),
.Y(n_3382)
);

OAI22xp5_ASAP7_75t_L g3383 ( 
.A1(n_3166),
.A2(n_3096),
.B1(n_3078),
.B2(n_2926),
.Y(n_3383)
);

AOI22xp33_ASAP7_75t_L g3384 ( 
.A1(n_3286),
.A2(n_3019),
.B1(n_3023),
.B2(n_2994),
.Y(n_3384)
);

BUFx6f_ASAP7_75t_L g3385 ( 
.A(n_3187),
.Y(n_3385)
);

BUFx6f_ASAP7_75t_L g3386 ( 
.A(n_3278),
.Y(n_3386)
);

INVx3_ASAP7_75t_SL g3387 ( 
.A(n_3161),
.Y(n_3387)
);

BUFx8_ASAP7_75t_SL g3388 ( 
.A(n_3242),
.Y(n_3388)
);

CKINVDCx5p33_ASAP7_75t_R g3389 ( 
.A(n_3201),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3303),
.B(n_2994),
.Y(n_3390)
);

BUFx3_ASAP7_75t_L g3391 ( 
.A(n_3177),
.Y(n_3391)
);

AOI21xp5_ASAP7_75t_L g3392 ( 
.A1(n_3162),
.A2(n_2923),
.B(n_2924),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_SL g3393 ( 
.A(n_3264),
.B(n_3131),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3251),
.Y(n_3394)
);

AOI22xp33_ASAP7_75t_L g3395 ( 
.A1(n_3288),
.A2(n_2994),
.B1(n_3023),
.B2(n_3019),
.Y(n_3395)
);

INVx2_ASAP7_75t_L g3396 ( 
.A(n_3256),
.Y(n_3396)
);

AOI22xp33_ASAP7_75t_L g3397 ( 
.A1(n_3275),
.A2(n_3019),
.B1(n_3023),
.B2(n_2924),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3252),
.Y(n_3398)
);

INVx2_ASAP7_75t_L g3399 ( 
.A(n_3280),
.Y(n_3399)
);

NAND3xp33_ASAP7_75t_SL g3400 ( 
.A(n_3268),
.B(n_3027),
.C(n_3031),
.Y(n_3400)
);

NOR2xp33_ASAP7_75t_L g3401 ( 
.A(n_3283),
.B(n_2965),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3308),
.B(n_3131),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3156),
.B(n_2970),
.Y(n_3403)
);

AOI22xp33_ASAP7_75t_L g3404 ( 
.A1(n_3295),
.A2(n_3073),
.B1(n_2988),
.B2(n_1606),
.Y(n_3404)
);

NOR2xp33_ASAP7_75t_L g3405 ( 
.A(n_3209),
.B(n_3041),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3253),
.Y(n_3406)
);

OR2x4_ASAP7_75t_L g3407 ( 
.A(n_3294),
.B(n_3082),
.Y(n_3407)
);

HB1xp67_ASAP7_75t_L g3408 ( 
.A(n_3299),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_SL g3409 ( 
.A(n_3312),
.B(n_3082),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3223),
.B(n_3111),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3287),
.Y(n_3411)
);

INVx2_ASAP7_75t_SL g3412 ( 
.A(n_3182),
.Y(n_3412)
);

AOI21xp5_ASAP7_75t_L g3413 ( 
.A1(n_3192),
.A2(n_1567),
.B(n_3113),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3226),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3237),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_3239),
.B(n_3114),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3171),
.B(n_3135),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_SL g3418 ( 
.A(n_3289),
.B(n_3144),
.Y(n_3418)
);

AOI22xp33_ASAP7_75t_L g3419 ( 
.A1(n_3297),
.A2(n_1613),
.B1(n_1619),
.B2(n_1598),
.Y(n_3419)
);

OAI21xp33_ASAP7_75t_SL g3420 ( 
.A1(n_3236),
.A2(n_1623),
.B(n_1621),
.Y(n_3420)
);

BUFx6f_ASAP7_75t_L g3421 ( 
.A(n_3214),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_SL g3422 ( 
.A(n_3291),
.B(n_2998),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3257),
.Y(n_3423)
);

AND2x4_ASAP7_75t_L g3424 ( 
.A(n_3313),
.B(n_2999),
.Y(n_3424)
);

INVx2_ASAP7_75t_L g3425 ( 
.A(n_3258),
.Y(n_3425)
);

BUFx6f_ASAP7_75t_L g3426 ( 
.A(n_3212),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3262),
.Y(n_3427)
);

AND2x2_ASAP7_75t_L g3428 ( 
.A(n_3274),
.B(n_3034),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3244),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3246),
.Y(n_3430)
);

AOI22xp5_ASAP7_75t_L g3431 ( 
.A1(n_3199),
.A2(n_3142),
.B1(n_3068),
.B2(n_3083),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_3298),
.B(n_3043),
.Y(n_3432)
);

AND2x6_ASAP7_75t_SL g3433 ( 
.A(n_3230),
.B(n_3093),
.Y(n_3433)
);

INVxp67_ASAP7_75t_SL g3434 ( 
.A(n_3197),
.Y(n_3434)
);

AND2x2_ASAP7_75t_L g3435 ( 
.A(n_3231),
.B(n_3021),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3185),
.B(n_3026),
.Y(n_3436)
);

OAI22xp5_ASAP7_75t_L g3437 ( 
.A1(n_3174),
.A2(n_3097),
.B1(n_3085),
.B2(n_1521),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_3296),
.B(n_1518),
.Y(n_3438)
);

OR2x4_ASAP7_75t_L g3439 ( 
.A(n_3314),
.B(n_1626),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_3307),
.B(n_3155),
.Y(n_3440)
);

BUFx6f_ASAP7_75t_L g3441 ( 
.A(n_3270),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3248),
.Y(n_3442)
);

INVx2_ASAP7_75t_L g3443 ( 
.A(n_3249),
.Y(n_3443)
);

AND2x2_ASAP7_75t_L g3444 ( 
.A(n_3309),
.B(n_2052),
.Y(n_3444)
);

INVx2_ASAP7_75t_L g3445 ( 
.A(n_3157),
.Y(n_3445)
);

AND2x4_ASAP7_75t_L g3446 ( 
.A(n_3230),
.B(n_3222),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3279),
.Y(n_3447)
);

OAI22xp5_ASAP7_75t_SL g3448 ( 
.A1(n_3200),
.A2(n_1526),
.B1(n_1531),
.B2(n_1523),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_SL g3449 ( 
.A(n_3217),
.B(n_1532),
.Y(n_3449)
);

BUFx2_ASAP7_75t_L g3450 ( 
.A(n_3302),
.Y(n_3450)
);

AOI22xp5_ASAP7_75t_L g3451 ( 
.A1(n_3169),
.A2(n_1534),
.B1(n_1536),
.B2(n_1533),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_SL g3452 ( 
.A(n_3389),
.B(n_3271),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_SL g3453 ( 
.A(n_3321),
.B(n_3292),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_SL g3454 ( 
.A(n_3405),
.B(n_3160),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_SL g3455 ( 
.A(n_3328),
.B(n_3300),
.Y(n_3455)
);

NAND2xp33_ASAP7_75t_SL g3456 ( 
.A(n_3317),
.B(n_3333),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_SL g3457 ( 
.A(n_3374),
.B(n_3435),
.Y(n_3457)
);

NAND2xp33_ASAP7_75t_SL g3458 ( 
.A(n_3385),
.B(n_3178),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_SL g3459 ( 
.A(n_3376),
.B(n_3173),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_3414),
.B(n_3307),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_SL g3461 ( 
.A(n_3415),
.B(n_3311),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_SL g3462 ( 
.A(n_3341),
.B(n_3215),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3337),
.B(n_3307),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_SL g3464 ( 
.A(n_3375),
.B(n_3213),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_SL g3465 ( 
.A(n_3325),
.B(n_3194),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_SL g3466 ( 
.A(n_3401),
.B(n_3293),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_SL g3467 ( 
.A(n_3324),
.B(n_3204),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_SL g3468 ( 
.A(n_3410),
.B(n_3207),
.Y(n_3468)
);

AND2x2_ASAP7_75t_L g3469 ( 
.A(n_3443),
.B(n_3224),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3411),
.B(n_3259),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_SL g3471 ( 
.A(n_3416),
.B(n_3219),
.Y(n_3471)
);

NAND2xp33_ASAP7_75t_SL g3472 ( 
.A(n_3385),
.B(n_3205),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3423),
.B(n_3265),
.Y(n_3473)
);

AND2x2_ASAP7_75t_L g3474 ( 
.A(n_3425),
.B(n_3188),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_SL g3475 ( 
.A(n_3347),
.B(n_3304),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_SL g3476 ( 
.A(n_3336),
.B(n_3285),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_SL g3477 ( 
.A(n_3329),
.B(n_3290),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_SL g3478 ( 
.A(n_3346),
.B(n_3180),
.Y(n_3478)
);

AND2x2_ASAP7_75t_L g3479 ( 
.A(n_3427),
.B(n_3281),
.Y(n_3479)
);

NAND2xp33_ASAP7_75t_SL g3480 ( 
.A(n_3350),
.B(n_3255),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_SL g3481 ( 
.A(n_3340),
.B(n_3228),
.Y(n_3481)
);

NAND2xp33_ASAP7_75t_SL g3482 ( 
.A(n_3350),
.B(n_3238),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_SL g3483 ( 
.A(n_3340),
.B(n_2052),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_SL g3484 ( 
.A(n_3319),
.B(n_2072),
.Y(n_3484)
);

NAND2xp33_ASAP7_75t_SL g3485 ( 
.A(n_3316),
.B(n_3208),
.Y(n_3485)
);

AND2x4_ASAP7_75t_L g3486 ( 
.A(n_3446),
.B(n_1628),
.Y(n_3486)
);

AND2x2_ASAP7_75t_L g3487 ( 
.A(n_3428),
.B(n_2072),
.Y(n_3487)
);

OR2x2_ASAP7_75t_L g3488 ( 
.A(n_3330),
.B(n_1539),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_3447),
.B(n_3240),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_SL g3490 ( 
.A(n_3431),
.B(n_1541),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_SL g3491 ( 
.A(n_3370),
.B(n_1543),
.Y(n_3491)
);

AND2x2_ASAP7_75t_L g3492 ( 
.A(n_3429),
.B(n_1544),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3430),
.B(n_1638),
.Y(n_3493)
);

NAND2xp33_ASAP7_75t_SL g3494 ( 
.A(n_3316),
.B(n_3339),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_SL g3495 ( 
.A(n_3368),
.B(n_1548),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_SL g3496 ( 
.A(n_3440),
.B(n_1549),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3442),
.B(n_1645),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_SL g3498 ( 
.A(n_3402),
.B(n_1551),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_SL g3499 ( 
.A(n_3450),
.B(n_1552),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3334),
.B(n_1647),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_SL g3501 ( 
.A(n_3338),
.B(n_1555),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_SL g3502 ( 
.A(n_3352),
.B(n_1556),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_SL g3503 ( 
.A(n_3369),
.B(n_3345),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_SL g3504 ( 
.A(n_3379),
.B(n_1558),
.Y(n_3504)
);

NAND2xp33_ASAP7_75t_SL g3505 ( 
.A(n_3339),
.B(n_1559),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_SL g3506 ( 
.A(n_3424),
.B(n_1566),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_SL g3507 ( 
.A(n_3351),
.B(n_1569),
.Y(n_3507)
);

NAND2xp33_ASAP7_75t_SL g3508 ( 
.A(n_3421),
.B(n_1572),
.Y(n_3508)
);

AND2x4_ASAP7_75t_L g3509 ( 
.A(n_3372),
.B(n_3320),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_SL g3510 ( 
.A(n_3386),
.B(n_1573),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_SL g3511 ( 
.A(n_3386),
.B(n_1577),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_SL g3512 ( 
.A(n_3421),
.B(n_1578),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_SL g3513 ( 
.A(n_3403),
.B(n_1583),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_SL g3514 ( 
.A(n_3343),
.B(n_3331),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3327),
.B(n_1652),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_SL g3516 ( 
.A(n_3438),
.B(n_1585),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_SL g3517 ( 
.A(n_3366),
.B(n_3408),
.Y(n_3517)
);

NAND2xp33_ASAP7_75t_SL g3518 ( 
.A(n_3426),
.B(n_1586),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_SL g3519 ( 
.A(n_3377),
.B(n_1587),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_SL g3520 ( 
.A(n_3357),
.B(n_1588),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_SL g3521 ( 
.A(n_3348),
.B(n_1592),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_SL g3522 ( 
.A(n_3335),
.B(n_1593),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_SL g3523 ( 
.A(n_3349),
.B(n_1603),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_SL g3524 ( 
.A(n_3354),
.B(n_3358),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_SL g3525 ( 
.A(n_3365),
.B(n_1604),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_L g3526 ( 
.A(n_3381),
.B(n_1654),
.Y(n_3526)
);

NOR2xp33_ASAP7_75t_L g3527 ( 
.A(n_3407),
.B(n_1609),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3394),
.B(n_1658),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_SL g3529 ( 
.A(n_3432),
.B(n_3398),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_SL g3530 ( 
.A(n_3406),
.B(n_1610),
.Y(n_3530)
);

NAND2xp33_ASAP7_75t_SL g3531 ( 
.A(n_3426),
.B(n_1614),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_SL g3532 ( 
.A(n_3363),
.B(n_1620),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_SL g3533 ( 
.A(n_3363),
.B(n_3436),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_SL g3534 ( 
.A(n_3404),
.B(n_1624),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_SL g3535 ( 
.A(n_3367),
.B(n_1625),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_SL g3536 ( 
.A(n_3322),
.B(n_1627),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_3373),
.B(n_1659),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_SL g3538 ( 
.A(n_3323),
.B(n_3332),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_SL g3539 ( 
.A(n_3342),
.B(n_1631),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_3419),
.B(n_1660),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_SL g3541 ( 
.A(n_3344),
.B(n_1634),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_SL g3542 ( 
.A(n_3371),
.B(n_1635),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_SL g3543 ( 
.A(n_3380),
.B(n_3382),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_SL g3544 ( 
.A(n_3396),
.B(n_1636),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_SL g3545 ( 
.A(n_3399),
.B(n_3361),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_SL g3546 ( 
.A(n_3417),
.B(n_3441),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3409),
.B(n_1665),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_SL g3548 ( 
.A(n_3441),
.B(n_1639),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3434),
.B(n_1683),
.Y(n_3549)
);

NAND2xp33_ASAP7_75t_SL g3550 ( 
.A(n_3387),
.B(n_1643),
.Y(n_3550)
);

NAND2xp33_ASAP7_75t_SL g3551 ( 
.A(n_3393),
.B(n_1644),
.Y(n_3551)
);

NAND2xp33_ASAP7_75t_SL g3552 ( 
.A(n_3362),
.B(n_1650),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_SL g3553 ( 
.A(n_3390),
.B(n_1651),
.Y(n_3553)
);

AND2x4_ASAP7_75t_L g3554 ( 
.A(n_3391),
.B(n_3412),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_SL g3555 ( 
.A(n_3448),
.B(n_1653),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_3418),
.B(n_1697),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_SL g3557 ( 
.A(n_3444),
.B(n_1655),
.Y(n_3557)
);

OR2x2_ASAP7_75t_L g3558 ( 
.A(n_3437),
.B(n_1667),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3422),
.B(n_1704),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_3383),
.B(n_1707),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_SL g3561 ( 
.A(n_3451),
.B(n_1668),
.Y(n_3561)
);

NAND2xp33_ASAP7_75t_SL g3562 ( 
.A(n_3359),
.B(n_3353),
.Y(n_3562)
);

AOI22xp5_ASAP7_75t_L g3563 ( 
.A1(n_3452),
.A2(n_3400),
.B1(n_3449),
.B2(n_3439),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3457),
.B(n_3378),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3524),
.Y(n_3565)
);

NOR2x1p5_ASAP7_75t_SL g3566 ( 
.A(n_3558),
.B(n_3445),
.Y(n_3566)
);

AOI22xp33_ASAP7_75t_L g3567 ( 
.A1(n_3514),
.A2(n_3364),
.B1(n_3420),
.B2(n_3360),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3479),
.B(n_3433),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_3538),
.Y(n_3569)
);

NAND2xp33_ASAP7_75t_SL g3570 ( 
.A(n_3453),
.B(n_3384),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3492),
.B(n_3413),
.Y(n_3571)
);

OR2x6_ASAP7_75t_L g3572 ( 
.A(n_3554),
.B(n_3356),
.Y(n_3572)
);

INVx2_ASAP7_75t_L g3573 ( 
.A(n_3543),
.Y(n_3573)
);

BUFx4f_ASAP7_75t_L g3574 ( 
.A(n_3554),
.Y(n_3574)
);

BUFx6f_ASAP7_75t_L g3575 ( 
.A(n_3509),
.Y(n_3575)
);

NOR2xp33_ASAP7_75t_SL g3576 ( 
.A(n_3509),
.B(n_3388),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_SL g3577 ( 
.A(n_3463),
.B(n_3318),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3469),
.B(n_3326),
.Y(n_3578)
);

CKINVDCx5p33_ASAP7_75t_R g3579 ( 
.A(n_3562),
.Y(n_3579)
);

CKINVDCx5p33_ASAP7_75t_R g3580 ( 
.A(n_3527),
.Y(n_3580)
);

HB1xp67_ASAP7_75t_L g3581 ( 
.A(n_3517),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3537),
.B(n_1670),
.Y(n_3582)
);

AOI22xp5_ASAP7_75t_L g3583 ( 
.A1(n_3456),
.A2(n_3355),
.B1(n_3395),
.B2(n_1672),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3462),
.B(n_3473),
.Y(n_3584)
);

NAND2x1p5_ASAP7_75t_L g3585 ( 
.A(n_3503),
.B(n_3392),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3470),
.B(n_1671),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3474),
.B(n_1673),
.Y(n_3587)
);

AND2x4_ASAP7_75t_L g3588 ( 
.A(n_3486),
.B(n_3397),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3529),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3466),
.B(n_1678),
.Y(n_3590)
);

BUFx6f_ASAP7_75t_L g3591 ( 
.A(n_3486),
.Y(n_3591)
);

BUFx6f_ASAP7_75t_L g3592 ( 
.A(n_3487),
.Y(n_3592)
);

AND2x2_ASAP7_75t_L g3593 ( 
.A(n_3465),
.B(n_1708),
.Y(n_3593)
);

NOR2xp33_ASAP7_75t_L g3594 ( 
.A(n_3460),
.B(n_1682),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_3478),
.B(n_3493),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_3461),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3497),
.B(n_1686),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3515),
.Y(n_3598)
);

HB1xp67_ASAP7_75t_L g3599 ( 
.A(n_3488),
.Y(n_3599)
);

NAND2x1p5_ASAP7_75t_L g3600 ( 
.A(n_3546),
.B(n_1714),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3526),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_SL g3602 ( 
.A(n_3489),
.B(n_1687),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3528),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_SL g3604 ( 
.A(n_3458),
.B(n_1688),
.Y(n_3604)
);

OR2x2_ASAP7_75t_L g3605 ( 
.A(n_3500),
.B(n_1719),
.Y(n_3605)
);

CKINVDCx16_ASAP7_75t_R g3606 ( 
.A(n_3518),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3464),
.B(n_3549),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3547),
.B(n_1694),
.Y(n_3608)
);

INVx2_ASAP7_75t_L g3609 ( 
.A(n_3533),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3560),
.B(n_1696),
.Y(n_3610)
);

CKINVDCx5p33_ASAP7_75t_R g3611 ( 
.A(n_3531),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_3459),
.B(n_1703),
.Y(n_3612)
);

BUFx4f_ASAP7_75t_L g3613 ( 
.A(n_3494),
.Y(n_3613)
);

NAND2x1p5_ASAP7_75t_L g3614 ( 
.A(n_3477),
.B(n_1721),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3559),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3481),
.Y(n_3616)
);

INVxp67_ASAP7_75t_SL g3617 ( 
.A(n_3545),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3490),
.B(n_1730),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_3557),
.B(n_1731),
.Y(n_3619)
);

INVx2_ASAP7_75t_L g3620 ( 
.A(n_3556),
.Y(n_3620)
);

NOR2xp33_ASAP7_75t_R g3621 ( 
.A(n_3472),
.B(n_1116),
.Y(n_3621)
);

AND2x2_ASAP7_75t_L g3622 ( 
.A(n_3455),
.B(n_1733),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_3475),
.B(n_3521),
.Y(n_3623)
);

CKINVDCx5p33_ASAP7_75t_R g3624 ( 
.A(n_3550),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_3454),
.B(n_3516),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_3502),
.B(n_1710),
.Y(n_3626)
);

BUFx4f_ASAP7_75t_SL g3627 ( 
.A(n_3548),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3501),
.B(n_1713),
.Y(n_3628)
);

INVxp33_ASAP7_75t_L g3629 ( 
.A(n_3495),
.Y(n_3629)
);

INVxp67_ASAP7_75t_L g3630 ( 
.A(n_3499),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_3507),
.B(n_1715),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3498),
.B(n_1716),
.Y(n_3632)
);

AND2x2_ASAP7_75t_L g3633 ( 
.A(n_3561),
.B(n_1735),
.Y(n_3633)
);

INVx2_ASAP7_75t_L g3634 ( 
.A(n_3471),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_L g3635 ( 
.A(n_3540),
.B(n_1722),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3476),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3484),
.B(n_1723),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_SL g3638 ( 
.A(n_3496),
.B(n_1724),
.Y(n_3638)
);

NAND2x1p5_ASAP7_75t_L g3639 ( 
.A(n_3512),
.B(n_1736),
.Y(n_3639)
);

OR2x2_ASAP7_75t_L g3640 ( 
.A(n_3522),
.B(n_1737),
.Y(n_3640)
);

BUFx8_ASAP7_75t_L g3641 ( 
.A(n_3505),
.Y(n_3641)
);

AND2x2_ASAP7_75t_L g3642 ( 
.A(n_3555),
.B(n_1743),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3468),
.B(n_1726),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3513),
.B(n_1727),
.Y(n_3644)
);

AND2x2_ASAP7_75t_L g3645 ( 
.A(n_3534),
.B(n_1752),
.Y(n_3645)
);

INVx2_ASAP7_75t_L g3646 ( 
.A(n_3536),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_3539),
.Y(n_3647)
);

CKINVDCx5p33_ASAP7_75t_R g3648 ( 
.A(n_3508),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3541),
.Y(n_3649)
);

AND3x1_ASAP7_75t_SL g3650 ( 
.A(n_3483),
.B(n_1758),
.C(n_1756),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_L g3651 ( 
.A(n_3523),
.B(n_1728),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3542),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3525),
.B(n_1732),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3530),
.B(n_1734),
.Y(n_3654)
);

AND2x2_ASAP7_75t_L g3655 ( 
.A(n_3506),
.B(n_3520),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3544),
.Y(n_3656)
);

BUFx6f_ASAP7_75t_L g3657 ( 
.A(n_3510),
.Y(n_3657)
);

INVx3_ASAP7_75t_L g3658 ( 
.A(n_3485),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3467),
.B(n_1740),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3553),
.B(n_1742),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3535),
.B(n_1745),
.Y(n_3661)
);

BUFx12f_ASAP7_75t_L g3662 ( 
.A(n_3532),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3519),
.B(n_1750),
.Y(n_3663)
);

BUFx12f_ASAP7_75t_L g3664 ( 
.A(n_3511),
.Y(n_3664)
);

AND2x2_ASAP7_75t_L g3665 ( 
.A(n_3491),
.B(n_1771),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3480),
.Y(n_3666)
);

AOI22xp33_ASAP7_75t_L g3667 ( 
.A1(n_3552),
.A2(n_1786),
.B1(n_1798),
.B2(n_1782),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3504),
.B(n_3551),
.Y(n_3668)
);

AND2x4_ASAP7_75t_L g3669 ( 
.A(n_3482),
.B(n_1799),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_SL g3670 ( 
.A(n_3463),
.B(n_1753),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3524),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_SL g3672 ( 
.A(n_3463),
.B(n_1755),
.Y(n_3672)
);

INVx2_ASAP7_75t_L g3673 ( 
.A(n_3524),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_L g3674 ( 
.A(n_3457),
.B(n_1757),
.Y(n_3674)
);

AND2x2_ASAP7_75t_L g3675 ( 
.A(n_3492),
.B(n_1803),
.Y(n_3675)
);

INVx2_ASAP7_75t_SL g3676 ( 
.A(n_3574),
.Y(n_3676)
);

NOR2xp33_ASAP7_75t_L g3677 ( 
.A(n_3629),
.B(n_1761),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_L g3678 ( 
.A(n_3595),
.B(n_1763),
.Y(n_3678)
);

AO21x2_ASAP7_75t_L g3679 ( 
.A1(n_3616),
.A2(n_3577),
.B(n_3623),
.Y(n_3679)
);

INVx5_ASAP7_75t_L g3680 ( 
.A(n_3592),
.Y(n_3680)
);

AO21x2_ASAP7_75t_L g3681 ( 
.A1(n_3571),
.A2(n_3607),
.B(n_3636),
.Y(n_3681)
);

AOI22xp33_ASAP7_75t_L g3682 ( 
.A1(n_3570),
.A2(n_1809),
.B1(n_1812),
.B2(n_1806),
.Y(n_3682)
);

NOR2xp67_ASAP7_75t_SL g3683 ( 
.A(n_3606),
.B(n_1768),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3569),
.Y(n_3684)
);

OAI21x1_ASAP7_75t_L g3685 ( 
.A1(n_3585),
.A2(n_1826),
.B(n_1815),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3589),
.Y(n_3686)
);

BUFx6f_ASAP7_75t_L g3687 ( 
.A(n_3592),
.Y(n_3687)
);

BUFx2_ASAP7_75t_L g3688 ( 
.A(n_3575),
.Y(n_3688)
);

AND2x2_ASAP7_75t_L g3689 ( 
.A(n_3593),
.B(n_3622),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3565),
.Y(n_3690)
);

INVx6_ASAP7_75t_L g3691 ( 
.A(n_3572),
.Y(n_3691)
);

OAI21x1_ASAP7_75t_L g3692 ( 
.A1(n_3634),
.A2(n_1842),
.B(n_1839),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3671),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3673),
.Y(n_3694)
);

INVx1_ASAP7_75t_SL g3695 ( 
.A(n_3599),
.Y(n_3695)
);

NAND2xp5_ASAP7_75t_L g3696 ( 
.A(n_3584),
.B(n_1770),
.Y(n_3696)
);

OA21x2_ASAP7_75t_L g3697 ( 
.A1(n_3567),
.A2(n_1869),
.B(n_1861),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3609),
.Y(n_3698)
);

BUFx4f_ASAP7_75t_L g3699 ( 
.A(n_3575),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3581),
.Y(n_3700)
);

OAI21x1_ASAP7_75t_L g3701 ( 
.A1(n_3573),
.A2(n_1881),
.B(n_1874),
.Y(n_3701)
);

AO21x2_ASAP7_75t_L g3702 ( 
.A1(n_3625),
.A2(n_1892),
.B(n_1889),
.Y(n_3702)
);

AO21x2_ASAP7_75t_L g3703 ( 
.A1(n_3659),
.A2(n_3672),
.B(n_3670),
.Y(n_3703)
);

AOI22x1_ASAP7_75t_L g3704 ( 
.A1(n_3666),
.A2(n_1785),
.B1(n_1788),
.B2(n_1784),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3596),
.Y(n_3705)
);

AND2x4_ASAP7_75t_L g3706 ( 
.A(n_3572),
.B(n_1117),
.Y(n_3706)
);

INVx3_ASAP7_75t_L g3707 ( 
.A(n_3613),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3620),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_3598),
.Y(n_3709)
);

INVx8_ASAP7_75t_L g3710 ( 
.A(n_3591),
.Y(n_3710)
);

BUFx3_ASAP7_75t_L g3711 ( 
.A(n_3591),
.Y(n_3711)
);

INVx5_ASAP7_75t_L g3712 ( 
.A(n_3662),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3578),
.Y(n_3713)
);

NAND2x1p5_ASAP7_75t_L g3714 ( 
.A(n_3658),
.B(n_1900),
.Y(n_3714)
);

OAI21x1_ASAP7_75t_L g3715 ( 
.A1(n_3600),
.A2(n_1907),
.B(n_1902),
.Y(n_3715)
);

OAI21xp5_ASAP7_75t_L g3716 ( 
.A1(n_3610),
.A2(n_1918),
.B(n_1914),
.Y(n_3716)
);

INVx2_ASAP7_75t_SL g3717 ( 
.A(n_3657),
.Y(n_3717)
);

BUFx3_ASAP7_75t_L g3718 ( 
.A(n_3657),
.Y(n_3718)
);

CKINVDCx16_ASAP7_75t_R g3719 ( 
.A(n_3576),
.Y(n_3719)
);

INVxp67_ASAP7_75t_L g3720 ( 
.A(n_3568),
.Y(n_3720)
);

AOI21x1_ASAP7_75t_L g3721 ( 
.A1(n_3643),
.A2(n_1932),
.B(n_1931),
.Y(n_3721)
);

INVx2_ASAP7_75t_L g3722 ( 
.A(n_3601),
.Y(n_3722)
);

INVx2_ASAP7_75t_SL g3723 ( 
.A(n_3641),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3617),
.Y(n_3724)
);

BUFx2_ASAP7_75t_R g3725 ( 
.A(n_3580),
.Y(n_3725)
);

OA21x2_ASAP7_75t_L g3726 ( 
.A1(n_3563),
.A2(n_1942),
.B(n_1935),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3603),
.B(n_1791),
.Y(n_3727)
);

INVx1_ASAP7_75t_L g3728 ( 
.A(n_3566),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3615),
.B(n_1795),
.Y(n_3729)
);

CKINVDCx6p67_ASAP7_75t_R g3730 ( 
.A(n_3664),
.Y(n_3730)
);

BUFx5_ASAP7_75t_L g3731 ( 
.A(n_3647),
.Y(n_3731)
);

INVx2_ASAP7_75t_L g3732 ( 
.A(n_3646),
.Y(n_3732)
);

INVx1_ASAP7_75t_SL g3733 ( 
.A(n_3564),
.Y(n_3733)
);

INVx2_ASAP7_75t_L g3734 ( 
.A(n_3656),
.Y(n_3734)
);

INVx4_ASAP7_75t_L g3735 ( 
.A(n_3611),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3649),
.Y(n_3736)
);

BUFx2_ASAP7_75t_L g3737 ( 
.A(n_3655),
.Y(n_3737)
);

BUFx4f_ASAP7_75t_L g3738 ( 
.A(n_3614),
.Y(n_3738)
);

BUFx6f_ASAP7_75t_L g3739 ( 
.A(n_3648),
.Y(n_3739)
);

OAI21x1_ASAP7_75t_L g3740 ( 
.A1(n_3602),
.A2(n_1945),
.B(n_1944),
.Y(n_3740)
);

BUFx3_ASAP7_75t_L g3741 ( 
.A(n_3627),
.Y(n_3741)
);

OAI21x1_ASAP7_75t_L g3742 ( 
.A1(n_3668),
.A2(n_3652),
.B(n_3612),
.Y(n_3742)
);

INVx4_ASAP7_75t_L g3743 ( 
.A(n_3624),
.Y(n_3743)
);

BUFx12f_ASAP7_75t_L g3744 ( 
.A(n_3579),
.Y(n_3744)
);

OAI21xp5_ASAP7_75t_L g3745 ( 
.A1(n_3594),
.A2(n_3582),
.B(n_3587),
.Y(n_3745)
);

NAND2x1p5_ASAP7_75t_L g3746 ( 
.A(n_3588),
.B(n_1946),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3618),
.Y(n_3747)
);

CKINVDCx20_ASAP7_75t_R g3748 ( 
.A(n_3650),
.Y(n_3748)
);

BUFx3_ASAP7_75t_L g3749 ( 
.A(n_3675),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_3645),
.Y(n_3750)
);

BUFx6f_ASAP7_75t_L g3751 ( 
.A(n_3665),
.Y(n_3751)
);

INVx2_ASAP7_75t_L g3752 ( 
.A(n_3633),
.Y(n_3752)
);

NAND2x1p5_ASAP7_75t_L g3753 ( 
.A(n_3604),
.B(n_1953),
.Y(n_3753)
);

INVx1_ASAP7_75t_SL g3754 ( 
.A(n_3619),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_3586),
.B(n_1796),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_3674),
.B(n_1797),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_L g3757 ( 
.A(n_3590),
.B(n_1800),
.Y(n_3757)
);

BUFx3_ASAP7_75t_L g3758 ( 
.A(n_3642),
.Y(n_3758)
);

OA21x2_ASAP7_75t_L g3759 ( 
.A1(n_3669),
.A2(n_1971),
.B(n_1957),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3605),
.Y(n_3760)
);

BUFx2_ASAP7_75t_L g3761 ( 
.A(n_3630),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3640),
.Y(n_3762)
);

BUFx12f_ASAP7_75t_L g3763 ( 
.A(n_3639),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3608),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3626),
.Y(n_3765)
);

OAI21x1_ASAP7_75t_L g3766 ( 
.A1(n_3638),
.A2(n_1977),
.B(n_1973),
.Y(n_3766)
);

HB1xp67_ASAP7_75t_L g3767 ( 
.A(n_3621),
.Y(n_3767)
);

CKINVDCx6p67_ASAP7_75t_R g3768 ( 
.A(n_3661),
.Y(n_3768)
);

AO21x2_ASAP7_75t_L g3769 ( 
.A1(n_3637),
.A2(n_1994),
.B(n_1992),
.Y(n_3769)
);

OAI21x1_ASAP7_75t_L g3770 ( 
.A1(n_3628),
.A2(n_2002),
.B(n_2000),
.Y(n_3770)
);

NAND2x1p5_ASAP7_75t_L g3771 ( 
.A(n_3583),
.B(n_2008),
.Y(n_3771)
);

INVx4_ASAP7_75t_L g3772 ( 
.A(n_3667),
.Y(n_3772)
);

INVx8_ASAP7_75t_L g3773 ( 
.A(n_3631),
.Y(n_3773)
);

OAI21xp5_ASAP7_75t_L g3774 ( 
.A1(n_3597),
.A2(n_2016),
.B(n_2013),
.Y(n_3774)
);

OAI21xp5_ASAP7_75t_SL g3775 ( 
.A1(n_3682),
.A2(n_3771),
.B(n_3745),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3690),
.Y(n_3776)
);

INVx2_ASAP7_75t_L g3777 ( 
.A(n_3686),
.Y(n_3777)
);

AOI22xp33_ASAP7_75t_L g3778 ( 
.A1(n_3772),
.A2(n_3660),
.B1(n_3644),
.B2(n_3663),
.Y(n_3778)
);

AOI22xp33_ASAP7_75t_L g3779 ( 
.A1(n_3758),
.A2(n_2030),
.B1(n_2032),
.B2(n_2029),
.Y(n_3779)
);

INVx4_ASAP7_75t_L g3780 ( 
.A(n_3707),
.Y(n_3780)
);

CKINVDCx5p33_ASAP7_75t_R g3781 ( 
.A(n_3725),
.Y(n_3781)
);

BUFx12f_ASAP7_75t_L g3782 ( 
.A(n_3739),
.Y(n_3782)
);

BUFx2_ASAP7_75t_L g3783 ( 
.A(n_3737),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3693),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3713),
.B(n_3635),
.Y(n_3785)
);

AOI22xp33_ASAP7_75t_L g3786 ( 
.A1(n_3749),
.A2(n_2038),
.B1(n_2044),
.B2(n_2036),
.Y(n_3786)
);

BUFx12f_ASAP7_75t_L g3787 ( 
.A(n_3723),
.Y(n_3787)
);

OAI22xp5_ASAP7_75t_L g3788 ( 
.A1(n_3748),
.A2(n_3632),
.B1(n_3653),
.B2(n_3651),
.Y(n_3788)
);

CKINVDCx20_ASAP7_75t_R g3789 ( 
.A(n_3719),
.Y(n_3789)
);

CKINVDCx20_ASAP7_75t_R g3790 ( 
.A(n_3768),
.Y(n_3790)
);

AOI22xp33_ASAP7_75t_SL g3791 ( 
.A1(n_3726),
.A2(n_3654),
.B1(n_2059),
.B2(n_2064),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_3709),
.Y(n_3792)
);

BUFx6f_ASAP7_75t_L g3793 ( 
.A(n_3687),
.Y(n_3793)
);

BUFx12f_ASAP7_75t_L g3794 ( 
.A(n_3751),
.Y(n_3794)
);

OAI22xp33_ASAP7_75t_L g3795 ( 
.A1(n_3746),
.A2(n_2065),
.B1(n_2066),
.B2(n_2047),
.Y(n_3795)
);

OAI22xp5_ASAP7_75t_L g3796 ( 
.A1(n_3714),
.A2(n_1802),
.B1(n_1805),
.B2(n_1801),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3700),
.B(n_1807),
.Y(n_3797)
);

INVx3_ASAP7_75t_L g3798 ( 
.A(n_3718),
.Y(n_3798)
);

INVxp33_ASAP7_75t_L g3799 ( 
.A(n_3767),
.Y(n_3799)
);

BUFx12f_ASAP7_75t_L g3800 ( 
.A(n_3735),
.Y(n_3800)
);

AOI22xp5_ASAP7_75t_L g3801 ( 
.A1(n_3689),
.A2(n_1813),
.B1(n_1816),
.B2(n_1811),
.Y(n_3801)
);

OAI22xp5_ASAP7_75t_L g3802 ( 
.A1(n_3720),
.A2(n_1819),
.B1(n_1821),
.B2(n_1818),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3736),
.Y(n_3803)
);

CKINVDCx11_ASAP7_75t_R g3804 ( 
.A(n_3744),
.Y(n_3804)
);

INVx3_ASAP7_75t_SL g3805 ( 
.A(n_3730),
.Y(n_3805)
);

INVx2_ASAP7_75t_SL g3806 ( 
.A(n_3680),
.Y(n_3806)
);

AOI22xp33_ASAP7_75t_SL g3807 ( 
.A1(n_3702),
.A2(n_2076),
.B1(n_2079),
.B2(n_2074),
.Y(n_3807)
);

OAI22xp33_ASAP7_75t_L g3808 ( 
.A1(n_3754),
.A2(n_1824),
.B1(n_1832),
.B2(n_1822),
.Y(n_3808)
);

AOI22xp33_ASAP7_75t_SL g3809 ( 
.A1(n_3716),
.A2(n_1834),
.B1(n_1836),
.B2(n_1833),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3695),
.B(n_1837),
.Y(n_3810)
);

INVx1_ASAP7_75t_SL g3811 ( 
.A(n_3761),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3724),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3694),
.Y(n_3813)
);

AOI22xp33_ASAP7_75t_L g3814 ( 
.A1(n_3703),
.A2(n_1844),
.B1(n_1845),
.B2(n_1840),
.Y(n_3814)
);

HB1xp67_ASAP7_75t_L g3815 ( 
.A(n_3681),
.Y(n_3815)
);

OAI22xp5_ASAP7_75t_L g3816 ( 
.A1(n_3738),
.A2(n_1851),
.B1(n_1852),
.B2(n_1849),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3722),
.Y(n_3817)
);

AOI22xp33_ASAP7_75t_SL g3818 ( 
.A1(n_3769),
.A2(n_1857),
.B1(n_1859),
.B2(n_1854),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3698),
.Y(n_3819)
);

BUFx12f_ASAP7_75t_L g3820 ( 
.A(n_3763),
.Y(n_3820)
);

INVx2_ASAP7_75t_L g3821 ( 
.A(n_3705),
.Y(n_3821)
);

BUFx2_ASAP7_75t_SL g3822 ( 
.A(n_3680),
.Y(n_3822)
);

AOI22xp33_ASAP7_75t_L g3823 ( 
.A1(n_3774),
.A2(n_1864),
.B1(n_1865),
.B2(n_1862),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_3684),
.Y(n_3824)
);

AOI22xp33_ASAP7_75t_SL g3825 ( 
.A1(n_3697),
.A2(n_1868),
.B1(n_1870),
.B2(n_1867),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_3764),
.B(n_3708),
.Y(n_3826)
);

INVx8_ASAP7_75t_L g3827 ( 
.A(n_3710),
.Y(n_3827)
);

INVx6_ASAP7_75t_L g3828 ( 
.A(n_3743),
.Y(n_3828)
);

AOI22xp5_ASAP7_75t_L g3829 ( 
.A1(n_3759),
.A2(n_1875),
.B1(n_1876),
.B2(n_1872),
.Y(n_3829)
);

OAI21xp33_ASAP7_75t_L g3830 ( 
.A1(n_3677),
.A2(n_1883),
.B(n_1879),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3731),
.Y(n_3831)
);

INVx5_ASAP7_75t_L g3832 ( 
.A(n_3773),
.Y(n_3832)
);

INVx2_ASAP7_75t_L g3833 ( 
.A(n_3732),
.Y(n_3833)
);

BUFx3_ASAP7_75t_L g3834 ( 
.A(n_3741),
.Y(n_3834)
);

BUFx8_ASAP7_75t_L g3835 ( 
.A(n_3688),
.Y(n_3835)
);

CKINVDCx5p33_ASAP7_75t_R g3836 ( 
.A(n_3711),
.Y(n_3836)
);

BUFx3_ASAP7_75t_L g3837 ( 
.A(n_3717),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_3733),
.B(n_1884),
.Y(n_3838)
);

AOI22xp33_ASAP7_75t_L g3839 ( 
.A1(n_3765),
.A2(n_1891),
.B1(n_1893),
.B2(n_1888),
.Y(n_3839)
);

INVx5_ASAP7_75t_L g3840 ( 
.A(n_3691),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3731),
.Y(n_3841)
);

AOI22xp33_ASAP7_75t_L g3842 ( 
.A1(n_3752),
.A2(n_1895),
.B1(n_1896),
.B2(n_1894),
.Y(n_3842)
);

BUFx2_ASAP7_75t_SL g3843 ( 
.A(n_3712),
.Y(n_3843)
);

INVx2_ASAP7_75t_L g3844 ( 
.A(n_3734),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3731),
.Y(n_3845)
);

CKINVDCx11_ASAP7_75t_R g3846 ( 
.A(n_3750),
.Y(n_3846)
);

AOI22xp33_ASAP7_75t_SL g3847 ( 
.A1(n_3747),
.A2(n_1899),
.B1(n_1901),
.B2(n_1898),
.Y(n_3847)
);

OAI21xp5_ASAP7_75t_SL g3848 ( 
.A1(n_3753),
.A2(n_1906),
.B(n_1903),
.Y(n_3848)
);

CKINVDCx6p67_ASAP7_75t_R g3849 ( 
.A(n_3712),
.Y(n_3849)
);

BUFx8_ASAP7_75t_L g3850 ( 
.A(n_3676),
.Y(n_3850)
);

OAI22xp33_ASAP7_75t_L g3851 ( 
.A1(n_3762),
.A2(n_1909),
.B1(n_1910),
.B2(n_1908),
.Y(n_3851)
);

BUFx8_ASAP7_75t_L g3852 ( 
.A(n_3760),
.Y(n_3852)
);

OAI21xp5_ASAP7_75t_SL g3853 ( 
.A1(n_3721),
.A2(n_1917),
.B(n_1916),
.Y(n_3853)
);

AOI22xp33_ASAP7_75t_L g3854 ( 
.A1(n_3742),
.A2(n_1920),
.B1(n_1922),
.B2(n_1919),
.Y(n_3854)
);

BUFx2_ASAP7_75t_L g3855 ( 
.A(n_3699),
.Y(n_3855)
);

OAI22xp5_ASAP7_75t_L g3856 ( 
.A1(n_3678),
.A2(n_1925),
.B1(n_1928),
.B2(n_1923),
.Y(n_3856)
);

INVx2_ASAP7_75t_L g3857 ( 
.A(n_3777),
.Y(n_3857)
);

AO21x1_ASAP7_75t_L g3858 ( 
.A1(n_3775),
.A2(n_3826),
.B(n_3819),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3776),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3812),
.B(n_3679),
.Y(n_3860)
);

INVx2_ASAP7_75t_L g3861 ( 
.A(n_3784),
.Y(n_3861)
);

OA21x2_ASAP7_75t_L g3862 ( 
.A1(n_3831),
.A2(n_3728),
.B(n_3685),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3803),
.Y(n_3863)
);

AO31x2_ASAP7_75t_L g3864 ( 
.A1(n_3841),
.A2(n_3696),
.A3(n_3729),
.B(n_3727),
.Y(n_3864)
);

AND2x2_ASAP7_75t_L g3865 ( 
.A(n_3783),
.B(n_3706),
.Y(n_3865)
);

AOI21xp5_ASAP7_75t_L g3866 ( 
.A1(n_3785),
.A2(n_3770),
.B(n_3755),
.Y(n_3866)
);

AOI22xp33_ASAP7_75t_SL g3867 ( 
.A1(n_3788),
.A2(n_3715),
.B1(n_3740),
.B2(n_3766),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_L g3868 ( 
.A(n_3817),
.B(n_3757),
.Y(n_3868)
);

OAI22xp5_ASAP7_75t_L g3869 ( 
.A1(n_3778),
.A2(n_3756),
.B1(n_3704),
.B2(n_1943),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3813),
.B(n_3692),
.Y(n_3870)
);

AOI21xp5_ASAP7_75t_L g3871 ( 
.A1(n_3815),
.A2(n_3814),
.B(n_3854),
.Y(n_3871)
);

INVx2_ASAP7_75t_L g3872 ( 
.A(n_3792),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3824),
.B(n_3701),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3821),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3833),
.Y(n_3875)
);

BUFx8_ASAP7_75t_L g3876 ( 
.A(n_3787),
.Y(n_3876)
);

AOI22xp33_ASAP7_75t_SL g3877 ( 
.A1(n_3852),
.A2(n_1947),
.B1(n_1949),
.B2(n_1939),
.Y(n_3877)
);

INVx2_ASAP7_75t_L g3878 ( 
.A(n_3844),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3845),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3811),
.B(n_3683),
.Y(n_3880)
);

OAI221xp5_ASAP7_75t_L g3881 ( 
.A1(n_3853),
.A2(n_1958),
.B1(n_1960),
.B2(n_1956),
.C(n_1952),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3797),
.Y(n_3882)
);

NOR2xp33_ASAP7_75t_L g3883 ( 
.A(n_3799),
.B(n_1963),
.Y(n_3883)
);

OA21x2_ASAP7_75t_L g3884 ( 
.A1(n_3829),
.A2(n_1972),
.B(n_1968),
.Y(n_3884)
);

OR2x2_ASAP7_75t_L g3885 ( 
.A(n_3798),
.B(n_0),
.Y(n_3885)
);

INVx2_ASAP7_75t_L g3886 ( 
.A(n_3837),
.Y(n_3886)
);

A2O1A1Ixp33_ASAP7_75t_L g3887 ( 
.A1(n_3848),
.A2(n_2088),
.B(n_2090),
.C(n_2087),
.Y(n_3887)
);

AOI22xp33_ASAP7_75t_L g3888 ( 
.A1(n_3818),
.A2(n_1976),
.B1(n_1978),
.B2(n_1975),
.Y(n_3888)
);

AOI22xp33_ASAP7_75t_L g3889 ( 
.A1(n_3791),
.A2(n_1983),
.B1(n_1989),
.B2(n_1981),
.Y(n_3889)
);

AND2x2_ASAP7_75t_L g3890 ( 
.A(n_3846),
.B(n_0),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_L g3891 ( 
.A(n_3838),
.B(n_1991),
.Y(n_3891)
);

AOI21xp5_ASAP7_75t_L g3892 ( 
.A1(n_3795),
.A2(n_1997),
.B(n_1995),
.Y(n_3892)
);

OA21x2_ASAP7_75t_L g3893 ( 
.A1(n_3810),
.A2(n_2001),
.B(n_1999),
.Y(n_3893)
);

AOI21x1_ASAP7_75t_L g3894 ( 
.A1(n_3856),
.A2(n_2006),
.B(n_2004),
.Y(n_3894)
);

AOI21xp5_ASAP7_75t_L g3895 ( 
.A1(n_3807),
.A2(n_2010),
.B(n_2009),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3843),
.Y(n_3896)
);

AO22x1_ASAP7_75t_L g3897 ( 
.A1(n_3832),
.A2(n_2014),
.B1(n_2017),
.B2(n_2012),
.Y(n_3897)
);

OAI21x1_ASAP7_75t_L g3898 ( 
.A1(n_3779),
.A2(n_1119),
.B(n_1118),
.Y(n_3898)
);

NAND2xp5_ASAP7_75t_L g3899 ( 
.A(n_3840),
.B(n_2018),
.Y(n_3899)
);

AND2x2_ASAP7_75t_L g3900 ( 
.A(n_3840),
.B(n_1),
.Y(n_3900)
);

AO21x2_ASAP7_75t_L g3901 ( 
.A1(n_3808),
.A2(n_3),
.B(n_4),
.Y(n_3901)
);

OA21x2_ASAP7_75t_L g3902 ( 
.A1(n_3806),
.A2(n_3786),
.B(n_3801),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3822),
.Y(n_3903)
);

OR2x2_ASAP7_75t_L g3904 ( 
.A(n_3780),
.B(n_3),
.Y(n_3904)
);

INVx2_ASAP7_75t_L g3905 ( 
.A(n_3832),
.Y(n_3905)
);

OA21x2_ASAP7_75t_L g3906 ( 
.A1(n_3830),
.A2(n_2020),
.B(n_2019),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_SL g3907 ( 
.A(n_3790),
.B(n_2023),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3849),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3851),
.B(n_2026),
.Y(n_3909)
);

HB1xp67_ASAP7_75t_L g3910 ( 
.A(n_3835),
.Y(n_3910)
);

HB1xp67_ASAP7_75t_L g3911 ( 
.A(n_3836),
.Y(n_3911)
);

OAI221xp5_ASAP7_75t_SL g3912 ( 
.A1(n_3823),
.A2(n_2033),
.B1(n_2035),
.B2(n_2031),
.C(n_2028),
.Y(n_3912)
);

OA21x2_ASAP7_75t_L g3913 ( 
.A1(n_3842),
.A2(n_2040),
.B(n_2039),
.Y(n_3913)
);

BUFx2_ASAP7_75t_L g3914 ( 
.A(n_3800),
.Y(n_3914)
);

AOI22xp33_ASAP7_75t_L g3915 ( 
.A1(n_3825),
.A2(n_2042),
.B1(n_2043),
.B2(n_2041),
.Y(n_3915)
);

AND2x2_ASAP7_75t_L g3916 ( 
.A(n_3834),
.B(n_4),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3855),
.Y(n_3917)
);

INVxp67_ASAP7_75t_L g3918 ( 
.A(n_3793),
.Y(n_3918)
);

AND2x2_ASAP7_75t_L g3919 ( 
.A(n_3789),
.B(n_5),
.Y(n_3919)
);

AOI21xp5_ASAP7_75t_L g3920 ( 
.A1(n_3809),
.A2(n_2050),
.B(n_2046),
.Y(n_3920)
);

AOI221xp5_ASAP7_75t_L g3921 ( 
.A1(n_3802),
.A2(n_2078),
.B1(n_2080),
.B2(n_2075),
.C(n_2073),
.Y(n_3921)
);

BUFx8_ASAP7_75t_L g3922 ( 
.A(n_3820),
.Y(n_3922)
);

AOI21xp5_ASAP7_75t_L g3923 ( 
.A1(n_3796),
.A2(n_2053),
.B(n_2051),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_3793),
.Y(n_3924)
);

AOI21xp5_ASAP7_75t_L g3925 ( 
.A1(n_3839),
.A2(n_2058),
.B(n_2057),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3828),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_L g3927 ( 
.A(n_3847),
.B(n_2060),
.Y(n_3927)
);

OAI21xp5_ASAP7_75t_L g3928 ( 
.A1(n_3816),
.A2(n_2062),
.B(n_2061),
.Y(n_3928)
);

INVx2_ASAP7_75t_L g3929 ( 
.A(n_3794),
.Y(n_3929)
);

OAI21xp5_ASAP7_75t_L g3930 ( 
.A1(n_3781),
.A2(n_2069),
.B(n_2067),
.Y(n_3930)
);

OAI22xp5_ASAP7_75t_L g3931 ( 
.A1(n_3805),
.A2(n_2081),
.B1(n_2083),
.B2(n_2070),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3850),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3827),
.B(n_2084),
.Y(n_3933)
);

AOI22xp33_ASAP7_75t_L g3934 ( 
.A1(n_3782),
.A2(n_2096),
.B1(n_2101),
.B2(n_2085),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_3827),
.B(n_2104),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3804),
.Y(n_3936)
);

AND2x4_ASAP7_75t_L g3937 ( 
.A(n_3783),
.B(n_1120),
.Y(n_3937)
);

AOI21xp5_ASAP7_75t_L g3938 ( 
.A1(n_3775),
.A2(n_5),
.B(n_6),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3776),
.Y(n_3939)
);

BUFx6f_ASAP7_75t_L g3940 ( 
.A(n_3924),
.Y(n_3940)
);

AND2x4_ASAP7_75t_L g3941 ( 
.A(n_3896),
.B(n_7),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3874),
.B(n_8),
.Y(n_3942)
);

OR2x2_ASAP7_75t_L g3943 ( 
.A(n_3860),
.B(n_9),
.Y(n_3943)
);

O2A1O1Ixp33_ASAP7_75t_L g3944 ( 
.A1(n_3938),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3859),
.Y(n_3945)
);

OAI22xp33_ASAP7_75t_L g3946 ( 
.A1(n_3871),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_3946)
);

AOI22xp33_ASAP7_75t_L g3947 ( 
.A1(n_3858),
.A2(n_18),
.B1(n_14),
.B2(n_17),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3863),
.Y(n_3948)
);

AND2x2_ASAP7_75t_L g3949 ( 
.A(n_3879),
.B(n_14),
.Y(n_3949)
);

AOI21xp5_ASAP7_75t_L g3950 ( 
.A1(n_3866),
.A2(n_1124),
.B(n_1123),
.Y(n_3950)
);

AOI221xp5_ASAP7_75t_L g3951 ( 
.A1(n_3869),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.C(n_21),
.Y(n_3951)
);

AOI22xp33_ASAP7_75t_L g3952 ( 
.A1(n_3884),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3861),
.Y(n_3953)
);

INVx2_ASAP7_75t_L g3954 ( 
.A(n_3939),
.Y(n_3954)
);

AOI222xp33_ASAP7_75t_L g3955 ( 
.A1(n_3928),
.A2(n_24),
.B1(n_26),
.B2(n_22),
.C1(n_23),
.C2(n_25),
.Y(n_3955)
);

AOI22xp5_ASAP7_75t_L g3956 ( 
.A1(n_3901),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_3956)
);

AOI22xp5_ASAP7_75t_L g3957 ( 
.A1(n_3902),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_3957)
);

INVx2_ASAP7_75t_L g3958 ( 
.A(n_3857),
.Y(n_3958)
);

AOI22xp33_ASAP7_75t_L g3959 ( 
.A1(n_3913),
.A2(n_3867),
.B1(n_3893),
.B2(n_3906),
.Y(n_3959)
);

BUFx6f_ASAP7_75t_L g3960 ( 
.A(n_3914),
.Y(n_3960)
);

AOI22xp33_ASAP7_75t_L g3961 ( 
.A1(n_3881),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_3961)
);

AOI22xp33_ASAP7_75t_L g3962 ( 
.A1(n_3882),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_3962)
);

NAND3xp33_ASAP7_75t_L g3963 ( 
.A(n_3909),
.B(n_35),
.C(n_36),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3875),
.Y(n_3964)
);

NOR2xp33_ASAP7_75t_L g3965 ( 
.A(n_3908),
.B(n_36),
.Y(n_3965)
);

OAI22xp33_ASAP7_75t_L g3966 ( 
.A1(n_3903),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3872),
.Y(n_3967)
);

OAI22xp5_ASAP7_75t_L g3968 ( 
.A1(n_3917),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_3968)
);

OAI22xp33_ASAP7_75t_L g3969 ( 
.A1(n_3905),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_3969)
);

AND2x2_ASAP7_75t_L g3970 ( 
.A(n_3865),
.B(n_42),
.Y(n_3970)
);

OAI221xp5_ASAP7_75t_L g3971 ( 
.A1(n_3877),
.A2(n_46),
.B1(n_43),
.B2(n_45),
.C(n_47),
.Y(n_3971)
);

AOI21xp5_ASAP7_75t_L g3972 ( 
.A1(n_3873),
.A2(n_1128),
.B(n_1125),
.Y(n_3972)
);

AND2x4_ASAP7_75t_L g3973 ( 
.A(n_3886),
.B(n_45),
.Y(n_3973)
);

OAI22xp5_ASAP7_75t_L g3974 ( 
.A1(n_3918),
.A2(n_49),
.B1(n_46),
.B2(n_48),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_3878),
.B(n_48),
.Y(n_3975)
);

OAI221xp5_ASAP7_75t_L g3976 ( 
.A1(n_3930),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.C(n_53),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3870),
.Y(n_3977)
);

AOI22xp33_ASAP7_75t_L g3978 ( 
.A1(n_3880),
.A2(n_55),
.B1(n_50),
.B2(n_51),
.Y(n_3978)
);

INVx2_ASAP7_75t_SL g3979 ( 
.A(n_3932),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3936),
.B(n_55),
.Y(n_3980)
);

NAND2xp5_ASAP7_75t_L g3981 ( 
.A(n_3868),
.B(n_56),
.Y(n_3981)
);

AOI222xp33_ASAP7_75t_L g3982 ( 
.A1(n_3915),
.A2(n_59),
.B1(n_62),
.B2(n_56),
.C1(n_57),
.C2(n_61),
.Y(n_3982)
);

OAI22xp5_ASAP7_75t_L g3983 ( 
.A1(n_3912),
.A2(n_61),
.B1(n_57),
.B2(n_59),
.Y(n_3983)
);

AOI22xp33_ASAP7_75t_L g3984 ( 
.A1(n_3919),
.A2(n_65),
.B1(n_62),
.B2(n_63),
.Y(n_3984)
);

BUFx3_ASAP7_75t_L g3985 ( 
.A(n_3876),
.Y(n_3985)
);

INVx4_ASAP7_75t_L g3986 ( 
.A(n_3911),
.Y(n_3986)
);

OAI221xp5_ASAP7_75t_L g3987 ( 
.A1(n_3927),
.A2(n_67),
.B1(n_63),
.B2(n_66),
.C(n_68),
.Y(n_3987)
);

AOI22xp33_ASAP7_75t_L g3988 ( 
.A1(n_3889),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_3988)
);

AOI21xp5_ASAP7_75t_L g3989 ( 
.A1(n_3887),
.A2(n_1132),
.B(n_1130),
.Y(n_3989)
);

OAI221xp5_ASAP7_75t_L g3990 ( 
.A1(n_3934),
.A2(n_3888),
.B1(n_3923),
.B2(n_3921),
.C(n_3891),
.Y(n_3990)
);

AND2x2_ASAP7_75t_L g3991 ( 
.A(n_3926),
.B(n_69),
.Y(n_3991)
);

AOI22xp33_ASAP7_75t_L g3992 ( 
.A1(n_3883),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_3992)
);

OA21x2_ASAP7_75t_L g3993 ( 
.A1(n_3929),
.A2(n_3899),
.B(n_3910),
.Y(n_3993)
);

CKINVDCx6p67_ASAP7_75t_R g3994 ( 
.A(n_3890),
.Y(n_3994)
);

OAI21x1_ASAP7_75t_L g3995 ( 
.A1(n_3862),
.A2(n_71),
.B(n_72),
.Y(n_3995)
);

OR2x2_ASAP7_75t_L g3996 ( 
.A(n_3864),
.B(n_73),
.Y(n_3996)
);

OAI211xp5_ASAP7_75t_L g3997 ( 
.A1(n_3920),
.A2(n_3925),
.B(n_3894),
.C(n_3892),
.Y(n_3997)
);

INVxp67_ASAP7_75t_L g3998 ( 
.A(n_3904),
.Y(n_3998)
);

AOI22xp33_ASAP7_75t_SL g3999 ( 
.A1(n_3937),
.A2(n_76),
.B1(n_77),
.B2(n_74),
.Y(n_3999)
);

INVx1_ASAP7_75t_SL g4000 ( 
.A(n_3916),
.Y(n_4000)
);

AOI22xp33_ASAP7_75t_L g4001 ( 
.A1(n_3898),
.A2(n_3907),
.B1(n_3900),
.B2(n_3933),
.Y(n_4001)
);

AOI22xp33_ASAP7_75t_L g4002 ( 
.A1(n_3935),
.A2(n_79),
.B1(n_73),
.B2(n_76),
.Y(n_4002)
);

OAI21x1_ASAP7_75t_SL g4003 ( 
.A1(n_3885),
.A2(n_80),
.B(n_82),
.Y(n_4003)
);

AOI22xp33_ASAP7_75t_L g4004 ( 
.A1(n_3922),
.A2(n_83),
.B1(n_80),
.B2(n_82),
.Y(n_4004)
);

AOI22xp33_ASAP7_75t_SL g4005 ( 
.A1(n_3931),
.A2(n_87),
.B1(n_88),
.B2(n_85),
.Y(n_4005)
);

OAI22xp33_ASAP7_75t_L g4006 ( 
.A1(n_3895),
.A2(n_87),
.B1(n_83),
.B2(n_85),
.Y(n_4006)
);

AOI22xp33_ASAP7_75t_SL g4007 ( 
.A1(n_3864),
.A2(n_93),
.B1(n_94),
.B2(n_91),
.Y(n_4007)
);

AND2x4_ASAP7_75t_L g4008 ( 
.A(n_3986),
.B(n_90),
.Y(n_4008)
);

AND2x2_ASAP7_75t_L g4009 ( 
.A(n_3998),
.B(n_3897),
.Y(n_4009)
);

INVx2_ASAP7_75t_L g4010 ( 
.A(n_3954),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3945),
.Y(n_4011)
);

AND2x2_ASAP7_75t_L g4012 ( 
.A(n_3993),
.B(n_91),
.Y(n_4012)
);

AND2x2_ASAP7_75t_L g4013 ( 
.A(n_3940),
.B(n_93),
.Y(n_4013)
);

INVx2_ASAP7_75t_L g4014 ( 
.A(n_3953),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_3948),
.Y(n_4015)
);

AND2x2_ASAP7_75t_L g4016 ( 
.A(n_3940),
.B(n_95),
.Y(n_4016)
);

AND2x2_ASAP7_75t_L g4017 ( 
.A(n_4000),
.B(n_95),
.Y(n_4017)
);

BUFx2_ASAP7_75t_L g4018 ( 
.A(n_3960),
.Y(n_4018)
);

AND2x2_ASAP7_75t_L g4019 ( 
.A(n_3979),
.B(n_96),
.Y(n_4019)
);

AND2x4_ASAP7_75t_L g4020 ( 
.A(n_3960),
.B(n_3964),
.Y(n_4020)
);

INVx2_ASAP7_75t_SL g4021 ( 
.A(n_3985),
.Y(n_4021)
);

AND2x4_ASAP7_75t_L g4022 ( 
.A(n_3958),
.B(n_96),
.Y(n_4022)
);

OA222x2_ASAP7_75t_L g4023 ( 
.A1(n_3996),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.C1(n_101),
.C2(n_103),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3977),
.Y(n_4024)
);

AND2x2_ASAP7_75t_L g4025 ( 
.A(n_3967),
.B(n_98),
.Y(n_4025)
);

BUFx3_ASAP7_75t_L g4026 ( 
.A(n_3994),
.Y(n_4026)
);

HB1xp67_ASAP7_75t_L g4027 ( 
.A(n_3943),
.Y(n_4027)
);

INVx2_ASAP7_75t_L g4028 ( 
.A(n_3949),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_3942),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_3975),
.Y(n_4030)
);

INVx2_ASAP7_75t_L g4031 ( 
.A(n_3995),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3981),
.B(n_98),
.Y(n_4032)
);

HB1xp67_ASAP7_75t_L g4033 ( 
.A(n_3970),
.Y(n_4033)
);

AND2x2_ASAP7_75t_L g4034 ( 
.A(n_3980),
.B(n_101),
.Y(n_4034)
);

AND2x2_ASAP7_75t_L g4035 ( 
.A(n_3941),
.B(n_103),
.Y(n_4035)
);

OAI21xp5_ASAP7_75t_L g4036 ( 
.A1(n_3957),
.A2(n_104),
.B(n_106),
.Y(n_4036)
);

AND2x2_ASAP7_75t_L g4037 ( 
.A(n_4001),
.B(n_3991),
.Y(n_4037)
);

OA21x2_ASAP7_75t_L g4038 ( 
.A1(n_3959),
.A2(n_106),
.B(n_107),
.Y(n_4038)
);

AND2x2_ASAP7_75t_L g4039 ( 
.A(n_3973),
.B(n_107),
.Y(n_4039)
);

OR2x6_ASAP7_75t_SL g4040 ( 
.A(n_3963),
.B(n_108),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_4007),
.B(n_110),
.Y(n_4041)
);

BUFx2_ASAP7_75t_L g4042 ( 
.A(n_3956),
.Y(n_4042)
);

AND2x2_ASAP7_75t_L g4043 ( 
.A(n_3965),
.B(n_111),
.Y(n_4043)
);

INVx3_ASAP7_75t_L g4044 ( 
.A(n_4003),
.Y(n_4044)
);

INVx2_ASAP7_75t_L g4045 ( 
.A(n_3987),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3968),
.Y(n_4046)
);

BUFx2_ASAP7_75t_L g4047 ( 
.A(n_3946),
.Y(n_4047)
);

AO31x2_ASAP7_75t_L g4048 ( 
.A1(n_3950),
.A2(n_113),
.A3(n_111),
.B(n_112),
.Y(n_4048)
);

INVx2_ASAP7_75t_SL g4049 ( 
.A(n_3974),
.Y(n_4049)
);

HB1xp67_ASAP7_75t_L g4050 ( 
.A(n_3947),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_3966),
.Y(n_4051)
);

INVx2_ASAP7_75t_L g4052 ( 
.A(n_3976),
.Y(n_4052)
);

HB1xp67_ASAP7_75t_L g4053 ( 
.A(n_3972),
.Y(n_4053)
);

OR2x2_ASAP7_75t_L g4054 ( 
.A(n_3984),
.B(n_112),
.Y(n_4054)
);

OR2x6_ASAP7_75t_L g4055 ( 
.A(n_3944),
.B(n_116),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_3952),
.B(n_116),
.Y(n_4056)
);

AND2x2_ASAP7_75t_L g4057 ( 
.A(n_3999),
.B(n_3955),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3969),
.Y(n_4058)
);

NOR2xp33_ASAP7_75t_L g4059 ( 
.A(n_3990),
.B(n_117),
.Y(n_4059)
);

AND2x2_ASAP7_75t_L g4060 ( 
.A(n_4004),
.B(n_118),
.Y(n_4060)
);

AND2x2_ASAP7_75t_L g4061 ( 
.A(n_3978),
.B(n_118),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_4006),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_3983),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3962),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_3971),
.Y(n_4065)
);

INVx2_ASAP7_75t_L g4066 ( 
.A(n_3997),
.Y(n_4066)
);

AND2x4_ASAP7_75t_L g4067 ( 
.A(n_3989),
.B(n_119),
.Y(n_4067)
);

OR2x2_ASAP7_75t_L g4068 ( 
.A(n_4002),
.B(n_3992),
.Y(n_4068)
);

AO31x2_ASAP7_75t_L g4069 ( 
.A1(n_3982),
.A2(n_124),
.A3(n_121),
.B(n_122),
.Y(n_4069)
);

AND2x4_ASAP7_75t_SL g4070 ( 
.A(n_3961),
.B(n_121),
.Y(n_4070)
);

AND2x2_ASAP7_75t_L g4071 ( 
.A(n_4005),
.B(n_122),
.Y(n_4071)
);

HB1xp67_ASAP7_75t_L g4072 ( 
.A(n_3951),
.Y(n_4072)
);

OR2x2_ASAP7_75t_L g4073 ( 
.A(n_3988),
.B(n_125),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_L g4074 ( 
.A(n_3943),
.B(n_125),
.Y(n_4074)
);

AND2x4_ASAP7_75t_L g4075 ( 
.A(n_3986),
.B(n_126),
.Y(n_4075)
);

INVx2_ASAP7_75t_L g4076 ( 
.A(n_3954),
.Y(n_4076)
);

OR2x2_ASAP7_75t_L g4077 ( 
.A(n_3977),
.B(n_126),
.Y(n_4077)
);

AND2x2_ASAP7_75t_L g4078 ( 
.A(n_3998),
.B(n_127),
.Y(n_4078)
);

OR2x2_ASAP7_75t_L g4079 ( 
.A(n_3977),
.B(n_128),
.Y(n_4079)
);

CKINVDCx5p33_ASAP7_75t_R g4080 ( 
.A(n_3985),
.Y(n_4080)
);

AOI22xp33_ASAP7_75t_L g4081 ( 
.A1(n_3955),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_4081)
);

INVx1_ASAP7_75t_SL g4082 ( 
.A(n_3994),
.Y(n_4082)
);

AND2x4_ASAP7_75t_L g4083 ( 
.A(n_3986),
.B(n_129),
.Y(n_4083)
);

INVx3_ASAP7_75t_L g4084 ( 
.A(n_3960),
.Y(n_4084)
);

OR2x2_ASAP7_75t_L g4085 ( 
.A(n_3977),
.B(n_130),
.Y(n_4085)
);

AND2x2_ASAP7_75t_L g4086 ( 
.A(n_3998),
.B(n_131),
.Y(n_4086)
);

HB1xp67_ASAP7_75t_L g4087 ( 
.A(n_3977),
.Y(n_4087)
);

OR2x2_ASAP7_75t_L g4088 ( 
.A(n_3977),
.B(n_132),
.Y(n_4088)
);

OR2x2_ASAP7_75t_L g4089 ( 
.A(n_3977),
.B(n_133),
.Y(n_4089)
);

AND2x2_ASAP7_75t_L g4090 ( 
.A(n_3998),
.B(n_133),
.Y(n_4090)
);

AND2x2_ASAP7_75t_L g4091 ( 
.A(n_3998),
.B(n_135),
.Y(n_4091)
);

AND2x2_ASAP7_75t_L g4092 ( 
.A(n_3998),
.B(n_135),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_3945),
.Y(n_4093)
);

INVx2_ASAP7_75t_L g4094 ( 
.A(n_3954),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_3945),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_3945),
.Y(n_4096)
);

BUFx2_ASAP7_75t_L g4097 ( 
.A(n_3993),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_3945),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_3945),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_3943),
.B(n_136),
.Y(n_4100)
);

OR2x2_ASAP7_75t_L g4101 ( 
.A(n_3977),
.B(n_137),
.Y(n_4101)
);

AND2x2_ASAP7_75t_L g4102 ( 
.A(n_3998),
.B(n_137),
.Y(n_4102)
);

OR2x2_ASAP7_75t_SL g4103 ( 
.A(n_3993),
.B(n_138),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3945),
.Y(n_4104)
);

AND2x2_ASAP7_75t_L g4105 ( 
.A(n_3998),
.B(n_140),
.Y(n_4105)
);

AND2x2_ASAP7_75t_L g4106 ( 
.A(n_3998),
.B(n_140),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_3945),
.Y(n_4107)
);

AND2x2_ASAP7_75t_L g4108 ( 
.A(n_3998),
.B(n_141),
.Y(n_4108)
);

AND2x4_ASAP7_75t_SL g4109 ( 
.A(n_3986),
.B(n_141),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_3945),
.Y(n_4110)
);

INVx2_ASAP7_75t_L g4111 ( 
.A(n_3954),
.Y(n_4111)
);

INVx3_ASAP7_75t_L g4112 ( 
.A(n_3960),
.Y(n_4112)
);

OR2x2_ASAP7_75t_L g4113 ( 
.A(n_3977),
.B(n_143),
.Y(n_4113)
);

INVx4_ASAP7_75t_L g4114 ( 
.A(n_3960),
.Y(n_4114)
);

CKINVDCx20_ASAP7_75t_R g4115 ( 
.A(n_3985),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3945),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_L g4117 ( 
.A(n_3943),
.B(n_144),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_SL g4118 ( 
.A(n_3960),
.B(n_144),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_3945),
.Y(n_4119)
);

AND2x2_ASAP7_75t_L g4120 ( 
.A(n_3998),
.B(n_145),
.Y(n_4120)
);

HB1xp67_ASAP7_75t_SL g4121 ( 
.A(n_3985),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_3945),
.Y(n_4122)
);

INVx2_ASAP7_75t_L g4123 ( 
.A(n_3954),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_3945),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_3945),
.Y(n_4125)
);

BUFx2_ASAP7_75t_L g4126 ( 
.A(n_3993),
.Y(n_4126)
);

INVx5_ASAP7_75t_L g4127 ( 
.A(n_4012),
.Y(n_4127)
);

AOI21xp5_ASAP7_75t_L g4128 ( 
.A1(n_4053),
.A2(n_145),
.B(n_146),
.Y(n_4128)
);

OR2x2_ASAP7_75t_L g4129 ( 
.A(n_4027),
.B(n_146),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_4011),
.Y(n_4130)
);

HB1xp67_ASAP7_75t_L g4131 ( 
.A(n_4087),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_4015),
.Y(n_4132)
);

INVx2_ASAP7_75t_L g4133 ( 
.A(n_4018),
.Y(n_4133)
);

INVx2_ASAP7_75t_SL g4134 ( 
.A(n_4026),
.Y(n_4134)
);

OAI211xp5_ASAP7_75t_L g4135 ( 
.A1(n_4072),
.A2(n_4047),
.B(n_4042),
.C(n_4036),
.Y(n_4135)
);

AO21x2_ASAP7_75t_L g4136 ( 
.A1(n_4009),
.A2(n_4059),
.B(n_4078),
.Y(n_4136)
);

INVx4_ASAP7_75t_SL g4137 ( 
.A(n_4021),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_4093),
.Y(n_4138)
);

INVx2_ASAP7_75t_L g4139 ( 
.A(n_4014),
.Y(n_4139)
);

OAI21x1_ASAP7_75t_L g4140 ( 
.A1(n_4031),
.A2(n_147),
.B(n_148),
.Y(n_4140)
);

INVx2_ASAP7_75t_L g4141 ( 
.A(n_4010),
.Y(n_4141)
);

OAI21x1_ASAP7_75t_L g4142 ( 
.A1(n_4024),
.A2(n_147),
.B(n_148),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_4095),
.Y(n_4143)
);

AOI22xp33_ASAP7_75t_L g4144 ( 
.A1(n_4057),
.A2(n_152),
.B1(n_149),
.B2(n_150),
.Y(n_4144)
);

AND2x2_ASAP7_75t_L g4145 ( 
.A(n_4084),
.B(n_149),
.Y(n_4145)
);

CKINVDCx5p33_ASAP7_75t_R g4146 ( 
.A(n_4080),
.Y(n_4146)
);

BUFx12f_ASAP7_75t_L g4147 ( 
.A(n_4008),
.Y(n_4147)
);

A2O1A1Ixp33_ASAP7_75t_L g4148 ( 
.A1(n_4052),
.A2(n_153),
.B(n_150),
.C(n_152),
.Y(n_4148)
);

OR2x2_ASAP7_75t_L g4149 ( 
.A(n_4029),
.B(n_154),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_4096),
.Y(n_4150)
);

HB1xp67_ASAP7_75t_L g4151 ( 
.A(n_4097),
.Y(n_4151)
);

INVxp67_ASAP7_75t_L g4152 ( 
.A(n_4126),
.Y(n_4152)
);

NOR2xp33_ASAP7_75t_L g4153 ( 
.A(n_4121),
.B(n_4066),
.Y(n_4153)
);

AO211x2_ASAP7_75t_L g4154 ( 
.A1(n_4051),
.A2(n_158),
.B(n_155),
.C(n_156),
.Y(n_4154)
);

AO31x2_ASAP7_75t_L g4155 ( 
.A1(n_4114),
.A2(n_159),
.A3(n_155),
.B(n_158),
.Y(n_4155)
);

AND2x2_ASAP7_75t_L g4156 ( 
.A(n_4112),
.B(n_160),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_4098),
.Y(n_4157)
);

OAI21xp33_ASAP7_75t_L g4158 ( 
.A1(n_4055),
.A2(n_160),
.B(n_162),
.Y(n_4158)
);

BUFx3_ASAP7_75t_L g4159 ( 
.A(n_4115),
.Y(n_4159)
);

AOI22xp33_ASAP7_75t_L g4160 ( 
.A1(n_4045),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_4160)
);

AND2x2_ASAP7_75t_L g4161 ( 
.A(n_4033),
.B(n_163),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_4099),
.Y(n_4162)
);

AND2x2_ASAP7_75t_L g4163 ( 
.A(n_4028),
.B(n_164),
.Y(n_4163)
);

INVx1_ASAP7_75t_SL g4164 ( 
.A(n_4082),
.Y(n_4164)
);

HB1xp67_ASAP7_75t_L g4165 ( 
.A(n_4104),
.Y(n_4165)
);

INVxp67_ASAP7_75t_SL g4166 ( 
.A(n_4044),
.Y(n_4166)
);

AO31x2_ASAP7_75t_L g4167 ( 
.A1(n_4062),
.A2(n_167),
.A3(n_165),
.B(n_166),
.Y(n_4167)
);

O2A1O1Ixp33_ASAP7_75t_L g4168 ( 
.A1(n_4050),
.A2(n_168),
.B(n_169),
.C(n_166),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_4107),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_4110),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_4116),
.Y(n_4171)
);

AND2x2_ASAP7_75t_L g4172 ( 
.A(n_4020),
.B(n_165),
.Y(n_4172)
);

BUFx2_ASAP7_75t_L g4173 ( 
.A(n_4103),
.Y(n_4173)
);

INVx2_ASAP7_75t_L g4174 ( 
.A(n_4076),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_4119),
.Y(n_4175)
);

AOI221xp5_ASAP7_75t_L g4176 ( 
.A1(n_4065),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.C(n_171),
.Y(n_4176)
);

AND2x2_ASAP7_75t_L g4177 ( 
.A(n_4037),
.B(n_171),
.Y(n_4177)
);

AOI221xp5_ASAP7_75t_L g4178 ( 
.A1(n_4063),
.A2(n_176),
.B1(n_173),
.B2(n_174),
.C(n_177),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_4122),
.Y(n_4179)
);

INVxp67_ASAP7_75t_L g4180 ( 
.A(n_4040),
.Y(n_4180)
);

OR2x2_ASAP7_75t_L g4181 ( 
.A(n_4030),
.B(n_173),
.Y(n_4181)
);

OAI22xp5_ASAP7_75t_L g4182 ( 
.A1(n_4055),
.A2(n_4081),
.B1(n_4046),
.B2(n_4058),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_4124),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_4125),
.Y(n_4184)
);

BUFx2_ASAP7_75t_L g4185 ( 
.A(n_4075),
.Y(n_4185)
);

NAND3xp33_ASAP7_75t_L g4186 ( 
.A(n_4038),
.B(n_177),
.C(n_178),
.Y(n_4186)
);

AND2x2_ASAP7_75t_L g4187 ( 
.A(n_4094),
.B(n_178),
.Y(n_4187)
);

AND2x4_ASAP7_75t_L g4188 ( 
.A(n_4025),
.B(n_179),
.Y(n_4188)
);

OAI21x1_ASAP7_75t_L g4189 ( 
.A1(n_4111),
.A2(n_179),
.B(n_180),
.Y(n_4189)
);

INVx2_ASAP7_75t_L g4190 ( 
.A(n_4123),
.Y(n_4190)
);

BUFx6f_ASAP7_75t_L g4191 ( 
.A(n_4083),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_4077),
.B(n_180),
.Y(n_4192)
);

INVx2_ASAP7_75t_L g4193 ( 
.A(n_4013),
.Y(n_4193)
);

HB1xp67_ASAP7_75t_L g4194 ( 
.A(n_4079),
.Y(n_4194)
);

NOR2x1p5_ASAP7_75t_L g4195 ( 
.A(n_4041),
.B(n_181),
.Y(n_4195)
);

BUFx2_ASAP7_75t_L g4196 ( 
.A(n_4022),
.Y(n_4196)
);

AND2x2_ASAP7_75t_L g4197 ( 
.A(n_4086),
.B(n_181),
.Y(n_4197)
);

BUFx3_ASAP7_75t_L g4198 ( 
.A(n_4019),
.Y(n_4198)
);

AOI22xp33_ASAP7_75t_SL g4199 ( 
.A1(n_4067),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4085),
.Y(n_4200)
);

INVx2_ASAP7_75t_L g4201 ( 
.A(n_4016),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_4088),
.Y(n_4202)
);

AND2x2_ASAP7_75t_L g4203 ( 
.A(n_4090),
.B(n_182),
.Y(n_4203)
);

AND2x4_ASAP7_75t_L g4204 ( 
.A(n_4091),
.B(n_183),
.Y(n_4204)
);

OR2x6_ASAP7_75t_L g4205 ( 
.A(n_4118),
.B(n_185),
.Y(n_4205)
);

OAI21x1_ASAP7_75t_L g4206 ( 
.A1(n_4089),
.A2(n_185),
.B(n_186),
.Y(n_4206)
);

INVx2_ASAP7_75t_L g4207 ( 
.A(n_4101),
.Y(n_4207)
);

OAI22xp5_ASAP7_75t_L g4208 ( 
.A1(n_4068),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_4208)
);

INVx2_ASAP7_75t_L g4209 ( 
.A(n_4113),
.Y(n_4209)
);

OAI21xp33_ASAP7_75t_L g4210 ( 
.A1(n_4056),
.A2(n_187),
.B(n_189),
.Y(n_4210)
);

INVx2_ASAP7_75t_L g4211 ( 
.A(n_4049),
.Y(n_4211)
);

HB1xp67_ASAP7_75t_L g4212 ( 
.A(n_4092),
.Y(n_4212)
);

AO31x2_ASAP7_75t_L g4213 ( 
.A1(n_4023),
.A2(n_193),
.A3(n_190),
.B(n_192),
.Y(n_4213)
);

OAI221xp5_ASAP7_75t_L g4214 ( 
.A1(n_4064),
.A2(n_193),
.B1(n_190),
.B2(n_192),
.C(n_194),
.Y(n_4214)
);

OAI21x1_ASAP7_75t_L g4215 ( 
.A1(n_4074),
.A2(n_195),
.B(n_196),
.Y(n_4215)
);

OAI21x1_ASAP7_75t_L g4216 ( 
.A1(n_4100),
.A2(n_196),
.B(n_197),
.Y(n_4216)
);

OA21x2_ASAP7_75t_L g4217 ( 
.A1(n_4117),
.A2(n_197),
.B(n_199),
.Y(n_4217)
);

HB1xp67_ASAP7_75t_L g4218 ( 
.A(n_4102),
.Y(n_4218)
);

INVx2_ASAP7_75t_L g4219 ( 
.A(n_4105),
.Y(n_4219)
);

AOI221xp5_ASAP7_75t_L g4220 ( 
.A1(n_4071),
.A2(n_4060),
.B1(n_4061),
.B2(n_4032),
.C(n_4043),
.Y(n_4220)
);

NOR2xp33_ASAP7_75t_SL g4221 ( 
.A(n_4109),
.B(n_200),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_4106),
.B(n_200),
.Y(n_4222)
);

INVx2_ASAP7_75t_L g4223 ( 
.A(n_4108),
.Y(n_4223)
);

INVx2_ASAP7_75t_L g4224 ( 
.A(n_4120),
.Y(n_4224)
);

AO21x2_ASAP7_75t_L g4225 ( 
.A1(n_4017),
.A2(n_201),
.B(n_202),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4048),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_4048),
.Y(n_4227)
);

BUFx6f_ASAP7_75t_L g4228 ( 
.A(n_4035),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_4039),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4069),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4069),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_4034),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_4054),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_4073),
.Y(n_4234)
);

AO31x2_ASAP7_75t_L g4235 ( 
.A1(n_4070),
.A2(n_204),
.A3(n_201),
.B(n_203),
.Y(n_4235)
);

BUFx3_ASAP7_75t_L g4236 ( 
.A(n_4115),
.Y(n_4236)
);

INVx2_ASAP7_75t_L g4237 ( 
.A(n_4018),
.Y(n_4237)
);

BUFx2_ASAP7_75t_L g4238 ( 
.A(n_4026),
.Y(n_4238)
);

INVx2_ASAP7_75t_L g4239 ( 
.A(n_4018),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_4011),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_L g4241 ( 
.A(n_4066),
.B(n_204),
.Y(n_4241)
);

INVxp67_ASAP7_75t_L g4242 ( 
.A(n_4097),
.Y(n_4242)
);

AND2x2_ASAP7_75t_L g4243 ( 
.A(n_4018),
.B(n_205),
.Y(n_4243)
);

AOI22xp33_ASAP7_75t_SL g4244 ( 
.A1(n_4042),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_4244)
);

AO31x2_ASAP7_75t_L g4245 ( 
.A1(n_4097),
.A2(n_208),
.A3(n_206),
.B(n_207),
.Y(n_4245)
);

INVx1_ASAP7_75t_SL g4246 ( 
.A(n_4121),
.Y(n_4246)
);

AND2x2_ASAP7_75t_L g4247 ( 
.A(n_4018),
.B(n_208),
.Y(n_4247)
);

AO21x2_ASAP7_75t_L g4248 ( 
.A1(n_4012),
.A2(n_209),
.B(n_210),
.Y(n_4248)
);

INVx2_ASAP7_75t_L g4249 ( 
.A(n_4018),
.Y(n_4249)
);

INVx2_ASAP7_75t_L g4250 ( 
.A(n_4018),
.Y(n_4250)
);

AND2x2_ASAP7_75t_L g4251 ( 
.A(n_4018),
.B(n_211),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_4011),
.Y(n_4252)
);

AOI21xp33_ASAP7_75t_L g4253 ( 
.A1(n_4072),
.A2(n_211),
.B(n_212),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_4018),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_L g4255 ( 
.A(n_4066),
.B(n_212),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4011),
.Y(n_4256)
);

AND2x4_ASAP7_75t_L g4257 ( 
.A(n_4114),
.B(n_213),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_4011),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_4011),
.Y(n_4259)
);

AND2x2_ASAP7_75t_L g4260 ( 
.A(n_4018),
.B(n_214),
.Y(n_4260)
);

AND2x2_ASAP7_75t_L g4261 ( 
.A(n_4018),
.B(n_215),
.Y(n_4261)
);

INVx2_ASAP7_75t_L g4262 ( 
.A(n_4018),
.Y(n_4262)
);

HB1xp67_ASAP7_75t_L g4263 ( 
.A(n_4087),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_L g4264 ( 
.A(n_4066),
.B(n_215),
.Y(n_4264)
);

AND2x2_ASAP7_75t_L g4265 ( 
.A(n_4018),
.B(n_216),
.Y(n_4265)
);

OAI22xp5_ASAP7_75t_L g4266 ( 
.A1(n_4103),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_4266)
);

INVx2_ASAP7_75t_L g4267 ( 
.A(n_4018),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4011),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_4066),
.B(n_218),
.Y(n_4269)
);

INVxp67_ASAP7_75t_L g4270 ( 
.A(n_4097),
.Y(n_4270)
);

AO21x2_ASAP7_75t_L g4271 ( 
.A1(n_4012),
.A2(n_219),
.B(n_220),
.Y(n_4271)
);

INVx2_ASAP7_75t_L g4272 ( 
.A(n_4018),
.Y(n_4272)
);

INVx2_ASAP7_75t_L g4273 ( 
.A(n_4018),
.Y(n_4273)
);

INVx2_ASAP7_75t_L g4274 ( 
.A(n_4018),
.Y(n_4274)
);

NOR2xp67_ASAP7_75t_L g4275 ( 
.A(n_4044),
.B(n_220),
.Y(n_4275)
);

OA21x2_ASAP7_75t_L g4276 ( 
.A1(n_4097),
.A2(n_221),
.B(n_222),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4011),
.Y(n_4277)
);

NOR2xp33_ASAP7_75t_R g4278 ( 
.A(n_4121),
.B(n_222),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_4066),
.B(n_221),
.Y(n_4279)
);

BUFx2_ASAP7_75t_L g4280 ( 
.A(n_4026),
.Y(n_4280)
);

AND2x2_ASAP7_75t_L g4281 ( 
.A(n_4018),
.B(n_223),
.Y(n_4281)
);

AOI22xp33_ASAP7_75t_SL g4282 ( 
.A1(n_4042),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_4282)
);

HB1xp67_ASAP7_75t_L g4283 ( 
.A(n_4087),
.Y(n_4283)
);

AND2x4_ASAP7_75t_L g4284 ( 
.A(n_4114),
.B(n_224),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_4018),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_SL g4286 ( 
.A(n_4066),
.B(n_225),
.Y(n_4286)
);

OR2x2_ASAP7_75t_L g4287 ( 
.A(n_4027),
.B(n_226),
.Y(n_4287)
);

BUFx3_ASAP7_75t_L g4288 ( 
.A(n_4115),
.Y(n_4288)
);

INVxp33_ASAP7_75t_L g4289 ( 
.A(n_4278),
.Y(n_4289)
);

BUFx3_ASAP7_75t_L g4290 ( 
.A(n_4159),
.Y(n_4290)
);

AND2x2_ASAP7_75t_L g4291 ( 
.A(n_4137),
.B(n_226),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4165),
.Y(n_4292)
);

INVx2_ASAP7_75t_L g4293 ( 
.A(n_4238),
.Y(n_4293)
);

AND2x4_ASAP7_75t_L g4294 ( 
.A(n_4280),
.B(n_227),
.Y(n_4294)
);

OR2x2_ASAP7_75t_L g4295 ( 
.A(n_4230),
.B(n_227),
.Y(n_4295)
);

OAI221xp5_ASAP7_75t_L g4296 ( 
.A1(n_4135),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.C(n_231),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_4173),
.B(n_4231),
.Y(n_4297)
);

INVx1_ASAP7_75t_SL g4298 ( 
.A(n_4246),
.Y(n_4298)
);

AND2x2_ASAP7_75t_L g4299 ( 
.A(n_4211),
.B(n_228),
.Y(n_4299)
);

AND2x2_ASAP7_75t_L g4300 ( 
.A(n_4133),
.B(n_229),
.Y(n_4300)
);

INVx1_ASAP7_75t_SL g4301 ( 
.A(n_4164),
.Y(n_4301)
);

AND2x4_ASAP7_75t_L g4302 ( 
.A(n_4134),
.B(n_230),
.Y(n_4302)
);

AND2x2_ASAP7_75t_L g4303 ( 
.A(n_4237),
.B(n_232),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4130),
.Y(n_4304)
);

OAI211xp5_ASAP7_75t_SL g4305 ( 
.A1(n_4180),
.A2(n_235),
.B(n_233),
.C(n_234),
.Y(n_4305)
);

AND2x4_ASAP7_75t_L g4306 ( 
.A(n_4239),
.B(n_235),
.Y(n_4306)
);

AND2x2_ASAP7_75t_L g4307 ( 
.A(n_4249),
.B(n_237),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_L g4308 ( 
.A(n_4127),
.B(n_4136),
.Y(n_4308)
);

AND2x2_ASAP7_75t_L g4309 ( 
.A(n_4250),
.B(n_4254),
.Y(n_4309)
);

HB1xp67_ASAP7_75t_L g4310 ( 
.A(n_4151),
.Y(n_4310)
);

AND2x2_ASAP7_75t_L g4311 ( 
.A(n_4262),
.B(n_237),
.Y(n_4311)
);

INVx3_ASAP7_75t_L g4312 ( 
.A(n_4191),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4132),
.Y(n_4313)
);

NAND3xp33_ASAP7_75t_L g4314 ( 
.A(n_4176),
.B(n_4178),
.C(n_4186),
.Y(n_4314)
);

OR2x2_ASAP7_75t_L g4315 ( 
.A(n_4207),
.B(n_238),
.Y(n_4315)
);

AND2x2_ASAP7_75t_L g4316 ( 
.A(n_4267),
.B(n_238),
.Y(n_4316)
);

BUFx3_ASAP7_75t_L g4317 ( 
.A(n_4236),
.Y(n_4317)
);

OAI22xp5_ASAP7_75t_L g4318 ( 
.A1(n_4127),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_4138),
.Y(n_4319)
);

INVx2_ASAP7_75t_L g4320 ( 
.A(n_4185),
.Y(n_4320)
);

OAI22xp5_ASAP7_75t_SL g4321 ( 
.A1(n_4205),
.A2(n_242),
.B1(n_239),
.B2(n_241),
.Y(n_4321)
);

NOR2x1_ASAP7_75t_L g4322 ( 
.A(n_4276),
.B(n_242),
.Y(n_4322)
);

INVx2_ASAP7_75t_SL g4323 ( 
.A(n_4191),
.Y(n_4323)
);

INVx2_ASAP7_75t_L g4324 ( 
.A(n_4228),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_4143),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4150),
.Y(n_4326)
);

OR2x2_ASAP7_75t_L g4327 ( 
.A(n_4209),
.B(n_243),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4157),
.Y(n_4328)
);

AND2x2_ASAP7_75t_L g4329 ( 
.A(n_4272),
.B(n_243),
.Y(n_4329)
);

OR2x2_ASAP7_75t_L g4330 ( 
.A(n_4212),
.B(n_244),
.Y(n_4330)
);

AOI221xp5_ASAP7_75t_L g4331 ( 
.A1(n_4182),
.A2(n_4266),
.B1(n_4168),
.B2(n_4242),
.C(n_4152),
.Y(n_4331)
);

HB1xp67_ASAP7_75t_L g4332 ( 
.A(n_4131),
.Y(n_4332)
);

BUFx3_ASAP7_75t_L g4333 ( 
.A(n_4288),
.Y(n_4333)
);

AND2x2_ASAP7_75t_L g4334 ( 
.A(n_4273),
.B(n_245),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_4162),
.Y(n_4335)
);

AND2x2_ASAP7_75t_L g4336 ( 
.A(n_4274),
.B(n_4285),
.Y(n_4336)
);

OR2x2_ASAP7_75t_L g4337 ( 
.A(n_4218),
.B(n_246),
.Y(n_4337)
);

BUFx3_ASAP7_75t_L g4338 ( 
.A(n_4147),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_4169),
.Y(n_4339)
);

HB1xp67_ASAP7_75t_L g4340 ( 
.A(n_4263),
.Y(n_4340)
);

INVx5_ASAP7_75t_L g4341 ( 
.A(n_4205),
.Y(n_4341)
);

AOI22xp33_ASAP7_75t_L g4342 ( 
.A1(n_4158),
.A2(n_249),
.B1(n_247),
.B2(n_248),
.Y(n_4342)
);

AND2x2_ASAP7_75t_L g4343 ( 
.A(n_4194),
.B(n_249),
.Y(n_4343)
);

INVx4_ASAP7_75t_L g4344 ( 
.A(n_4146),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_4170),
.Y(n_4345)
);

INVx3_ASAP7_75t_L g4346 ( 
.A(n_4228),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4171),
.Y(n_4347)
);

BUFx3_ASAP7_75t_L g4348 ( 
.A(n_4257),
.Y(n_4348)
);

NAND3xp33_ASAP7_75t_L g4349 ( 
.A(n_4128),
.B(n_250),
.C(n_251),
.Y(n_4349)
);

HB1xp67_ASAP7_75t_L g4350 ( 
.A(n_4283),
.Y(n_4350)
);

NOR2xp33_ASAP7_75t_SL g4351 ( 
.A(n_4153),
.B(n_250),
.Y(n_4351)
);

BUFx2_ASAP7_75t_L g4352 ( 
.A(n_4166),
.Y(n_4352)
);

NAND4xp25_ASAP7_75t_L g4353 ( 
.A(n_4144),
.B(n_254),
.C(n_255),
.D(n_253),
.Y(n_4353)
);

OR2x2_ASAP7_75t_L g4354 ( 
.A(n_4200),
.B(n_252),
.Y(n_4354)
);

NAND2x1_ASAP7_75t_L g4355 ( 
.A(n_4275),
.B(n_252),
.Y(n_4355)
);

AND2x2_ASAP7_75t_L g4356 ( 
.A(n_4234),
.B(n_255),
.Y(n_4356)
);

AOI21xp5_ASAP7_75t_L g4357 ( 
.A1(n_4154),
.A2(n_256),
.B(n_257),
.Y(n_4357)
);

NOR2x1_ASAP7_75t_L g4358 ( 
.A(n_4225),
.B(n_256),
.Y(n_4358)
);

AND2x2_ASAP7_75t_L g4359 ( 
.A(n_4233),
.B(n_258),
.Y(n_4359)
);

INVxp67_ASAP7_75t_SL g4360 ( 
.A(n_4270),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4175),
.Y(n_4361)
);

OAI221xp5_ASAP7_75t_L g4362 ( 
.A1(n_4244),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.C(n_261),
.Y(n_4362)
);

INVx2_ASAP7_75t_L g4363 ( 
.A(n_4198),
.Y(n_4363)
);

AND2x2_ASAP7_75t_L g4364 ( 
.A(n_4219),
.B(n_4223),
.Y(n_4364)
);

OAI21xp33_ASAP7_75t_L g4365 ( 
.A1(n_4282),
.A2(n_259),
.B(n_260),
.Y(n_4365)
);

INVxp67_ASAP7_75t_SL g4366 ( 
.A(n_4226),
.Y(n_4366)
);

AND2x2_ASAP7_75t_L g4367 ( 
.A(n_4224),
.B(n_261),
.Y(n_4367)
);

AOI22xp5_ASAP7_75t_L g4368 ( 
.A1(n_4208),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_4368)
);

OR2x2_ASAP7_75t_L g4369 ( 
.A(n_4202),
.B(n_262),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4179),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_4183),
.Y(n_4371)
);

NOR2xp33_ASAP7_75t_L g4372 ( 
.A(n_4193),
.B(n_264),
.Y(n_4372)
);

INVx2_ASAP7_75t_L g4373 ( 
.A(n_4196),
.Y(n_4373)
);

OAI21xp5_ASAP7_75t_L g4374 ( 
.A1(n_4148),
.A2(n_265),
.B(n_266),
.Y(n_4374)
);

OAI221xp5_ASAP7_75t_L g4375 ( 
.A1(n_4210),
.A2(n_4214),
.B1(n_4160),
.B2(n_4227),
.C(n_4220),
.Y(n_4375)
);

INVx2_ASAP7_75t_L g4376 ( 
.A(n_4201),
.Y(n_4376)
);

NAND2xp5_ASAP7_75t_L g4377 ( 
.A(n_4248),
.B(n_266),
.Y(n_4377)
);

OR2x2_ASAP7_75t_L g4378 ( 
.A(n_4141),
.B(n_267),
.Y(n_4378)
);

AND2x4_ASAP7_75t_L g4379 ( 
.A(n_4229),
.B(n_4232),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4184),
.Y(n_4380)
);

OR2x2_ASAP7_75t_L g4381 ( 
.A(n_4174),
.B(n_267),
.Y(n_4381)
);

BUFx2_ASAP7_75t_L g4382 ( 
.A(n_4213),
.Y(n_4382)
);

AND2x2_ASAP7_75t_L g4383 ( 
.A(n_4139),
.B(n_269),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_4190),
.Y(n_4384)
);

AND2x2_ASAP7_75t_L g4385 ( 
.A(n_4161),
.B(n_270),
.Y(n_4385)
);

INVx2_ASAP7_75t_L g4386 ( 
.A(n_4240),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4252),
.Y(n_4387)
);

INVx2_ASAP7_75t_SL g4388 ( 
.A(n_4284),
.Y(n_4388)
);

OR2x2_ASAP7_75t_L g4389 ( 
.A(n_4256),
.B(n_271),
.Y(n_4389)
);

AO21x2_ASAP7_75t_L g4390 ( 
.A1(n_4241),
.A2(n_4264),
.B(n_4255),
.Y(n_4390)
);

NAND2xp5_ASAP7_75t_L g4391 ( 
.A(n_4271),
.B(n_271),
.Y(n_4391)
);

AND2x2_ASAP7_75t_L g4392 ( 
.A(n_4172),
.B(n_272),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_4258),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_4259),
.Y(n_4394)
);

OR2x2_ASAP7_75t_L g4395 ( 
.A(n_4268),
.B(n_272),
.Y(n_4395)
);

AO21x2_ASAP7_75t_L g4396 ( 
.A1(n_4269),
.A2(n_274),
.B(n_275),
.Y(n_4396)
);

OR2x2_ASAP7_75t_L g4397 ( 
.A(n_4277),
.B(n_275),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4245),
.Y(n_4398)
);

AND2x2_ASAP7_75t_L g4399 ( 
.A(n_4177),
.B(n_276),
.Y(n_4399)
);

NAND2xp5_ASAP7_75t_L g4400 ( 
.A(n_4217),
.B(n_277),
.Y(n_4400)
);

BUFx3_ASAP7_75t_L g4401 ( 
.A(n_4188),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4245),
.Y(n_4402)
);

AND2x2_ASAP7_75t_L g4403 ( 
.A(n_4243),
.B(n_277),
.Y(n_4403)
);

OAI31xp33_ASAP7_75t_L g4404 ( 
.A1(n_4195),
.A2(n_280),
.A3(n_278),
.B(n_279),
.Y(n_4404)
);

OAI211xp5_ASAP7_75t_L g4405 ( 
.A1(n_4253),
.A2(n_282),
.B(n_278),
.C(n_280),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_4187),
.Y(n_4406)
);

INVxp67_ASAP7_75t_SL g4407 ( 
.A(n_4286),
.Y(n_4407)
);

OAI221xp5_ASAP7_75t_L g4408 ( 
.A1(n_4199),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.C(n_285),
.Y(n_4408)
);

OA21x2_ASAP7_75t_L g4409 ( 
.A1(n_4279),
.A2(n_283),
.B(n_285),
.Y(n_4409)
);

OAI21xp33_ASAP7_75t_L g4410 ( 
.A1(n_4221),
.A2(n_286),
.B(n_287),
.Y(n_4410)
);

AOI22xp33_ASAP7_75t_L g4411 ( 
.A1(n_4204),
.A2(n_289),
.B1(n_286),
.B2(n_288),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4149),
.Y(n_4412)
);

BUFx3_ASAP7_75t_L g4413 ( 
.A(n_4247),
.Y(n_4413)
);

AOI22xp5_ASAP7_75t_L g4414 ( 
.A1(n_4251),
.A2(n_291),
.B1(n_288),
.B2(n_290),
.Y(n_4414)
);

HB1xp67_ASAP7_75t_L g4415 ( 
.A(n_4213),
.Y(n_4415)
);

AND2x2_ASAP7_75t_L g4416 ( 
.A(n_4260),
.B(n_290),
.Y(n_4416)
);

INVx2_ASAP7_75t_L g4417 ( 
.A(n_4145),
.Y(n_4417)
);

AND2x2_ASAP7_75t_L g4418 ( 
.A(n_4261),
.B(n_292),
.Y(n_4418)
);

INVx2_ASAP7_75t_L g4419 ( 
.A(n_4156),
.Y(n_4419)
);

OA21x2_ASAP7_75t_L g4420 ( 
.A1(n_4140),
.A2(n_4142),
.B(n_4206),
.Y(n_4420)
);

INVx2_ASAP7_75t_L g4421 ( 
.A(n_4181),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_L g4422 ( 
.A(n_4265),
.B(n_292),
.Y(n_4422)
);

AND2x2_ASAP7_75t_L g4423 ( 
.A(n_4281),
.B(n_4163),
.Y(n_4423)
);

INVx2_ASAP7_75t_L g4424 ( 
.A(n_4129),
.Y(n_4424)
);

INVx3_ASAP7_75t_L g4425 ( 
.A(n_4287),
.Y(n_4425)
);

AOI21xp5_ASAP7_75t_L g4426 ( 
.A1(n_4192),
.A2(n_293),
.B(n_294),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_4167),
.Y(n_4427)
);

AOI33xp33_ASAP7_75t_L g4428 ( 
.A1(n_4197),
.A2(n_296),
.A3(n_298),
.B1(n_293),
.B2(n_295),
.B3(n_297),
.Y(n_4428)
);

BUFx2_ASAP7_75t_L g4429 ( 
.A(n_4155),
.Y(n_4429)
);

AND2x4_ASAP7_75t_L g4430 ( 
.A(n_4203),
.B(n_295),
.Y(n_4430)
);

AND2x2_ASAP7_75t_L g4431 ( 
.A(n_4215),
.B(n_297),
.Y(n_4431)
);

AND2x2_ASAP7_75t_L g4432 ( 
.A(n_4216),
.B(n_298),
.Y(n_4432)
);

NOR2xp33_ASAP7_75t_L g4433 ( 
.A(n_4222),
.B(n_4189),
.Y(n_4433)
);

AND2x2_ASAP7_75t_L g4434 ( 
.A(n_4167),
.B(n_4155),
.Y(n_4434)
);

AND2x2_ASAP7_75t_L g4435 ( 
.A(n_4235),
.B(n_299),
.Y(n_4435)
);

OR2x2_ASAP7_75t_L g4436 ( 
.A(n_4235),
.B(n_299),
.Y(n_4436)
);

AND2x2_ASAP7_75t_L g4437 ( 
.A(n_4137),
.B(n_300),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_L g4438 ( 
.A(n_4173),
.B(n_300),
.Y(n_4438)
);

OR2x2_ASAP7_75t_L g4439 ( 
.A(n_4230),
.B(n_301),
.Y(n_4439)
);

AOI21xp33_ASAP7_75t_L g4440 ( 
.A1(n_4135),
.A2(n_302),
.B(n_303),
.Y(n_4440)
);

AND2x2_ASAP7_75t_L g4441 ( 
.A(n_4137),
.B(n_302),
.Y(n_4441)
);

AND2x2_ASAP7_75t_L g4442 ( 
.A(n_4137),
.B(n_303),
.Y(n_4442)
);

AOI22xp33_ASAP7_75t_SL g4443 ( 
.A1(n_4135),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_4443)
);

OR2x2_ASAP7_75t_L g4444 ( 
.A(n_4230),
.B(n_305),
.Y(n_4444)
);

INVxp67_ASAP7_75t_R g4445 ( 
.A(n_4206),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_4165),
.Y(n_4446)
);

HB1xp67_ASAP7_75t_L g4447 ( 
.A(n_4151),
.Y(n_4447)
);

INVx2_ASAP7_75t_L g4448 ( 
.A(n_4238),
.Y(n_4448)
);

BUFx6f_ASAP7_75t_L g4449 ( 
.A(n_4159),
.Y(n_4449)
);

AND2x2_ASAP7_75t_L g4450 ( 
.A(n_4137),
.B(n_306),
.Y(n_4450)
);

INVx3_ASAP7_75t_L g4451 ( 
.A(n_4191),
.Y(n_4451)
);

INVx2_ASAP7_75t_SL g4452 ( 
.A(n_4137),
.Y(n_4452)
);

HB1xp67_ASAP7_75t_L g4453 ( 
.A(n_4151),
.Y(n_4453)
);

INVx2_ASAP7_75t_L g4454 ( 
.A(n_4238),
.Y(n_4454)
);

INVx1_ASAP7_75t_SL g4455 ( 
.A(n_4246),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_4165),
.Y(n_4456)
);

OR2x2_ASAP7_75t_L g4457 ( 
.A(n_4230),
.B(n_307),
.Y(n_4457)
);

INVx4_ASAP7_75t_L g4458 ( 
.A(n_4146),
.Y(n_4458)
);

OR2x2_ASAP7_75t_L g4459 ( 
.A(n_4230),
.B(n_308),
.Y(n_4459)
);

AND2x2_ASAP7_75t_L g4460 ( 
.A(n_4137),
.B(n_309),
.Y(n_4460)
);

OR2x2_ASAP7_75t_L g4461 ( 
.A(n_4230),
.B(n_309),
.Y(n_4461)
);

NOR2x1_ASAP7_75t_SL g4462 ( 
.A(n_4127),
.B(n_310),
.Y(n_4462)
);

INVxp67_ASAP7_75t_L g4463 ( 
.A(n_4173),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_L g4464 ( 
.A(n_4173),
.B(n_310),
.Y(n_4464)
);

BUFx2_ASAP7_75t_L g4465 ( 
.A(n_4137),
.Y(n_4465)
);

AOI221xp5_ASAP7_75t_L g4466 ( 
.A1(n_4135),
.A2(n_314),
.B1(n_312),
.B2(n_313),
.C(n_315),
.Y(n_4466)
);

INVx1_ASAP7_75t_L g4467 ( 
.A(n_4165),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_4165),
.Y(n_4468)
);

AND2x2_ASAP7_75t_L g4469 ( 
.A(n_4137),
.B(n_313),
.Y(n_4469)
);

AND2x2_ASAP7_75t_L g4470 ( 
.A(n_4137),
.B(n_316),
.Y(n_4470)
);

AND2x2_ASAP7_75t_L g4471 ( 
.A(n_4137),
.B(n_317),
.Y(n_4471)
);

AO21x2_ASAP7_75t_L g4472 ( 
.A1(n_4151),
.A2(n_317),
.B(n_318),
.Y(n_4472)
);

NOR2x1_ASAP7_75t_L g4473 ( 
.A(n_4276),
.B(n_319),
.Y(n_4473)
);

AND2x2_ASAP7_75t_L g4474 ( 
.A(n_4137),
.B(n_319),
.Y(n_4474)
);

INVx2_ASAP7_75t_L g4475 ( 
.A(n_4238),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4165),
.Y(n_4476)
);

NAND4xp25_ASAP7_75t_L g4477 ( 
.A(n_4135),
.B(n_324),
.C(n_325),
.D(n_323),
.Y(n_4477)
);

INVx2_ASAP7_75t_L g4478 ( 
.A(n_4238),
.Y(n_4478)
);

INVx1_ASAP7_75t_L g4479 ( 
.A(n_4165),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_4165),
.Y(n_4480)
);

AOI221xp5_ASAP7_75t_L g4481 ( 
.A1(n_4135),
.A2(n_325),
.B1(n_322),
.B2(n_323),
.C(n_326),
.Y(n_4481)
);

INVx1_ASAP7_75t_L g4482 ( 
.A(n_4165),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4165),
.Y(n_4483)
);

BUFx2_ASAP7_75t_L g4484 ( 
.A(n_4137),
.Y(n_4484)
);

CKINVDCx20_ASAP7_75t_R g4485 ( 
.A(n_4338),
.Y(n_4485)
);

OR2x2_ASAP7_75t_L g4486 ( 
.A(n_4463),
.B(n_322),
.Y(n_4486)
);

OR2x2_ASAP7_75t_L g4487 ( 
.A(n_4297),
.B(n_327),
.Y(n_4487)
);

OR2x2_ASAP7_75t_L g4488 ( 
.A(n_4373),
.B(n_327),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_4332),
.Y(n_4489)
);

INVx2_ASAP7_75t_L g4490 ( 
.A(n_4484),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_L g4491 ( 
.A(n_4382),
.B(n_328),
.Y(n_4491)
);

INVx1_ASAP7_75t_SL g4492 ( 
.A(n_4465),
.Y(n_4492)
);

AND2x2_ASAP7_75t_L g4493 ( 
.A(n_4452),
.B(n_329),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_SL g4494 ( 
.A(n_4301),
.B(n_331),
.Y(n_4494)
);

AOI321xp33_ASAP7_75t_L g4495 ( 
.A1(n_4375),
.A2(n_333),
.A3(n_335),
.B1(n_331),
.B2(n_332),
.C(n_334),
.Y(n_4495)
);

AND2x2_ASAP7_75t_SL g4496 ( 
.A(n_4415),
.B(n_4434),
.Y(n_4496)
);

AND2x4_ASAP7_75t_SL g4497 ( 
.A(n_4449),
.B(n_333),
.Y(n_4497)
);

INVx3_ASAP7_75t_L g4498 ( 
.A(n_4449),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_4340),
.Y(n_4499)
);

CKINVDCx5p33_ASAP7_75t_R g4500 ( 
.A(n_4290),
.Y(n_4500)
);

NAND2xp5_ASAP7_75t_L g4501 ( 
.A(n_4298),
.B(n_334),
.Y(n_4501)
);

INVx2_ASAP7_75t_L g4502 ( 
.A(n_4348),
.Y(n_4502)
);

AND2x2_ASAP7_75t_L g4503 ( 
.A(n_4455),
.B(n_336),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_4350),
.Y(n_4504)
);

NAND2xp5_ASAP7_75t_L g4505 ( 
.A(n_4407),
.B(n_338),
.Y(n_4505)
);

HB1xp67_ASAP7_75t_L g4506 ( 
.A(n_4352),
.Y(n_4506)
);

INVx1_ASAP7_75t_SL g4507 ( 
.A(n_4291),
.Y(n_4507)
);

NOR2xp33_ASAP7_75t_L g4508 ( 
.A(n_4289),
.B(n_339),
.Y(n_4508)
);

AND2x2_ASAP7_75t_L g4509 ( 
.A(n_4312),
.B(n_339),
.Y(n_4509)
);

INVx2_ASAP7_75t_L g4510 ( 
.A(n_4451),
.Y(n_4510)
);

INVx1_ASAP7_75t_SL g4511 ( 
.A(n_4437),
.Y(n_4511)
);

AND2x2_ASAP7_75t_L g4512 ( 
.A(n_4293),
.B(n_340),
.Y(n_4512)
);

AND2x4_ASAP7_75t_L g4513 ( 
.A(n_4323),
.B(n_341),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4310),
.Y(n_4514)
);

AND2x2_ASAP7_75t_L g4515 ( 
.A(n_4448),
.B(n_342),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_4447),
.Y(n_4516)
);

AOI22xp33_ASAP7_75t_SL g4517 ( 
.A1(n_4308),
.A2(n_345),
.B1(n_342),
.B2(n_343),
.Y(n_4517)
);

NAND2xp5_ASAP7_75t_SL g4518 ( 
.A(n_4341),
.B(n_343),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_4341),
.B(n_345),
.Y(n_4519)
);

NOR2x1_ASAP7_75t_L g4520 ( 
.A(n_4322),
.B(n_346),
.Y(n_4520)
);

NAND2xp5_ASAP7_75t_L g4521 ( 
.A(n_4454),
.B(n_346),
.Y(n_4521)
);

INVx1_ASAP7_75t_L g4522 ( 
.A(n_4453),
.Y(n_4522)
);

AND2x4_ASAP7_75t_L g4523 ( 
.A(n_4475),
.B(n_347),
.Y(n_4523)
);

INVx2_ASAP7_75t_L g4524 ( 
.A(n_4478),
.Y(n_4524)
);

AND2x4_ASAP7_75t_L g4525 ( 
.A(n_4388),
.B(n_347),
.Y(n_4525)
);

NOR2xp33_ASAP7_75t_R g4526 ( 
.A(n_4351),
.B(n_4317),
.Y(n_4526)
);

INVx2_ASAP7_75t_L g4527 ( 
.A(n_4401),
.Y(n_4527)
);

INVxp67_ASAP7_75t_SL g4528 ( 
.A(n_4462),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4386),
.Y(n_4529)
);

AND2x4_ASAP7_75t_SL g4530 ( 
.A(n_4344),
.B(n_348),
.Y(n_4530)
);

OR2x2_ASAP7_75t_L g4531 ( 
.A(n_4320),
.B(n_348),
.Y(n_4531)
);

NAND2xp5_ASAP7_75t_L g4532 ( 
.A(n_4473),
.B(n_4425),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_L g4533 ( 
.A(n_4417),
.B(n_4419),
.Y(n_4533)
);

AND2x2_ASAP7_75t_L g4534 ( 
.A(n_4346),
.B(n_349),
.Y(n_4534)
);

AND2x2_ASAP7_75t_L g4535 ( 
.A(n_4324),
.B(n_349),
.Y(n_4535)
);

HB1xp67_ASAP7_75t_L g4536 ( 
.A(n_4413),
.Y(n_4536)
);

HB1xp67_ASAP7_75t_L g4537 ( 
.A(n_4420),
.Y(n_4537)
);

NOR2xp33_ASAP7_75t_L g4538 ( 
.A(n_4458),
.B(n_350),
.Y(n_4538)
);

BUFx2_ASAP7_75t_L g4539 ( 
.A(n_4360),
.Y(n_4539)
);

INVx2_ASAP7_75t_SL g4540 ( 
.A(n_4441),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_L g4541 ( 
.A(n_4443),
.B(n_350),
.Y(n_4541)
);

AND2x2_ASAP7_75t_L g4542 ( 
.A(n_4309),
.B(n_351),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_L g4543 ( 
.A(n_4409),
.B(n_351),
.Y(n_4543)
);

AND2x2_ASAP7_75t_L g4544 ( 
.A(n_4336),
.B(n_352),
.Y(n_4544)
);

AND2x2_ASAP7_75t_L g4545 ( 
.A(n_4363),
.B(n_353),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_L g4546 ( 
.A(n_4406),
.B(n_353),
.Y(n_4546)
);

HB1xp67_ASAP7_75t_L g4547 ( 
.A(n_4429),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_4390),
.B(n_354),
.Y(n_4548)
);

AND2x2_ASAP7_75t_L g4549 ( 
.A(n_4445),
.B(n_354),
.Y(n_4549)
);

INVx2_ASAP7_75t_L g4550 ( 
.A(n_4333),
.Y(n_4550)
);

INVx2_ASAP7_75t_L g4551 ( 
.A(n_4378),
.Y(n_4551)
);

AND2x4_ASAP7_75t_L g4552 ( 
.A(n_4423),
.B(n_355),
.Y(n_4552)
);

AND2x2_ASAP7_75t_L g4553 ( 
.A(n_4364),
.B(n_356),
.Y(n_4553)
);

AND2x2_ASAP7_75t_L g4554 ( 
.A(n_4424),
.B(n_356),
.Y(n_4554)
);

INVx2_ASAP7_75t_L g4555 ( 
.A(n_4381),
.Y(n_4555)
);

AND2x2_ASAP7_75t_L g4556 ( 
.A(n_4421),
.B(n_357),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_4393),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_4304),
.Y(n_4558)
);

INVx1_ASAP7_75t_L g4559 ( 
.A(n_4313),
.Y(n_4559)
);

AND2x2_ASAP7_75t_L g4560 ( 
.A(n_4412),
.B(n_358),
.Y(n_4560)
);

AND2x4_ASAP7_75t_L g4561 ( 
.A(n_4379),
.B(n_358),
.Y(n_4561)
);

AND2x2_ASAP7_75t_L g4562 ( 
.A(n_4376),
.B(n_359),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4319),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_4325),
.Y(n_4564)
);

NAND4xp25_ASAP7_75t_L g4565 ( 
.A(n_4331),
.B(n_362),
.C(n_359),
.D(n_360),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_4326),
.Y(n_4566)
);

OR2x2_ASAP7_75t_L g4567 ( 
.A(n_4292),
.B(n_363),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4328),
.Y(n_4568)
);

AND2x4_ASAP7_75t_SL g4569 ( 
.A(n_4442),
.B(n_363),
.Y(n_4569)
);

AND2x2_ASAP7_75t_L g4570 ( 
.A(n_4433),
.B(n_364),
.Y(n_4570)
);

OR2x2_ASAP7_75t_L g4571 ( 
.A(n_4446),
.B(n_364),
.Y(n_4571)
);

NAND2xp5_ASAP7_75t_L g4572 ( 
.A(n_4396),
.B(n_365),
.Y(n_4572)
);

BUFx2_ASAP7_75t_L g4573 ( 
.A(n_4450),
.Y(n_4573)
);

AND2x2_ASAP7_75t_L g4574 ( 
.A(n_4460),
.B(n_366),
.Y(n_4574)
);

INVx2_ASAP7_75t_L g4575 ( 
.A(n_4355),
.Y(n_4575)
);

INVx1_ASAP7_75t_SL g4576 ( 
.A(n_4469),
.Y(n_4576)
);

AND2x2_ASAP7_75t_L g4577 ( 
.A(n_4470),
.B(n_366),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_4335),
.Y(n_4578)
);

CKINVDCx16_ASAP7_75t_R g4579 ( 
.A(n_4321),
.Y(n_4579)
);

NAND2xp5_ASAP7_75t_L g4580 ( 
.A(n_4358),
.B(n_367),
.Y(n_4580)
);

NAND4xp25_ASAP7_75t_L g4581 ( 
.A(n_4466),
.B(n_4481),
.C(n_4314),
.D(n_4477),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4339),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_4345),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4347),
.Y(n_4584)
);

NAND2x1p5_ASAP7_75t_L g4585 ( 
.A(n_4471),
.B(n_368),
.Y(n_4585)
);

NOR2xp33_ASAP7_75t_R g4586 ( 
.A(n_4474),
.B(n_369),
.Y(n_4586)
);

INVx2_ASAP7_75t_L g4587 ( 
.A(n_4315),
.Y(n_4587)
);

AND2x2_ASAP7_75t_L g4588 ( 
.A(n_4356),
.B(n_369),
.Y(n_4588)
);

NAND2xp5_ASAP7_75t_L g4589 ( 
.A(n_4398),
.B(n_370),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4361),
.Y(n_4590)
);

INVx2_ASAP7_75t_L g4591 ( 
.A(n_4327),
.Y(n_4591)
);

AND2x2_ASAP7_75t_L g4592 ( 
.A(n_4359),
.B(n_370),
.Y(n_4592)
);

AND2x2_ASAP7_75t_L g4593 ( 
.A(n_4300),
.B(n_371),
.Y(n_4593)
);

AND2x2_ASAP7_75t_L g4594 ( 
.A(n_4303),
.B(n_372),
.Y(n_4594)
);

BUFx3_ASAP7_75t_L g4595 ( 
.A(n_4302),
.Y(n_4595)
);

OR2x2_ASAP7_75t_L g4596 ( 
.A(n_4456),
.B(n_372),
.Y(n_4596)
);

AND2x4_ASAP7_75t_L g4597 ( 
.A(n_4307),
.B(n_373),
.Y(n_4597)
);

AND2x2_ASAP7_75t_L g4598 ( 
.A(n_4311),
.B(n_373),
.Y(n_4598)
);

AND2x2_ASAP7_75t_L g4599 ( 
.A(n_4316),
.B(n_374),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_L g4600 ( 
.A(n_4402),
.B(n_374),
.Y(n_4600)
);

AND2x2_ASAP7_75t_L g4601 ( 
.A(n_4329),
.B(n_375),
.Y(n_4601)
);

OR2x2_ASAP7_75t_L g4602 ( 
.A(n_4467),
.B(n_376),
.Y(n_4602)
);

AND2x2_ASAP7_75t_L g4603 ( 
.A(n_4334),
.B(n_4399),
.Y(n_4603)
);

OR2x2_ASAP7_75t_L g4604 ( 
.A(n_4468),
.B(n_376),
.Y(n_4604)
);

INVx1_ASAP7_75t_L g4605 ( 
.A(n_4370),
.Y(n_4605)
);

NAND2xp5_ASAP7_75t_L g4606 ( 
.A(n_4427),
.B(n_377),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_4440),
.B(n_378),
.Y(n_4607)
);

NOR2xp33_ASAP7_75t_L g4608 ( 
.A(n_4438),
.B(n_378),
.Y(n_4608)
);

AND2x2_ASAP7_75t_L g4609 ( 
.A(n_4299),
.B(n_379),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4371),
.Y(n_4610)
);

INVx2_ASAP7_75t_L g4611 ( 
.A(n_4384),
.Y(n_4611)
);

AND2x2_ASAP7_75t_L g4612 ( 
.A(n_4343),
.B(n_379),
.Y(n_4612)
);

AND2x2_ASAP7_75t_L g4613 ( 
.A(n_4403),
.B(n_380),
.Y(n_4613)
);

INVx1_ASAP7_75t_SL g4614 ( 
.A(n_4294),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_4380),
.Y(n_4615)
);

OR2x6_ASAP7_75t_L g4616 ( 
.A(n_4426),
.B(n_381),
.Y(n_4616)
);

AND2x2_ASAP7_75t_L g4617 ( 
.A(n_4416),
.B(n_381),
.Y(n_4617)
);

INVx1_ASAP7_75t_L g4618 ( 
.A(n_4387),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4394),
.Y(n_4619)
);

AND2x4_ASAP7_75t_L g4620 ( 
.A(n_4306),
.B(n_382),
.Y(n_4620)
);

NAND2xp5_ASAP7_75t_SL g4621 ( 
.A(n_4357),
.B(n_382),
.Y(n_4621)
);

NAND2xp5_ASAP7_75t_L g4622 ( 
.A(n_4472),
.B(n_383),
.Y(n_4622)
);

AND2x2_ASAP7_75t_L g4623 ( 
.A(n_4492),
.B(n_4476),
.Y(n_4623)
);

NAND2xp5_ASAP7_75t_L g4624 ( 
.A(n_4579),
.B(n_4479),
.Y(n_4624)
);

INVx2_ASAP7_75t_L g4625 ( 
.A(n_4485),
.Y(n_4625)
);

INVx2_ASAP7_75t_SL g4626 ( 
.A(n_4595),
.Y(n_4626)
);

INVx1_ASAP7_75t_SL g4627 ( 
.A(n_4526),
.Y(n_4627)
);

INVx1_ASAP7_75t_SL g4628 ( 
.A(n_4586),
.Y(n_4628)
);

AND2x2_ASAP7_75t_L g4629 ( 
.A(n_4573),
.B(n_4480),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_L g4630 ( 
.A(n_4507),
.B(n_4482),
.Y(n_4630)
);

OR2x2_ASAP7_75t_L g4631 ( 
.A(n_4539),
.B(n_4464),
.Y(n_4631)
);

AOI211xp5_ASAP7_75t_SL g4632 ( 
.A1(n_4528),
.A2(n_4296),
.B(n_4506),
.C(n_4537),
.Y(n_4632)
);

AND4x2_ASAP7_75t_L g4633 ( 
.A(n_4520),
.B(n_4366),
.C(n_4404),
.D(n_4428),
.Y(n_4633)
);

INVx1_ASAP7_75t_L g4634 ( 
.A(n_4547),
.Y(n_4634)
);

INVx2_ASAP7_75t_SL g4635 ( 
.A(n_4490),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4489),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_4499),
.Y(n_4637)
);

NAND2xp5_ASAP7_75t_L g4638 ( 
.A(n_4511),
.B(n_4483),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_L g4639 ( 
.A(n_4576),
.B(n_4400),
.Y(n_4639)
);

HB1xp67_ASAP7_75t_L g4640 ( 
.A(n_4536),
.Y(n_4640)
);

INVx4_ASAP7_75t_L g4641 ( 
.A(n_4500),
.Y(n_4641)
);

NAND2xp5_ASAP7_75t_L g4642 ( 
.A(n_4540),
.B(n_4435),
.Y(n_4642)
);

XOR2x2_ASAP7_75t_L g4643 ( 
.A(n_4621),
.B(n_4349),
.Y(n_4643)
);

NAND4xp75_ASAP7_75t_SL g4644 ( 
.A(n_4549),
.B(n_4372),
.C(n_4432),
.D(n_4431),
.Y(n_4644)
);

AND2x2_ASAP7_75t_L g4645 ( 
.A(n_4498),
.B(n_4550),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4504),
.Y(n_4646)
);

AND2x2_ASAP7_75t_L g4647 ( 
.A(n_4603),
.B(n_4418),
.Y(n_4647)
);

OAI21xp5_ASAP7_75t_SL g4648 ( 
.A1(n_4581),
.A2(n_4374),
.B(n_4353),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_4514),
.Y(n_4649)
);

XNOR2xp5_ASAP7_75t_L g4650 ( 
.A(n_4565),
.B(n_4414),
.Y(n_4650)
);

OR2x2_ASAP7_75t_L g4651 ( 
.A(n_4532),
.B(n_4516),
.Y(n_4651)
);

NOR2xp33_ASAP7_75t_L g4652 ( 
.A(n_4614),
.B(n_4354),
.Y(n_4652)
);

BUFx5_ASAP7_75t_L g4653 ( 
.A(n_4493),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4522),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_4575),
.Y(n_4655)
);

NOR2x1_ASAP7_75t_L g4656 ( 
.A(n_4518),
.B(n_4295),
.Y(n_4656)
);

NAND2xp5_ASAP7_75t_L g4657 ( 
.A(n_4570),
.B(n_4502),
.Y(n_4657)
);

INVx2_ASAP7_75t_L g4658 ( 
.A(n_4527),
.Y(n_4658)
);

HB1xp67_ASAP7_75t_L g4659 ( 
.A(n_4519),
.Y(n_4659)
);

AND2x2_ASAP7_75t_L g4660 ( 
.A(n_4510),
.B(n_4385),
.Y(n_4660)
);

NOR3xp33_ASAP7_75t_SL g4661 ( 
.A(n_4533),
.B(n_4410),
.C(n_4362),
.Y(n_4661)
);

OR2x2_ASAP7_75t_L g4662 ( 
.A(n_4524),
.B(n_4439),
.Y(n_4662)
);

HB1xp67_ASAP7_75t_L g4663 ( 
.A(n_4496),
.Y(n_4663)
);

NOR2x1p5_ASAP7_75t_L g4664 ( 
.A(n_4587),
.B(n_4422),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4556),
.Y(n_4665)
);

AOI21xp5_ASAP7_75t_L g4666 ( 
.A1(n_4548),
.A2(n_4391),
.B(n_4377),
.Y(n_4666)
);

AND2x2_ASAP7_75t_L g4667 ( 
.A(n_4591),
.B(n_4392),
.Y(n_4667)
);

NAND4xp75_ASAP7_75t_L g4668 ( 
.A(n_4494),
.B(n_4368),
.C(n_4367),
.D(n_4383),
.Y(n_4668)
);

INVx2_ASAP7_75t_L g4669 ( 
.A(n_4585),
.Y(n_4669)
);

INVx2_ASAP7_75t_L g4670 ( 
.A(n_4512),
.Y(n_4670)
);

NAND4xp75_ASAP7_75t_SL g4671 ( 
.A(n_4508),
.B(n_4365),
.C(n_4305),
.D(n_4405),
.Y(n_4671)
);

NAND2xp5_ASAP7_75t_L g4672 ( 
.A(n_4551),
.B(n_4444),
.Y(n_4672)
);

OAI22xp33_ASAP7_75t_L g4673 ( 
.A1(n_4616),
.A2(n_4408),
.B1(n_4459),
.B2(n_4457),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_4554),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_4560),
.Y(n_4675)
);

NAND4xp75_ASAP7_75t_L g4676 ( 
.A(n_4622),
.B(n_4318),
.C(n_4342),
.D(n_4436),
.Y(n_4676)
);

INVx2_ASAP7_75t_SL g4677 ( 
.A(n_4569),
.Y(n_4677)
);

INVx3_ASAP7_75t_R g4678 ( 
.A(n_4523),
.Y(n_4678)
);

INVx1_ASAP7_75t_L g4679 ( 
.A(n_4567),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4571),
.Y(n_4680)
);

INVx2_ASAP7_75t_SL g4681 ( 
.A(n_4513),
.Y(n_4681)
);

OR2x2_ASAP7_75t_L g4682 ( 
.A(n_4487),
.B(n_4461),
.Y(n_4682)
);

INVx2_ASAP7_75t_L g4683 ( 
.A(n_4515),
.Y(n_4683)
);

XOR2xp5_ASAP7_75t_L g4684 ( 
.A(n_4517),
.B(n_4430),
.Y(n_4684)
);

XOR2xp5_ASAP7_75t_L g4685 ( 
.A(n_4597),
.B(n_4552),
.Y(n_4685)
);

NAND2xp5_ASAP7_75t_L g4686 ( 
.A(n_4555),
.B(n_4369),
.Y(n_4686)
);

AND2x2_ASAP7_75t_L g4687 ( 
.A(n_4503),
.B(n_4330),
.Y(n_4687)
);

INVxp67_ASAP7_75t_L g4688 ( 
.A(n_4616),
.Y(n_4688)
);

NAND4xp75_ASAP7_75t_SL g4689 ( 
.A(n_4538),
.B(n_4608),
.C(n_4542),
.D(n_4544),
.Y(n_4689)
);

XNOR2xp5_ASAP7_75t_L g4690 ( 
.A(n_4574),
.B(n_4411),
.Y(n_4690)
);

INVx2_ASAP7_75t_SL g4691 ( 
.A(n_4530),
.Y(n_4691)
);

AND2x2_ASAP7_75t_L g4692 ( 
.A(n_4553),
.B(n_4337),
.Y(n_4692)
);

AOI22xp5_ASAP7_75t_L g4693 ( 
.A1(n_4541),
.A2(n_4389),
.B1(n_4397),
.B2(n_4395),
.Y(n_4693)
);

XOR2x2_ASAP7_75t_L g4694 ( 
.A(n_4607),
.B(n_383),
.Y(n_4694)
);

AND2x2_ASAP7_75t_L g4695 ( 
.A(n_4613),
.B(n_384),
.Y(n_4695)
);

OR2x2_ASAP7_75t_L g4696 ( 
.A(n_4488),
.B(n_384),
.Y(n_4696)
);

NAND4xp75_ASAP7_75t_SL g4697 ( 
.A(n_4509),
.B(n_387),
.C(n_385),
.D(n_386),
.Y(n_4697)
);

XOR2x2_ASAP7_75t_L g4698 ( 
.A(n_4572),
.B(n_385),
.Y(n_4698)
);

AND2x2_ASAP7_75t_L g4699 ( 
.A(n_4617),
.B(n_387),
.Y(n_4699)
);

INVx1_ASAP7_75t_SL g4700 ( 
.A(n_4497),
.Y(n_4700)
);

INVx2_ASAP7_75t_L g4701 ( 
.A(n_4525),
.Y(n_4701)
);

OR2x2_ASAP7_75t_L g4702 ( 
.A(n_4531),
.B(n_389),
.Y(n_4702)
);

NAND2xp5_ASAP7_75t_L g4703 ( 
.A(n_4611),
.B(n_389),
.Y(n_4703)
);

AOI21xp5_ASAP7_75t_L g4704 ( 
.A1(n_4491),
.A2(n_390),
.B(n_391),
.Y(n_4704)
);

INVx1_ASAP7_75t_L g4705 ( 
.A(n_4596),
.Y(n_4705)
);

NOR4xp25_ASAP7_75t_L g4706 ( 
.A(n_4495),
.B(n_393),
.C(n_391),
.D(n_392),
.Y(n_4706)
);

AND2x2_ASAP7_75t_L g4707 ( 
.A(n_4612),
.B(n_393),
.Y(n_4707)
);

XOR2x2_ASAP7_75t_L g4708 ( 
.A(n_4580),
.B(n_394),
.Y(n_4708)
);

INVx5_ASAP7_75t_L g4709 ( 
.A(n_4545),
.Y(n_4709)
);

INVx2_ASAP7_75t_L g4710 ( 
.A(n_4562),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_4543),
.B(n_394),
.Y(n_4711)
);

BUFx3_ASAP7_75t_L g4712 ( 
.A(n_4620),
.Y(n_4712)
);

OAI22xp5_ASAP7_75t_L g4713 ( 
.A1(n_4505),
.A2(n_397),
.B1(n_398),
.B2(n_396),
.Y(n_4713)
);

AND2x2_ASAP7_75t_L g4714 ( 
.A(n_4588),
.B(n_395),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4602),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_4640),
.Y(n_4716)
);

AND2x4_ASAP7_75t_SL g4717 ( 
.A(n_4625),
.B(n_4561),
.Y(n_4717)
);

AOI22xp5_ASAP7_75t_L g4718 ( 
.A1(n_4648),
.A2(n_4529),
.B1(n_4557),
.B2(n_4521),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4629),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_4630),
.Y(n_4720)
);

INVxp67_ASAP7_75t_SL g4721 ( 
.A(n_4656),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4638),
.Y(n_4722)
);

NAND2xp5_ASAP7_75t_L g4723 ( 
.A(n_4706),
.B(n_4486),
.Y(n_4723)
);

AND2x2_ASAP7_75t_L g4724 ( 
.A(n_4628),
.B(n_4577),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_L g4725 ( 
.A(n_4681),
.B(n_4589),
.Y(n_4725)
);

INVxp33_ASAP7_75t_L g4726 ( 
.A(n_4684),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4634),
.Y(n_4727)
);

INVx1_ASAP7_75t_L g4728 ( 
.A(n_4696),
.Y(n_4728)
);

INVx1_ASAP7_75t_L g4729 ( 
.A(n_4702),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4667),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_L g4731 ( 
.A(n_4677),
.B(n_4600),
.Y(n_4731)
);

OR2x2_ASAP7_75t_L g4732 ( 
.A(n_4631),
.B(n_4546),
.Y(n_4732)
);

AND2x2_ASAP7_75t_L g4733 ( 
.A(n_4691),
.B(n_4534),
.Y(n_4733)
);

INVx2_ASAP7_75t_L g4734 ( 
.A(n_4653),
.Y(n_4734)
);

NAND2xp5_ASAP7_75t_L g4735 ( 
.A(n_4626),
.B(n_4606),
.Y(n_4735)
);

NAND2x1_ASAP7_75t_L g4736 ( 
.A(n_4669),
.B(n_4558),
.Y(n_4736)
);

INVx2_ASAP7_75t_SL g4737 ( 
.A(n_4709),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4675),
.Y(n_4738)
);

OAI21xp5_ASAP7_75t_L g4739 ( 
.A1(n_4632),
.A2(n_4501),
.B(n_4604),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4703),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4679),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4680),
.Y(n_4742)
);

INVxp67_ASAP7_75t_SL g4743 ( 
.A(n_4663),
.Y(n_4743)
);

AOI21xp33_ASAP7_75t_SL g4744 ( 
.A1(n_4673),
.A2(n_4650),
.B(n_4624),
.Y(n_4744)
);

INVx2_ASAP7_75t_L g4745 ( 
.A(n_4653),
.Y(n_4745)
);

AND2x2_ASAP7_75t_L g4746 ( 
.A(n_4700),
.B(n_4535),
.Y(n_4746)
);

NAND2x1_ASAP7_75t_L g4747 ( 
.A(n_4701),
.B(n_4559),
.Y(n_4747)
);

OR2x2_ASAP7_75t_L g4748 ( 
.A(n_4642),
.B(n_4563),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4705),
.Y(n_4749)
);

NAND4xp25_ASAP7_75t_SL g4750 ( 
.A(n_4666),
.B(n_4566),
.C(n_4568),
.D(n_4564),
.Y(n_4750)
);

NOR2xp33_ASAP7_75t_L g4751 ( 
.A(n_4641),
.B(n_4593),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4715),
.Y(n_4752)
);

AND2x2_ASAP7_75t_L g4753 ( 
.A(n_4645),
.B(n_4592),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4659),
.Y(n_4754)
);

INVx3_ASAP7_75t_L g4755 ( 
.A(n_4712),
.Y(n_4755)
);

NOR2xp67_ASAP7_75t_L g4756 ( 
.A(n_4709),
.B(n_4578),
.Y(n_4756)
);

AND2x2_ASAP7_75t_L g4757 ( 
.A(n_4627),
.B(n_4609),
.Y(n_4757)
);

INVx1_ASAP7_75t_L g4758 ( 
.A(n_4623),
.Y(n_4758)
);

AND2x2_ASAP7_75t_L g4759 ( 
.A(n_4647),
.B(n_4594),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_L g4760 ( 
.A(n_4635),
.B(n_4598),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4665),
.Y(n_4761)
);

OR2x2_ASAP7_75t_L g4762 ( 
.A(n_4651),
.B(n_4582),
.Y(n_4762)
);

NAND2xp5_ASAP7_75t_L g4763 ( 
.A(n_4709),
.B(n_4653),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4674),
.Y(n_4764)
);

INVx2_ASAP7_75t_L g4765 ( 
.A(n_4653),
.Y(n_4765)
);

AND2x2_ASAP7_75t_L g4766 ( 
.A(n_4687),
.B(n_4660),
.Y(n_4766)
);

OR2x2_ASAP7_75t_L g4767 ( 
.A(n_4662),
.B(n_4583),
.Y(n_4767)
);

INVx2_ASAP7_75t_L g4768 ( 
.A(n_4655),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4672),
.Y(n_4769)
);

INVx3_ASAP7_75t_L g4770 ( 
.A(n_4658),
.Y(n_4770)
);

INVx1_ASAP7_75t_SL g4771 ( 
.A(n_4697),
.Y(n_4771)
);

AND2x2_ASAP7_75t_L g4772 ( 
.A(n_4688),
.B(n_4599),
.Y(n_4772)
);

NAND2xp5_ASAP7_75t_L g4773 ( 
.A(n_4692),
.B(n_4601),
.Y(n_4773)
);

NAND3xp33_ASAP7_75t_L g4774 ( 
.A(n_4661),
.B(n_4590),
.C(n_4584),
.Y(n_4774)
);

OR2x2_ASAP7_75t_L g4775 ( 
.A(n_4682),
.B(n_4605),
.Y(n_4775)
);

HB1xp67_ASAP7_75t_L g4776 ( 
.A(n_4756),
.Y(n_4776)
);

AOI21xp33_ASAP7_75t_SL g4777 ( 
.A1(n_4723),
.A2(n_4652),
.B(n_4657),
.Y(n_4777)
);

INVxp67_ASAP7_75t_SL g4778 ( 
.A(n_4721),
.Y(n_4778)
);

AO22x1_ASAP7_75t_L g4779 ( 
.A1(n_4743),
.A2(n_4670),
.B1(n_4683),
.B2(n_4633),
.Y(n_4779)
);

XNOR2x1_ASAP7_75t_SL g4780 ( 
.A(n_4737),
.B(n_4707),
.Y(n_4780)
);

INVx2_ASAP7_75t_L g4781 ( 
.A(n_4755),
.Y(n_4781)
);

OAI211xp5_ASAP7_75t_SL g4782 ( 
.A1(n_4739),
.A2(n_4639),
.B(n_4637),
.C(n_4636),
.Y(n_4782)
);

NAND2xp5_ASAP7_75t_L g4783 ( 
.A(n_4724),
.B(n_4690),
.Y(n_4783)
);

OAI22xp5_ASAP7_75t_L g4784 ( 
.A1(n_4726),
.A2(n_4676),
.B1(n_4668),
.B2(n_4693),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_4716),
.Y(n_4785)
);

INVxp67_ASAP7_75t_L g4786 ( 
.A(n_4763),
.Y(n_4786)
);

XOR2xp5_ASAP7_75t_L g4787 ( 
.A(n_4733),
.B(n_4685),
.Y(n_4787)
);

INVx1_ASAP7_75t_SL g4788 ( 
.A(n_4717),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4772),
.Y(n_4789)
);

AOI21xp5_ASAP7_75t_L g4790 ( 
.A1(n_4744),
.A2(n_4643),
.B(n_4704),
.Y(n_4790)
);

NAND3xp33_ASAP7_75t_L g4791 ( 
.A(n_4774),
.B(n_4649),
.C(n_4646),
.Y(n_4791)
);

OAI22xp5_ASAP7_75t_L g4792 ( 
.A1(n_4758),
.A2(n_4710),
.B1(n_4664),
.B2(n_4686),
.Y(n_4792)
);

INVxp67_ASAP7_75t_L g4793 ( 
.A(n_4757),
.Y(n_4793)
);

OAI22xp5_ASAP7_75t_L g4794 ( 
.A1(n_4719),
.A2(n_4654),
.B1(n_4711),
.B2(n_4713),
.Y(n_4794)
);

INVx1_ASAP7_75t_L g4795 ( 
.A(n_4730),
.Y(n_4795)
);

INVxp67_ASAP7_75t_L g4796 ( 
.A(n_4746),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_L g4797 ( 
.A(n_4766),
.B(n_4708),
.Y(n_4797)
);

NAND3xp33_ASAP7_75t_SL g4798 ( 
.A(n_4771),
.B(n_4678),
.C(n_4671),
.Y(n_4798)
);

XOR2x2_ASAP7_75t_L g4799 ( 
.A(n_4751),
.B(n_4689),
.Y(n_4799)
);

AOI22xp33_ASAP7_75t_L g4800 ( 
.A1(n_4753),
.A2(n_4698),
.B1(n_4694),
.B2(n_4615),
.Y(n_4800)
);

OAI21xp5_ASAP7_75t_SL g4801 ( 
.A1(n_4718),
.A2(n_4618),
.B(n_4610),
.Y(n_4801)
);

AOI22xp33_ASAP7_75t_L g4802 ( 
.A1(n_4759),
.A2(n_4619),
.B1(n_4714),
.B2(n_4699),
.Y(n_4802)
);

NAND2xp5_ASAP7_75t_L g4803 ( 
.A(n_4770),
.B(n_4695),
.Y(n_4803)
);

XOR2x2_ASAP7_75t_L g4804 ( 
.A(n_4773),
.B(n_4644),
.Y(n_4804)
);

AOI21xp5_ASAP7_75t_L g4805 ( 
.A1(n_4736),
.A2(n_399),
.B(n_400),
.Y(n_4805)
);

OAI22xp5_ASAP7_75t_L g4806 ( 
.A1(n_4760),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_4806)
);

HB1xp67_ASAP7_75t_L g4807 ( 
.A(n_4747),
.Y(n_4807)
);

INVxp67_ASAP7_75t_L g4808 ( 
.A(n_4731),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4775),
.Y(n_4809)
);

OAI21xp5_ASAP7_75t_L g4810 ( 
.A1(n_4750),
.A2(n_401),
.B(n_402),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4767),
.Y(n_4811)
);

OAI21xp5_ASAP7_75t_L g4812 ( 
.A1(n_4735),
.A2(n_403),
.B(n_404),
.Y(n_4812)
);

OAI21xp33_ASAP7_75t_SL g4813 ( 
.A1(n_4734),
.A2(n_403),
.B(n_404),
.Y(n_4813)
);

AOI211xp5_ASAP7_75t_L g4814 ( 
.A1(n_4720),
.A2(n_407),
.B(n_405),
.C(n_406),
.Y(n_4814)
);

OAI22xp5_ASAP7_75t_L g4815 ( 
.A1(n_4722),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_4815)
);

INVx2_ASAP7_75t_L g4816 ( 
.A(n_4745),
.Y(n_4816)
);

AOI21xp33_ASAP7_75t_SL g4817 ( 
.A1(n_4762),
.A2(n_408),
.B(n_409),
.Y(n_4817)
);

INVx1_ASAP7_75t_L g4818 ( 
.A(n_4725),
.Y(n_4818)
);

INVx2_ASAP7_75t_L g4819 ( 
.A(n_4765),
.Y(n_4819)
);

AOI21xp5_ASAP7_75t_L g4820 ( 
.A1(n_4728),
.A2(n_408),
.B(n_409),
.Y(n_4820)
);

OAI21xp5_ASAP7_75t_L g4821 ( 
.A1(n_4754),
.A2(n_410),
.B(n_411),
.Y(n_4821)
);

OAI21xp33_ASAP7_75t_L g4822 ( 
.A1(n_4800),
.A2(n_4769),
.B(n_4727),
.Y(n_4822)
);

INVxp67_ASAP7_75t_L g4823 ( 
.A(n_4807),
.Y(n_4823)
);

OAI221xp5_ASAP7_75t_L g4824 ( 
.A1(n_4810),
.A2(n_4764),
.B1(n_4761),
.B2(n_4738),
.C(n_4749),
.Y(n_4824)
);

AND2x2_ASAP7_75t_L g4825 ( 
.A(n_4788),
.B(n_4729),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4789),
.Y(n_4826)
);

AOI21xp33_ASAP7_75t_L g4827 ( 
.A1(n_4784),
.A2(n_4732),
.B(n_4748),
.Y(n_4827)
);

OAI222xp33_ASAP7_75t_L g4828 ( 
.A1(n_4790),
.A2(n_4752),
.B1(n_4741),
.B2(n_4742),
.C1(n_4768),
.C2(n_4740),
.Y(n_4828)
);

NOR2x1_ASAP7_75t_L g4829 ( 
.A(n_4798),
.B(n_410),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4778),
.Y(n_4830)
);

OAI32xp33_ASAP7_75t_L g4831 ( 
.A1(n_4780),
.A2(n_430),
.A3(n_439),
.B1(n_420),
.B2(n_411),
.Y(n_4831)
);

INVx2_ASAP7_75t_L g4832 ( 
.A(n_4776),
.Y(n_4832)
);

INVx1_ASAP7_75t_L g4833 ( 
.A(n_4796),
.Y(n_4833)
);

NOR2xp33_ASAP7_75t_L g4834 ( 
.A(n_4787),
.B(n_412),
.Y(n_4834)
);

INVx1_ASAP7_75t_L g4835 ( 
.A(n_4793),
.Y(n_4835)
);

OAI22xp5_ASAP7_75t_L g4836 ( 
.A1(n_4791),
.A2(n_416),
.B1(n_413),
.B2(n_414),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4777),
.B(n_4781),
.Y(n_4837)
);

OAI322xp33_ASAP7_75t_L g4838 ( 
.A1(n_4786),
.A2(n_421),
.A3(n_419),
.B1(n_417),
.B2(n_414),
.C1(n_416),
.C2(n_418),
.Y(n_4838)
);

HB1xp67_ASAP7_75t_L g4839 ( 
.A(n_4809),
.Y(n_4839)
);

NAND2xp5_ASAP7_75t_L g4840 ( 
.A(n_4779),
.B(n_417),
.Y(n_4840)
);

AOI21xp5_ASAP7_75t_L g4841 ( 
.A1(n_4797),
.A2(n_419),
.B(n_421),
.Y(n_4841)
);

NAND2xp5_ASAP7_75t_SL g4842 ( 
.A(n_4813),
.B(n_4817),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_4811),
.Y(n_4843)
);

NAND2xp5_ASAP7_75t_L g4844 ( 
.A(n_4802),
.B(n_422),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4803),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4792),
.Y(n_4846)
);

NAND4xp25_ASAP7_75t_L g4847 ( 
.A(n_4783),
.B(n_4782),
.C(n_4794),
.D(n_4808),
.Y(n_4847)
);

AOI221xp5_ASAP7_75t_L g4848 ( 
.A1(n_4801),
.A2(n_425),
.B1(n_423),
.B2(n_424),
.C(n_426),
.Y(n_4848)
);

AOI211xp5_ASAP7_75t_L g4849 ( 
.A1(n_4805),
.A2(n_436),
.B(n_444),
.C(n_425),
.Y(n_4849)
);

INVx2_ASAP7_75t_L g4850 ( 
.A(n_4816),
.Y(n_4850)
);

INVx2_ASAP7_75t_L g4851 ( 
.A(n_4819),
.Y(n_4851)
);

AND2x2_ASAP7_75t_L g4852 ( 
.A(n_4818),
.B(n_426),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_4785),
.Y(n_4853)
);

OAI21xp5_ASAP7_75t_SL g4854 ( 
.A1(n_4795),
.A2(n_428),
.B(n_430),
.Y(n_4854)
);

AOI22xp5_ASAP7_75t_L g4855 ( 
.A1(n_4804),
.A2(n_434),
.B1(n_432),
.B2(n_433),
.Y(n_4855)
);

NAND2xp5_ASAP7_75t_L g4856 ( 
.A(n_4820),
.B(n_432),
.Y(n_4856)
);

NAND2xp5_ASAP7_75t_L g4857 ( 
.A(n_4814),
.B(n_433),
.Y(n_4857)
);

A2O1A1Ixp33_ASAP7_75t_L g4858 ( 
.A1(n_4821),
.A2(n_437),
.B(n_435),
.C(n_436),
.Y(n_4858)
);

OAI21xp5_ASAP7_75t_L g4859 ( 
.A1(n_4812),
.A2(n_439),
.B(n_438),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_4815),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_4806),
.Y(n_4861)
);

AOI21xp5_ASAP7_75t_L g4862 ( 
.A1(n_4799),
.A2(n_435),
.B(n_438),
.Y(n_4862)
);

INVx1_ASAP7_75t_L g4863 ( 
.A(n_4789),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4789),
.Y(n_4864)
);

INVx1_ASAP7_75t_SL g4865 ( 
.A(n_4788),
.Y(n_4865)
);

INVx2_ASAP7_75t_L g4866 ( 
.A(n_4776),
.Y(n_4866)
);

NAND2xp33_ASAP7_75t_L g4867 ( 
.A(n_4788),
.B(n_440),
.Y(n_4867)
);

NAND2xp5_ASAP7_75t_SL g4868 ( 
.A(n_4865),
.B(n_4829),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4825),
.Y(n_4869)
);

NOR2xp33_ASAP7_75t_L g4870 ( 
.A(n_4828),
.B(n_440),
.Y(n_4870)
);

AND2x2_ASAP7_75t_SL g4871 ( 
.A(n_4867),
.B(n_441),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_4832),
.Y(n_4872)
);

OAI21xp33_ASAP7_75t_L g4873 ( 
.A1(n_4822),
.A2(n_441),
.B(n_442),
.Y(n_4873)
);

AOI22xp5_ASAP7_75t_L g4874 ( 
.A1(n_4834),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.Y(n_4874)
);

NOR2xp33_ASAP7_75t_L g4875 ( 
.A(n_4842),
.B(n_4831),
.Y(n_4875)
);

AOI22xp5_ASAP7_75t_L g4876 ( 
.A1(n_4846),
.A2(n_446),
.B1(n_443),
.B2(n_445),
.Y(n_4876)
);

AND2x2_ASAP7_75t_L g4877 ( 
.A(n_4866),
.B(n_446),
.Y(n_4877)
);

INVx2_ASAP7_75t_L g4878 ( 
.A(n_4830),
.Y(n_4878)
);

AOI22xp5_ASAP7_75t_L g4879 ( 
.A1(n_4847),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_4879)
);

NOR2xp33_ASAP7_75t_L g4880 ( 
.A(n_4824),
.B(n_448),
.Y(n_4880)
);

NAND2xp5_ASAP7_75t_L g4881 ( 
.A(n_4823),
.B(n_450),
.Y(n_4881)
);

AND2x2_ASAP7_75t_L g4882 ( 
.A(n_4839),
.B(n_450),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4837),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4852),
.Y(n_4884)
);

O2A1O1Ixp33_ASAP7_75t_SL g4885 ( 
.A1(n_4840),
.A2(n_453),
.B(n_451),
.C(n_452),
.Y(n_4885)
);

OR2x2_ASAP7_75t_L g4886 ( 
.A(n_4844),
.B(n_4843),
.Y(n_4886)
);

AOI211x1_ASAP7_75t_L g4887 ( 
.A1(n_4862),
.A2(n_455),
.B(n_453),
.C(n_454),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4826),
.Y(n_4888)
);

INVx2_ASAP7_75t_L g4889 ( 
.A(n_4850),
.Y(n_4889)
);

O2A1O1Ixp5_ASAP7_75t_L g4890 ( 
.A1(n_4827),
.A2(n_457),
.B(n_454),
.C(n_456),
.Y(n_4890)
);

AOI21xp5_ASAP7_75t_L g4891 ( 
.A1(n_4841),
.A2(n_457),
.B(n_458),
.Y(n_4891)
);

OAI221xp5_ASAP7_75t_L g4892 ( 
.A1(n_4855),
.A2(n_4848),
.B1(n_4835),
.B2(n_4833),
.C(n_4860),
.Y(n_4892)
);

INVxp33_ASAP7_75t_L g4893 ( 
.A(n_4857),
.Y(n_4893)
);

NAND2xp5_ASAP7_75t_L g4894 ( 
.A(n_4849),
.B(n_458),
.Y(n_4894)
);

INVx1_ASAP7_75t_L g4895 ( 
.A(n_4863),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4864),
.Y(n_4896)
);

NAND2xp5_ASAP7_75t_L g4897 ( 
.A(n_4854),
.B(n_459),
.Y(n_4897)
);

AOI322xp5_ASAP7_75t_L g4898 ( 
.A1(n_4861),
.A2(n_466),
.A3(n_465),
.B1(n_462),
.B2(n_460),
.C1(n_461),
.C2(n_463),
.Y(n_4898)
);

BUFx2_ASAP7_75t_L g4899 ( 
.A(n_4851),
.Y(n_4899)
);

NAND2x1p5_ASAP7_75t_L g4900 ( 
.A(n_4853),
.B(n_461),
.Y(n_4900)
);

OAI21xp33_ASAP7_75t_SL g4901 ( 
.A1(n_4845),
.A2(n_462),
.B(n_463),
.Y(n_4901)
);

AOI22xp5_ASAP7_75t_L g4902 ( 
.A1(n_4836),
.A2(n_467),
.B1(n_465),
.B2(n_466),
.Y(n_4902)
);

NAND2xp5_ASAP7_75t_L g4903 ( 
.A(n_4858),
.B(n_467),
.Y(n_4903)
);

INVx2_ASAP7_75t_SL g4904 ( 
.A(n_4856),
.Y(n_4904)
);

OR2x2_ASAP7_75t_L g4905 ( 
.A(n_4859),
.B(n_468),
.Y(n_4905)
);

OAI22xp5_ASAP7_75t_L g4906 ( 
.A1(n_4838),
.A2(n_471),
.B1(n_469),
.B2(n_470),
.Y(n_4906)
);

AND2x2_ASAP7_75t_L g4907 ( 
.A(n_4865),
.B(n_472),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_4825),
.Y(n_4908)
);

AOI21xp5_ASAP7_75t_L g4909 ( 
.A1(n_4831),
.A2(n_473),
.B(n_474),
.Y(n_4909)
);

NAND2xp5_ASAP7_75t_L g4910 ( 
.A(n_4865),
.B(n_473),
.Y(n_4910)
);

INVxp67_ASAP7_75t_L g4911 ( 
.A(n_4829),
.Y(n_4911)
);

AOI21xp5_ASAP7_75t_L g4912 ( 
.A1(n_4831),
.A2(n_475),
.B(n_477),
.Y(n_4912)
);

INVx2_ASAP7_75t_L g4913 ( 
.A(n_4832),
.Y(n_4913)
);

INVx1_ASAP7_75t_SL g4914 ( 
.A(n_4865),
.Y(n_4914)
);

AOI22xp5_ASAP7_75t_L g4915 ( 
.A1(n_4865),
.A2(n_478),
.B1(n_475),
.B2(n_477),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4825),
.Y(n_4916)
);

AOI21xp5_ASAP7_75t_L g4917 ( 
.A1(n_4831),
.A2(n_478),
.B(n_480),
.Y(n_4917)
);

NAND3xp33_ASAP7_75t_L g4918 ( 
.A(n_4829),
.B(n_480),
.C(n_481),
.Y(n_4918)
);

NAND2xp5_ASAP7_75t_L g4919 ( 
.A(n_4865),
.B(n_481),
.Y(n_4919)
);

OR2x2_ASAP7_75t_L g4920 ( 
.A(n_4865),
.B(n_482),
.Y(n_4920)
);

A2O1A1Ixp33_ASAP7_75t_L g4921 ( 
.A1(n_4831),
.A2(n_492),
.B(n_501),
.C(n_482),
.Y(n_4921)
);

NOR2x1_ASAP7_75t_L g4922 ( 
.A(n_4918),
.B(n_484),
.Y(n_4922)
);

AOI221xp5_ASAP7_75t_L g4923 ( 
.A1(n_4870),
.A2(n_487),
.B1(n_489),
.B2(n_485),
.C(n_488),
.Y(n_4923)
);

OR2x2_ASAP7_75t_L g4924 ( 
.A(n_4914),
.B(n_484),
.Y(n_4924)
);

NOR2xp33_ASAP7_75t_L g4925 ( 
.A(n_4911),
.B(n_487),
.Y(n_4925)
);

NOR2xp33_ASAP7_75t_L g4926 ( 
.A(n_4868),
.B(n_488),
.Y(n_4926)
);

NAND2xp33_ASAP7_75t_L g4927 ( 
.A(n_4921),
.B(n_489),
.Y(n_4927)
);

INVx2_ASAP7_75t_SL g4928 ( 
.A(n_4920),
.Y(n_4928)
);

INVx1_ASAP7_75t_L g4929 ( 
.A(n_4907),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4882),
.Y(n_4930)
);

NOR3xp33_ASAP7_75t_L g4931 ( 
.A(n_4892),
.B(n_500),
.C(n_490),
.Y(n_4931)
);

AOI221xp5_ASAP7_75t_L g4932 ( 
.A1(n_4880),
.A2(n_4875),
.B1(n_4890),
.B2(n_4906),
.C(n_4883),
.Y(n_4932)
);

NAND3xp33_ASAP7_75t_SL g4933 ( 
.A(n_4909),
.B(n_491),
.C(n_493),
.Y(n_4933)
);

OAI21xp5_ASAP7_75t_L g4934 ( 
.A1(n_4912),
.A2(n_491),
.B(n_493),
.Y(n_4934)
);

NAND3xp33_ASAP7_75t_L g4935 ( 
.A(n_4901),
.B(n_494),
.C(n_495),
.Y(n_4935)
);

NOR3xp33_ASAP7_75t_L g4936 ( 
.A(n_4873),
.B(n_4908),
.C(n_4869),
.Y(n_4936)
);

NOR3x1_ASAP7_75t_L g4937 ( 
.A(n_4899),
.B(n_494),
.C(n_495),
.Y(n_4937)
);

NAND2xp5_ASAP7_75t_L g4938 ( 
.A(n_4871),
.B(n_497),
.Y(n_4938)
);

NOR2xp33_ASAP7_75t_L g4939 ( 
.A(n_4916),
.B(n_498),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4910),
.Y(n_4940)
);

NAND3xp33_ASAP7_75t_SL g4941 ( 
.A(n_4917),
.B(n_499),
.C(n_500),
.Y(n_4941)
);

AOI221xp5_ASAP7_75t_L g4942 ( 
.A1(n_4872),
.A2(n_502),
.B1(n_504),
.B2(n_501),
.C(n_503),
.Y(n_4942)
);

INVx1_ASAP7_75t_L g4943 ( 
.A(n_4919),
.Y(n_4943)
);

AOI21xp33_ASAP7_75t_SL g4944 ( 
.A1(n_4900),
.A2(n_505),
.B(n_503),
.Y(n_4944)
);

NOR3x1_ASAP7_75t_L g4945 ( 
.A(n_4904),
.B(n_499),
.C(n_505),
.Y(n_4945)
);

AOI221xp5_ASAP7_75t_L g4946 ( 
.A1(n_4879),
.A2(n_508),
.B1(n_510),
.B2(n_507),
.C(n_509),
.Y(n_4946)
);

NAND2xp5_ASAP7_75t_L g4947 ( 
.A(n_4887),
.B(n_506),
.Y(n_4947)
);

CKINVDCx5p33_ASAP7_75t_R g4948 ( 
.A(n_4877),
.Y(n_4948)
);

OR2x2_ASAP7_75t_L g4949 ( 
.A(n_4913),
.B(n_507),
.Y(n_4949)
);

NOR3xp33_ASAP7_75t_SL g4950 ( 
.A(n_4884),
.B(n_509),
.C(n_510),
.Y(n_4950)
);

OAI21xp5_ASAP7_75t_SL g4951 ( 
.A1(n_4893),
.A2(n_4878),
.B(n_4891),
.Y(n_4951)
);

NOR3xp33_ASAP7_75t_L g4952 ( 
.A(n_4886),
.B(n_521),
.C(n_511),
.Y(n_4952)
);

NAND2xp5_ASAP7_75t_SL g4953 ( 
.A(n_4889),
.B(n_512),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_4885),
.Y(n_4954)
);

INVx1_ASAP7_75t_L g4955 ( 
.A(n_4881),
.Y(n_4955)
);

INVx2_ASAP7_75t_SL g4956 ( 
.A(n_4888),
.Y(n_4956)
);

INVxp33_ASAP7_75t_SL g4957 ( 
.A(n_4915),
.Y(n_4957)
);

NAND3xp33_ASAP7_75t_L g4958 ( 
.A(n_4895),
.B(n_512),
.C(n_513),
.Y(n_4958)
);

AND2x2_ASAP7_75t_L g4959 ( 
.A(n_4905),
.B(n_513),
.Y(n_4959)
);

INVx2_ASAP7_75t_SL g4960 ( 
.A(n_4896),
.Y(n_4960)
);

AOI211xp5_ASAP7_75t_L g4961 ( 
.A1(n_4897),
.A2(n_516),
.B(n_514),
.C(n_515),
.Y(n_4961)
);

INVxp67_ASAP7_75t_L g4962 ( 
.A(n_4903),
.Y(n_4962)
);

AOI221xp5_ASAP7_75t_L g4963 ( 
.A1(n_4894),
.A2(n_520),
.B1(n_523),
.B2(n_519),
.C(n_522),
.Y(n_4963)
);

CKINVDCx6p67_ASAP7_75t_R g4964 ( 
.A(n_4898),
.Y(n_4964)
);

OA22x2_ASAP7_75t_L g4965 ( 
.A1(n_4902),
.A2(n_522),
.B1(n_523),
.B2(n_519),
.Y(n_4965)
);

OA22x2_ASAP7_75t_L g4966 ( 
.A1(n_4876),
.A2(n_526),
.B1(n_527),
.B2(n_525),
.Y(n_4966)
);

OAI22xp5_ASAP7_75t_L g4967 ( 
.A1(n_4874),
.A2(n_526),
.B1(n_515),
.B2(n_525),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4907),
.Y(n_4968)
);

NAND2xp5_ASAP7_75t_L g4969 ( 
.A(n_4914),
.B(n_527),
.Y(n_4969)
);

NAND2xp5_ASAP7_75t_SL g4970 ( 
.A(n_4871),
.B(n_528),
.Y(n_4970)
);

INVx1_ASAP7_75t_L g4971 ( 
.A(n_4907),
.Y(n_4971)
);

NAND2xp5_ASAP7_75t_SL g4972 ( 
.A(n_4871),
.B(n_528),
.Y(n_4972)
);

INVx2_ASAP7_75t_L g4973 ( 
.A(n_4920),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4907),
.Y(n_4974)
);

NOR2xp33_ASAP7_75t_SL g4975 ( 
.A(n_4914),
.B(n_529),
.Y(n_4975)
);

NAND3xp33_ASAP7_75t_SL g4976 ( 
.A(n_4914),
.B(n_529),
.C(n_530),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_L g4977 ( 
.A(n_4914),
.B(n_530),
.Y(n_4977)
);

AND2x2_ASAP7_75t_L g4978 ( 
.A(n_4914),
.B(n_531),
.Y(n_4978)
);

OR2x2_ASAP7_75t_L g4979 ( 
.A(n_4914),
.B(n_531),
.Y(n_4979)
);

NAND2xp5_ASAP7_75t_SL g4980 ( 
.A(n_4871),
.B(n_532),
.Y(n_4980)
);

INVx1_ASAP7_75t_L g4981 ( 
.A(n_4907),
.Y(n_4981)
);

AOI22xp5_ASAP7_75t_L g4982 ( 
.A1(n_4914),
.A2(n_535),
.B1(n_533),
.B2(n_534),
.Y(n_4982)
);

NOR2x1_ASAP7_75t_L g4983 ( 
.A(n_4918),
.B(n_534),
.Y(n_4983)
);

NAND2xp5_ASAP7_75t_L g4984 ( 
.A(n_4914),
.B(n_535),
.Y(n_4984)
);

NAND2xp5_ASAP7_75t_L g4985 ( 
.A(n_4914),
.B(n_536),
.Y(n_4985)
);

NOR2xp33_ASAP7_75t_L g4986 ( 
.A(n_4914),
.B(n_536),
.Y(n_4986)
);

OAI22xp5_ASAP7_75t_SL g4987 ( 
.A1(n_4871),
.A2(n_539),
.B1(n_537),
.B2(n_538),
.Y(n_4987)
);

NOR2x1_ASAP7_75t_L g4988 ( 
.A(n_4918),
.B(n_537),
.Y(n_4988)
);

XNOR2xp5_ASAP7_75t_L g4989 ( 
.A(n_4914),
.B(n_539),
.Y(n_4989)
);

NAND2xp5_ASAP7_75t_L g4990 ( 
.A(n_4914),
.B(n_538),
.Y(n_4990)
);

XNOR2x1_ASAP7_75t_L g4991 ( 
.A(n_4914),
.B(n_540),
.Y(n_4991)
);

NOR2xp33_ASAP7_75t_L g4992 ( 
.A(n_4914),
.B(n_541),
.Y(n_4992)
);

NAND2xp5_ASAP7_75t_SL g4993 ( 
.A(n_4871),
.B(n_542),
.Y(n_4993)
);

NAND2xp5_ASAP7_75t_SL g4994 ( 
.A(n_4871),
.B(n_542),
.Y(n_4994)
);

OAI21xp5_ASAP7_75t_L g4995 ( 
.A1(n_4911),
.A2(n_544),
.B(n_545),
.Y(n_4995)
);

O2A1O1Ixp5_ASAP7_75t_L g4996 ( 
.A1(n_4868),
.A2(n_546),
.B(n_544),
.C(n_545),
.Y(n_4996)
);

NAND2xp33_ASAP7_75t_L g4997 ( 
.A(n_4914),
.B(n_547),
.Y(n_4997)
);

OAI21xp33_ASAP7_75t_L g4998 ( 
.A1(n_4914),
.A2(n_556),
.B(n_548),
.Y(n_4998)
);

OAI22x1_ASAP7_75t_L g4999 ( 
.A1(n_4911),
.A2(n_551),
.B1(n_549),
.B2(n_550),
.Y(n_4999)
);

OAI211xp5_ASAP7_75t_SL g5000 ( 
.A1(n_4914),
.A2(n_551),
.B(n_549),
.C(n_550),
.Y(n_5000)
);

INVx1_ASAP7_75t_L g5001 ( 
.A(n_4907),
.Y(n_5001)
);

NAND3xp33_ASAP7_75t_SL g5002 ( 
.A(n_4914),
.B(n_552),
.C(n_553),
.Y(n_5002)
);

NOR2xp33_ASAP7_75t_SL g5003 ( 
.A(n_4914),
.B(n_552),
.Y(n_5003)
);

OR2x2_ASAP7_75t_L g5004 ( 
.A(n_4914),
.B(n_553),
.Y(n_5004)
);

AOI21xp5_ASAP7_75t_L g5005 ( 
.A1(n_4868),
.A2(n_554),
.B(n_555),
.Y(n_5005)
);

INVx2_ASAP7_75t_SL g5006 ( 
.A(n_4920),
.Y(n_5006)
);

INVx1_ASAP7_75t_L g5007 ( 
.A(n_4907),
.Y(n_5007)
);

AOI22xp5_ASAP7_75t_L g5008 ( 
.A1(n_4957),
.A2(n_556),
.B1(n_554),
.B2(n_555),
.Y(n_5008)
);

AOI211xp5_ASAP7_75t_L g5009 ( 
.A1(n_4933),
.A2(n_559),
.B(n_557),
.C(n_558),
.Y(n_5009)
);

AOI221xp5_ASAP7_75t_L g5010 ( 
.A1(n_4931),
.A2(n_560),
.B1(n_557),
.B2(n_559),
.C(n_562),
.Y(n_5010)
);

NOR3x1_ASAP7_75t_L g5011 ( 
.A(n_4935),
.B(n_563),
.C(n_562),
.Y(n_5011)
);

AOI21xp5_ASAP7_75t_L g5012 ( 
.A1(n_4970),
.A2(n_560),
.B(n_564),
.Y(n_5012)
);

OAI221xp5_ASAP7_75t_L g5013 ( 
.A1(n_4951),
.A2(n_567),
.B1(n_565),
.B2(n_566),
.C(n_568),
.Y(n_5013)
);

OAI21xp5_ASAP7_75t_SL g5014 ( 
.A1(n_4932),
.A2(n_565),
.B(n_566),
.Y(n_5014)
);

OAI211xp5_ASAP7_75t_SL g5015 ( 
.A1(n_4962),
.A2(n_569),
.B(n_567),
.C(n_568),
.Y(n_5015)
);

OAI22xp5_ASAP7_75t_L g5016 ( 
.A1(n_4964),
.A2(n_572),
.B1(n_569),
.B2(n_570),
.Y(n_5016)
);

AOI22xp5_ASAP7_75t_L g5017 ( 
.A1(n_4936),
.A2(n_573),
.B1(n_570),
.B2(n_572),
.Y(n_5017)
);

OAI21xp33_ASAP7_75t_L g5018 ( 
.A1(n_4929),
.A2(n_573),
.B(n_574),
.Y(n_5018)
);

AOI221xp5_ASAP7_75t_L g5019 ( 
.A1(n_4926),
.A2(n_577),
.B1(n_574),
.B2(n_575),
.C(n_578),
.Y(n_5019)
);

NAND2xp5_ASAP7_75t_L g5020 ( 
.A(n_4954),
.B(n_577),
.Y(n_5020)
);

OAI21xp5_ASAP7_75t_SL g5021 ( 
.A1(n_4941),
.A2(n_578),
.B(n_579),
.Y(n_5021)
);

NAND4xp25_ASAP7_75t_SL g5022 ( 
.A(n_4923),
.B(n_581),
.C(n_579),
.D(n_580),
.Y(n_5022)
);

OAI211xp5_ASAP7_75t_SL g5023 ( 
.A1(n_4968),
.A2(n_583),
.B(n_580),
.C(n_582),
.Y(n_5023)
);

AOI221xp5_ASAP7_75t_L g5024 ( 
.A1(n_4934),
.A2(n_585),
.B1(n_582),
.B2(n_584),
.C(n_586),
.Y(n_5024)
);

AOI222xp33_ASAP7_75t_L g5025 ( 
.A1(n_4927),
.A2(n_586),
.B1(n_588),
.B2(n_584),
.C1(n_585),
.C2(n_587),
.Y(n_5025)
);

NAND2xp5_ASAP7_75t_L g5026 ( 
.A(n_4978),
.B(n_4989),
.Y(n_5026)
);

NAND2x1_ASAP7_75t_L g5027 ( 
.A(n_4928),
.B(n_588),
.Y(n_5027)
);

NOR3xp33_ASAP7_75t_L g5028 ( 
.A(n_4972),
.B(n_589),
.C(n_590),
.Y(n_5028)
);

OAI221xp5_ASAP7_75t_L g5029 ( 
.A1(n_4956),
.A2(n_591),
.B1(n_589),
.B2(n_590),
.C(n_592),
.Y(n_5029)
);

AOI22xp5_ASAP7_75t_L g5030 ( 
.A1(n_4986),
.A2(n_594),
.B1(n_592),
.B2(n_593),
.Y(n_5030)
);

NAND3xp33_ASAP7_75t_L g5031 ( 
.A(n_4997),
.B(n_593),
.C(n_594),
.Y(n_5031)
);

OAI21xp5_ASAP7_75t_SL g5032 ( 
.A1(n_4991),
.A2(n_595),
.B(n_596),
.Y(n_5032)
);

AOI21xp5_ASAP7_75t_L g5033 ( 
.A1(n_4980),
.A2(n_595),
.B(n_596),
.Y(n_5033)
);

OAI211xp5_ASAP7_75t_SL g5034 ( 
.A1(n_4971),
.A2(n_599),
.B(n_597),
.C(n_598),
.Y(n_5034)
);

NOR2xp33_ASAP7_75t_L g5035 ( 
.A(n_4975),
.B(n_598),
.Y(n_5035)
);

OAI222xp33_ASAP7_75t_R g5036 ( 
.A1(n_5006),
.A2(n_602),
.B1(n_604),
.B2(n_600),
.C1(n_601),
.C2(n_603),
.Y(n_5036)
);

AOI21xp5_ASAP7_75t_L g5037 ( 
.A1(n_4993),
.A2(n_600),
.B(n_601),
.Y(n_5037)
);

AOI221x1_ASAP7_75t_L g5038 ( 
.A1(n_5005),
.A2(n_604),
.B1(n_602),
.B2(n_603),
.C(n_605),
.Y(n_5038)
);

NOR3xp33_ASAP7_75t_L g5039 ( 
.A(n_4994),
.B(n_605),
.C(n_606),
.Y(n_5039)
);

NOR4xp25_ASAP7_75t_L g5040 ( 
.A(n_4960),
.B(n_608),
.C(n_606),
.D(n_607),
.Y(n_5040)
);

NAND2xp5_ASAP7_75t_L g5041 ( 
.A(n_4930),
.B(n_607),
.Y(n_5041)
);

OAI21xp5_ASAP7_75t_SL g5042 ( 
.A1(n_5007),
.A2(n_608),
.B(n_609),
.Y(n_5042)
);

OAI211xp5_ASAP7_75t_L g5043 ( 
.A1(n_4922),
.A2(n_618),
.B(n_626),
.C(n_609),
.Y(n_5043)
);

OAI21xp5_ASAP7_75t_SL g5044 ( 
.A1(n_4974),
.A2(n_5001),
.B(n_4981),
.Y(n_5044)
);

OAI221xp5_ASAP7_75t_L g5045 ( 
.A1(n_4996),
.A2(n_613),
.B1(n_611),
.B2(n_612),
.C(n_614),
.Y(n_5045)
);

NOR2xp33_ASAP7_75t_L g5046 ( 
.A(n_5003),
.B(n_612),
.Y(n_5046)
);

NAND3xp33_ASAP7_75t_L g5047 ( 
.A(n_4950),
.B(n_614),
.C(n_615),
.Y(n_5047)
);

AOI21xp33_ASAP7_75t_L g5048 ( 
.A1(n_4983),
.A2(n_616),
.B(n_617),
.Y(n_5048)
);

AOI22xp5_ASAP7_75t_L g5049 ( 
.A1(n_4992),
.A2(n_619),
.B1(n_616),
.B2(n_617),
.Y(n_5049)
);

INVx1_ASAP7_75t_L g5050 ( 
.A(n_4987),
.Y(n_5050)
);

AOI211x1_ASAP7_75t_SL g5051 ( 
.A1(n_4976),
.A2(n_5002),
.B(n_5000),
.C(n_4973),
.Y(n_5051)
);

AOI22xp5_ASAP7_75t_L g5052 ( 
.A1(n_4948),
.A2(n_621),
.B1(n_619),
.B2(n_620),
.Y(n_5052)
);

AOI211x1_ASAP7_75t_L g5053 ( 
.A1(n_4995),
.A2(n_622),
.B(n_620),
.C(n_621),
.Y(n_5053)
);

AOI22xp5_ASAP7_75t_L g5054 ( 
.A1(n_4925),
.A2(n_4952),
.B1(n_4977),
.B2(n_4969),
.Y(n_5054)
);

INVx1_ASAP7_75t_L g5055 ( 
.A(n_4924),
.Y(n_5055)
);

AOI21xp5_ASAP7_75t_L g5056 ( 
.A1(n_4938),
.A2(n_622),
.B(n_623),
.Y(n_5056)
);

AOI22xp5_ASAP7_75t_L g5057 ( 
.A1(n_4984),
.A2(n_627),
.B1(n_624),
.B2(n_625),
.Y(n_5057)
);

OAI211xp5_ASAP7_75t_SL g5058 ( 
.A1(n_4940),
.A2(n_4943),
.B(n_4955),
.C(n_4988),
.Y(n_5058)
);

O2A1O1Ixp33_ASAP7_75t_L g5059 ( 
.A1(n_4947),
.A2(n_4944),
.B(n_4953),
.C(n_4985),
.Y(n_5059)
);

AOI321xp33_ASAP7_75t_L g5060 ( 
.A1(n_4961),
.A2(n_628),
.A3(n_633),
.B1(n_625),
.B2(n_627),
.C(n_629),
.Y(n_5060)
);

AOI221xp5_ASAP7_75t_L g5061 ( 
.A1(n_4963),
.A2(n_4946),
.B1(n_4967),
.B2(n_4990),
.C(n_4998),
.Y(n_5061)
);

AOI221x1_ASAP7_75t_L g5062 ( 
.A1(n_4999),
.A2(n_634),
.B1(n_628),
.B2(n_633),
.C(n_635),
.Y(n_5062)
);

A2O1A1Ixp33_ASAP7_75t_L g5063 ( 
.A1(n_4939),
.A2(n_638),
.B(n_635),
.C(n_637),
.Y(n_5063)
);

AOI21xp5_ASAP7_75t_L g5064 ( 
.A1(n_4959),
.A2(n_639),
.B(n_640),
.Y(n_5064)
);

AOI21xp5_ASAP7_75t_L g5065 ( 
.A1(n_4979),
.A2(n_639),
.B(n_640),
.Y(n_5065)
);

OAI321xp33_ASAP7_75t_L g5066 ( 
.A1(n_5004),
.A2(n_644),
.A3(n_646),
.B1(n_642),
.B2(n_643),
.C(n_645),
.Y(n_5066)
);

OAI21xp33_ASAP7_75t_L g5067 ( 
.A1(n_4965),
.A2(n_642),
.B(n_643),
.Y(n_5067)
);

AO21x1_ASAP7_75t_L g5068 ( 
.A1(n_4949),
.A2(n_645),
.B(n_648),
.Y(n_5068)
);

AOI211xp5_ASAP7_75t_L g5069 ( 
.A1(n_4958),
.A2(n_650),
.B(n_648),
.C(n_649),
.Y(n_5069)
);

NOR3xp33_ASAP7_75t_L g5070 ( 
.A(n_4942),
.B(n_651),
.C(n_653),
.Y(n_5070)
);

AOI22xp5_ASAP7_75t_L g5071 ( 
.A1(n_4966),
.A2(n_654),
.B1(n_651),
.B2(n_653),
.Y(n_5071)
);

OAI211xp5_ASAP7_75t_L g5072 ( 
.A1(n_4982),
.A2(n_663),
.B(n_671),
.C(n_655),
.Y(n_5072)
);

AOI21xp5_ASAP7_75t_L g5073 ( 
.A1(n_4945),
.A2(n_655),
.B(n_656),
.Y(n_5073)
);

AOI221xp5_ASAP7_75t_L g5074 ( 
.A1(n_4937),
.A2(n_658),
.B1(n_656),
.B2(n_657),
.C(n_659),
.Y(n_5074)
);

NAND2xp5_ASAP7_75t_SL g5075 ( 
.A(n_4954),
.B(n_657),
.Y(n_5075)
);

AOI22xp5_ASAP7_75t_L g5076 ( 
.A1(n_4957),
.A2(n_660),
.B1(n_658),
.B2(n_659),
.Y(n_5076)
);

NOR2xp33_ASAP7_75t_L g5077 ( 
.A(n_4957),
.B(n_660),
.Y(n_5077)
);

O2A1O1Ixp33_ASAP7_75t_L g5078 ( 
.A1(n_4976),
.A2(n_663),
.B(n_661),
.C(n_662),
.Y(n_5078)
);

NOR4xp25_ASAP7_75t_L g5079 ( 
.A(n_4951),
.B(n_664),
.C(n_661),
.D(n_662),
.Y(n_5079)
);

AOI222xp33_ASAP7_75t_L g5080 ( 
.A1(n_4932),
.A2(n_666),
.B1(n_668),
.B2(n_664),
.C1(n_665),
.C2(n_667),
.Y(n_5080)
);

NAND3xp33_ASAP7_75t_L g5081 ( 
.A(n_4997),
.B(n_665),
.C(n_667),
.Y(n_5081)
);

NOR2xp33_ASAP7_75t_SL g5082 ( 
.A(n_4954),
.B(n_668),
.Y(n_5082)
);

AOI21xp5_ASAP7_75t_L g5083 ( 
.A1(n_4970),
.A2(n_669),
.B(n_670),
.Y(n_5083)
);

OAI221xp5_ASAP7_75t_SL g5084 ( 
.A1(n_4951),
.A2(n_673),
.B1(n_671),
.B2(n_672),
.C(n_674),
.Y(n_5084)
);

NAND3xp33_ASAP7_75t_L g5085 ( 
.A(n_4997),
.B(n_672),
.C(n_675),
.Y(n_5085)
);

AOI21xp5_ASAP7_75t_L g5086 ( 
.A1(n_4970),
.A2(n_675),
.B(n_676),
.Y(n_5086)
);

OAI31xp33_ASAP7_75t_L g5087 ( 
.A1(n_5000),
.A2(n_678),
.A3(n_676),
.B(n_677),
.Y(n_5087)
);

AOI221xp5_ASAP7_75t_L g5088 ( 
.A1(n_4931),
.A2(n_679),
.B1(n_677),
.B2(n_678),
.C(n_680),
.Y(n_5088)
);

AOI222xp33_ASAP7_75t_L g5089 ( 
.A1(n_4932),
.A2(n_681),
.B1(n_684),
.B2(n_679),
.C1(n_680),
.C2(n_683),
.Y(n_5089)
);

AOI221xp5_ASAP7_75t_L g5090 ( 
.A1(n_4931),
.A2(n_686),
.B1(n_683),
.B2(n_685),
.C(n_687),
.Y(n_5090)
);

AOI222xp33_ASAP7_75t_L g5091 ( 
.A1(n_4932),
.A2(n_688),
.B1(n_690),
.B2(n_685),
.C1(n_687),
.C2(n_689),
.Y(n_5091)
);

AOI21xp5_ASAP7_75t_L g5092 ( 
.A1(n_4970),
.A2(n_688),
.B(n_690),
.Y(n_5092)
);

INVx2_ASAP7_75t_L g5093 ( 
.A(n_5027),
.Y(n_5093)
);

INVx1_ASAP7_75t_L g5094 ( 
.A(n_5068),
.Y(n_5094)
);

INVx1_ASAP7_75t_L g5095 ( 
.A(n_5020),
.Y(n_5095)
);

INVx1_ASAP7_75t_L g5096 ( 
.A(n_5026),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_5050),
.Y(n_5097)
);

INVx1_ASAP7_75t_L g5098 ( 
.A(n_5016),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_5071),
.Y(n_5099)
);

OA22x2_ASAP7_75t_L g5100 ( 
.A1(n_5014),
.A2(n_5032),
.B1(n_5021),
.B2(n_5044),
.Y(n_5100)
);

INVx1_ASAP7_75t_L g5101 ( 
.A(n_5041),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_5035),
.Y(n_5102)
);

INVx2_ASAP7_75t_L g5103 ( 
.A(n_5011),
.Y(n_5103)
);

INVxp67_ASAP7_75t_L g5104 ( 
.A(n_5082),
.Y(n_5104)
);

OAI22x1_ASAP7_75t_L g5105 ( 
.A1(n_5017),
.A2(n_693),
.B1(n_691),
.B2(n_692),
.Y(n_5105)
);

INVx1_ASAP7_75t_L g5106 ( 
.A(n_5046),
.Y(n_5106)
);

INVx2_ASAP7_75t_SL g5107 ( 
.A(n_5055),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_5077),
.Y(n_5108)
);

INVx1_ASAP7_75t_L g5109 ( 
.A(n_5031),
.Y(n_5109)
);

INVx1_ASAP7_75t_L g5110 ( 
.A(n_5081),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_5085),
.Y(n_5111)
);

INVxp67_ASAP7_75t_L g5112 ( 
.A(n_5075),
.Y(n_5112)
);

INVx1_ASAP7_75t_L g5113 ( 
.A(n_5062),
.Y(n_5113)
);

AO22x2_ASAP7_75t_L g5114 ( 
.A1(n_5053),
.A2(n_693),
.B1(n_691),
.B2(n_692),
.Y(n_5114)
);

OAI22x1_ASAP7_75t_L g5115 ( 
.A1(n_5054),
.A2(n_696),
.B1(n_694),
.B2(n_695),
.Y(n_5115)
);

INVxp67_ASAP7_75t_SL g5116 ( 
.A(n_5078),
.Y(n_5116)
);

INVx1_ASAP7_75t_L g5117 ( 
.A(n_5047),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_5067),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_5008),
.Y(n_5119)
);

AO22x2_ASAP7_75t_L g5120 ( 
.A1(n_5043),
.A2(n_5073),
.B1(n_5042),
.B2(n_5038),
.Y(n_5120)
);

INVx1_ASAP7_75t_L g5121 ( 
.A(n_5076),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_5059),
.Y(n_5122)
);

OAI22xp5_ASAP7_75t_L g5123 ( 
.A1(n_5084),
.A2(n_697),
.B1(n_695),
.B2(n_696),
.Y(n_5123)
);

OAI22xp33_ASAP7_75t_L g5124 ( 
.A1(n_5045),
.A2(n_700),
.B1(n_698),
.B2(n_699),
.Y(n_5124)
);

OAI221xp5_ASAP7_75t_SL g5125 ( 
.A1(n_5061),
.A2(n_5087),
.B1(n_5079),
.B2(n_5009),
.C(n_5070),
.Y(n_5125)
);

AOI22xp5_ASAP7_75t_L g5126 ( 
.A1(n_5022),
.A2(n_701),
.B1(n_698),
.B2(n_699),
.Y(n_5126)
);

INVx1_ASAP7_75t_L g5127 ( 
.A(n_5018),
.Y(n_5127)
);

OAI22x1_ASAP7_75t_L g5128 ( 
.A1(n_5030),
.A2(n_704),
.B1(n_702),
.B2(n_703),
.Y(n_5128)
);

INVx1_ASAP7_75t_L g5129 ( 
.A(n_5057),
.Y(n_5129)
);

AOI31xp33_ASAP7_75t_L g5130 ( 
.A1(n_5048),
.A2(n_713),
.A3(n_721),
.B(n_704),
.Y(n_5130)
);

A2O1A1Ixp33_ASAP7_75t_SL g5131 ( 
.A1(n_5058),
.A2(n_707),
.B(n_705),
.C(n_706),
.Y(n_5131)
);

NAND2xp5_ASAP7_75t_SL g5132 ( 
.A(n_5040),
.B(n_705),
.Y(n_5132)
);

AO22x1_ASAP7_75t_L g5133 ( 
.A1(n_5028),
.A2(n_709),
.B1(n_706),
.B2(n_708),
.Y(n_5133)
);

BUFx2_ASAP7_75t_L g5134 ( 
.A(n_5063),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_5049),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_5060),
.Y(n_5136)
);

A2O1A1Ixp33_ASAP7_75t_L g5137 ( 
.A1(n_5065),
.A2(n_5064),
.B(n_5012),
.C(n_5037),
.Y(n_5137)
);

OAI22xp5_ASAP7_75t_L g5138 ( 
.A1(n_5013),
.A2(n_712),
.B1(n_708),
.B2(n_711),
.Y(n_5138)
);

AOI22xp5_ASAP7_75t_L g5139 ( 
.A1(n_5039),
.A2(n_714),
.B1(n_711),
.B2(n_712),
.Y(n_5139)
);

AOI22xp5_ASAP7_75t_L g5140 ( 
.A1(n_5072),
.A2(n_716),
.B1(n_714),
.B2(n_715),
.Y(n_5140)
);

AOI22x1_ASAP7_75t_L g5141 ( 
.A1(n_5080),
.A2(n_719),
.B1(n_717),
.B2(n_718),
.Y(n_5141)
);

INVx1_ASAP7_75t_L g5142 ( 
.A(n_5052),
.Y(n_5142)
);

AO22x1_ASAP7_75t_L g5143 ( 
.A1(n_5036),
.A2(n_719),
.B1(n_717),
.B2(n_718),
.Y(n_5143)
);

INVx1_ASAP7_75t_L g5144 ( 
.A(n_5029),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_5023),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_5034),
.Y(n_5146)
);

OA22x2_ASAP7_75t_L g5147 ( 
.A1(n_5051),
.A2(n_723),
.B1(n_720),
.B2(n_722),
.Y(n_5147)
);

INVx1_ASAP7_75t_L g5148 ( 
.A(n_5025),
.Y(n_5148)
);

A2O1A1Ixp33_ASAP7_75t_SL g5149 ( 
.A1(n_5066),
.A2(n_5069),
.B(n_5056),
.C(n_5033),
.Y(n_5149)
);

AOI22xp5_ASAP7_75t_L g5150 ( 
.A1(n_5074),
.A2(n_725),
.B1(n_723),
.B2(n_724),
.Y(n_5150)
);

BUFx6f_ASAP7_75t_L g5151 ( 
.A(n_5089),
.Y(n_5151)
);

INVx1_ASAP7_75t_L g5152 ( 
.A(n_5015),
.Y(n_5152)
);

AOI22xp5_ASAP7_75t_L g5153 ( 
.A1(n_5091),
.A2(n_726),
.B1(n_724),
.B2(n_725),
.Y(n_5153)
);

INVx1_ASAP7_75t_L g5154 ( 
.A(n_5083),
.Y(n_5154)
);

O2A1O1Ixp33_ASAP7_75t_L g5155 ( 
.A1(n_5086),
.A2(n_728),
.B(n_726),
.C(n_727),
.Y(n_5155)
);

AOI22xp5_ASAP7_75t_L g5156 ( 
.A1(n_5010),
.A2(n_731),
.B1(n_728),
.B2(n_729),
.Y(n_5156)
);

INVx1_ASAP7_75t_L g5157 ( 
.A(n_5092),
.Y(n_5157)
);

AOI22xp33_ASAP7_75t_L g5158 ( 
.A1(n_5024),
.A2(n_733),
.B1(n_731),
.B2(n_732),
.Y(n_5158)
);

AOI221xp5_ASAP7_75t_L g5159 ( 
.A1(n_5090),
.A2(n_734),
.B1(n_732),
.B2(n_733),
.C(n_735),
.Y(n_5159)
);

INVx2_ASAP7_75t_L g5160 ( 
.A(n_5019),
.Y(n_5160)
);

A2O1A1Ixp33_ASAP7_75t_L g5161 ( 
.A1(n_5088),
.A2(n_737),
.B(n_735),
.C(n_736),
.Y(n_5161)
);

AO22x2_ASAP7_75t_L g5162 ( 
.A1(n_5016),
.A2(n_739),
.B1(n_737),
.B2(n_738),
.Y(n_5162)
);

OAI22xp5_ASAP7_75t_L g5163 ( 
.A1(n_5047),
.A2(n_740),
.B1(n_738),
.B2(n_739),
.Y(n_5163)
);

AOI22x1_ASAP7_75t_L g5164 ( 
.A1(n_5080),
.A2(n_742),
.B1(n_740),
.B2(n_741),
.Y(n_5164)
);

INVx1_ASAP7_75t_L g5165 ( 
.A(n_5027),
.Y(n_5165)
);

AOI22xp5_ASAP7_75t_L g5166 ( 
.A1(n_5016),
.A2(n_744),
.B1(n_741),
.B2(n_743),
.Y(n_5166)
);

INVx1_ASAP7_75t_L g5167 ( 
.A(n_5027),
.Y(n_5167)
);

INVx1_ASAP7_75t_L g5168 ( 
.A(n_5027),
.Y(n_5168)
);

INVx1_ASAP7_75t_L g5169 ( 
.A(n_5027),
.Y(n_5169)
);

INVxp67_ASAP7_75t_L g5170 ( 
.A(n_5082),
.Y(n_5170)
);

AO22x2_ASAP7_75t_L g5171 ( 
.A1(n_5016),
.A2(n_748),
.B1(n_745),
.B2(n_746),
.Y(n_5171)
);

OAI22xp5_ASAP7_75t_L g5172 ( 
.A1(n_5047),
.A2(n_749),
.B1(n_745),
.B2(n_748),
.Y(n_5172)
);

OAI22xp5_ASAP7_75t_L g5173 ( 
.A1(n_5047),
.A2(n_751),
.B1(n_749),
.B2(n_750),
.Y(n_5173)
);

HB1xp67_ASAP7_75t_L g5174 ( 
.A(n_5027),
.Y(n_5174)
);

OAI22xp5_ASAP7_75t_L g5175 ( 
.A1(n_5047),
.A2(n_752),
.B1(n_750),
.B2(n_751),
.Y(n_5175)
);

OAI22xp5_ASAP7_75t_L g5176 ( 
.A1(n_5047),
.A2(n_754),
.B1(n_752),
.B2(n_753),
.Y(n_5176)
);

AOI22xp5_ASAP7_75t_L g5177 ( 
.A1(n_5016),
.A2(n_755),
.B1(n_753),
.B2(n_754),
.Y(n_5177)
);

OAI22xp5_ASAP7_75t_L g5178 ( 
.A1(n_5047),
.A2(n_760),
.B1(n_756),
.B2(n_759),
.Y(n_5178)
);

OAI22xp5_ASAP7_75t_L g5179 ( 
.A1(n_5126),
.A2(n_761),
.B1(n_756),
.B2(n_760),
.Y(n_5179)
);

INVxp67_ASAP7_75t_SL g5180 ( 
.A(n_5174),
.Y(n_5180)
);

AOI211x1_ASAP7_75t_SL g5181 ( 
.A1(n_5137),
.A2(n_764),
.B(n_762),
.C(n_763),
.Y(n_5181)
);

AOI22xp33_ASAP7_75t_L g5182 ( 
.A1(n_5097),
.A2(n_764),
.B1(n_762),
.B2(n_763),
.Y(n_5182)
);

NOR2xp33_ASAP7_75t_SL g5183 ( 
.A(n_5093),
.B(n_767),
.Y(n_5183)
);

OAI21xp5_ASAP7_75t_SL g5184 ( 
.A1(n_5153),
.A2(n_768),
.B(n_767),
.Y(n_5184)
);

NAND4xp25_ASAP7_75t_L g5185 ( 
.A(n_5125),
.B(n_769),
.C(n_765),
.D(n_768),
.Y(n_5185)
);

AND2x2_ASAP7_75t_L g5186 ( 
.A(n_5120),
.B(n_765),
.Y(n_5186)
);

OAI22xp5_ASAP7_75t_L g5187 ( 
.A1(n_5158),
.A2(n_772),
.B1(n_770),
.B2(n_771),
.Y(n_5187)
);

NOR3xp33_ASAP7_75t_L g5188 ( 
.A(n_5122),
.B(n_771),
.C(n_772),
.Y(n_5188)
);

NAND4xp25_ASAP7_75t_L g5189 ( 
.A(n_5149),
.B(n_775),
.C(n_773),
.D(n_774),
.Y(n_5189)
);

OAI221xp5_ASAP7_75t_L g5190 ( 
.A1(n_5131),
.A2(n_5094),
.B1(n_5164),
.B2(n_5141),
.C(n_5104),
.Y(n_5190)
);

AOI221xp5_ASAP7_75t_L g5191 ( 
.A1(n_5143),
.A2(n_777),
.B1(n_774),
.B2(n_776),
.C(n_778),
.Y(n_5191)
);

A2O1A1Ixp33_ASAP7_75t_L g5192 ( 
.A1(n_5155),
.A2(n_779),
.B(n_777),
.C(n_778),
.Y(n_5192)
);

OAI21xp5_ASAP7_75t_L g5193 ( 
.A1(n_5170),
.A2(n_779),
.B(n_780),
.Y(n_5193)
);

OAI211xp5_ASAP7_75t_L g5194 ( 
.A1(n_5132),
.A2(n_5167),
.B(n_5168),
.C(n_5165),
.Y(n_5194)
);

NAND2xp5_ASAP7_75t_L g5195 ( 
.A(n_5169),
.B(n_780),
.Y(n_5195)
);

AOI221xp5_ASAP7_75t_SL g5196 ( 
.A1(n_5112),
.A2(n_783),
.B1(n_781),
.B2(n_782),
.C(n_784),
.Y(n_5196)
);

NOR2xp33_ASAP7_75t_L g5197 ( 
.A(n_5113),
.B(n_781),
.Y(n_5197)
);

AOI221xp5_ASAP7_75t_L g5198 ( 
.A1(n_5124),
.A2(n_785),
.B1(n_782),
.B2(n_783),
.C(n_786),
.Y(n_5198)
);

XOR2x2_ASAP7_75t_L g5199 ( 
.A(n_5100),
.B(n_785),
.Y(n_5199)
);

AOI211xp5_ASAP7_75t_L g5200 ( 
.A1(n_5123),
.A2(n_789),
.B(n_786),
.C(n_787),
.Y(n_5200)
);

AOI221xp5_ASAP7_75t_L g5201 ( 
.A1(n_5120),
.A2(n_791),
.B1(n_787),
.B2(n_790),
.C(n_793),
.Y(n_5201)
);

INVx1_ASAP7_75t_L g5202 ( 
.A(n_5162),
.Y(n_5202)
);

AOI211xp5_ASAP7_75t_L g5203 ( 
.A1(n_5163),
.A2(n_794),
.B(n_790),
.C(n_791),
.Y(n_5203)
);

AOI221xp5_ASAP7_75t_L g5204 ( 
.A1(n_5116),
.A2(n_797),
.B1(n_794),
.B2(n_796),
.C(n_798),
.Y(n_5204)
);

AND2x2_ASAP7_75t_L g5205 ( 
.A(n_5103),
.B(n_796),
.Y(n_5205)
);

AOI222xp33_ASAP7_75t_L g5206 ( 
.A1(n_5136),
.A2(n_802),
.B1(n_804),
.B2(n_799),
.C1(n_800),
.C2(n_803),
.Y(n_5206)
);

AOI221xp5_ASAP7_75t_L g5207 ( 
.A1(n_5098),
.A2(n_803),
.B1(n_799),
.B2(n_802),
.C(n_805),
.Y(n_5207)
);

NAND2xp5_ASAP7_75t_L g5208 ( 
.A(n_5133),
.B(n_805),
.Y(n_5208)
);

OAI22xp33_ASAP7_75t_L g5209 ( 
.A1(n_5140),
.A2(n_808),
.B1(n_806),
.B2(n_807),
.Y(n_5209)
);

O2A1O1Ixp33_ASAP7_75t_L g5210 ( 
.A1(n_5130),
.A2(n_811),
.B(n_809),
.C(n_810),
.Y(n_5210)
);

OAI221xp5_ASAP7_75t_L g5211 ( 
.A1(n_5150),
.A2(n_811),
.B1(n_809),
.B2(n_810),
.C(n_812),
.Y(n_5211)
);

AOI211xp5_ASAP7_75t_L g5212 ( 
.A1(n_5172),
.A2(n_815),
.B(n_813),
.C(n_814),
.Y(n_5212)
);

INVx1_ASAP7_75t_L g5213 ( 
.A(n_5162),
.Y(n_5213)
);

AOI221xp5_ASAP7_75t_L g5214 ( 
.A1(n_5145),
.A2(n_816),
.B1(n_813),
.B2(n_815),
.C(n_817),
.Y(n_5214)
);

O2A1O1Ixp5_ASAP7_75t_L g5215 ( 
.A1(n_5146),
.A2(n_5152),
.B(n_5118),
.C(n_5117),
.Y(n_5215)
);

OAI221xp5_ASAP7_75t_L g5216 ( 
.A1(n_5161),
.A2(n_820),
.B1(n_817),
.B2(n_819),
.C(n_821),
.Y(n_5216)
);

AOI221xp5_ASAP7_75t_L g5217 ( 
.A1(n_5173),
.A2(n_5175),
.B1(n_5178),
.B2(n_5176),
.C(n_5114),
.Y(n_5217)
);

NOR2xp33_ASAP7_75t_L g5218 ( 
.A(n_5107),
.B(n_820),
.Y(n_5218)
);

OAI21xp33_ASAP7_75t_L g5219 ( 
.A1(n_5099),
.A2(n_822),
.B(n_823),
.Y(n_5219)
);

NAND2xp33_ASAP7_75t_L g5220 ( 
.A(n_5115),
.B(n_823),
.Y(n_5220)
);

NAND2xp5_ASAP7_75t_L g5221 ( 
.A(n_5171),
.B(n_824),
.Y(n_5221)
);

NOR2x1_ASAP7_75t_L g5222 ( 
.A(n_5154),
.B(n_5157),
.Y(n_5222)
);

NAND2xp5_ASAP7_75t_L g5223 ( 
.A(n_5171),
.B(n_825),
.Y(n_5223)
);

AOI22xp5_ASAP7_75t_L g5224 ( 
.A1(n_5148),
.A2(n_828),
.B1(n_826),
.B2(n_827),
.Y(n_5224)
);

OAI211xp5_ASAP7_75t_L g5225 ( 
.A1(n_5156),
.A2(n_829),
.B(n_826),
.C(n_827),
.Y(n_5225)
);

OAI211xp5_ASAP7_75t_L g5226 ( 
.A1(n_5159),
.A2(n_831),
.B(n_829),
.C(n_830),
.Y(n_5226)
);

NOR2xp33_ASAP7_75t_L g5227 ( 
.A(n_5151),
.B(n_830),
.Y(n_5227)
);

OAI221xp5_ASAP7_75t_L g5228 ( 
.A1(n_5144),
.A2(n_835),
.B1(n_833),
.B2(n_834),
.C(n_836),
.Y(n_5228)
);

INVx1_ASAP7_75t_SL g5229 ( 
.A(n_5147),
.Y(n_5229)
);

OAI211xp5_ASAP7_75t_L g5230 ( 
.A1(n_5139),
.A2(n_836),
.B(n_834),
.C(n_835),
.Y(n_5230)
);

OAI21xp5_ASAP7_75t_L g5231 ( 
.A1(n_5138),
.A2(n_837),
.B(n_838),
.Y(n_5231)
);

OAI22xp5_ASAP7_75t_L g5232 ( 
.A1(n_5166),
.A2(n_839),
.B1(n_837),
.B2(n_838),
.Y(n_5232)
);

OAI211xp5_ASAP7_75t_SL g5233 ( 
.A1(n_5096),
.A2(n_844),
.B(n_841),
.C(n_842),
.Y(n_5233)
);

NAND3xp33_ASAP7_75t_SL g5234 ( 
.A(n_5134),
.B(n_841),
.C(n_844),
.Y(n_5234)
);

NAND3xp33_ASAP7_75t_L g5235 ( 
.A(n_5151),
.B(n_846),
.C(n_847),
.Y(n_5235)
);

INVx3_ASAP7_75t_L g5236 ( 
.A(n_5114),
.Y(n_5236)
);

NOR2xp33_ASAP7_75t_L g5237 ( 
.A(n_5177),
.B(n_846),
.Y(n_5237)
);

OAI22xp5_ASAP7_75t_L g5238 ( 
.A1(n_5109),
.A2(n_849),
.B1(n_847),
.B2(n_848),
.Y(n_5238)
);

OAI21xp33_ASAP7_75t_SL g5239 ( 
.A1(n_5110),
.A2(n_850),
.B(n_851),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_5105),
.Y(n_5240)
);

OAI221xp5_ASAP7_75t_SL g5241 ( 
.A1(n_5111),
.A2(n_854),
.B1(n_850),
.B2(n_853),
.C(n_855),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_5128),
.Y(n_5242)
);

AOI221xp5_ASAP7_75t_L g5243 ( 
.A1(n_5127),
.A2(n_5142),
.B1(n_5121),
.B2(n_5119),
.C(n_5129),
.Y(n_5243)
);

A2O1A1Ixp33_ASAP7_75t_SL g5244 ( 
.A1(n_5108),
.A2(n_856),
.B(n_853),
.C(n_855),
.Y(n_5244)
);

AOI211xp5_ASAP7_75t_L g5245 ( 
.A1(n_5135),
.A2(n_858),
.B(n_856),
.C(n_857),
.Y(n_5245)
);

AOI221xp5_ASAP7_75t_L g5246 ( 
.A1(n_5102),
.A2(n_859),
.B1(n_857),
.B2(n_858),
.C(n_860),
.Y(n_5246)
);

OAI21xp33_ASAP7_75t_L g5247 ( 
.A1(n_5160),
.A2(n_859),
.B(n_861),
.Y(n_5247)
);

NOR4xp25_ASAP7_75t_L g5248 ( 
.A(n_5106),
.B(n_864),
.C(n_862),
.D(n_863),
.Y(n_5248)
);

INVx2_ASAP7_75t_L g5249 ( 
.A(n_5095),
.Y(n_5249)
);

NOR3xp33_ASAP7_75t_SL g5250 ( 
.A(n_5101),
.B(n_862),
.C(n_864),
.Y(n_5250)
);

NAND2xp5_ASAP7_75t_L g5251 ( 
.A(n_5143),
.B(n_866),
.Y(n_5251)
);

AOI221xp5_ASAP7_75t_L g5252 ( 
.A1(n_5143),
.A2(n_871),
.B1(n_867),
.B2(n_870),
.C(n_872),
.Y(n_5252)
);

NOR2x1_ASAP7_75t_L g5253 ( 
.A(n_5094),
.B(n_871),
.Y(n_5253)
);

OAI211xp5_ASAP7_75t_SL g5254 ( 
.A1(n_5122),
.A2(n_874),
.B(n_872),
.C(n_873),
.Y(n_5254)
);

NAND2xp5_ASAP7_75t_SL g5255 ( 
.A(n_5093),
.B(n_873),
.Y(n_5255)
);

AOI221xp5_ASAP7_75t_L g5256 ( 
.A1(n_5180),
.A2(n_876),
.B1(n_874),
.B2(n_875),
.C(n_877),
.Y(n_5256)
);

OAI22xp33_ASAP7_75t_L g5257 ( 
.A1(n_5224),
.A2(n_877),
.B1(n_875),
.B2(n_876),
.Y(n_5257)
);

AOI22xp5_ASAP7_75t_L g5258 ( 
.A1(n_5229),
.A2(n_880),
.B1(n_878),
.B2(n_879),
.Y(n_5258)
);

AOI21x1_ASAP7_75t_L g5259 ( 
.A1(n_5202),
.A2(n_879),
.B(n_880),
.Y(n_5259)
);

OAI211xp5_ASAP7_75t_L g5260 ( 
.A1(n_5239),
.A2(n_884),
.B(n_881),
.C(n_882),
.Y(n_5260)
);

O2A1O1Ixp33_ASAP7_75t_L g5261 ( 
.A1(n_5244),
.A2(n_886),
.B(n_881),
.C(n_885),
.Y(n_5261)
);

AOI222xp33_ASAP7_75t_L g5262 ( 
.A1(n_5186),
.A2(n_889),
.B1(n_891),
.B2(n_886),
.C1(n_888),
.C2(n_890),
.Y(n_5262)
);

NOR3xp33_ASAP7_75t_L g5263 ( 
.A(n_5194),
.B(n_898),
.C(n_888),
.Y(n_5263)
);

OAI221xp5_ASAP7_75t_L g5264 ( 
.A1(n_5191),
.A2(n_908),
.B1(n_917),
.B2(n_899),
.C(n_889),
.Y(n_5264)
);

INVx2_ASAP7_75t_SL g5265 ( 
.A(n_5253),
.Y(n_5265)
);

OAI21x1_ASAP7_75t_SL g5266 ( 
.A1(n_5210),
.A2(n_890),
.B(n_891),
.Y(n_5266)
);

OAI21xp33_ASAP7_75t_L g5267 ( 
.A1(n_5251),
.A2(n_892),
.B(n_894),
.Y(n_5267)
);

OAI211xp5_ASAP7_75t_SL g5268 ( 
.A1(n_5243),
.A2(n_897),
.B(n_892),
.C(n_895),
.Y(n_5268)
);

CKINVDCx16_ASAP7_75t_R g5269 ( 
.A(n_5183),
.Y(n_5269)
);

OAI22x1_ASAP7_75t_L g5270 ( 
.A1(n_5242),
.A2(n_898),
.B1(n_895),
.B2(n_897),
.Y(n_5270)
);

INVx1_ASAP7_75t_L g5271 ( 
.A(n_5221),
.Y(n_5271)
);

NAND4xp25_ASAP7_75t_SL g5272 ( 
.A(n_5252),
.B(n_902),
.C(n_900),
.D(n_901),
.Y(n_5272)
);

OR2x2_ASAP7_75t_L g5273 ( 
.A(n_5248),
.B(n_900),
.Y(n_5273)
);

AOI222xp33_ASAP7_75t_L g5274 ( 
.A1(n_5220),
.A2(n_904),
.B1(n_906),
.B2(n_902),
.C1(n_903),
.C2(n_905),
.Y(n_5274)
);

NAND3xp33_ASAP7_75t_L g5275 ( 
.A(n_5200),
.B(n_903),
.C(n_904),
.Y(n_5275)
);

AOI22xp33_ASAP7_75t_L g5276 ( 
.A1(n_5240),
.A2(n_5227),
.B1(n_5236),
.B2(n_5197),
.Y(n_5276)
);

NOR3xp33_ASAP7_75t_L g5277 ( 
.A(n_5215),
.B(n_916),
.C(n_905),
.Y(n_5277)
);

A2O1A1Ixp33_ASAP7_75t_L g5278 ( 
.A1(n_5218),
.A2(n_911),
.B(n_908),
.C(n_909),
.Y(n_5278)
);

AOI222xp33_ASAP7_75t_L g5279 ( 
.A1(n_5213),
.A2(n_912),
.B1(n_914),
.B2(n_909),
.C1(n_911),
.C2(n_913),
.Y(n_5279)
);

HB1xp67_ASAP7_75t_L g5280 ( 
.A(n_5236),
.Y(n_5280)
);

AOI31xp33_ASAP7_75t_L g5281 ( 
.A1(n_5203),
.A2(n_923),
.A3(n_932),
.B(n_914),
.Y(n_5281)
);

OAI211xp5_ASAP7_75t_SL g5282 ( 
.A1(n_5217),
.A2(n_918),
.B(n_915),
.C(n_917),
.Y(n_5282)
);

AOI322xp5_ASAP7_75t_L g5283 ( 
.A1(n_5222),
.A2(n_922),
.A3(n_921),
.B1(n_919),
.B2(n_915),
.C1(n_918),
.C2(n_920),
.Y(n_5283)
);

AOI22xp5_ASAP7_75t_L g5284 ( 
.A1(n_5199),
.A2(n_923),
.B1(n_921),
.B2(n_922),
.Y(n_5284)
);

AOI211xp5_ASAP7_75t_L g5285 ( 
.A1(n_5190),
.A2(n_926),
.B(n_924),
.C(n_925),
.Y(n_5285)
);

O2A1O1Ixp5_ASAP7_75t_SL g5286 ( 
.A1(n_5255),
.A2(n_935),
.B(n_944),
.C(n_925),
.Y(n_5286)
);

BUFx6f_ASAP7_75t_L g5287 ( 
.A(n_5249),
.Y(n_5287)
);

AOI221xp5_ASAP7_75t_L g5288 ( 
.A1(n_5189),
.A2(n_929),
.B1(n_927),
.B2(n_928),
.C(n_930),
.Y(n_5288)
);

AOI221xp5_ASAP7_75t_SL g5289 ( 
.A1(n_5185),
.A2(n_929),
.B1(n_927),
.B2(n_928),
.C(n_930),
.Y(n_5289)
);

NAND2xp5_ASAP7_75t_L g5290 ( 
.A(n_5201),
.B(n_932),
.Y(n_5290)
);

AOI31xp33_ASAP7_75t_L g5291 ( 
.A1(n_5212),
.A2(n_5208),
.A3(n_5196),
.B(n_5223),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_5195),
.Y(n_5292)
);

NOR3xp33_ASAP7_75t_L g5293 ( 
.A(n_5234),
.B(n_942),
.C(n_933),
.Y(n_5293)
);

AOI21xp33_ASAP7_75t_SL g5294 ( 
.A1(n_5209),
.A2(n_935),
.B(n_934),
.Y(n_5294)
);

INVx1_ASAP7_75t_SL g5295 ( 
.A(n_5205),
.Y(n_5295)
);

AOI221xp5_ASAP7_75t_L g5296 ( 
.A1(n_5184),
.A2(n_937),
.B1(n_933),
.B2(n_934),
.C(n_938),
.Y(n_5296)
);

AOI222xp33_ASAP7_75t_L g5297 ( 
.A1(n_5231),
.A2(n_940),
.B1(n_942),
.B2(n_937),
.C1(n_939),
.C2(n_941),
.Y(n_5297)
);

NOR3xp33_ASAP7_75t_SL g5298 ( 
.A(n_5226),
.B(n_940),
.C(n_941),
.Y(n_5298)
);

NAND4xp25_ASAP7_75t_L g5299 ( 
.A(n_5181),
.B(n_945),
.C(n_943),
.D(n_944),
.Y(n_5299)
);

AOI321xp33_ASAP7_75t_L g5300 ( 
.A1(n_5187),
.A2(n_946),
.A3(n_948),
.B1(n_943),
.B2(n_945),
.C(n_947),
.Y(n_5300)
);

OAI222xp33_ASAP7_75t_L g5301 ( 
.A1(n_5216),
.A2(n_949),
.B1(n_951),
.B2(n_947),
.C1(n_948),
.C2(n_950),
.Y(n_5301)
);

INVx1_ASAP7_75t_L g5302 ( 
.A(n_5235),
.Y(n_5302)
);

OAI211xp5_ASAP7_75t_L g5303 ( 
.A1(n_5225),
.A2(n_951),
.B(n_949),
.C(n_950),
.Y(n_5303)
);

AOI221xp5_ASAP7_75t_L g5304 ( 
.A1(n_5188),
.A2(n_5179),
.B1(n_5254),
.B2(n_5192),
.C(n_5247),
.Y(n_5304)
);

NAND2xp5_ASAP7_75t_L g5305 ( 
.A(n_5245),
.B(n_952),
.Y(n_5305)
);

AOI221xp5_ASAP7_75t_L g5306 ( 
.A1(n_5237),
.A2(n_954),
.B1(n_952),
.B2(n_953),
.C(n_955),
.Y(n_5306)
);

OAI221xp5_ASAP7_75t_L g5307 ( 
.A1(n_5198),
.A2(n_956),
.B1(n_954),
.B2(n_955),
.C(n_957),
.Y(n_5307)
);

AOI211xp5_ASAP7_75t_SL g5308 ( 
.A1(n_5230),
.A2(n_959),
.B(n_956),
.C(n_958),
.Y(n_5308)
);

AOI22xp5_ASAP7_75t_L g5309 ( 
.A1(n_5219),
.A2(n_961),
.B1(n_958),
.B2(n_960),
.Y(n_5309)
);

O2A1O1Ixp33_ASAP7_75t_L g5310 ( 
.A1(n_5233),
.A2(n_963),
.B(n_961),
.C(n_962),
.Y(n_5310)
);

AOI222xp33_ASAP7_75t_L g5311 ( 
.A1(n_5204),
.A2(n_964),
.B1(n_966),
.B2(n_962),
.C1(n_963),
.C2(n_965),
.Y(n_5311)
);

OAI221xp5_ASAP7_75t_SL g5312 ( 
.A1(n_5276),
.A2(n_5211),
.B1(n_5228),
.B2(n_5207),
.C(n_5182),
.Y(n_5312)
);

XOR2xp5_ASAP7_75t_L g5313 ( 
.A(n_5284),
.B(n_5232),
.Y(n_5313)
);

AOI22xp33_ASAP7_75t_L g5314 ( 
.A1(n_5263),
.A2(n_5193),
.B1(n_5214),
.B2(n_5206),
.Y(n_5314)
);

INVx1_ASAP7_75t_L g5315 ( 
.A(n_5259),
.Y(n_5315)
);

AOI21xp5_ASAP7_75t_L g5316 ( 
.A1(n_5280),
.A2(n_5241),
.B(n_5238),
.Y(n_5316)
);

INVx1_ASAP7_75t_L g5317 ( 
.A(n_5270),
.Y(n_5317)
);

NOR2x1_ASAP7_75t_L g5318 ( 
.A(n_5260),
.B(n_5250),
.Y(n_5318)
);

INVx1_ASAP7_75t_L g5319 ( 
.A(n_5273),
.Y(n_5319)
);

OR2x2_ASAP7_75t_L g5320 ( 
.A(n_5299),
.B(n_5246),
.Y(n_5320)
);

NOR2x1p5_ASAP7_75t_L g5321 ( 
.A(n_5305),
.B(n_964),
.Y(n_5321)
);

OAI22xp5_ASAP7_75t_L g5322 ( 
.A1(n_5258),
.A2(n_969),
.B1(n_965),
.B2(n_967),
.Y(n_5322)
);

AOI222xp33_ASAP7_75t_L g5323 ( 
.A1(n_5265),
.A2(n_5304),
.B1(n_5302),
.B2(n_5295),
.C1(n_5287),
.C2(n_5271),
.Y(n_5323)
);

NOR3xp33_ASAP7_75t_L g5324 ( 
.A(n_5269),
.B(n_967),
.C(n_969),
.Y(n_5324)
);

INVx1_ASAP7_75t_SL g5325 ( 
.A(n_5287),
.Y(n_5325)
);

NAND2xp5_ASAP7_75t_SL g5326 ( 
.A(n_5287),
.B(n_970),
.Y(n_5326)
);

NAND2x1p5_ASAP7_75t_L g5327 ( 
.A(n_5292),
.B(n_5309),
.Y(n_5327)
);

OAI32xp33_ASAP7_75t_L g5328 ( 
.A1(n_5277),
.A2(n_972),
.A3(n_970),
.B1(n_971),
.B2(n_973),
.Y(n_5328)
);

INVxp67_ASAP7_75t_L g5329 ( 
.A(n_5262),
.Y(n_5329)
);

NOR4xp75_ASAP7_75t_L g5330 ( 
.A(n_5266),
.B(n_974),
.C(n_972),
.D(n_973),
.Y(n_5330)
);

AND2x4_ASAP7_75t_L g5331 ( 
.A(n_5293),
.B(n_975),
.Y(n_5331)
);

AOI21xp5_ASAP7_75t_L g5332 ( 
.A1(n_5261),
.A2(n_975),
.B(n_977),
.Y(n_5332)
);

AOI221xp5_ASAP7_75t_L g5333 ( 
.A1(n_5294),
.A2(n_979),
.B1(n_977),
.B2(n_978),
.C(n_980),
.Y(n_5333)
);

OAI211xp5_ASAP7_75t_L g5334 ( 
.A1(n_5285),
.A2(n_980),
.B(n_978),
.C(n_979),
.Y(n_5334)
);

NOR3xp33_ASAP7_75t_L g5335 ( 
.A(n_5267),
.B(n_981),
.C(n_982),
.Y(n_5335)
);

O2A1O1Ixp33_ASAP7_75t_L g5336 ( 
.A1(n_5281),
.A2(n_985),
.B(n_983),
.C(n_984),
.Y(n_5336)
);

AOI22xp5_ASAP7_75t_L g5337 ( 
.A1(n_5272),
.A2(n_985),
.B1(n_983),
.B2(n_984),
.Y(n_5337)
);

INVx2_ASAP7_75t_SL g5338 ( 
.A(n_5290),
.Y(n_5338)
);

OAI21xp5_ASAP7_75t_L g5339 ( 
.A1(n_5310),
.A2(n_986),
.B(n_988),
.Y(n_5339)
);

AND2x2_ASAP7_75t_L g5340 ( 
.A(n_5298),
.B(n_986),
.Y(n_5340)
);

NAND3xp33_ASAP7_75t_L g5341 ( 
.A(n_5274),
.B(n_989),
.C(n_990),
.Y(n_5341)
);

INVx1_ASAP7_75t_SL g5342 ( 
.A(n_5275),
.Y(n_5342)
);

NAND2xp33_ASAP7_75t_L g5343 ( 
.A(n_5278),
.B(n_990),
.Y(n_5343)
);

AND2x4_ASAP7_75t_L g5344 ( 
.A(n_5308),
.B(n_991),
.Y(n_5344)
);

NAND2xp5_ASAP7_75t_L g5345 ( 
.A(n_5283),
.B(n_991),
.Y(n_5345)
);

NAND2xp5_ASAP7_75t_SL g5346 ( 
.A(n_5300),
.B(n_992),
.Y(n_5346)
);

NAND2xp5_ASAP7_75t_L g5347 ( 
.A(n_5344),
.B(n_5289),
.Y(n_5347)
);

INVx1_ASAP7_75t_L g5348 ( 
.A(n_5340),
.Y(n_5348)
);

INVx1_ASAP7_75t_L g5349 ( 
.A(n_5344),
.Y(n_5349)
);

AOI221xp5_ASAP7_75t_L g5350 ( 
.A1(n_5328),
.A2(n_5291),
.B1(n_5268),
.B2(n_5282),
.C(n_5264),
.Y(n_5350)
);

INVx2_ASAP7_75t_SL g5351 ( 
.A(n_5315),
.Y(n_5351)
);

NOR3xp33_ASAP7_75t_L g5352 ( 
.A(n_5329),
.B(n_5307),
.C(n_5288),
.Y(n_5352)
);

AOI22xp5_ASAP7_75t_L g5353 ( 
.A1(n_5317),
.A2(n_5303),
.B1(n_5296),
.B2(n_5311),
.Y(n_5353)
);

NOR3xp33_ASAP7_75t_L g5354 ( 
.A(n_5325),
.B(n_5301),
.C(n_5257),
.Y(n_5354)
);

INVx1_ASAP7_75t_L g5355 ( 
.A(n_5345),
.Y(n_5355)
);

AOI21xp5_ASAP7_75t_SL g5356 ( 
.A1(n_5336),
.A2(n_5256),
.B(n_5306),
.Y(n_5356)
);

AOI21xp33_ASAP7_75t_SL g5357 ( 
.A1(n_5324),
.A2(n_5297),
.B(n_5279),
.Y(n_5357)
);

NOR2xp33_ASAP7_75t_L g5358 ( 
.A(n_5334),
.B(n_5286),
.Y(n_5358)
);

NOR3xp33_ASAP7_75t_SL g5359 ( 
.A(n_5316),
.B(n_992),
.C(n_993),
.Y(n_5359)
);

CKINVDCx5p33_ASAP7_75t_R g5360 ( 
.A(n_5319),
.Y(n_5360)
);

AOI211xp5_ASAP7_75t_SL g5361 ( 
.A1(n_5312),
.A2(n_5343),
.B(n_5332),
.C(n_5335),
.Y(n_5361)
);

OAI31xp33_ASAP7_75t_L g5362 ( 
.A1(n_5341),
.A2(n_996),
.A3(n_994),
.B(n_995),
.Y(n_5362)
);

NOR2x1p5_ASAP7_75t_L g5363 ( 
.A(n_5320),
.B(n_5331),
.Y(n_5363)
);

NAND2xp5_ASAP7_75t_SL g5364 ( 
.A(n_5350),
.B(n_5333),
.Y(n_5364)
);

INVx1_ASAP7_75t_L g5365 ( 
.A(n_5347),
.Y(n_5365)
);

AOI22xp33_ASAP7_75t_L g5366 ( 
.A1(n_5354),
.A2(n_5352),
.B1(n_5349),
.B2(n_5318),
.Y(n_5366)
);

AOI22xp33_ASAP7_75t_SL g5367 ( 
.A1(n_5351),
.A2(n_5342),
.B1(n_5338),
.B2(n_5339),
.Y(n_5367)
);

NOR2xp33_ASAP7_75t_L g5368 ( 
.A(n_5357),
.B(n_5346),
.Y(n_5368)
);

AO22x2_ASAP7_75t_L g5369 ( 
.A1(n_5348),
.A2(n_5322),
.B1(n_5326),
.B2(n_5313),
.Y(n_5369)
);

NAND3xp33_ASAP7_75t_SL g5370 ( 
.A(n_5362),
.B(n_5330),
.C(n_5323),
.Y(n_5370)
);

INVx1_ASAP7_75t_L g5371 ( 
.A(n_5359),
.Y(n_5371)
);

OAI211xp5_ASAP7_75t_L g5372 ( 
.A1(n_5353),
.A2(n_5337),
.B(n_5361),
.C(n_5356),
.Y(n_5372)
);

NOR2x1_ASAP7_75t_L g5373 ( 
.A(n_5363),
.B(n_5321),
.Y(n_5373)
);

AOI211x1_ASAP7_75t_L g5374 ( 
.A1(n_5355),
.A2(n_5314),
.B(n_5327),
.C(n_997),
.Y(n_5374)
);

XOR2xp5_ASAP7_75t_L g5375 ( 
.A(n_5366),
.B(n_5360),
.Y(n_5375)
);

OAI22xp5_ASAP7_75t_L g5376 ( 
.A1(n_5367),
.A2(n_5358),
.B1(n_998),
.B2(n_995),
.Y(n_5376)
);

INVx2_ASAP7_75t_L g5377 ( 
.A(n_5369),
.Y(n_5377)
);

NOR2x2_ASAP7_75t_L g5378 ( 
.A(n_5370),
.B(n_5374),
.Y(n_5378)
);

INVx1_ASAP7_75t_L g5379 ( 
.A(n_5373),
.Y(n_5379)
);

INVx1_ASAP7_75t_L g5380 ( 
.A(n_5371),
.Y(n_5380)
);

INVx2_ASAP7_75t_L g5381 ( 
.A(n_5365),
.Y(n_5381)
);

INVx1_ASAP7_75t_L g5382 ( 
.A(n_5376),
.Y(n_5382)
);

AOI22xp33_ASAP7_75t_L g5383 ( 
.A1(n_5377),
.A2(n_5368),
.B1(n_5364),
.B2(n_5372),
.Y(n_5383)
);

INVx1_ASAP7_75t_L g5384 ( 
.A(n_5375),
.Y(n_5384)
);

AOI22xp5_ASAP7_75t_L g5385 ( 
.A1(n_5379),
.A2(n_1000),
.B1(n_996),
.B2(n_999),
.Y(n_5385)
);

INVx3_ASAP7_75t_L g5386 ( 
.A(n_5381),
.Y(n_5386)
);

AOI22xp5_ASAP7_75t_L g5387 ( 
.A1(n_5386),
.A2(n_5380),
.B1(n_5378),
.B2(n_1001),
.Y(n_5387)
);

OAI22xp5_ASAP7_75t_L g5388 ( 
.A1(n_5383),
.A2(n_1001),
.B1(n_999),
.B2(n_1000),
.Y(n_5388)
);

AOI22xp33_ASAP7_75t_SL g5389 ( 
.A1(n_5388),
.A2(n_5384),
.B1(n_5382),
.B2(n_5385),
.Y(n_5389)
);

AOI22xp33_ASAP7_75t_L g5390 ( 
.A1(n_5389),
.A2(n_5387),
.B1(n_1004),
.B2(n_1002),
.Y(n_5390)
);

OAI21x1_ASAP7_75t_SL g5391 ( 
.A1(n_5390),
.A2(n_1002),
.B(n_1003),
.Y(n_5391)
);

OAI21xp5_ASAP7_75t_SL g5392 ( 
.A1(n_5391),
.A2(n_1003),
.B(n_1004),
.Y(n_5392)
);

NAND3xp33_ASAP7_75t_L g5393 ( 
.A(n_5392),
.B(n_1005),
.C(n_1006),
.Y(n_5393)
);

HB1xp67_ASAP7_75t_L g5394 ( 
.A(n_5393),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_5393),
.Y(n_5395)
);

OR2x6_ASAP7_75t_L g5396 ( 
.A(n_5395),
.B(n_1005),
.Y(n_5396)
);

OA21x2_ASAP7_75t_L g5397 ( 
.A1(n_5394),
.A2(n_1006),
.B(n_1007),
.Y(n_5397)
);

AOI21xp5_ASAP7_75t_L g5398 ( 
.A1(n_5396),
.A2(n_1008),
.B(n_1009),
.Y(n_5398)
);

AOI211xp5_ASAP7_75t_L g5399 ( 
.A1(n_5398),
.A2(n_5397),
.B(n_1010),
.C(n_1008),
.Y(n_5399)
);


endmodule