module fake_jpeg_15885_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_R g33 ( 
.A(n_23),
.B(n_32),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_24),
.Y(n_44)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_16),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_31),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_44),
.A2(n_64),
.B(n_38),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_29),
.C(n_18),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_41),
.C(n_38),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_30),
.B1(n_21),
.B2(n_28),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_51),
.B1(n_21),
.B2(n_25),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_30),
.B1(n_21),
.B2(n_31),
.Y(n_51)
);

HAxp5_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_29),
.CON(n_52),
.SN(n_52)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_58),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_59),
.Y(n_81)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_64),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_66),
.B(n_77),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_17),
.B1(n_26),
.B2(n_22),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_82),
.C(n_53),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_74),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_40),
.B1(n_39),
.B2(n_36),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_71),
.A2(n_41),
.B1(n_54),
.B2(n_34),
.Y(n_100)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_42),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_42),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_83),
.Y(n_107)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_40),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_80),
.A2(n_78),
.B(n_86),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_40),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_39),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_0),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_90),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

AOI32xp33_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_34),
.A3(n_59),
.B1(n_36),
.B2(n_47),
.Y(n_91)
);

OAI32xp33_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_53),
.A3(n_37),
.B1(n_34),
.B2(n_43),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_80),
.B1(n_84),
.B2(n_66),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_92),
.A2(n_97),
.B1(n_100),
.B2(n_82),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_61),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_82),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_38),
.B1(n_57),
.B2(n_46),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_119),
.B1(n_65),
.B2(n_85),
.Y(n_122)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_89),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_96),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_115),
.C(n_116),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_106),
.B1(n_76),
.B2(n_65),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_17),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_109),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_41),
.B1(n_58),
.B2(n_37),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_26),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_88),
.B(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_24),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_0),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_43),
.C(n_49),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_22),
.Y(n_118)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_79),
.A2(n_37),
.B1(n_54),
.B2(n_58),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_120),
.B(n_128),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_133),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_127),
.B1(n_132),
.B2(n_138),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_140),
.B1(n_114),
.B2(n_102),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_124),
.Y(n_159)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_126),
.A2(n_134),
.B1(n_136),
.B2(n_142),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_130),
.B(n_143),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_92),
.A2(n_90),
.B1(n_72),
.B2(n_69),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_69),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_73),
.B(n_75),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_0),
.Y(n_135)
);

XNOR2x1_ASAP7_75t_SL g170 ( 
.A(n_135),
.B(n_24),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_75),
.B(n_49),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_99),
.A2(n_37),
.B1(n_55),
.B2(n_14),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_97),
.A2(n_55),
.B1(n_87),
.B2(n_19),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_75),
.B(n_18),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_19),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_106),
.A2(n_87),
.B1(n_19),
.B2(n_29),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_113),
.B1(n_24),
.B2(n_29),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_95),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_149),
.C(n_160),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_145),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_148),
.B(n_162),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_133),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_95),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_152),
.B(n_156),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_169),
.B1(n_171),
.B2(n_137),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_112),
.A3(n_102),
.B1(n_114),
.B2(n_118),
.C1(n_104),
.C2(n_101),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g194 ( 
.A1(n_155),
.A2(n_170),
.B(n_18),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_93),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_121),
.B(n_93),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_164),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_100),
.C(n_98),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_129),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_119),
.C(n_111),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_108),
.B1(n_117),
.B2(n_96),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_165),
.A2(n_137),
.B1(n_144),
.B2(n_129),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_125),
.B(n_109),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_27),
.Y(n_193)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_96),
.B1(n_111),
.B2(n_29),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_123),
.B1(n_135),
.B2(n_141),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_172),
.A2(n_179),
.B1(n_182),
.B2(n_188),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_175),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_154),
.A2(n_139),
.B(n_125),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_174),
.A2(n_1),
.B(n_2),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_128),
.Y(n_176)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_138),
.Y(n_177)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_122),
.B1(n_126),
.B2(n_120),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_162),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_190),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_159),
.B1(n_156),
.B2(n_157),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_153),
.A2(n_145),
.B1(n_129),
.B2(n_113),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_165),
.A2(n_124),
.B1(n_18),
.B2(n_110),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_168),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_159),
.Y(n_191)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_196),
.Y(n_212)
);

XNOR2x2_ASAP7_75t_SL g216 ( 
.A(n_194),
.B(n_7),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_151),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_152),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_7),
.Y(n_218)
);

OAI22x1_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_170),
.B1(n_161),
.B2(n_171),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_201),
.A2(n_209),
.B1(n_186),
.B2(n_194),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_149),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_217),
.Y(n_228)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_146),
.C(n_163),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_208),
.C(n_185),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_195),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_210),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_110),
.C(n_27),
.Y(n_208)
);

XOR2x2_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_27),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_192),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_189),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_197),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_218),
.B(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_184),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_174),
.Y(n_223)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_223),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_179),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_224),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_232),
.C(n_234),
.Y(n_246)
);

AND2x4_ASAP7_75t_SL g226 ( 
.A(n_201),
.B(n_175),
.Y(n_226)
);

INVx13_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_202),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_240),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_177),
.B1(n_188),
.B2(n_172),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_231),
.A2(n_206),
.B1(n_204),
.B2(n_214),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_176),
.C(n_183),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_184),
.C(n_181),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_215),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_238),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_7),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_216),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_14),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_1),
.C(n_2),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_219),
.C(n_220),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_230),
.A2(n_200),
.B(n_220),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_243),
.A2(n_8),
.B(n_14),
.Y(n_271)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_224),
.A2(n_214),
.B1(n_199),
.B2(n_198),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_259),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_232),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_254),
.C(n_255),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_212),
.Y(n_251)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_198),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_226),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_239),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_238),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_242),
.Y(n_261)
);

BUFx12_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_1),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_274),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_222),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_257),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_227),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_267),
.Y(n_279)
);

OA21x2_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_199),
.B(n_233),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_260),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_258),
.A2(n_211),
.B1(n_2),
.B2(n_3),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_270),
.B(n_272),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_271),
.A2(n_256),
.B(n_11),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_15),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_3),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_260),
.A2(n_8),
.B(n_12),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_277),
.B(n_278),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_275),
.A2(n_253),
.B1(n_246),
.B2(n_248),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_281),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_286),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_288),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_266),
.B(n_246),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_285),
.B(n_284),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_255),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_287),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_273),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_269),
.C(n_261),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_296),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_249),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_291),
.B(n_289),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_283),
.A2(n_268),
.B1(n_253),
.B2(n_274),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_279),
.B(n_264),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g299 ( 
.A(n_284),
.B(n_248),
.CI(n_263),
.CON(n_299),
.SN(n_299)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_303),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_290),
.B(n_276),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_268),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_307),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_305),
.A2(n_294),
.B(n_299),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_297),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_301),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_311),
.C(n_312),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_15),
.B1(n_4),
.B2(n_5),
.Y(n_313)
);

AOI321xp33_ASAP7_75t_SL g314 ( 
.A1(n_313),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_310),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_315),
.Y(n_317)
);

AOI321xp33_ASAP7_75t_L g315 ( 
.A1(n_308),
.A2(n_3),
.A3(n_4),
.B1(n_6),
.B2(n_311),
.C(n_312),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_316),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_318),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_4),
.Y(n_320)
);


endmodule