module fake_jpeg_16572_n_249 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_12),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_11),
.B(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_1),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_41),
.Y(n_53)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_17),
.Y(n_39)
);

HAxp5_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_17),
.CON(n_61),
.SN(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_28),
.B(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_25),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_48),
.Y(n_75)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_35),
.Y(n_78)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_26),
.B1(n_31),
.B2(n_20),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_50),
.A2(n_51),
.B1(n_63),
.B2(n_39),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_26),
.B1(n_31),
.B2(n_20),
.Y(n_51)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_26),
.B1(n_20),
.B2(n_31),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_35),
.B1(n_15),
.B2(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_18),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_33),
.A2(n_23),
.B(n_30),
.C(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_23),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

AND2x4_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_39),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_23),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_22),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_35),
.A2(n_26),
.B1(n_42),
.B2(n_24),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_53),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_69),
.A2(n_72),
.B1(n_43),
.B2(n_46),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_50),
.B1(n_64),
.B2(n_60),
.Y(n_98)
);

NOR3xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_41),
.C(n_36),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_81),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_76),
.B(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_44),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_49),
.Y(n_94)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_32),
.C(n_17),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_17),
.C(n_51),
.Y(n_93)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_90),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_48),
.B1(n_54),
.B2(n_52),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_89),
.A2(n_98),
.B1(n_71),
.B2(n_43),
.Y(n_122)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_80),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_100),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_58),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_103),
.C(n_69),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_58),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_64),
.B1(n_47),
.B2(n_46),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_84),
.B1(n_43),
.B2(n_67),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_63),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_105),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_68),
.B1(n_85),
.B2(n_76),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_55),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_55),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_69),
.B1(n_68),
.B2(n_70),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_117),
.B1(n_121),
.B2(n_122),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_113),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_69),
.C(n_79),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_115),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_68),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_27),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_131),
.Y(n_145)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_104),
.B(n_27),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_88),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_97),
.Y(n_138)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_32),
.B1(n_55),
.B2(n_24),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_128),
.A2(n_86),
.B1(n_90),
.B2(n_21),
.Y(n_134)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_92),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_87),
.B(n_92),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_143),
.B(n_153),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_147),
.B1(n_129),
.B2(n_19),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_113),
.A2(n_93),
.B1(n_95),
.B2(n_103),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_137),
.A2(n_148),
.B1(n_119),
.B2(n_112),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_116),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_140),
.B(n_141),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_124),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_88),
.B(n_22),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_144),
.B(n_118),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_105),
.B1(n_30),
.B2(n_22),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_130),
.A2(n_30),
.B1(n_21),
.B2(n_19),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_17),
.Y(n_152)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_115),
.A2(n_111),
.B(n_119),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_147),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_118),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_153),
.C(n_137),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_142),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_161),
.Y(n_180)
);

NAND2xp33_ASAP7_75t_SL g160 ( 
.A(n_136),
.B(n_109),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_160),
.A2(n_174),
.B1(n_25),
.B2(n_18),
.Y(n_192)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_135),
.A2(n_109),
.B1(n_122),
.B2(n_121),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_165),
.A2(n_169),
.B1(n_172),
.B2(n_139),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_128),
.C(n_32),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_170),
.Y(n_189)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_168),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_140),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_171),
.B(n_173),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_135),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_19),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_146),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_177),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_132),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_165),
.A2(n_149),
.B1(n_141),
.B2(n_150),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_184),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_152),
.C(n_143),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_148),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_185),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_160),
.A2(n_164),
.B1(n_163),
.B2(n_172),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_134),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_192),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_164),
.A2(n_144),
.B1(n_14),
.B2(n_6),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_156),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_191),
.Y(n_195)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_194),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_163),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_203),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_186),
.A2(n_166),
.B1(n_187),
.B2(n_185),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_201),
.A2(n_176),
.B1(n_177),
.B2(n_25),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_SL g202 ( 
.A(n_180),
.B(n_155),
.C(n_158),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_202),
.A2(n_5),
.B(n_7),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_158),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_182),
.B(n_3),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_206),
.Y(n_219)
);

BUFx12_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_206),
.Y(n_223)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_18),
.C(n_7),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_211),
.C(n_216),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_5),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_206),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_204),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_200),
.B1(n_204),
.B2(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_198),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_7),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_8),
.C(n_9),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_218),
.B(n_201),
.Y(n_220)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_220),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_222),
.B(n_217),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_223),
.B(n_227),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_214),
.B(n_8),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_228),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_9),
.Y(n_228)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_230),
.Y(n_238)
);

NOR2xp67_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_210),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_232),
.A2(n_213),
.B(n_225),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_219),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_233),
.B(n_235),
.Y(n_239)
);

NOR2x1_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_212),
.Y(n_235)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_236),
.Y(n_244)
);

AOI21xp33_ASAP7_75t_L g237 ( 
.A1(n_231),
.A2(n_225),
.B(n_216),
.Y(n_237)
);

O2A1O1Ixp33_ASAP7_75t_SL g242 ( 
.A1(n_237),
.A2(n_240),
.B(n_10),
.C(n_13),
.Y(n_242)
);

AOI21xp33_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_10),
.B(n_12),
.Y(n_240)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_238),
.B(n_230),
.CI(n_229),
.CON(n_241),
.SN(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_242),
.A2(n_243),
.B(n_10),
.Y(n_245)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_239),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_245),
.B(n_243),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_246),
.B1(n_244),
.B2(n_13),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_13),
.Y(n_249)
);


endmodule