module real_aes_18120_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_1102;
wire n_661;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1457;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_578;
wire n_372;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_0), .A2(n_1), .B1(n_1177), .B2(n_1180), .Y(n_1190) );
INVx1_ASAP7_75t_L g409 ( .A(n_2), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g840 ( .A1(n_3), .A2(n_256), .B1(n_738), .B2(n_841), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_3), .A2(n_174), .B1(n_681), .B2(n_852), .Y(n_851) );
OAI211xp5_ASAP7_75t_L g758 ( .A1(n_4), .A2(n_423), .B(n_600), .C(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g769 ( .A(n_4), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_5), .A2(n_263), .B1(n_844), .B2(n_1104), .Y(n_1103) );
INVxp33_ASAP7_75t_SL g1136 ( .A(n_5), .Y(n_1136) );
INVx1_ASAP7_75t_L g648 ( .A(n_6), .Y(n_648) );
AOI22xp33_ASAP7_75t_SL g832 ( .A1(n_7), .A2(n_238), .B1(n_738), .B2(n_833), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_7), .A2(n_216), .B1(n_675), .B2(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g341 ( .A(n_8), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_8), .B(n_303), .Y(n_407) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_8), .B(n_224), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_8), .B(n_324), .Y(n_1406) );
OAI22xp33_ASAP7_75t_L g573 ( .A1(n_9), .A2(n_203), .B1(n_332), .B2(n_574), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_9), .A2(n_203), .B1(n_385), .B2(n_512), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g1411 ( .A1(n_10), .A2(n_77), .B1(n_738), .B2(n_1076), .Y(n_1411) );
AOI22xp33_ASAP7_75t_L g1457 ( .A1(n_10), .A2(n_128), .B1(n_854), .B2(n_1458), .Y(n_1457) );
INVx1_ASAP7_75t_L g774 ( .A(n_11), .Y(n_774) );
INVx1_ASAP7_75t_L g707 ( .A(n_12), .Y(n_707) );
INVx2_ASAP7_75t_L g1173 ( .A(n_13), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_13), .B(n_102), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_13), .B(n_1179), .Y(n_1181) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_14), .A2(n_123), .B1(n_511), .B2(n_512), .Y(n_510) );
OAI22xp33_ASAP7_75t_L g527 ( .A1(n_14), .A2(n_123), .B1(n_332), .B2(n_528), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g1206 ( .A1(n_15), .A2(n_231), .B1(n_1177), .B2(n_1180), .Y(n_1206) );
INVx1_ASAP7_75t_L g645 ( .A(n_16), .Y(n_645) );
OAI22xp33_ASAP7_75t_L g982 ( .A1(n_17), .A2(n_150), .B1(n_334), .B2(n_608), .Y(n_982) );
OAI22xp33_ASAP7_75t_L g984 ( .A1(n_17), .A2(n_271), .B1(n_387), .B2(n_709), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_18), .A2(n_204), .B1(n_1078), .B2(n_1082), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_18), .A2(n_235), .B1(n_702), .B2(n_854), .Y(n_1090) );
CKINVDCx5p33_ASAP7_75t_R g963 ( .A(n_19), .Y(n_963) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_20), .A2(n_134), .B1(n_574), .B2(n_611), .Y(n_610) );
OAI22xp33_ASAP7_75t_SL g613 ( .A1(n_20), .A2(n_134), .B1(n_387), .B2(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g431 ( .A(n_21), .Y(n_431) );
OAI22xp33_ASAP7_75t_L g946 ( .A1(n_22), .A2(n_197), .B1(n_326), .B2(n_611), .Y(n_946) );
OAI22xp33_ASAP7_75t_L g949 ( .A1(n_22), .A2(n_98), .B1(n_387), .B2(n_709), .Y(n_949) );
AOI22xp5_ASAP7_75t_L g1195 ( .A1(n_23), .A2(n_268), .B1(n_1170), .B2(n_1196), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_24), .A2(n_108), .B1(n_767), .B2(n_1111), .Y(n_1110) );
INVx1_ASAP7_75t_L g1143 ( .A(n_24), .Y(n_1143) );
INVx1_ASAP7_75t_L g430 ( .A(n_25), .Y(n_430) );
INVx1_ASAP7_75t_L g862 ( .A(n_26), .Y(n_862) );
INVx1_ASAP7_75t_L g945 ( .A(n_27), .Y(n_945) );
OAI211xp5_ASAP7_75t_L g950 ( .A1(n_27), .A2(n_570), .B(n_616), .C(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g1008 ( .A(n_28), .Y(n_1008) );
INVx1_ASAP7_75t_L g1494 ( .A(n_29), .Y(n_1494) );
INVx1_ASAP7_75t_L g479 ( .A(n_30), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g968 ( .A(n_31), .Y(n_968) );
CKINVDCx5p33_ASAP7_75t_R g960 ( .A(n_32), .Y(n_960) );
OAI22xp33_ASAP7_75t_L g757 ( .A1(n_33), .A2(n_119), .B1(n_608), .B2(n_609), .Y(n_757) );
OAI22xp33_ASAP7_75t_L g770 ( .A1(n_33), .A2(n_47), .B1(n_359), .B2(n_709), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g1199 ( .A1(n_34), .A2(n_247), .B1(n_1177), .B2(n_1180), .Y(n_1199) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_35), .A2(n_168), .B1(n_359), .B2(n_709), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_35), .A2(n_36), .B1(n_608), .B2(n_609), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_36), .A2(n_278), .B1(n_349), .B2(n_387), .Y(n_698) );
AO22x1_ASAP7_75t_L g1203 ( .A1(n_37), .A2(n_61), .B1(n_1170), .B2(n_1185), .Y(n_1203) );
INVx1_ASAP7_75t_L g1486 ( .A(n_38), .Y(n_1486) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_39), .A2(n_139), .B1(n_868), .B2(n_869), .Y(n_867) );
INVxp67_ASAP7_75t_SL g880 ( .A(n_39), .Y(n_880) );
INVx1_ASAP7_75t_L g812 ( .A(n_40), .Y(n_812) );
INVx1_ASAP7_75t_L g606 ( .A(n_41), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_42), .A2(n_76), .B1(n_1078), .B2(n_1080), .Y(n_1077) );
AOI22xp33_ASAP7_75t_SL g1091 ( .A1(n_42), .A2(n_89), .B1(n_901), .B2(n_928), .Y(n_1091) );
INVx1_ASAP7_75t_L g356 ( .A(n_43), .Y(n_356) );
INVx1_ASAP7_75t_L g362 ( .A(n_43), .Y(n_362) );
AOI221xp5_ASAP7_75t_L g1408 ( .A1(n_44), .A2(n_122), .B1(n_878), .B2(n_890), .C(n_1409), .Y(n_1408) );
AOI22xp33_ASAP7_75t_SL g1459 ( .A1(n_44), .A2(n_195), .B1(n_637), .B2(n_901), .Y(n_1459) );
INVx1_ASAP7_75t_L g1512 ( .A(n_45), .Y(n_1512) );
OAI211xp5_ASAP7_75t_L g1518 ( .A1(n_45), .A2(n_616), .B(n_1519), .C(n_1520), .Y(n_1518) );
INVx1_ASAP7_75t_L g1063 ( .A(n_46), .Y(n_1063) );
OAI221xp5_ASAP7_75t_L g1070 ( .A1(n_46), .A2(n_101), .B1(n_452), .B2(n_869), .C(n_1071), .Y(n_1070) );
OAI22xp33_ASAP7_75t_L g762 ( .A1(n_47), .A2(n_201), .B1(n_574), .B2(n_611), .Y(n_762) );
INVx1_ASAP7_75t_L g556 ( .A(n_48), .Y(n_556) );
XOR2x2_ASAP7_75t_L g858 ( .A(n_49), .B(n_859), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_50), .A2(n_74), .B1(n_738), .B2(n_893), .Y(n_892) );
AOI22xp33_ASAP7_75t_SL g907 ( .A1(n_50), .A2(n_246), .B1(n_623), .B2(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g549 ( .A(n_51), .Y(n_549) );
INVx1_ASAP7_75t_L g1036 ( .A(n_52), .Y(n_1036) );
OAI22xp33_ASAP7_75t_L g1047 ( .A1(n_52), .A2(n_152), .B1(n_334), .B2(n_611), .Y(n_1047) );
OAI211xp5_ASAP7_75t_L g941 ( .A1(n_53), .A2(n_600), .B(n_942), .C(n_943), .Y(n_941) );
INVx1_ASAP7_75t_L g952 ( .A(n_53), .Y(n_952) );
INVx1_ASAP7_75t_L g1156 ( .A(n_54), .Y(n_1156) );
OAI22xp33_ASAP7_75t_L g1123 ( .A1(n_55), .A2(n_219), .B1(n_534), .B2(n_1124), .Y(n_1123) );
OAI22xp5_ASAP7_75t_L g1132 ( .A1(n_55), .A2(n_219), .B1(n_523), .B2(n_1133), .Y(n_1132) );
INVx2_ASAP7_75t_L g352 ( .A(n_56), .Y(n_352) );
XNOR2x2_ASAP7_75t_L g539 ( .A(n_57), .B(n_540), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_58), .A2(n_244), .B1(n_675), .B2(n_676), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_58), .A2(n_172), .B1(n_741), .B2(n_743), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_59), .A2(n_223), .B1(n_318), .B2(n_583), .Y(n_582) );
OAI22xp33_ASAP7_75t_L g590 ( .A1(n_59), .A2(n_223), .B1(n_522), .B2(n_591), .Y(n_590) );
INVxp67_ASAP7_75t_SL g865 ( .A(n_60), .Y(n_865) );
OAI22xp33_ASAP7_75t_L g881 ( .A1(n_60), .A2(n_139), .B1(n_579), .B2(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g705 ( .A(n_62), .Y(n_705) );
INVx1_ASAP7_75t_L g761 ( .A(n_63), .Y(n_761) );
INVx1_ASAP7_75t_L g701 ( .A(n_64), .Y(n_701) );
INVx1_ASAP7_75t_L g1005 ( .A(n_65), .Y(n_1005) );
AOI22xp5_ASAP7_75t_L g1200 ( .A1(n_66), .A2(n_170), .B1(n_1170), .B2(n_1185), .Y(n_1200) );
INVx1_ASAP7_75t_L g1108 ( .A(n_67), .Y(n_1108) );
INVx1_ASAP7_75t_L g550 ( .A(n_68), .Y(n_550) );
INVx1_ASAP7_75t_L g779 ( .A(n_69), .Y(n_779) );
AO221x2_ASAP7_75t_L g1242 ( .A1(n_70), .A2(n_213), .B1(n_1177), .B2(n_1180), .C(n_1243), .Y(n_1242) );
OAI22xp33_ASAP7_75t_L g947 ( .A1(n_71), .A2(n_98), .B1(n_319), .B2(n_334), .Y(n_947) );
OAI22xp33_ASAP7_75t_L g953 ( .A1(n_71), .A2(n_197), .B1(n_349), .B2(n_359), .Y(n_953) );
OAI211xp5_ASAP7_75t_L g513 ( .A1(n_72), .A2(n_370), .B(n_514), .C(n_517), .Y(n_513) );
INVx1_ASAP7_75t_L g532 ( .A(n_72), .Y(n_532) );
INVx1_ASAP7_75t_L g635 ( .A(n_73), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_74), .A2(n_86), .B1(n_623), .B2(n_854), .Y(n_902) );
CKINVDCx5p33_ASAP7_75t_R g926 ( .A(n_75), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_76), .A2(n_183), .B1(n_901), .B2(n_1088), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g1463 ( .A1(n_77), .A2(n_275), .B1(n_854), .B2(n_1464), .Y(n_1463) );
INVx1_ASAP7_75t_L g417 ( .A(n_78), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_79), .A2(n_277), .B1(n_455), .B2(n_681), .C(n_685), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_79), .A2(n_127), .B1(n_746), .B2(n_749), .Y(n_745) );
XOR2xp5_ASAP7_75t_L g1478 ( .A(n_80), .B(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g1120 ( .A(n_81), .Y(n_1120) );
INVx1_ASAP7_75t_L g497 ( .A(n_82), .Y(n_497) );
INVx1_ASAP7_75t_L g605 ( .A(n_83), .Y(n_605) );
INVx1_ASAP7_75t_L g820 ( .A(n_84), .Y(n_820) );
OAI221xp5_ASAP7_75t_L g825 ( .A1(n_84), .A2(n_245), .B1(n_633), .B2(n_826), .C(n_827), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_85), .A2(n_149), .B1(n_608), .B2(n_609), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_85), .A2(n_149), .B1(n_349), .B2(n_359), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_86), .A2(n_246), .B1(n_741), .B2(n_891), .Y(n_896) );
XOR2x2_ASAP7_75t_L g594 ( .A(n_87), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g1009 ( .A(n_88), .Y(n_1009) );
AOI22xp33_ASAP7_75t_SL g1083 ( .A1(n_89), .A2(n_183), .B1(n_1084), .B2(n_1085), .Y(n_1083) );
INVx1_ASAP7_75t_L g545 ( .A(n_90), .Y(n_545) );
OAI211xp5_ASAP7_75t_L g575 ( .A1(n_91), .A2(n_292), .B(n_576), .C(n_581), .Y(n_575) );
INVx1_ASAP7_75t_L g589 ( .A(n_91), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g1511 ( .A(n_92), .Y(n_1511) );
INVx1_ASAP7_75t_L g476 ( .A(n_93), .Y(n_476) );
INVx1_ASAP7_75t_L g913 ( .A(n_94), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_95), .A2(n_162), .B1(n_608), .B2(n_609), .Y(n_607) );
OAI22xp33_ASAP7_75t_L g624 ( .A1(n_95), .A2(n_162), .B1(n_349), .B2(n_359), .Y(n_624) );
OAI22xp33_ASAP7_75t_L g1515 ( .A1(n_96), .A2(n_156), .B1(n_334), .B2(n_611), .Y(n_1515) );
OAI22xp5_ASAP7_75t_L g1517 ( .A1(n_96), .A2(n_117), .B1(n_387), .B2(n_522), .Y(n_1517) );
OAI22xp5_ASAP7_75t_L g1066 ( .A1(n_97), .A2(n_206), .B1(n_608), .B2(n_609), .Y(n_1066) );
OAI22xp5_ASAP7_75t_L g1072 ( .A1(n_97), .A2(n_206), .B1(n_349), .B2(n_359), .Y(n_1072) );
HB1xp67_ASAP7_75t_L g1158 ( .A(n_99), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_99), .B(n_1156), .Y(n_1171) );
AOI22xp33_ASAP7_75t_SL g838 ( .A1(n_100), .A2(n_216), .B1(n_835), .B2(n_839), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_100), .A2(n_238), .B1(n_844), .B2(n_846), .Y(n_843) );
INVx1_ASAP7_75t_L g1065 ( .A(n_101), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_102), .B(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1179 ( .A(n_102), .Y(n_1179) );
INVx1_ASAP7_75t_L g1493 ( .A(n_103), .Y(n_1493) );
AOI22xp5_ASAP7_75t_L g1419 ( .A1(n_104), .A2(n_195), .B1(n_1076), .B2(n_1420), .Y(n_1419) );
AOI22xp5_ASAP7_75t_L g1460 ( .A1(n_104), .A2(n_122), .B1(n_901), .B2(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1415 ( .A(n_105), .Y(n_1415) );
INVx1_ASAP7_75t_L g871 ( .A(n_106), .Y(n_871) );
CKINVDCx5p33_ASAP7_75t_R g965 ( .A(n_107), .Y(n_965) );
INVx1_ASAP7_75t_L g1137 ( .A(n_108), .Y(n_1137) );
INVx1_ASAP7_75t_L g1426 ( .A(n_109), .Y(n_1426) );
INVx2_ASAP7_75t_L g397 ( .A(n_110), .Y(n_397) );
INVx1_ASAP7_75t_L g464 ( .A(n_110), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g1390 ( .A(n_110), .B(n_352), .Y(n_1390) );
CKINVDCx5p33_ASAP7_75t_R g919 ( .A(n_111), .Y(n_919) );
INVx1_ASAP7_75t_L g783 ( .A(n_112), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_113), .A2(n_209), .B1(n_1170), .B2(n_1185), .Y(n_1189) );
XOR2xp5_ASAP7_75t_L g470 ( .A(n_114), .B(n_471), .Y(n_470) );
AOI22xp33_ASAP7_75t_SL g897 ( .A1(n_115), .A2(n_261), .B1(n_738), .B2(n_893), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_115), .A2(n_182), .B1(n_900), .B2(n_901), .Y(n_904) );
INVx1_ASAP7_75t_L g632 ( .A(n_116), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g1513 ( .A1(n_117), .A2(n_120), .B1(n_318), .B2(n_1514), .Y(n_1513) );
CKINVDCx5p33_ASAP7_75t_R g924 ( .A(n_118), .Y(n_924) );
OAI22xp5_ASAP7_75t_SL g764 ( .A1(n_119), .A2(n_201), .B1(n_349), .B2(n_387), .Y(n_764) );
OAI22xp5_ASAP7_75t_L g1522 ( .A1(n_120), .A2(n_156), .B1(n_388), .B2(n_1523), .Y(n_1522) );
INVx1_ASAP7_75t_L g787 ( .A(n_121), .Y(n_787) );
INVx1_ASAP7_75t_L g647 ( .A(n_124), .Y(n_647) );
INVx1_ASAP7_75t_L g1011 ( .A(n_125), .Y(n_1011) );
INVx1_ASAP7_75t_L g490 ( .A(n_126), .Y(n_490) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_127), .A2(n_215), .B1(n_455), .B2(n_681), .C(n_689), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g1416 ( .A1(n_128), .A2(n_275), .B1(n_743), .B2(n_1417), .C(n_1418), .Y(n_1416) );
INVx1_ASAP7_75t_L g1423 ( .A(n_129), .Y(n_1423) );
OAI21xp5_ASAP7_75t_L g1428 ( .A1(n_130), .A2(n_1429), .B(n_1433), .Y(n_1428) );
CKINVDCx5p33_ASAP7_75t_R g979 ( .A(n_131), .Y(n_979) );
INVx1_ASAP7_75t_L g1101 ( .A(n_132), .Y(n_1101) );
INVx1_ASAP7_75t_L g1484 ( .A(n_133), .Y(n_1484) );
INVx1_ASAP7_75t_L g784 ( .A(n_135), .Y(n_784) );
AOI31xp33_ASAP7_75t_L g672 ( .A1(n_136), .A2(n_673), .A3(n_697), .B(n_712), .Y(n_672) );
NAND2xp33_ASAP7_75t_SL g730 ( .A(n_136), .B(n_731), .Y(n_730) );
INVxp67_ASAP7_75t_SL g752 ( .A(n_136), .Y(n_752) );
AO22x1_ASAP7_75t_L g1204 ( .A1(n_136), .A2(n_228), .B1(n_1177), .B2(n_1180), .Y(n_1204) );
INVx1_ASAP7_75t_L g1057 ( .A(n_137), .Y(n_1057) );
INVx1_ASAP7_75t_L g1034 ( .A(n_138), .Y(n_1034) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_138), .A2(n_262), .B1(n_318), .B2(n_583), .Y(n_1043) );
BUFx3_ASAP7_75t_L g354 ( .A(n_140), .Y(n_354) );
INVx1_ASAP7_75t_L g1030 ( .A(n_141), .Y(n_1030) );
OA211x2_ASAP7_75t_L g1044 ( .A1(n_141), .A2(n_299), .B(n_423), .C(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_L g777 ( .A(n_142), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g932 ( .A(n_143), .Y(n_932) );
CKINVDCx5p33_ASAP7_75t_R g969 ( .A(n_144), .Y(n_969) );
OAI22xp33_ASAP7_75t_L g1114 ( .A1(n_145), .A2(n_254), .B1(n_332), .B2(n_334), .Y(n_1114) );
OAI22xp33_ASAP7_75t_L g1126 ( .A1(n_145), .A2(n_254), .B1(n_388), .B2(n_1127), .Y(n_1126) );
OAI22xp5_ASAP7_75t_SL g993 ( .A1(n_146), .A2(n_994), .B1(n_1041), .B2(n_1049), .Y(n_993) );
NAND4xp25_ASAP7_75t_L g994 ( .A(n_146), .B(n_995), .C(n_1013), .D(n_1024), .Y(n_994) );
INVx1_ASAP7_75t_L g520 ( .A(n_147), .Y(n_520) );
OAI211xp5_ASAP7_75t_L g529 ( .A1(n_147), .A2(n_292), .B(n_530), .C(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g547 ( .A(n_148), .Y(n_547) );
OAI22xp33_ASAP7_75t_L g988 ( .A1(n_150), .A2(n_276), .B1(n_349), .B2(n_359), .Y(n_988) );
CKINVDCx5p33_ASAP7_75t_R g966 ( .A(n_151), .Y(n_966) );
INVx1_ASAP7_75t_L g1033 ( .A(n_152), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1186 ( .A1(n_153), .A2(n_166), .B1(n_1177), .B2(n_1180), .Y(n_1186) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_154), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g959 ( .A(n_155), .Y(n_959) );
INVx1_ASAP7_75t_L g1109 ( .A(n_157), .Y(n_1109) );
INVx1_ASAP7_75t_L g1496 ( .A(n_158), .Y(n_1496) );
XOR2x2_ASAP7_75t_L g754 ( .A(n_159), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g1122 ( .A(n_160), .Y(n_1122) );
OAI211xp5_ASAP7_75t_L g1128 ( .A1(n_160), .A2(n_370), .B(n_1129), .C(n_1130), .Y(n_1128) );
OAI22xp33_ASAP7_75t_L g331 ( .A1(n_161), .A2(n_191), .B1(n_332), .B2(n_334), .Y(n_331) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_161), .A2(n_191), .B1(n_385), .B2(n_388), .Y(n_384) );
INVx1_ASAP7_75t_L g694 ( .A(n_163), .Y(n_694) );
AOI22xp33_ASAP7_75t_SL g733 ( .A1(n_163), .A2(n_244), .B1(n_734), .B2(n_738), .Y(n_733) );
INVx1_ASAP7_75t_L g554 ( .A(n_164), .Y(n_554) );
OAI211xp5_ASAP7_75t_L g1508 ( .A1(n_165), .A2(n_299), .B(n_1509), .C(n_1510), .Y(n_1508) );
INVx1_ASAP7_75t_L g1521 ( .A(n_165), .Y(n_1521) );
INVx1_ASAP7_75t_L g1385 ( .A(n_167), .Y(n_1385) );
INVxp67_ASAP7_75t_SL g716 ( .A(n_168), .Y(n_716) );
INVx1_ASAP7_75t_L g1498 ( .A(n_169), .Y(n_1498) );
AOI22xp5_ASAP7_75t_L g1207 ( .A1(n_171), .A2(n_249), .B1(n_1170), .B2(n_1185), .Y(n_1207) );
INVx1_ASAP7_75t_L g691 ( .A(n_172), .Y(n_691) );
INVx1_ASAP7_75t_L g1488 ( .A(n_173), .Y(n_1488) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_174), .A2(n_248), .B1(n_835), .B2(n_837), .Y(n_834) );
INVx1_ASAP7_75t_L g1001 ( .A(n_175), .Y(n_1001) );
XNOR2xp5_ASAP7_75t_L g288 ( .A(n_176), .B(n_289), .Y(n_288) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_177), .Y(n_444) );
INVx1_ASAP7_75t_L g863 ( .A(n_178), .Y(n_863) );
INVx1_ASAP7_75t_L g789 ( .A(n_179), .Y(n_789) );
OAI211xp5_ASAP7_75t_SL g291 ( .A1(n_180), .A2(n_292), .B(n_299), .C(n_306), .Y(n_291) );
INVx1_ASAP7_75t_L g380 ( .A(n_180), .Y(n_380) );
INVx1_ASAP7_75t_L g412 ( .A(n_181), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_182), .A2(n_189), .B1(n_888), .B2(n_891), .Y(n_887) );
INVx1_ASAP7_75t_L g810 ( .A(n_184), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g962 ( .A(n_185), .Y(n_962) );
INVx1_ASAP7_75t_L g1004 ( .A(n_186), .Y(n_1004) );
INVx1_ASAP7_75t_L g495 ( .A(n_187), .Y(n_495) );
INVx1_ASAP7_75t_L g488 ( .A(n_188), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_189), .A2(n_261), .B1(n_900), .B2(n_901), .Y(n_899) );
CKINVDCx5p33_ASAP7_75t_R g923 ( .A(n_190), .Y(n_923) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_192), .Y(n_297) );
INVx1_ASAP7_75t_L g1000 ( .A(n_193), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1184 ( .A1(n_194), .A2(n_240), .B1(n_1170), .B2(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g817 ( .A(n_196), .Y(n_817) );
INVx1_ASAP7_75t_L g980 ( .A(n_198), .Y(n_980) );
OAI211xp5_ASAP7_75t_L g985 ( .A1(n_198), .A2(n_570), .B(n_616), .C(n_986), .Y(n_985) );
CKINVDCx5p33_ASAP7_75t_R g918 ( .A(n_199), .Y(n_918) );
INVx1_ASAP7_75t_L g760 ( .A(n_200), .Y(n_760) );
AO22x1_ASAP7_75t_L g1169 ( .A1(n_202), .A2(n_230), .B1(n_1170), .B2(n_1174), .Y(n_1169) );
AOI221xp5_ASAP7_75t_L g1092 ( .A1(n_204), .A2(n_265), .B1(n_623), .B2(n_685), .C(n_854), .Y(n_1092) );
CKINVDCx16_ASAP7_75t_R g1244 ( .A(n_205), .Y(n_1244) );
OAI211xp5_ASAP7_75t_L g1115 ( .A1(n_207), .A2(n_530), .B(n_1116), .C(n_1119), .Y(n_1115) );
INVx1_ASAP7_75t_L g1131 ( .A(n_207), .Y(n_1131) );
INVx1_ASAP7_75t_L g642 ( .A(n_208), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g1381 ( .A1(n_209), .A2(n_1382), .B1(n_1383), .B2(n_1467), .Y(n_1381) );
INVxp67_ASAP7_75t_SL g1467 ( .A(n_209), .Y(n_1467) );
AOI22xp33_ASAP7_75t_L g1473 ( .A1(n_209), .A2(n_1474), .B1(n_1477), .B2(n_1524), .Y(n_1473) );
INVx1_ASAP7_75t_L g580 ( .A(n_210), .Y(n_580) );
OAI211xp5_ASAP7_75t_L g587 ( .A1(n_210), .A2(n_364), .B(n_370), .C(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g781 ( .A(n_211), .Y(n_781) );
INVx1_ASAP7_75t_L g311 ( .A(n_212), .Y(n_311) );
OA22x2_ASAP7_75t_L g806 ( .A1(n_213), .A2(n_807), .B1(n_856), .B2(n_857), .Y(n_806) );
INVxp67_ASAP7_75t_SL g857 ( .A(n_213), .Y(n_857) );
INVx1_ASAP7_75t_L g483 ( .A(n_214), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_215), .A2(n_277), .B1(n_741), .B2(n_743), .Y(n_740) );
INVx1_ASAP7_75t_L g1058 ( .A(n_217), .Y(n_1058) );
CKINVDCx5p33_ASAP7_75t_R g944 ( .A(n_218), .Y(n_944) );
INVx1_ASAP7_75t_L g422 ( .A(n_220), .Y(n_422) );
INVx1_ASAP7_75t_L g638 ( .A(n_221), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g1194 ( .A1(n_222), .A2(n_252), .B1(n_1177), .B2(n_1180), .Y(n_1194) );
BUFx3_ASAP7_75t_L g303 ( .A(n_224), .Y(n_303) );
INVx1_ASAP7_75t_L g324 ( .A(n_224), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_225), .A2(n_267), .B1(n_318), .B2(n_325), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_225), .A2(n_267), .B1(n_348), .B2(n_357), .Y(n_347) );
INVx1_ASAP7_75t_L g577 ( .A(n_226), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g1246 ( .A(n_227), .Y(n_1246) );
OAI22xp33_ASAP7_75t_L g521 ( .A1(n_229), .A2(n_260), .B1(n_522), .B2(n_523), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_229), .A2(n_260), .B1(n_318), .B2(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g1403 ( .A(n_232), .Y(n_1403) );
INVx1_ASAP7_75t_L g1029 ( .A(n_233), .Y(n_1029) );
INVx1_ASAP7_75t_L g1012 ( .A(n_234), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_235), .A2(n_265), .B1(n_749), .B2(n_1076), .Y(n_1075) );
OAI211xp5_ASAP7_75t_L g977 ( .A1(n_236), .A2(n_600), .B(n_942), .C(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g987 ( .A(n_236), .Y(n_987) );
INVx1_ASAP7_75t_L g630 ( .A(n_237), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g930 ( .A(n_239), .Y(n_930) );
OAI211xp5_ASAP7_75t_L g597 ( .A1(n_241), .A2(n_598), .B(n_600), .C(n_604), .Y(n_597) );
INVx1_ASAP7_75t_L g619 ( .A(n_241), .Y(n_619) );
INVx1_ASAP7_75t_L g345 ( .A(n_242), .Y(n_345) );
INVx2_ASAP7_75t_L g406 ( .A(n_242), .Y(n_406) );
INVx1_ASAP7_75t_L g463 ( .A(n_242), .Y(n_463) );
INVx1_ASAP7_75t_L g519 ( .A(n_243), .Y(n_519) );
OAI211xp5_ASAP7_75t_L g814 ( .A1(n_245), .A2(n_725), .B(n_815), .C(n_816), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_248), .A2(n_256), .B1(n_848), .B2(n_850), .Y(n_847) );
XNOR2x1_ASAP7_75t_L g1095 ( .A(n_250), .B(n_1096), .Y(n_1095) );
AO22x1_ASAP7_75t_L g1176 ( .A1(n_250), .A2(n_272), .B1(n_1177), .B2(n_1180), .Y(n_1176) );
INVx1_ASAP7_75t_L g1407 ( .A(n_251), .Y(n_1407) );
XNOR2xp5_ASAP7_75t_L g1053 ( .A(n_253), .B(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g312 ( .A(n_255), .Y(n_312) );
OAI211xp5_ASAP7_75t_L g363 ( .A1(n_255), .A2(n_364), .B(n_370), .C(n_374), .Y(n_363) );
INVx1_ASAP7_75t_L g557 ( .A(n_257), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g1062 ( .A(n_258), .Y(n_1062) );
INVx1_ASAP7_75t_L g1490 ( .A(n_259), .Y(n_1490) );
INVx1_ASAP7_75t_L g1038 ( .A(n_262), .Y(n_1038) );
INVxp67_ASAP7_75t_SL g1141 ( .A(n_263), .Y(n_1141) );
INVx1_ASAP7_75t_L g873 ( .A(n_264), .Y(n_873) );
INVx1_ASAP7_75t_L g1102 ( .A(n_266), .Y(n_1102) );
INVx1_ASAP7_75t_L g1031 ( .A(n_269), .Y(n_1031) );
XNOR2xp5_ASAP7_75t_L g954 ( .A(n_270), .B(n_955), .Y(n_954) );
OAI22xp33_ASAP7_75t_L g981 ( .A1(n_271), .A2(n_276), .B1(n_326), .B2(n_611), .Y(n_981) );
INVx1_ASAP7_75t_L g441 ( .A(n_273), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g933 ( .A(n_274), .Y(n_933) );
INVx1_ASAP7_75t_L g714 ( .A(n_278), .Y(n_714) );
INVx1_ASAP7_75t_L g552 ( .A(n_279), .Y(n_552) );
INVx1_ASAP7_75t_L g475 ( .A(n_280), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_1148), .B(n_1162), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_990), .B1(n_1146), .B2(n_1147), .Y(n_282) );
INVx1_ASAP7_75t_L g1146 ( .A(n_283), .Y(n_1146) );
XNOR2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_802), .Y(n_283) );
XNOR2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_537), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_288), .B1(n_469), .B2(n_470), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND3xp33_ASAP7_75t_L g289 ( .A(n_290), .B(n_346), .C(n_401), .Y(n_289) );
OAI31xp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_317), .A3(n_331), .B(n_338), .Y(n_290) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g1487 ( .A1(n_294), .A2(n_1488), .B1(n_1489), .B2(n_1490), .Y(n_1487) );
BUFx4f_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx4f_ASAP7_75t_L g506 ( .A(n_295), .Y(n_506) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_295), .Y(n_599) );
INVx4_ASAP7_75t_L g659 ( .A(n_295), .Y(n_659) );
BUFx4f_ASAP7_75t_L g1142 ( .A(n_295), .Y(n_1142) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
BUFx3_ASAP7_75t_L g425 ( .A(n_296), .Y(n_425) );
NAND2x1_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x2_ASAP7_75t_L g305 ( .A(n_297), .B(n_298), .Y(n_305) );
INVx1_ASAP7_75t_L g316 ( .A(n_297), .Y(n_316) );
OR2x2_ASAP7_75t_L g322 ( .A(n_297), .B(n_298), .Y(n_322) );
INVx2_ASAP7_75t_L g330 ( .A(n_297), .Y(n_330) );
AND2x2_ASAP7_75t_L g336 ( .A(n_297), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g421 ( .A(n_297), .Y(n_421) );
BUFx2_ASAP7_75t_L g310 ( .A(n_298), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_298), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g337 ( .A(n_298), .Y(n_337) );
OR2x2_ASAP7_75t_L g420 ( .A(n_298), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g737 ( .A(n_298), .Y(n_737) );
AND2x2_ASAP7_75t_L g739 ( .A(n_298), .B(n_330), .Y(n_739) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g530 ( .A(n_300), .Y(n_530) );
INVx1_ASAP7_75t_L g581 ( .A(n_300), .Y(n_581) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_304), .Y(n_300) );
AND2x2_ASAP7_75t_L g601 ( .A(n_301), .B(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g609 ( .A(n_301), .B(n_328), .Y(n_609) );
AND2x2_ASAP7_75t_L g721 ( .A(n_301), .B(n_310), .Y(n_721) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVxp67_ASAP7_75t_L g333 ( .A(n_302), .Y(n_333) );
AND2x4_ASAP7_75t_L g1410 ( .A(n_302), .B(n_341), .Y(n_1410) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx2_ASAP7_75t_L g309 ( .A(n_303), .Y(n_309) );
AND2x4_ASAP7_75t_L g314 ( .A(n_303), .B(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g434 ( .A(n_303), .B(n_341), .Y(n_434) );
BUFx3_ASAP7_75t_L g743 ( .A(n_304), .Y(n_743) );
BUFx6f_ASAP7_75t_L g837 ( .A(n_304), .Y(n_837) );
BUFx3_ASAP7_75t_L g839 ( .A(n_304), .Y(n_839) );
BUFx3_ASAP7_75t_L g891 ( .A(n_304), .Y(n_891) );
AND2x4_ASAP7_75t_SL g1405 ( .A(n_304), .B(n_1406), .Y(n_1405) );
AND2x6_ASAP7_75t_L g1421 ( .A(n_304), .B(n_1394), .Y(n_1421) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g603 ( .A(n_305), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_311), .B1(n_312), .B2(n_313), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_307), .A2(n_577), .B1(n_578), .B2(n_580), .Y(n_576) );
BUFx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_308), .A2(n_314), .B1(n_519), .B2(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_308), .A2(n_313), .B1(n_605), .B2(n_606), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_308), .A2(n_313), .B1(n_760), .B2(n_761), .Y(n_759) );
INVx1_ASAP7_75t_L g882 ( .A(n_308), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_308), .A2(n_578), .B1(n_1029), .B2(n_1031), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1510 ( .A1(n_308), .A2(n_818), .B1(n_1511), .B2(n_1512), .Y(n_1510) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
OR2x2_ASAP7_75t_L g327 ( .A(n_309), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g884 ( .A(n_309), .B(n_748), .Y(n_884) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_309), .B(n_310), .Y(n_1121) );
BUFx2_ASAP7_75t_L g1402 ( .A(n_310), .Y(n_1402) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_311), .A2(n_375), .B1(n_380), .B2(n_381), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g978 ( .A1(n_313), .A2(n_721), .B1(n_979), .B2(n_980), .Y(n_978) );
BUFx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g579 ( .A(n_314), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_314), .A2(n_701), .B1(n_705), .B2(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g819 ( .A(n_314), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_314), .A2(n_721), .B1(n_1062), .B2(n_1063), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_314), .A2(n_1120), .B1(n_1121), .B2(n_1122), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1432 ( .A(n_315), .B(n_1394), .Y(n_1432) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx2_ASAP7_75t_L g1124 ( .A(n_319), .Y(n_1124) );
OR2x6_ASAP7_75t_L g319 ( .A(n_320), .B(n_323), .Y(n_319) );
OR2x6_ASAP7_75t_L g332 ( .A(n_320), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g608 ( .A(n_320), .B(n_323), .Y(n_608) );
INVx1_ASAP7_75t_L g665 ( .A(n_320), .Y(n_665) );
BUFx4f_ASAP7_75t_L g1017 ( .A(n_320), .Y(n_1017) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx3_ASAP7_75t_L g411 ( .A(n_321), .Y(n_411) );
BUFx4f_ASAP7_75t_L g440 ( .A(n_321), .Y(n_440) );
INVx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g335 ( .A(n_323), .B(n_336), .Y(n_335) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g535 ( .A(n_327), .Y(n_535) );
INVx8_ASAP7_75t_L g415 ( .A(n_328), .Y(n_415) );
BUFx2_ASAP7_75t_L g1018 ( .A(n_328), .Y(n_1018) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx3_ASAP7_75t_L g811 ( .A(n_332), .Y(n_811) );
OR2x6_ASAP7_75t_L g611 ( .A(n_333), .B(n_411), .Y(n_611) );
CKINVDCx16_ASAP7_75t_R g334 ( .A(n_335), .Y(n_334) );
INVx3_ASAP7_75t_SL g528 ( .A(n_335), .Y(n_528) );
INVx4_ASAP7_75t_L g574 ( .A(n_335), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_335), .A2(n_714), .B1(n_715), .B2(n_716), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_335), .A2(n_810), .B1(n_811), .B2(n_812), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_335), .A2(n_862), .B1(n_863), .B2(n_876), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g1056 ( .A1(n_335), .A2(n_715), .B1(n_1057), .B2(n_1058), .Y(n_1056) );
BUFx6f_ASAP7_75t_L g742 ( .A(n_336), .Y(n_742) );
BUFx3_ASAP7_75t_L g890 ( .A(n_336), .Y(n_890) );
OAI31xp33_ASAP7_75t_L g940 ( .A1(n_338), .A2(n_941), .A3(n_946), .B(n_947), .Y(n_940) );
OAI31xp33_ASAP7_75t_L g976 ( .A1(n_338), .A2(n_977), .A3(n_981), .B(n_982), .Y(n_976) );
INVx1_ASAP7_75t_L g1048 ( .A(n_338), .Y(n_1048) );
OAI31xp33_ASAP7_75t_SL g1113 ( .A1(n_338), .A2(n_1114), .A3(n_1115), .B(n_1123), .Y(n_1113) );
OAI31xp33_ASAP7_75t_L g1507 ( .A1(n_338), .A2(n_1508), .A3(n_1513), .B(n_1515), .Y(n_1507) );
BUFx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx2_ASAP7_75t_SL g536 ( .A(n_339), .Y(n_536) );
BUFx3_ASAP7_75t_L g584 ( .A(n_339), .Y(n_584) );
INVx1_ASAP7_75t_L g726 ( .A(n_339), .Y(n_726) );
OAI31xp33_ASAP7_75t_L g756 ( .A1(n_339), .A2(n_757), .A3(n_758), .B(n_762), .Y(n_756) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
INVx1_ASAP7_75t_L g1161 ( .A(n_340), .Y(n_1161) );
NOR2xp33_ASAP7_75t_L g1472 ( .A(n_340), .B(n_1153), .Y(n_1472) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g1431 ( .A(n_343), .B(n_1432), .Y(n_1431) );
INVxp67_ASAP7_75t_L g1445 ( .A(n_343), .Y(n_1445) );
BUFx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g400 ( .A(n_344), .Y(n_400) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OAI31xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_363), .A3(n_384), .B(n_394), .Y(n_346) );
BUFx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx3_ASAP7_75t_L g522 ( .A(n_349), .Y(n_522) );
INVx2_ASAP7_75t_SL g872 ( .A(n_349), .Y(n_872) );
OR2x4_ASAP7_75t_L g349 ( .A(n_350), .B(n_353), .Y(n_349) );
AND2x4_ASAP7_75t_L g389 ( .A(n_350), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g710 ( .A(n_350), .B(n_390), .Y(n_710) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OR2x6_ASAP7_75t_L g359 ( .A(n_351), .B(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g371 ( .A(n_351), .B(n_372), .Y(n_371) );
OR2x4_ASAP7_75t_L g387 ( .A(n_351), .B(n_353), .Y(n_387) );
NAND3x1_ASAP7_75t_L g461 ( .A(n_351), .B(n_462), .C(n_464), .Y(n_461) );
NAND2x1p5_ASAP7_75t_L g650 ( .A(n_351), .B(n_464), .Y(n_650) );
AND2x4_ASAP7_75t_L g1443 ( .A(n_351), .B(n_1444), .Y(n_1443) );
INVx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx3_ASAP7_75t_L g378 ( .A(n_352), .Y(n_378) );
NAND2xp33_ASAP7_75t_SL g448 ( .A(n_352), .B(n_397), .Y(n_448) );
BUFx3_ASAP7_75t_L g450 ( .A(n_353), .Y(n_450) );
BUFx3_ASAP7_75t_L g468 ( .A(n_353), .Y(n_468) );
BUFx4f_ASAP7_75t_L g631 ( .A(n_353), .Y(n_631) );
INVx2_ASAP7_75t_L g793 ( .A(n_353), .Y(n_793) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_354), .B(n_362), .Y(n_361) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_354), .Y(n_369) );
AND2x4_ASAP7_75t_L g372 ( .A(n_354), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g393 ( .A(n_354), .Y(n_393) );
INVx1_ASAP7_75t_L g679 ( .A(n_355), .Y(n_679) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g392 ( .A(n_356), .Y(n_392) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g524 ( .A(n_359), .Y(n_524) );
INVx1_ASAP7_75t_L g592 ( .A(n_359), .Y(n_592) );
BUFx3_ASAP7_75t_L g1523 ( .A(n_359), .Y(n_1523) );
BUFx3_ASAP7_75t_L g456 ( .A(n_360), .Y(n_456) );
INVx1_ASAP7_75t_L g486 ( .A(n_360), .Y(n_486) );
BUFx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g493 ( .A(n_361), .Y(n_493) );
INVx1_ASAP7_75t_L g368 ( .A(n_362), .Y(n_368) );
INVx2_ASAP7_75t_L g373 ( .A(n_362), .Y(n_373) );
OAI22xp33_ASAP7_75t_L g465 ( .A1(n_364), .A2(n_412), .B1(n_431), .B2(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g496 ( .A(n_365), .Y(n_496) );
INVx1_ASAP7_75t_L g1129 ( .A(n_365), .Y(n_1129) );
INVx1_ASAP7_75t_L g1519 ( .A(n_365), .Y(n_1519) );
INVx4_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_366), .Y(n_633) );
INVx3_ASAP7_75t_L g921 ( .A(n_366), .Y(n_921) );
OR2x2_ASAP7_75t_L g1430 ( .A(n_366), .B(n_1389), .Y(n_1430) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx3_ASAP7_75t_L g452 ( .A(n_367), .Y(n_452) );
BUFx2_ASAP7_75t_L g516 ( .A(n_367), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
BUFx2_ASAP7_75t_L g383 ( .A(n_368), .Y(n_383) );
BUFx2_ASAP7_75t_L g379 ( .A(n_369), .Y(n_379) );
AND2x4_ASAP7_75t_L g683 ( .A(n_369), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g1451 ( .A(n_369), .Y(n_1451) );
CKINVDCx8_ASAP7_75t_R g370 ( .A(n_371), .Y(n_370) );
CKINVDCx8_ASAP7_75t_R g616 ( .A(n_371), .Y(n_616) );
NOR3xp33_ASAP7_75t_L g823 ( .A(n_371), .B(n_824), .C(n_825), .Y(n_823) );
AOI211xp5_ASAP7_75t_L g864 ( .A1(n_371), .A2(n_865), .B(n_866), .C(n_867), .Y(n_864) );
NOR2xp33_ASAP7_75t_L g1026 ( .A(n_371), .B(n_1027), .Y(n_1026) );
NOR3xp33_ASAP7_75t_L g1069 ( .A(n_371), .B(n_1070), .C(n_1072), .Y(n_1069) );
BUFx3_ASAP7_75t_L g623 ( .A(n_372), .Y(n_623) );
BUFx2_ASAP7_75t_L g675 ( .A(n_372), .Y(n_675) );
INVx2_ASAP7_75t_L g703 ( .A(n_372), .Y(n_703) );
BUFx2_ASAP7_75t_L g767 ( .A(n_372), .Y(n_767) );
BUFx2_ASAP7_75t_L g866 ( .A(n_372), .Y(n_866) );
BUFx2_ASAP7_75t_L g1104 ( .A(n_372), .Y(n_1104) );
BUFx2_ASAP7_75t_L g1458 ( .A(n_372), .Y(n_1458) );
INVx1_ASAP7_75t_L g684 ( .A(n_373), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_375), .A2(n_381), .B1(n_1120), .B2(n_1131), .Y(n_1130) );
BUFx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx3_ASAP7_75t_L g518 ( .A(n_376), .Y(n_518) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
AND2x4_ASAP7_75t_L g382 ( .A(n_377), .B(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g618 ( .A(n_377), .B(n_379), .Y(n_618) );
AND2x2_ASAP7_75t_L g620 ( .A(n_377), .B(n_383), .Y(n_620) );
AND2x4_ASAP7_75t_L g706 ( .A(n_377), .B(n_379), .Y(n_706) );
INVx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND3x4_ASAP7_75t_L g686 ( .A(n_378), .B(n_397), .C(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_381), .A2(n_518), .B1(n_519), .B2(n_520), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_381), .A2(n_518), .B1(n_577), .B2(n_589), .Y(n_588) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g826 ( .A(n_382), .Y(n_826) );
AOI222xp33_ASAP7_75t_L g1028 ( .A1(n_382), .A2(n_675), .B1(n_706), .B2(n_1029), .C1(n_1030), .C2(n_1031), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1520 ( .A1(n_382), .A2(n_618), .B1(n_1511), .B2(n_1521), .Y(n_1520) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_387), .Y(n_511) );
INVx2_ASAP7_75t_SL g829 ( .A(n_387), .Y(n_829) );
INVx1_ASAP7_75t_L g1037 ( .A(n_387), .Y(n_1037) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g512 ( .A(n_389), .Y(n_512) );
INVx1_ASAP7_75t_L g614 ( .A(n_389), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_389), .A2(n_810), .B1(n_812), .B2(n_829), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_389), .A2(n_829), .B1(n_862), .B2(n_863), .Y(n_861) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_390), .Y(n_455) );
INVx2_ASAP7_75t_L g458 ( .A(n_390), .Y(n_458) );
INVx1_ASAP7_75t_L g489 ( .A(n_390), .Y(n_489) );
INVx2_ASAP7_75t_L g849 ( .A(n_390), .Y(n_849) );
BUFx6f_ASAP7_75t_L g900 ( .A(n_390), .Y(n_900) );
INVx2_ASAP7_75t_L g1462 ( .A(n_390), .Y(n_1462) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_391), .Y(n_482) );
BUFx8_ASAP7_75t_L g637 ( .A(n_391), .Y(n_637) );
INVx2_ASAP7_75t_L g929 ( .A(n_391), .Y(n_929) );
AND2x4_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
AND2x4_ASAP7_75t_L g678 ( .A(n_393), .B(n_679), .Y(n_678) );
BUFx2_ASAP7_75t_L g593 ( .A(n_394), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g859 ( .A1(n_394), .A2(n_536), .B1(n_860), .B2(n_874), .C(n_885), .Y(n_859) );
OAI31xp33_ASAP7_75t_L g1125 ( .A1(n_394), .A2(n_1126), .A3(n_1128), .B(n_1132), .Y(n_1125) );
AND2x2_ASAP7_75t_SL g394 ( .A(n_395), .B(n_398), .Y(n_394) );
AND2x2_ASAP7_75t_L g525 ( .A(n_395), .B(n_398), .Y(n_525) );
AND2x2_ASAP7_75t_L g625 ( .A(n_395), .B(n_398), .Y(n_625) );
AND2x2_ASAP7_75t_L g711 ( .A(n_395), .B(n_398), .Y(n_711) );
AND2x4_ASAP7_75t_L g1040 ( .A(n_395), .B(n_398), .Y(n_1040) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g1444 ( .A(n_397), .Y(n_1444) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g436 ( .A(n_400), .Y(n_436) );
OR2x2_ASAP7_75t_L g447 ( .A(n_400), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_SL g662 ( .A(n_400), .B(n_434), .Y(n_662) );
OR2x2_ASAP7_75t_L g1389 ( .A(n_400), .B(n_1390), .Y(n_1389) );
NOR2xp33_ASAP7_75t_SL g401 ( .A(n_402), .B(n_445), .Y(n_401) );
OAI33xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_408), .A3(n_416), .B1(n_426), .B2(n_432), .B3(n_437), .Y(n_402) );
INVx2_ASAP7_75t_SL g732 ( .A(n_403), .Y(n_732) );
INVx2_ASAP7_75t_SL g1074 ( .A(n_403), .Y(n_1074) );
OAI33xp33_ASAP7_75t_L g1482 ( .A1(n_403), .A2(n_1145), .A3(n_1483), .B1(n_1487), .B2(n_1491), .B3(n_1495), .Y(n_1482) );
INVx4_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g500 ( .A(n_404), .Y(n_500) );
INVx2_ASAP7_75t_L g543 ( .A(n_404), .Y(n_543) );
INVx2_ASAP7_75t_L g654 ( .A(n_404), .Y(n_654) );
AND2x4_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
OR2x2_ASAP7_75t_L g649 ( .A(n_405), .B(n_650), .Y(n_649) );
OR2x6_ASAP7_75t_L g696 ( .A(n_405), .B(n_650), .Y(n_696) );
INVx1_ASAP7_75t_L g1398 ( .A(n_405), .Y(n_1398) );
BUFx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g687 ( .A(n_406), .Y(n_687) );
OAI22xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_412), .B2(n_413), .Y(n_408) );
OAI22xp33_ASAP7_75t_L g449 ( .A1(n_409), .A2(n_430), .B1(n_450), .B2(n_451), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_410), .A2(n_413), .B1(n_483), .B2(n_490), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_410), .A2(n_413), .B1(n_556), .B2(n_557), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g1144 ( .A1(n_410), .A2(n_413), .B1(n_1102), .B2(n_1109), .Y(n_1144) );
OAI22xp5_ASAP7_75t_L g1495 ( .A1(n_410), .A2(n_1496), .B1(n_1497), .B2(n_1498), .Y(n_1495) );
BUFx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OAI22xp5_ASAP7_75t_SL g544 ( .A1(n_413), .A2(n_545), .B1(n_546), .B2(n_547), .Y(n_544) );
INVx6_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx5_ASAP7_75t_L g1138 ( .A(n_414), .Y(n_1138) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g443 ( .A(n_415), .Y(n_443) );
INVx1_ASAP7_75t_L g503 ( .A(n_415), .Y(n_503) );
INVx4_ASAP7_75t_L g666 ( .A(n_415), .Y(n_666) );
INVx2_ASAP7_75t_L g776 ( .A(n_415), .Y(n_776) );
INVx2_ASAP7_75t_SL g788 ( .A(n_415), .Y(n_788) );
INVx2_ASAP7_75t_L g1497 ( .A(n_415), .Y(n_1497) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_422), .B2(n_423), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_417), .A2(n_441), .B1(n_454), .B2(n_456), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_418), .A2(n_425), .B1(n_549), .B2(n_550), .Y(n_548) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g780 ( .A(n_419), .Y(n_780) );
BUFx2_ASAP7_75t_L g1022 ( .A(n_419), .Y(n_1022) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx2_ASAP7_75t_L g429 ( .A(n_420), .Y(n_429) );
INVx1_ASAP7_75t_L g657 ( .A(n_420), .Y(n_657) );
BUFx2_ASAP7_75t_L g938 ( .A(n_420), .Y(n_938) );
AND2x2_ASAP7_75t_L g736 ( .A(n_421), .B(n_737), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_422), .A2(n_444), .B1(n_456), .B2(n_458), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g1491 ( .A1(n_423), .A2(n_1492), .B1(n_1493), .B2(n_1494), .Y(n_1491) );
INVx5_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_425), .A2(n_427), .B1(n_430), .B2(n_431), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_425), .A2(n_427), .B1(n_476), .B2(n_497), .Y(n_507) );
BUFx2_ASAP7_75t_SL g553 ( .A(n_425), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_425), .A2(n_632), .B1(n_648), .B2(n_656), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_425), .A2(n_919), .B1(n_933), .B2(n_938), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_425), .A2(n_780), .B1(n_962), .B2(n_963), .Y(n_961) );
BUFx3_ASAP7_75t_L g1118 ( .A(n_425), .Y(n_1118) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_427), .A2(n_552), .B1(n_553), .B2(n_554), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g1139 ( .A1(n_427), .A2(n_553), .B1(n_1101), .B2(n_1108), .Y(n_1139) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx4_ASAP7_75t_L g505 ( .A(n_428), .Y(n_505) );
INVx2_ASAP7_75t_L g1489 ( .A(n_428), .Y(n_1489) );
INVx4_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI33xp33_ASAP7_75t_L g498 ( .A1(n_432), .A2(n_499), .A3(n_501), .B1(n_504), .B2(n_507), .B3(n_508), .Y(n_498) );
OAI33xp33_ASAP7_75t_L g542 ( .A1(n_432), .A2(n_543), .A3(n_544), .B1(n_548), .B2(n_551), .B3(n_555), .Y(n_542) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND3xp33_ASAP7_75t_L g895 ( .A(n_433), .B(n_896), .C(n_897), .Y(n_895) );
CKINVDCx5p33_ASAP7_75t_R g1145 ( .A(n_433), .Y(n_1145) );
AND2x4_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx4_ASAP7_75t_L g1418 ( .A(n_434), .Y(n_1418) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_441), .B1(n_442), .B2(n_444), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g502 ( .A(n_439), .Y(n_502) );
INVx3_ASAP7_75t_L g1485 ( .A(n_439), .Y(n_1485) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx3_ASAP7_75t_L g546 ( .A(n_440), .Y(n_546) );
INVx4_ASAP7_75t_L g653 ( .A(n_440), .Y(n_653) );
BUFx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI33xp33_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_449), .A3(n_453), .B1(n_457), .B2(n_459), .B3(n_465), .Y(n_445) );
OAI33xp33_ASAP7_75t_L g473 ( .A1(n_446), .A2(n_459), .A3(n_474), .B1(n_478), .B2(n_487), .B3(n_494), .Y(n_473) );
OAI33xp33_ASAP7_75t_L g1499 ( .A1(n_446), .A2(n_1112), .A3(n_1500), .B1(n_1503), .B2(n_1504), .B3(n_1505), .Y(n_1499) );
BUFx8_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx4f_ASAP7_75t_L g559 ( .A(n_447), .Y(n_559) );
BUFx4f_ASAP7_75t_L g628 ( .A(n_447), .Y(n_628) );
BUFx2_ASAP7_75t_L g997 ( .A(n_447), .Y(n_997) );
OAI22xp33_ASAP7_75t_L g474 ( .A1(n_450), .A2(n_475), .B1(n_476), .B2(n_477), .Y(n_474) );
OAI22xp33_ASAP7_75t_L g494 ( .A1(n_450), .A2(n_495), .B1(n_496), .B2(n_497), .Y(n_494) );
OAI22xp33_ASAP7_75t_L g1010 ( .A1(n_450), .A2(n_633), .B1(n_1011), .B2(n_1012), .Y(n_1010) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_452), .Y(n_477) );
INVx2_ASAP7_75t_L g564 ( .A(n_452), .Y(n_564) );
OAI22xp33_ASAP7_75t_L g646 ( .A1(n_452), .A2(n_631), .B1(n_647), .B2(n_648), .Y(n_646) );
OAI22xp33_ASAP7_75t_L g791 ( .A1(n_452), .A2(n_774), .B1(n_783), .B2(n_792), .Y(n_791) );
OAI22xp33_ASAP7_75t_L g931 ( .A1(n_452), .A2(n_792), .B1(n_932), .B2(n_933), .Y(n_931) );
OAI22xp33_ASAP7_75t_L g975 ( .A1(n_452), .A2(n_792), .B1(n_960), .B2(n_966), .Y(n_975) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_456), .A2(n_550), .B1(n_557), .B2(n_567), .Y(n_566) );
OAI221xp5_ASAP7_75t_L g1099 ( .A1(n_456), .A2(n_1100), .B1(n_1101), .B2(n_1102), .C(n_1103), .Y(n_1099) );
OAI221xp5_ASAP7_75t_L g1106 ( .A1(n_456), .A2(n_1107), .B1(n_1108), .B2(n_1109), .C(n_1110), .Y(n_1106) );
OAI22xp5_ASAP7_75t_L g1503 ( .A1(n_456), .A2(n_1100), .B1(n_1488), .B2(n_1496), .Y(n_1503) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_458), .A2(n_781), .B1(n_789), .B2(n_798), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_458), .A2(n_796), .B1(n_923), .B2(n_924), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g972 ( .A1(n_458), .A2(n_796), .B1(n_962), .B2(n_968), .Y(n_972) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g568 ( .A(n_460), .Y(n_568) );
INVx2_ASAP7_75t_L g1112 ( .A(n_460), .Y(n_1112) );
INVx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx3_ASAP7_75t_L g906 ( .A(n_461), .Y(n_906) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g1392 ( .A(n_463), .Y(n_1392) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVxp67_ASAP7_75t_SL g562 ( .A(n_468), .Y(n_562) );
INVx1_ASAP7_75t_L g1502 ( .A(n_468), .Y(n_1502) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_509), .C(n_526), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_498), .Y(n_472) );
OAI22xp33_ASAP7_75t_L g501 ( .A1(n_475), .A2(n_495), .B1(n_502), .B2(n_503), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B1(n_483), .B2(n_484), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_479), .A2(n_488), .B1(n_505), .B2(n_506), .Y(n_504) );
BUFx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_481), .A2(n_491), .B1(n_549), .B2(n_556), .Y(n_565) );
INVx5_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_SL g567 ( .A(n_482), .Y(n_567) );
INVx3_ASAP7_75t_L g795 ( .A(n_482), .Y(n_795) );
INVx2_ASAP7_75t_SL g1089 ( .A(n_482), .Y(n_1089) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g639 ( .A(n_486), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B1(n_490), .B2(n_491), .Y(n_487) );
INVx1_ASAP7_75t_L g852 ( .A(n_489), .Y(n_852) );
OAI22xp33_ASAP7_75t_SL g1504 ( .A1(n_491), .A2(n_1462), .B1(n_1490), .B2(n_1498), .Y(n_1504) );
CKINVDCx8_ASAP7_75t_R g491 ( .A(n_492), .Y(n_491) );
INVx3_ASAP7_75t_L g796 ( .A(n_492), .Y(n_796) );
INVx3_ASAP7_75t_L g798 ( .A(n_492), .Y(n_798) );
INVx3_ASAP7_75t_L g974 ( .A(n_492), .Y(n_974) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g644 ( .A(n_493), .Y(n_644) );
OAI22xp33_ASAP7_75t_L g799 ( .A1(n_496), .A2(n_631), .B1(n_777), .B2(n_784), .Y(n_799) );
OA33x2_ASAP7_75t_L g1134 ( .A1(n_499), .A2(n_1135), .A3(n_1139), .B1(n_1140), .B2(n_1144), .B3(n_1145), .Y(n_1134) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI33xp33_ASAP7_75t_L g772 ( .A1(n_500), .A2(n_773), .A3(n_778), .B1(n_782), .B2(n_785), .B3(n_786), .Y(n_772) );
OAI33xp33_ASAP7_75t_L g957 ( .A1(n_500), .A2(n_785), .A3(n_958), .B1(n_961), .B2(n_964), .B3(n_967), .Y(n_957) );
OAI22xp33_ASAP7_75t_L g652 ( .A1(n_503), .A2(n_630), .B1(n_647), .B2(n_653), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_506), .A2(n_780), .B1(n_783), .B2(n_784), .Y(n_782) );
OAI31xp33_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_513), .A3(n_521), .B(n_525), .Y(n_509) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g571 ( .A(n_516), .Y(n_571) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_524), .A2(n_871), .B1(n_872), .B2(n_873), .Y(n_870) );
OAI31xp33_ASAP7_75t_L g1516 ( .A1(n_525), .A2(n_1517), .A3(n_1518), .B(n_1522), .Y(n_1516) );
OAI31xp33_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_529), .A3(n_533), .B(n_536), .Y(n_526) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g583 ( .A(n_535), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_535), .A2(n_871), .B1(n_873), .B2(n_884), .Y(n_883) );
INVxp67_ASAP7_75t_SL g1514 ( .A(n_535), .Y(n_1514) );
OAI31xp33_ASAP7_75t_SL g596 ( .A1(n_536), .A2(n_597), .A3(n_607), .B(n_610), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_669), .B1(n_800), .B2(n_801), .Y(n_537) );
INVx1_ASAP7_75t_L g800 ( .A(n_538), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_594), .B1(n_667), .B2(n_668), .Y(n_538) );
INVx1_ASAP7_75t_L g668 ( .A(n_539), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_572), .C(n_585), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_558), .Y(n_541) );
OAI22xp33_ASAP7_75t_L g560 ( .A1(n_545), .A2(n_552), .B1(n_561), .B2(n_563), .Y(n_560) );
OAI22xp33_ASAP7_75t_L g569 ( .A1(n_547), .A2(n_554), .B1(n_561), .B2(n_570), .Y(n_569) );
OAI33xp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .A3(n_565), .B1(n_566), .B2(n_568), .B3(n_569), .Y(n_558) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g973 ( .A1(n_567), .A2(n_963), .B1(n_969), .B2(n_974), .Y(n_973) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OAI31xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_575), .A3(n_582), .B(n_584), .Y(n_572) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI31xp33_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .A3(n_590), .B(n_593), .Y(n_585) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_592), .A2(n_710), .B1(n_1033), .B2(n_1034), .Y(n_1032) );
INVx2_ASAP7_75t_SL g667 ( .A(n_594), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_612), .C(n_626), .Y(n_595) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_599), .A2(n_779), .B1(n_780), .B2(n_781), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_599), .A2(n_780), .B1(n_965), .B2(n_966), .Y(n_964) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g725 ( .A(n_601), .Y(n_725) );
AOI211xp5_ASAP7_75t_L g877 ( .A1(n_601), .A2(n_878), .B(n_880), .C(n_881), .Y(n_877) );
INVx1_ASAP7_75t_L g724 ( .A(n_602), .Y(n_724) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
BUFx2_ASAP7_75t_L g879 ( .A(n_603), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_605), .A2(n_618), .B1(n_619), .B2(n_620), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_606), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g715 ( .A(n_611), .Y(n_715) );
INVx1_ASAP7_75t_L g876 ( .A(n_611), .Y(n_876) );
OAI31xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_615), .A3(n_624), .B(n_625), .Y(n_612) );
NAND3xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .C(n_621), .Y(n_615) );
NAND3xp33_ASAP7_75t_SL g699 ( .A(n_616), .B(n_700), .C(n_704), .Y(n_699) );
NAND3xp33_ASAP7_75t_SL g765 ( .A(n_616), .B(n_766), .C(n_768), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_620), .A2(n_705), .B1(n_706), .B2(n_707), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_620), .A2(n_706), .B1(n_760), .B2(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g869 ( .A(n_620), .Y(n_869) );
AOI22xp33_ASAP7_75t_SL g951 ( .A1(n_620), .A2(n_706), .B1(n_944), .B2(n_952), .Y(n_951) );
AOI22xp33_ASAP7_75t_SL g986 ( .A1(n_620), .A2(n_706), .B1(n_979), .B2(n_987), .Y(n_986) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g690 ( .A(n_623), .Y(n_690) );
OAI31xp33_ASAP7_75t_SL g948 ( .A1(n_625), .A2(n_949), .A3(n_950), .B(n_953), .Y(n_948) );
OAI31xp33_ASAP7_75t_SL g983 ( .A1(n_625), .A2(n_984), .A3(n_985), .B(n_988), .Y(n_983) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_651), .Y(n_626) );
OAI33xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .A3(n_634), .B1(n_640), .B2(n_646), .B3(n_649), .Y(n_627) );
OAI33xp33_ASAP7_75t_L g790 ( .A1(n_628), .A2(n_649), .A3(n_791), .B1(n_794), .B2(n_797), .B3(n_799), .Y(n_790) );
OAI33xp33_ASAP7_75t_L g916 ( .A1(n_628), .A2(n_649), .A3(n_917), .B1(n_922), .B2(n_925), .B3(n_931), .Y(n_916) );
OAI33xp33_ASAP7_75t_L g970 ( .A1(n_628), .A2(n_649), .A3(n_971), .B1(n_972), .B2(n_973), .B3(n_975), .Y(n_970) );
BUFx3_ASAP7_75t_L g1105 ( .A(n_628), .Y(n_1105) );
OAI22xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B1(n_632), .B2(n_633), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_631), .A2(n_918), .B1(n_919), .B2(n_920), .Y(n_917) );
OAI22xp33_ASAP7_75t_L g971 ( .A1(n_633), .A2(n_792), .B1(n_959), .B2(n_965), .Y(n_971) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .B1(n_638), .B2(n_639), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_635), .A2(n_642), .B1(n_656), .B2(n_658), .Y(n_655) );
INVx3_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_SL g641 ( .A(n_637), .Y(n_641) );
INVx3_ASAP7_75t_L g1007 ( .A(n_637), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_638), .A2(n_645), .B1(n_664), .B2(n_666), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_639), .A2(n_926), .B1(n_927), .B2(n_930), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_643), .B2(n_645), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_643), .A2(n_1003), .B1(n_1004), .B2(n_1005), .Y(n_1002) );
OAI22xp5_ASAP7_75t_L g1006 ( .A1(n_643), .A2(n_1007), .B1(n_1008), .B2(n_1009), .Y(n_1006) );
BUFx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g1388 ( .A(n_644), .B(n_1389), .Y(n_1388) );
OAI33xp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .A3(n_655), .B1(n_660), .B2(n_661), .B3(n_663), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g773 ( .A1(n_653), .A2(n_774), .B1(n_775), .B2(n_777), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_653), .A2(n_787), .B1(n_788), .B2(n_789), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g935 ( .A1(n_653), .A2(n_775), .B1(n_918), .B2(n_932), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_653), .A2(n_666), .B1(n_924), .B2(n_930), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g958 ( .A1(n_653), .A2(n_788), .B1(n_959), .B2(n_960), .Y(n_958) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_653), .A2(n_775), .B1(n_968), .B2(n_969), .Y(n_967) );
OAI33xp33_ASAP7_75t_L g934 ( .A1(n_654), .A2(n_785), .A3(n_935), .B1(n_936), .B2(n_937), .B3(n_939), .Y(n_934) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g1492 ( .A(n_657), .Y(n_1492) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_658), .A2(n_780), .B1(n_923), .B2(n_926), .Y(n_936) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g815 ( .A(n_659), .Y(n_815) );
INVx1_ASAP7_75t_L g942 ( .A(n_659), .Y(n_942) );
INVx2_ASAP7_75t_L g1509 ( .A(n_659), .Y(n_1509) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AOI33xp33_ASAP7_75t_L g731 ( .A1(n_662), .A2(n_732), .A3(n_733), .B1(n_740), .B2(n_744), .B3(n_745), .Y(n_731) );
INVx2_ASAP7_75t_L g785 ( .A(n_662), .Y(n_785) );
AOI33xp33_ASAP7_75t_L g831 ( .A1(n_662), .A2(n_732), .A3(n_832), .B1(n_834), .B2(n_838), .B3(n_840), .Y(n_831) );
AOI33xp33_ASAP7_75t_L g1073 ( .A1(n_662), .A2(n_1074), .A3(n_1075), .B1(n_1077), .B2(n_1081), .B3(n_1083), .Y(n_1073) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g801 ( .A(n_669), .Y(n_801) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
XNOR2x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_754), .Y(n_670) );
OR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_727), .Y(n_671) );
INVx1_ASAP7_75t_L g729 ( .A(n_673), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_680), .B(n_688), .Y(n_673) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx8_ASAP7_75t_L g854 ( .A(n_677), .Y(n_854) );
INVx2_ASAP7_75t_L g1435 ( .A(n_677), .Y(n_1435) );
INVx8_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
BUFx3_ASAP7_75t_L g693 ( .A(n_678), .Y(n_693) );
BUFx3_ASAP7_75t_L g845 ( .A(n_678), .Y(n_845) );
NAND2x1p5_ASAP7_75t_L g1442 ( .A(n_678), .B(n_1443), .Y(n_1442) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_R g850 ( .A(n_682), .Y(n_850) );
INVx5_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
BUFx12f_ASAP7_75t_L g901 ( .A(n_683), .Y(n_901) );
INVx1_ASAP7_75t_L g1455 ( .A(n_684), .Y(n_1455) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI33xp33_ASAP7_75t_L g842 ( .A1(n_686), .A2(n_843), .A3(n_847), .B1(n_851), .B2(n_853), .B3(n_855), .Y(n_842) );
NAND3xp33_ASAP7_75t_L g898 ( .A(n_686), .B(n_899), .C(n_902), .Y(n_898) );
AOI33xp33_ASAP7_75t_L g1456 ( .A1(n_686), .A2(n_1457), .A3(n_1459), .B1(n_1460), .B2(n_1463), .B3(n_1465), .Y(n_1456) );
OAI221xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_691), .B1(n_692), .B2(n_694), .C(n_695), .Y(n_689) );
INVx2_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
AOI32xp33_ASAP7_75t_L g1086 ( .A1(n_695), .A2(n_1087), .A3(n_1090), .B1(n_1091), .B2(n_1092), .Y(n_1086) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g855 ( .A(n_696), .Y(n_855) );
OAI33xp33_ASAP7_75t_L g996 ( .A1(n_696), .A2(n_997), .A3(n_998), .B1(n_1002), .B2(n_1006), .B3(n_1010), .Y(n_996) );
INVx1_ASAP7_75t_SL g1465 ( .A(n_696), .Y(n_1465) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_697), .B(n_712), .Y(n_728) );
OAI31xp33_ASAP7_75t_SL g697 ( .A1(n_698), .A2(n_699), .A3(n_708), .B(n_711), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g846 ( .A(n_703), .Y(n_846) );
INVx2_ASAP7_75t_L g1464 ( .A(n_703), .Y(n_1464) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_706), .B(n_817), .Y(n_827) );
INVx1_ASAP7_75t_L g868 ( .A(n_706), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_706), .B(n_1062), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_707), .B(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g1068 ( .A1(n_710), .A2(n_829), .B1(n_1057), .B2(n_1058), .Y(n_1068) );
OAI31xp33_ASAP7_75t_SL g763 ( .A1(n_711), .A2(n_764), .A3(n_765), .B(n_770), .Y(n_763) );
INVx1_ASAP7_75t_L g830 ( .A(n_711), .Y(n_830) );
AO21x1_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_717), .B(n_726), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_722), .C(n_725), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_721), .A2(n_817), .B1(n_818), .B2(n_820), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g943 ( .A1(n_721), .A2(n_818), .B1(n_944), .B2(n_945), .Y(n_943) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g1060 ( .A(n_725), .B(n_1061), .C(n_1064), .Y(n_1060) );
AO21x1_ASAP7_75t_L g808 ( .A1(n_726), .A2(n_809), .B(n_813), .Y(n_808) );
AO21x1_ASAP7_75t_L g1055 ( .A1(n_726), .A2(n_1056), .B(n_1059), .Y(n_1055) );
OAI31xp33_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .A3(n_730), .B(n_751), .Y(n_727) );
INVx1_ASAP7_75t_L g753 ( .A(n_731), .Y(n_753) );
HB1xp67_ASAP7_75t_L g894 ( .A(n_732), .Y(n_894) );
INVx1_ASAP7_75t_L g1015 ( .A(n_732), .Y(n_1015) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g893 ( .A(n_735), .Y(n_893) );
INVx2_ASAP7_75t_SL g1076 ( .A(n_735), .Y(n_1076) );
INVx1_ASAP7_75t_L g1084 ( .A(n_735), .Y(n_1084) );
INVx3_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
BUFx6f_ASAP7_75t_L g748 ( .A(n_736), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_736), .B(n_1394), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1425 ( .A(n_736), .B(n_1406), .Y(n_1425) );
BUFx3_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g750 ( .A(n_739), .Y(n_750) );
BUFx6f_ASAP7_75t_L g1085 ( .A(n_739), .Y(n_1085) );
BUFx3_ASAP7_75t_L g1420 ( .A(n_739), .Y(n_1420) );
BUFx6f_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g836 ( .A(n_742), .Y(n_836) );
INVx2_ASAP7_75t_L g1079 ( .A(n_742), .Y(n_1079) );
AND2x4_ASAP7_75t_L g1427 ( .A(n_742), .B(n_1406), .Y(n_1427) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_SL g841 ( .A(n_747), .Y(n_841) );
INVx3_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
BUFx6f_ASAP7_75t_L g833 ( .A(n_748), .Y(n_833) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx3_ASAP7_75t_L g1414 ( .A(n_750), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
NAND3xp33_ASAP7_75t_SL g755 ( .A(n_756), .B(n_763), .C(n_771), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_761), .B(n_767), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_790), .Y(n_771) );
BUFx6f_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_779), .A2(n_787), .B1(n_795), .B2(n_796), .Y(n_794) );
OAI33xp33_ASAP7_75t_L g1014 ( .A1(n_785), .A2(n_1015), .A3(n_1016), .B1(n_1019), .B2(n_1020), .B3(n_1023), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_788), .A2(n_1005), .B1(n_1009), .B2(n_1017), .Y(n_1023) );
OAI22xp33_ASAP7_75t_L g1483 ( .A1(n_788), .A2(n_1484), .B1(n_1485), .B2(n_1486), .Y(n_1483) );
INVx2_ASAP7_75t_SL g792 ( .A(n_793), .Y(n_792) );
INVx3_ASAP7_75t_L g999 ( .A(n_793), .Y(n_999) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_805), .B1(n_910), .B2(n_989), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
XNOR2xp5_ASAP7_75t_L g805 ( .A(n_806), .B(n_858), .Y(n_805) );
INVx1_ASAP7_75t_L g856 ( .A(n_807), .Y(n_856) );
NAND4xp75_ASAP7_75t_L g807 ( .A(n_808), .B(n_822), .C(n_831), .D(n_842), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_811), .B(n_1161), .Y(n_1160) );
AND2x4_ASAP7_75t_SL g1471 ( .A(n_811), .B(n_1472), .Y(n_1471) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_814), .B(n_821), .Y(n_813) );
OAI22xp5_ASAP7_75t_SL g1019 ( .A1(n_815), .A2(n_938), .B1(n_1004), .B2(n_1008), .Y(n_1019) );
OAI22xp5_ASAP7_75t_L g1020 ( .A1(n_815), .A2(n_1001), .B1(n_1012), .B2(n_1021), .Y(n_1020) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
AO21x1_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_828), .B(n_830), .Y(n_822) );
INVx2_ASAP7_75t_SL g1127 ( .A(n_829), .Y(n_1127) );
AO21x1_ASAP7_75t_L g1067 ( .A1(n_830), .A2(n_1068), .B(n_1069), .Y(n_1067) );
INVx2_ASAP7_75t_SL g835 ( .A(n_836), .Y(n_835) );
BUFx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g909 ( .A(n_845), .Y(n_909) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
BUFx2_ASAP7_75t_L g1111 ( .A(n_854), .Y(n_1111) );
NAND3xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_864), .C(n_870), .Y(n_860) );
AOI22xp5_ASAP7_75t_L g1035 ( .A1(n_872), .A2(n_1036), .B1(n_1037), .B2(n_1038), .Y(n_1035) );
INVx2_ASAP7_75t_L g1133 ( .A(n_872), .Y(n_1133) );
NAND3xp33_ASAP7_75t_L g874 ( .A(n_875), .B(n_877), .C(n_883), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_878), .B(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx2_ASAP7_75t_L g1080 ( .A(n_879), .Y(n_1080) );
INVx1_ASAP7_75t_L g1082 ( .A(n_879), .Y(n_1082) );
NAND4xp25_ASAP7_75t_L g885 ( .A(n_886), .B(n_895), .C(n_898), .D(n_903), .Y(n_885) );
NAND3xp33_ASAP7_75t_L g886 ( .A(n_887), .B(n_892), .C(n_894), .Y(n_886) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx2_ASAP7_75t_SL g1107 ( .A(n_900), .Y(n_1107) );
NAND3xp33_ASAP7_75t_L g903 ( .A(n_904), .B(n_905), .C(n_907), .Y(n_903) );
BUFx2_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
BUFx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g989 ( .A(n_911), .Y(n_989) );
XNOR2x1_ASAP7_75t_L g911 ( .A(n_912), .B(n_954), .Y(n_911) );
XNOR2xp5_ASAP7_75t_L g912 ( .A(n_913), .B(n_914), .Y(n_912) );
AND3x1_ASAP7_75t_L g914 ( .A(n_915), .B(n_940), .C(n_948), .Y(n_914) );
NOR2xp33_ASAP7_75t_SL g915 ( .A(n_916), .B(n_934), .Y(n_915) );
OAI22xp33_ASAP7_75t_L g998 ( .A1(n_920), .A2(n_999), .B1(n_1000), .B2(n_1001), .Y(n_998) );
INVx3_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx2_ASAP7_75t_L g1506 ( .A(n_921), .Y(n_1506) );
INVx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx2_ASAP7_75t_L g1100 ( .A(n_928), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1437 ( .A(n_928), .B(n_1438), .Y(n_1437) );
INVx3_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
BUFx2_ASAP7_75t_L g1003 ( .A(n_929), .Y(n_1003) );
AND3x1_ASAP7_75t_L g955 ( .A(n_956), .B(n_976), .C(n_983), .Y(n_955) );
NOR2xp33_ASAP7_75t_L g956 ( .A(n_957), .B(n_970), .Y(n_956) );
INVx1_ASAP7_75t_L g1147 ( .A(n_990), .Y(n_1147) );
XNOR2xp5_ASAP7_75t_L g990 ( .A(n_991), .B(n_1050), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
HB1xp67_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
INVxp67_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
NOR4xp25_ASAP7_75t_L g1049 ( .A(n_996), .B(n_1014), .C(n_1025), .D(n_1041), .Y(n_1049) );
OAI22xp33_ASAP7_75t_L g1016 ( .A1(n_1000), .A2(n_1011), .B1(n_1017), .B2(n_1018), .Y(n_1016) );
INVxp67_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
OAI22xp33_ASAP7_75t_L g1135 ( .A1(n_1017), .A2(n_1136), .B1(n_1137), .B2(n_1138), .Y(n_1135) );
OAI22xp5_ASAP7_75t_L g1140 ( .A1(n_1021), .A2(n_1141), .B1(n_1142), .B2(n_1143), .Y(n_1140) );
INVx4_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVxp67_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
AOI31xp33_ASAP7_75t_L g1025 ( .A1(n_1026), .A2(n_1032), .A3(n_1035), .B(n_1039), .Y(n_1025) );
INVxp67_ASAP7_75t_SL g1027 ( .A(n_1028), .Y(n_1027) );
CKINVDCx14_ASAP7_75t_R g1039 ( .A(n_1040), .Y(n_1039) );
AOI31xp67_ASAP7_75t_SL g1041 ( .A1(n_1042), .A2(n_1044), .A3(n_1046), .B(n_1048), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
INVxp67_ASAP7_75t_SL g1046 ( .A(n_1047), .Y(n_1046) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_1051), .A2(n_1052), .B1(n_1093), .B2(n_1094), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
HB1xp67_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
NAND4xp75_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1067), .C(n_1073), .D(n_1086), .Y(n_1054) );
NOR2xp33_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1066), .Y(n_1059) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx2_ASAP7_75t_L g1417 ( .A(n_1079), .Y(n_1417) );
INVx2_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
NAND4xp75_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1113), .C(n_1125), .D(n_1134), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_1099), .A2(n_1105), .B1(n_1106), .B2(n_1112), .Y(n_1098) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
OAI22xp33_ASAP7_75t_L g1500 ( .A1(n_1129), .A2(n_1484), .B1(n_1493), .B2(n_1501), .Y(n_1500) );
INVx2_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
BUFx4f_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
INVx3_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
OR2x2_ASAP7_75t_L g1152 ( .A(n_1153), .B(n_1159), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
NOR2xp33_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1157), .Y(n_1154) );
NOR2xp33_ASAP7_75t_L g1476 ( .A(n_1155), .B(n_1158), .Y(n_1476) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1155), .Y(n_1526) );
HB1xp67_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
NOR2xp33_ASAP7_75t_L g1528 ( .A(n_1158), .B(n_1526), .Y(n_1528) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
OAI221xp5_ASAP7_75t_L g1162 ( .A1(n_1163), .A2(n_1376), .B1(n_1378), .B2(n_1468), .C(n_1473), .Y(n_1162) );
NOR3xp33_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1313), .C(n_1352), .Y(n_1163) );
NAND3xp33_ASAP7_75t_L g1164 ( .A(n_1165), .B(n_1248), .C(n_1280), .Y(n_1164) );
AOI211xp5_ASAP7_75t_L g1165 ( .A1(n_1166), .A2(n_1191), .B(n_1208), .C(n_1227), .Y(n_1165) );
NAND2xp5_ASAP7_75t_L g1225 ( .A(n_1166), .B(n_1226), .Y(n_1225) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1166), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1182), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1167), .B(n_1188), .Y(n_1296) );
NAND3xp33_ASAP7_75t_L g1300 ( .A(n_1167), .B(n_1286), .C(n_1301), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1167), .B(n_1217), .Y(n_1306) );
OR2x2_ASAP7_75t_L g1324 ( .A(n_1167), .B(n_1188), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1338 ( .A(n_1167), .B(n_1281), .Y(n_1338) );
CKINVDCx6p67_ASAP7_75t_R g1167 ( .A(n_1168), .Y(n_1167) );
OR2x2_ASAP7_75t_L g1215 ( .A(n_1168), .B(n_1188), .Y(n_1215) );
OR2x2_ASAP7_75t_L g1287 ( .A(n_1168), .B(n_1288), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1168), .B(n_1217), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1168), .B(n_1188), .Y(n_1317) );
CKINVDCx5p33_ASAP7_75t_R g1340 ( .A(n_1168), .Y(n_1340) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1168), .B(n_1242), .Y(n_1345) );
OR2x6_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1176), .Y(n_1168) );
OR2x2_ASAP7_75t_L g1329 ( .A(n_1169), .B(n_1176), .Y(n_1329) );
INVx2_ASAP7_75t_L g1245 ( .A(n_1170), .Y(n_1245) );
AND2x6_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1172), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1171), .B(n_1175), .Y(n_1174) );
AND2x4_ASAP7_75t_L g1177 ( .A(n_1171), .B(n_1178), .Y(n_1177) );
AND2x6_ASAP7_75t_L g1180 ( .A(n_1171), .B(n_1181), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1171), .B(n_1175), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1171), .B(n_1175), .Y(n_1196) );
OAI21xp5_ASAP7_75t_L g1525 ( .A1(n_1172), .A2(n_1526), .B(n_1527), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1173), .B(n_1179), .Y(n_1178) );
AOI21xp33_ASAP7_75t_L g1265 ( .A1(n_1182), .A2(n_1241), .B(n_1266), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1364 ( .A(n_1182), .B(n_1212), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1187), .Y(n_1182) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1183), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1183), .B(n_1188), .Y(n_1229) );
OR2x2_ASAP7_75t_L g1279 ( .A(n_1183), .B(n_1188), .Y(n_1279) );
OR2x2_ASAP7_75t_L g1302 ( .A(n_1183), .B(n_1198), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1184), .B(n_1186), .Y(n_1183) );
INVxp67_ASAP7_75t_L g1247 ( .A(n_1185), .Y(n_1247) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
OAI221xp5_ASAP7_75t_L g1208 ( .A1(n_1188), .A2(n_1209), .B1(n_1213), .B2(n_1219), .C(n_1225), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1188), .B(n_1218), .Y(n_1240) );
A2O1A1Ixp33_ASAP7_75t_L g1248 ( .A1(n_1188), .A2(n_1249), .B(n_1263), .C(n_1264), .Y(n_1248) );
INVx3_ASAP7_75t_L g1309 ( .A(n_1188), .Y(n_1309) );
O2A1O1Ixp33_ASAP7_75t_L g1353 ( .A1(n_1188), .A2(n_1354), .B(n_1355), .C(n_1356), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1367 ( .A(n_1188), .B(n_1198), .Y(n_1367) );
AND2x4_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1190), .Y(n_1188) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
AOI21xp5_ASAP7_75t_L g1356 ( .A1(n_1192), .A2(n_1279), .B(n_1357), .Y(n_1356) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1197), .Y(n_1192) );
INVx2_ASAP7_75t_L g1210 ( .A(n_1193), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1193), .B(n_1222), .Y(n_1226) );
BUFx2_ASAP7_75t_L g1254 ( .A(n_1193), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1193), .B(n_1201), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1193), .B(n_1268), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1194), .B(n_1195), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1201), .Y(n_1197) );
INVx2_ASAP7_75t_L g1212 ( .A(n_1198), .Y(n_1212) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1198), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1198), .B(n_1254), .Y(n_1261) );
OR2x2_ASAP7_75t_L g1271 ( .A(n_1198), .B(n_1272), .Y(n_1271) );
NOR2xp33_ASAP7_75t_L g1321 ( .A(n_1198), .B(n_1322), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1328 ( .A(n_1198), .B(n_1222), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1199), .B(n_1200), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1201), .B(n_1212), .Y(n_1211) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1201), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1342 ( .A(n_1201), .B(n_1343), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1201), .B(n_1261), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1202), .B(n_1205), .Y(n_1201) );
INVx2_ASAP7_75t_L g1223 ( .A(n_1202), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1202), .B(n_1224), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1272 ( .A(n_1202), .B(n_1254), .Y(n_1272) );
OR2x2_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1204), .Y(n_1202) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1205), .Y(n_1224) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1205), .B(n_1210), .Y(n_1233) );
OR2x2_ASAP7_75t_L g1253 ( .A(n_1205), .B(n_1254), .Y(n_1253) );
AND3x1_ASAP7_75t_L g1257 ( .A(n_1205), .B(n_1210), .C(n_1223), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1205), .B(n_1254), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1205), .B(n_1223), .Y(n_1286) );
OAI21xp33_ASAP7_75t_L g1318 ( .A1(n_1205), .A2(n_1319), .B(n_1320), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1207), .Y(n_1205) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_1210), .B(n_1211), .Y(n_1209) );
OR2x2_ASAP7_75t_L g1219 ( .A(n_1210), .B(n_1220), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1210), .B(n_1222), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1210), .B(n_1268), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1210), .B(n_1223), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1210), .B(n_1212), .Y(n_1343) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1212), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_1212), .B(n_1268), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1212), .B(n_1275), .Y(n_1274) );
NOR2xp33_ASAP7_75t_L g1294 ( .A(n_1212), .B(n_1272), .Y(n_1294) );
O2A1O1Ixp33_ASAP7_75t_L g1303 ( .A1(n_1212), .A2(n_1236), .B(n_1304), .C(n_1305), .Y(n_1303) );
NOR2xp33_ASAP7_75t_L g1312 ( .A(n_1212), .B(n_1253), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_1212), .B(n_1217), .Y(n_1327) );
NOR2xp33_ASAP7_75t_L g1213 ( .A(n_1214), .B(n_1216), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
OAI21xp33_ASAP7_75t_L g1297 ( .A1(n_1215), .A2(n_1298), .B(n_1300), .Y(n_1297) );
OAI222xp33_ASAP7_75t_L g1346 ( .A1(n_1215), .A2(n_1305), .B1(n_1347), .B2(n_1348), .C1(n_1349), .C2(n_1351), .Y(n_1346) );
OAI211xp5_ASAP7_75t_L g1249 ( .A1(n_1216), .A2(n_1250), .B(n_1255), .C(n_1258), .Y(n_1249) );
INVx2_ASAP7_75t_L g1311 ( .A(n_1216), .Y(n_1311) );
O2A1O1Ixp33_ASAP7_75t_L g1332 ( .A1(n_1216), .A2(n_1273), .B(n_1299), .C(n_1333), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1374 ( .A(n_1216), .B(n_1375), .Y(n_1374) );
INVx2_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1217), .B(n_1259), .Y(n_1258) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
OAI211xp5_ASAP7_75t_SL g1323 ( .A1(n_1219), .A2(n_1281), .B(n_1324), .C(n_1325), .Y(n_1323) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1220), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_1221), .B(n_1222), .Y(n_1220) );
INVx2_ASAP7_75t_L g1252 ( .A(n_1221), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1221), .B(n_1278), .Y(n_1277) );
NAND2xp5_ASAP7_75t_SL g1319 ( .A(n_1221), .B(n_1229), .Y(n_1319) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1222), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_1222), .B(n_1277), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1222), .B(n_1343), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1223), .B(n_1224), .Y(n_1222) );
OR2x2_ASAP7_75t_L g1322 ( .A(n_1223), .B(n_1254), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1223), .B(n_1254), .Y(n_1350) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1226), .Y(n_1351) );
O2A1O1Ixp33_ASAP7_75t_SL g1227 ( .A1(n_1228), .A2(n_1230), .B(n_1234), .C(n_1241), .Y(n_1227) );
INVx2_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
OAI21xp5_ASAP7_75t_SL g1334 ( .A1(n_1229), .A2(n_1335), .B(n_1336), .Y(n_1334) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
NOR2xp33_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1233), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1232), .B(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
AOI21xp33_ASAP7_75t_L g1235 ( .A1(n_1236), .A2(n_1238), .B(n_1239), .Y(n_1235) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
AOI221xp5_ASAP7_75t_L g1325 ( .A1(n_1238), .A2(n_1261), .B1(n_1286), .B2(n_1326), .C(n_1328), .Y(n_1325) );
AOI21xp33_ASAP7_75t_L g1333 ( .A1(n_1238), .A2(n_1239), .B(n_1304), .Y(n_1333) );
OAI21xp5_ASAP7_75t_L g1269 ( .A1(n_1240), .A2(n_1270), .B(n_1273), .Y(n_1269) );
CKINVDCx6p67_ASAP7_75t_R g1288 ( .A(n_1240), .Y(n_1288) );
INVx3_ASAP7_75t_L g1263 ( .A(n_1241), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1241), .B(n_1309), .Y(n_1308) );
INVx2_ASAP7_75t_SL g1241 ( .A(n_1242), .Y(n_1241) );
INVx2_ASAP7_75t_SL g1281 ( .A(n_1242), .Y(n_1281) );
OAI22xp5_ASAP7_75t_SL g1243 ( .A1(n_1244), .A2(n_1245), .B1(n_1246), .B2(n_1247), .Y(n_1243) );
CKINVDCx20_ASAP7_75t_R g1377 ( .A(n_1245), .Y(n_1377) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
NOR2xp33_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1253), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1252), .B(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1252), .Y(n_1292) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
A2O1A1Ixp33_ASAP7_75t_L g1365 ( .A1(n_1256), .A2(n_1309), .B(n_1344), .C(n_1366), .Y(n_1365) );
AND2x2_ASAP7_75t_SL g1373 ( .A(n_1257), .B(n_1278), .Y(n_1373) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1258), .Y(n_1354) );
OR2x2_ASAP7_75t_L g1259 ( .A(n_1260), .B(n_1262), .Y(n_1259) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1261), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1261), .B(n_1268), .Y(n_1335) );
O2A1O1Ixp33_ASAP7_75t_L g1341 ( .A1(n_1263), .A2(n_1278), .B(n_1342), .C(n_1344), .Y(n_1341) );
NAND3xp33_ASAP7_75t_L g1264 ( .A(n_1265), .B(n_1269), .C(n_1276), .Y(n_1264) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
OAI211xp5_ASAP7_75t_L g1331 ( .A1(n_1271), .A2(n_1288), .B(n_1332), .C(n_1334), .Y(n_1331) );
AOI211xp5_ASAP7_75t_L g1295 ( .A1(n_1273), .A2(n_1296), .B(n_1297), .C(n_1303), .Y(n_1295) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1275), .Y(n_1371) );
OAI21xp5_ASAP7_75t_L g1289 ( .A1(n_1278), .A2(n_1290), .B(n_1294), .Y(n_1289) );
INVx2_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
AOI22xp5_ASAP7_75t_L g1280 ( .A1(n_1281), .A2(n_1282), .B1(n_1307), .B2(n_1310), .Y(n_1280) );
NAND3xp33_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1289), .C(n_1295), .Y(n_1282) );
INVxp67_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
NOR2xp33_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1287), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
AOI211xp5_ASAP7_75t_L g1359 ( .A1(n_1290), .A2(n_1309), .B(n_1360), .C(n_1362), .Y(n_1359) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1293), .Y(n_1291) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1293), .B(n_1326), .Y(n_1361) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1293), .Y(n_1370) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
INVxp33_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1311), .B(n_1312), .Y(n_1310) );
AOI21xp5_ASAP7_75t_L g1372 ( .A1(n_1311), .A2(n_1355), .B(n_1373), .Y(n_1372) );
AOI221xp5_ASAP7_75t_SL g1313 ( .A1(n_1314), .A2(n_1329), .B1(n_1330), .B2(n_1337), .C(n_1339), .Y(n_1313) );
O2A1O1Ixp33_ASAP7_75t_L g1314 ( .A1(n_1315), .A2(n_1317), .B(n_1318), .C(n_1323), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
INVxp67_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
AOI211xp5_ASAP7_75t_L g1339 ( .A1(n_1331), .A2(n_1340), .B(n_1341), .C(n_1346), .Y(n_1339) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1335), .Y(n_1347) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
A2O1A1Ixp33_ASAP7_75t_L g1352 ( .A1(n_1340), .A2(n_1353), .B(n_1359), .C(n_1365), .Y(n_1352) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
CKINVDCx14_ASAP7_75t_R g1349 ( .A(n_1350), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1350), .B(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
INVxp67_ASAP7_75t_SL g1362 ( .A(n_1363), .Y(n_1362) );
OAI211xp5_ASAP7_75t_SL g1366 ( .A1(n_1367), .A2(n_1368), .B(n_1372), .C(n_1374), .Y(n_1366) );
INVxp67_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
NAND2xp5_ASAP7_75t_SL g1369 ( .A(n_1370), .B(n_1371), .Y(n_1369) );
CKINVDCx20_ASAP7_75t_R g1376 ( .A(n_1377), .Y(n_1376) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
HB1xp67_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
NAND3xp33_ASAP7_75t_L g1383 ( .A(n_1384), .B(n_1395), .C(n_1439), .Y(n_1383) );
NAND2xp5_ASAP7_75t_L g1384 ( .A(n_1385), .B(n_1386), .Y(n_1384) );
INVx8_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
AND2x4_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1391), .Y(n_1387) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1389), .Y(n_1436) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1389), .Y(n_1438) );
OR2x2_ASAP7_75t_L g1391 ( .A(n_1392), .B(n_1393), .Y(n_1391) );
AND2x4_ASAP7_75t_L g1449 ( .A(n_1392), .B(n_1443), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1394), .B(n_1402), .Y(n_1401) );
AOI21xp5_ASAP7_75t_L g1395 ( .A1(n_1396), .A2(n_1399), .B(n_1428), .Y(n_1395) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
BUFx2_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
NAND3xp33_ASAP7_75t_L g1399 ( .A(n_1400), .B(n_1412), .C(n_1422), .Y(n_1399) );
AOI222xp33_ASAP7_75t_L g1400 ( .A1(n_1401), .A2(n_1403), .B1(n_1404), .B2(n_1407), .C1(n_1408), .C2(n_1411), .Y(n_1400) );
AOI22xp33_ASAP7_75t_L g1447 ( .A1(n_1403), .A2(n_1407), .B1(n_1448), .B2(n_1452), .Y(n_1447) );
BUFx3_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1406), .B(n_1414), .Y(n_1413) );
INVx3_ASAP7_75t_L g1409 ( .A(n_1410), .Y(n_1409) );
AOI221xp5_ASAP7_75t_L g1412 ( .A1(n_1413), .A2(n_1415), .B1(n_1416), .B2(n_1419), .C(n_1421), .Y(n_1412) );
AOI211xp5_ASAP7_75t_L g1439 ( .A1(n_1415), .A2(n_1440), .B(n_1446), .C(n_1466), .Y(n_1439) );
AOI22xp33_ASAP7_75t_L g1422 ( .A1(n_1423), .A2(n_1424), .B1(n_1426), .B2(n_1427), .Y(n_1422) );
AOI22xp33_ASAP7_75t_L g1433 ( .A1(n_1423), .A2(n_1426), .B1(n_1434), .B2(n_1437), .Y(n_1433) );
BUFx6f_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
AND2x4_ASAP7_75t_L g1429 ( .A(n_1430), .B(n_1431), .Y(n_1429) );
AND2x4_ASAP7_75t_L g1434 ( .A(n_1435), .B(n_1436), .Y(n_1434) );
INVx3_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
OR2x6_ASAP7_75t_L g1441 ( .A(n_1442), .B(n_1445), .Y(n_1441) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_1447), .B(n_1456), .Y(n_1446) );
AND2x4_ASAP7_75t_SL g1448 ( .A(n_1449), .B(n_1450), .Y(n_1448) );
AND2x4_ASAP7_75t_SL g1452 ( .A(n_1449), .B(n_1453), .Y(n_1452) );
AND2x4_ASAP7_75t_L g1466 ( .A(n_1449), .B(n_1458), .Y(n_1466) );
INVx3_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
INVx2_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
CKINVDCx20_ASAP7_75t_R g1468 ( .A(n_1469), .Y(n_1468) );
CKINVDCx20_ASAP7_75t_R g1469 ( .A(n_1470), .Y(n_1469) );
INVx3_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
HB1xp67_ASAP7_75t_SL g1474 ( .A(n_1475), .Y(n_1474) );
BUFx3_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
INVxp33_ASAP7_75t_SL g1477 ( .A(n_1478), .Y(n_1477) );
HB1xp67_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
NAND3xp33_ASAP7_75t_L g1480 ( .A(n_1481), .B(n_1507), .C(n_1516), .Y(n_1480) );
NOR2xp33_ASAP7_75t_L g1481 ( .A(n_1482), .B(n_1499), .Y(n_1481) );
OAI22xp33_ASAP7_75t_L g1505 ( .A1(n_1486), .A2(n_1494), .B1(n_1501), .B2(n_1506), .Y(n_1505) );
INVx2_ASAP7_75t_L g1501 ( .A(n_1502), .Y(n_1501) );
HB1xp67_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
endmodule