module fake_netlist_1_6183_n_652 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_652);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_652;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_73;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g72 ( .A(n_55), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_25), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_35), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_30), .Y(n_75) );
INVxp67_ASAP7_75t_SL g76 ( .A(n_70), .Y(n_76) );
INVx2_ASAP7_75t_L g77 ( .A(n_0), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_49), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_0), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_45), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_22), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_52), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_53), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_20), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_56), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_19), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_43), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_71), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_31), .Y(n_89) );
NAND2xp5_ASAP7_75t_L g90 ( .A(n_50), .B(n_44), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_65), .Y(n_91) );
HB1xp67_ASAP7_75t_L g92 ( .A(n_42), .Y(n_92) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_66), .Y(n_93) );
HB1xp67_ASAP7_75t_L g94 ( .A(n_58), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_4), .Y(n_95) );
BUFx3_ASAP7_75t_L g96 ( .A(n_9), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_27), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_4), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_62), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_59), .Y(n_100) );
INVxp33_ASAP7_75t_SL g101 ( .A(n_11), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_38), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_26), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_9), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_3), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_1), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_37), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_11), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_3), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_17), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_67), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_54), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_81), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_111), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_72), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_72), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_81), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_74), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_74), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_75), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_78), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_79), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_78), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_80), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_111), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_80), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_86), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_82), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_82), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_85), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_96), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_111), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_88), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_87), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_92), .B(n_2), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_96), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_94), .B(n_5), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_88), .Y(n_141) );
INVxp67_ASAP7_75t_SL g142 ( .A(n_77), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_111), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_86), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_100), .B(n_5), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_87), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_99), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_99), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_95), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_100), .Y(n_150) );
NAND2xp33_ASAP7_75t_L g151 ( .A(n_112), .B(n_34), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_142), .B(n_97), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_114), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_115), .B(n_77), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_133), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_114), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_138), .B(n_98), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_133), .Y(n_158) );
BUFx2_ASAP7_75t_L g159 ( .A(n_149), .Y(n_159) );
BUFx2_ASAP7_75t_L g160 ( .A(n_137), .Y(n_160) );
INVx4_ASAP7_75t_L g161 ( .A(n_133), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_133), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_139), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_114), .Y(n_164) );
OR2x2_ASAP7_75t_L g165 ( .A(n_146), .B(n_98), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_139), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_114), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_116), .B(n_106), .Y(n_168) );
INVx4_ASAP7_75t_L g169 ( .A(n_139), .Y(n_169) );
BUFx2_ASAP7_75t_L g170 ( .A(n_147), .Y(n_170) );
OR2x6_ASAP7_75t_L g171 ( .A(n_138), .B(n_110), .Y(n_171) );
INVxp67_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_116), .B(n_109), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_139), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_114), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_118), .B(n_108), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_118), .B(n_93), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_114), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_113), .Y(n_179) );
INVx4_ASAP7_75t_L g180 ( .A(n_119), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_113), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_117), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_117), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_119), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_120), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_125), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_120), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_129), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_129), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_121), .B(n_91), .Y(n_190) );
INVxp67_ASAP7_75t_SL g191 ( .A(n_123), .Y(n_191) );
AND2x6_ASAP7_75t_L g192 ( .A(n_123), .B(n_112), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_125), .Y(n_193) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_127), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_135), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_124), .Y(n_196) );
OR2x2_ASAP7_75t_SL g197 ( .A(n_140), .B(n_105), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_125), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_135), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_124), .Y(n_200) );
INVx5_ASAP7_75t_L g201 ( .A(n_125), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_125), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_125), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_144), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_126), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_141), .Y(n_206) );
OR2x2_ASAP7_75t_L g207 ( .A(n_126), .B(n_104), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_128), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_134), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_141), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_128), .B(n_102), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_130), .B(n_103), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_184), .Y(n_213) );
BUFx4f_ASAP7_75t_SL g214 ( .A(n_159), .Y(n_214) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_159), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_191), .B(n_136), .Y(n_216) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_160), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_171), .B(n_136), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_155), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_184), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_177), .B(n_130), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_155), .Y(n_222) );
BUFx8_ASAP7_75t_L g223 ( .A(n_160), .Y(n_223) );
INVx2_ASAP7_75t_SL g224 ( .A(n_196), .Y(n_224) );
BUFx3_ASAP7_75t_L g225 ( .A(n_196), .Y(n_225) );
OR2x6_ASAP7_75t_L g226 ( .A(n_171), .B(n_170), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_205), .B(n_131), .Y(n_227) );
NOR2xp33_ASAP7_75t_R g228 ( .A(n_204), .B(n_122), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_200), .A2(n_151), .B(n_150), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_171), .B(n_150), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_205), .B(n_131), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_185), .Y(n_232) );
OR2x6_ASAP7_75t_L g233 ( .A(n_171), .B(n_145), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_170), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_172), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_200), .B(n_132), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_185), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_165), .B(n_132), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_168), .A2(n_102), .B(n_107), .C(n_73), .Y(n_239) );
INVxp67_ASAP7_75t_L g240 ( .A(n_194), .Y(n_240) );
AND2x6_ASAP7_75t_SL g241 ( .A(n_157), .B(n_107), .Y(n_241) );
OR2x2_ASAP7_75t_L g242 ( .A(n_165), .B(n_6), .Y(n_242) );
INVxp67_ASAP7_75t_L g243 ( .A(n_157), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_208), .A2(n_101), .B1(n_89), .B2(n_84), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_187), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_192), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_155), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_168), .B(n_76), .Y(n_248) );
INVx4_ASAP7_75t_L g249 ( .A(n_180), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_158), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_192), .Y(n_251) );
INVx4_ASAP7_75t_L g252 ( .A(n_180), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_168), .B(n_90), .Y(n_253) );
BUFx2_ASAP7_75t_L g254 ( .A(n_192), .Y(n_254) );
NOR2xp33_ASAP7_75t_SL g255 ( .A(n_192), .B(n_143), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_187), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_158), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_168), .B(n_143), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_188), .Y(n_259) );
BUFx10_ASAP7_75t_L g260 ( .A(n_192), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_211), .A2(n_134), .B1(n_143), .B2(n_8), .Y(n_261) );
NOR2xp33_ASAP7_75t_R g262 ( .A(n_192), .B(n_6), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_173), .B(n_143), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_176), .B(n_7), .Y(n_264) );
NOR2xp33_ASAP7_75t_SL g265 ( .A(n_192), .B(n_143), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_162), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_211), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_162), .Y(n_268) );
NOR3xp33_ASAP7_75t_SL g269 ( .A(n_152), .B(n_7), .C(n_8), .Y(n_269) );
NOR2xp33_ASAP7_75t_R g270 ( .A(n_207), .B(n_10), .Y(n_270) );
INVxp67_ASAP7_75t_L g271 ( .A(n_176), .Y(n_271) );
INVx2_ASAP7_75t_SL g272 ( .A(n_173), .Y(n_272) );
OR2x2_ASAP7_75t_L g273 ( .A(n_197), .B(n_10), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_188), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_161), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_189), .Y(n_276) );
INVx6_ASAP7_75t_L g277 ( .A(n_180), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_163), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_173), .B(n_211), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_246), .Y(n_280) );
INVx4_ASAP7_75t_L g281 ( .A(n_226), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_218), .A2(n_211), .B1(n_173), .B2(n_154), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_249), .Y(n_283) );
BUFx4f_ASAP7_75t_L g284 ( .A(n_226), .Y(n_284) );
INVx5_ASAP7_75t_L g285 ( .A(n_249), .Y(n_285) );
NAND2x1p5_ASAP7_75t_L g286 ( .A(n_218), .B(n_154), .Y(n_286) );
OAI21xp33_ASAP7_75t_SL g287 ( .A1(n_279), .A2(n_212), .B(n_190), .Y(n_287) );
INVx2_ASAP7_75t_SL g288 ( .A(n_214), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_L g289 ( .A1(n_243), .A2(n_210), .B(n_189), .C(n_206), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_218), .Y(n_290) );
INVx4_ASAP7_75t_L g291 ( .A(n_226), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_230), .B(n_154), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_264), .Y(n_293) );
BUFx3_ASAP7_75t_L g294 ( .A(n_277), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_267), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_271), .B(n_154), .Y(n_296) );
INVx2_ASAP7_75t_SL g297 ( .A(n_214), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_250), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_260), .B(n_161), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_223), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_215), .Y(n_301) );
AOI22xp33_ASAP7_75t_SL g302 ( .A1(n_270), .A2(n_182), .B1(n_179), .B2(n_181), .Y(n_302) );
INVx3_ASAP7_75t_L g303 ( .A(n_249), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_272), .B(n_163), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_238), .B(n_169), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_267), .B(n_169), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_252), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_272), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_244), .A2(n_166), .B1(n_174), .B2(n_206), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_221), .A2(n_210), .B1(n_195), .B2(n_199), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_217), .B(n_181), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_277), .Y(n_312) );
INVx5_ASAP7_75t_L g313 ( .A(n_252), .Y(n_313) );
INVxp67_ASAP7_75t_L g314 ( .A(n_234), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_216), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_213), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_235), .B(n_182), .Y(n_317) );
INVx4_ASAP7_75t_SL g318 ( .A(n_246), .Y(n_318) );
NOR3xp33_ASAP7_75t_L g319 ( .A(n_240), .B(n_199), .C(n_195), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_251), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_220), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_236), .A2(n_166), .B(n_174), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_223), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_252), .B(n_179), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_248), .B(n_183), .Y(n_325) );
OAI21x1_ASAP7_75t_L g326 ( .A1(n_229), .A2(n_183), .B(n_203), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_253), .A2(n_209), .B(n_203), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_224), .A2(n_209), .B(n_202), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g329 ( .A1(n_242), .A2(n_197), .B1(n_134), .B2(n_143), .C(n_175), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_250), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_251), .B(n_12), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_232), .A2(n_134), .B1(n_202), .B2(n_167), .Y(n_332) );
OR2x6_ASAP7_75t_L g333 ( .A(n_281), .B(n_254), .Y(n_333) );
INVx6_ASAP7_75t_L g334 ( .A(n_285), .Y(n_334) );
OAI21xp5_ASAP7_75t_L g335 ( .A1(n_287), .A2(n_239), .B(n_257), .Y(n_335) );
OAI211xp5_ASAP7_75t_L g336 ( .A1(n_302), .A2(n_270), .B(n_269), .C(n_273), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_314), .B(n_241), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_298), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_298), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_286), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_285), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_315), .B(n_237), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_330), .Y(n_343) );
INVx4_ASAP7_75t_L g344 ( .A(n_285), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_319), .A2(n_223), .B1(n_233), .B2(n_277), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_330), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_316), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_302), .A2(n_239), .B1(n_276), .B2(n_259), .Y(n_348) );
AO31x2_ASAP7_75t_L g349 ( .A1(n_321), .A2(n_245), .A3(n_274), .B(n_256), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_319), .A2(n_233), .B1(n_278), .B2(n_228), .Y(n_350) );
AND2x4_ASAP7_75t_SL g351 ( .A(n_281), .B(n_260), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_286), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_282), .B(n_275), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_282), .B(n_227), .Y(n_354) );
INVxp67_ASAP7_75t_SL g355 ( .A(n_284), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_300), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_291), .B(n_275), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_285), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_292), .B(n_275), .Y(n_359) );
AO21x2_ASAP7_75t_L g360 ( .A1(n_326), .A2(n_262), .B(n_263), .Y(n_360) );
INVx4_ASAP7_75t_L g361 ( .A(n_313), .Y(n_361) );
NAND2xp33_ASAP7_75t_R g362 ( .A(n_323), .B(n_228), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_292), .A2(n_278), .B1(n_247), .B2(n_225), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_304), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_310), .A2(n_231), .B1(n_224), .B2(n_261), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_301), .Y(n_366) );
OAI322xp33_ASAP7_75t_L g367 ( .A1(n_337), .A2(n_293), .A3(n_314), .B1(n_309), .B2(n_291), .C1(n_300), .C2(n_295), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_342), .B(n_317), .Y(n_368) );
INVx2_ASAP7_75t_SL g369 ( .A(n_334), .Y(n_369) );
A2O1A1Ixp33_ASAP7_75t_L g370 ( .A1(n_335), .A2(n_289), .B(n_284), .C(n_310), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_338), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_338), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_339), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_342), .B(n_311), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_339), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_366), .A2(n_296), .B1(n_331), .B2(n_290), .Y(n_376) );
OAI22xp33_ASAP7_75t_L g377 ( .A1(n_366), .A2(n_297), .B1(n_288), .B2(n_305), .Y(n_377) );
OAI22xp33_ASAP7_75t_L g378 ( .A1(n_362), .A2(n_306), .B1(n_331), .B2(n_313), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_354), .A2(n_329), .B1(n_324), .B2(n_325), .Y(n_379) );
OA21x2_ASAP7_75t_L g380 ( .A1(n_335), .A2(n_327), .B(n_328), .Y(n_380) );
OAI221xp5_ASAP7_75t_L g381 ( .A1(n_345), .A2(n_308), .B1(n_247), .B2(n_283), .C(n_303), .Y(n_381) );
OA21x2_ASAP7_75t_L g382 ( .A1(n_348), .A2(n_332), .B(n_322), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_353), .A2(n_262), .B1(n_304), .B2(n_283), .Y(n_383) );
INVx2_ASAP7_75t_SL g384 ( .A(n_334), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_343), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_353), .A2(n_304), .B1(n_303), .B2(n_307), .Y(n_386) );
BUFx10_ASAP7_75t_L g387 ( .A(n_334), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_353), .A2(n_307), .B1(n_247), .B2(n_313), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_346), .B(n_313), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_346), .B(n_268), .Y(n_390) );
OR2x6_ASAP7_75t_L g391 ( .A(n_333), .B(n_280), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_350), .A2(n_312), .B1(n_294), .B2(n_225), .Y(n_392) );
OAI22xp33_ASAP7_75t_L g393 ( .A1(n_355), .A2(n_294), .B1(n_312), .B2(n_280), .Y(n_393) );
AOI222xp33_ASAP7_75t_L g394 ( .A1(n_347), .A2(n_318), .B1(n_266), .B2(n_257), .C1(n_268), .C2(n_219), .Y(n_394) );
AOI22xp33_ASAP7_75t_SL g395 ( .A1(n_374), .A2(n_336), .B1(n_340), .B2(n_352), .Y(n_395) );
INVx4_ASAP7_75t_L g396 ( .A(n_391), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_371), .Y(n_397) );
OAI21x1_ASAP7_75t_L g398 ( .A1(n_380), .A2(n_343), .B(n_341), .Y(n_398) );
AOI211xp5_ASAP7_75t_L g399 ( .A1(n_367), .A2(n_336), .B(n_340), .C(n_352), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_371), .B(n_343), .Y(n_400) );
OAI31xp33_ASAP7_75t_L g401 ( .A1(n_370), .A2(n_365), .A3(n_359), .B(n_347), .Y(n_401) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_367), .A2(n_359), .B1(n_356), .B2(n_365), .C(n_357), .Y(n_402) );
OAI211xp5_ASAP7_75t_L g403 ( .A1(n_368), .A2(n_376), .B(n_374), .C(n_392), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_372), .B(n_349), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_385), .Y(n_405) );
OAI33xp33_ASAP7_75t_L g406 ( .A1(n_377), .A2(n_372), .A3(n_373), .B1(n_375), .B2(n_378), .B3(n_379), .Y(n_406) );
NAND2x1p5_ASAP7_75t_L g407 ( .A(n_389), .B(n_344), .Y(n_407) );
OAI33xp33_ASAP7_75t_L g408 ( .A1(n_373), .A2(n_258), .A3(n_364), .B1(n_156), .B2(n_167), .B3(n_153), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_385), .Y(n_409) );
OAI211xp5_ASAP7_75t_SL g410 ( .A1(n_388), .A2(n_363), .B(n_358), .C(n_341), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_385), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_389), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_375), .Y(n_413) );
AO21x2_ASAP7_75t_L g414 ( .A1(n_393), .A2(n_360), .B(n_364), .Y(n_414) );
BUFx2_ASAP7_75t_L g415 ( .A(n_391), .Y(n_415) );
OAI21x1_ASAP7_75t_L g416 ( .A1(n_380), .A2(n_341), .B(n_358), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_390), .B(n_349), .Y(n_417) );
AOI31xp33_ASAP7_75t_L g418 ( .A1(n_383), .A2(n_357), .A3(n_361), .B(n_344), .Y(n_418) );
OR2x6_ASAP7_75t_L g419 ( .A(n_391), .B(n_361), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_390), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_380), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_387), .B(n_349), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_386), .A2(n_357), .B1(n_358), .B2(n_341), .C(n_344), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_381), .A2(n_358), .B1(n_344), .B2(n_361), .C(n_219), .Y(n_424) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_387), .A2(n_334), .B1(n_361), .B2(n_333), .Y(n_425) );
INVxp67_ASAP7_75t_L g426 ( .A(n_394), .Y(n_426) );
OAI31xp33_ASAP7_75t_SL g427 ( .A1(n_394), .A2(n_349), .A3(n_360), .B(n_334), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_369), .A2(n_222), .B1(n_266), .B2(n_332), .C(n_360), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_417), .B(n_349), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_397), .Y(n_430) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_401), .A2(n_333), .B1(n_391), .B2(n_384), .C(n_369), .Y(n_431) );
AND2x4_ASAP7_75t_L g432 ( .A(n_396), .B(n_391), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_417), .B(n_349), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_404), .B(n_349), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_404), .B(n_382), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_421), .Y(n_436) );
INVx3_ASAP7_75t_L g437 ( .A(n_416), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_396), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_422), .B(n_382), .Y(n_439) );
INVx2_ASAP7_75t_SL g440 ( .A(n_419), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_422), .B(n_382), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_397), .B(n_384), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_400), .B(n_382), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_400), .B(n_360), .Y(n_444) );
INVx5_ASAP7_75t_L g445 ( .A(n_419), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_413), .B(n_380), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_421), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_396), .B(n_61), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_396), .B(n_63), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_403), .B(n_333), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_413), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_405), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_405), .B(n_387), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_405), .Y(n_454) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_409), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_409), .B(n_387), .Y(n_456) );
OAI31xp33_ASAP7_75t_L g457 ( .A1(n_401), .A2(n_351), .A3(n_222), .B(n_15), .Y(n_457) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_399), .B(n_134), .C(n_198), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_411), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_411), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_411), .B(n_13), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_398), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_412), .B(n_13), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_398), .Y(n_464) );
NAND3xp33_ASAP7_75t_L g465 ( .A(n_399), .B(n_134), .C(n_198), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_415), .B(n_14), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_416), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_420), .Y(n_468) );
OAI221xp5_ASAP7_75t_SL g469 ( .A1(n_427), .A2(n_333), .B1(n_15), .B2(n_16), .C(n_17), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_415), .B(n_14), .Y(n_470) );
OAI31xp33_ASAP7_75t_SL g471 ( .A1(n_395), .A2(n_16), .A3(n_18), .B(n_333), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_420), .B(n_18), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_414), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_414), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_414), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_419), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_419), .Y(n_477) );
NAND3xp33_ASAP7_75t_L g478 ( .A(n_427), .B(n_198), .C(n_153), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_419), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_429), .B(n_426), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_430), .Y(n_481) );
BUFx12f_ASAP7_75t_L g482 ( .A(n_463), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_436), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_434), .B(n_407), .Y(n_484) );
NAND2x1_ASAP7_75t_L g485 ( .A(n_448), .B(n_418), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_439), .B(n_407), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_439), .B(n_428), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_433), .B(n_402), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_442), .B(n_418), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_442), .B(n_425), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_457), .A2(n_406), .B1(n_408), .B2(n_410), .Y(n_491) );
INVxp67_ASAP7_75t_L g492 ( .A(n_463), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_455), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_468), .B(n_423), .Y(n_494) );
AOI33xp33_ASAP7_75t_L g495 ( .A1(n_472), .A2(n_424), .A3(n_178), .B1(n_193), .B2(n_186), .B3(n_175), .Y(n_495) );
NAND2x1_ASAP7_75t_L g496 ( .A(n_448), .B(n_320), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_455), .Y(n_497) );
OAI31xp33_ASAP7_75t_L g498 ( .A1(n_469), .A2(n_351), .A3(n_299), .B(n_265), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_451), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_476), .B(n_21), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_468), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_441), .B(n_23), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_441), .B(n_24), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_435), .B(n_28), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_461), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_435), .B(n_29), .Y(n_506) );
NAND3xp33_ASAP7_75t_L g507 ( .A(n_471), .B(n_198), .C(n_156), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_443), .B(n_32), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_443), .B(n_33), .Y(n_509) );
NOR2xp33_ASAP7_75t_SL g510 ( .A(n_469), .B(n_320), .Y(n_510) );
NOR3xp33_ASAP7_75t_L g511 ( .A(n_458), .B(n_186), .C(n_178), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_436), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_452), .B(n_36), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_453), .B(n_39), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_461), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_452), .B(n_40), .Y(n_516) );
INVx1_ASAP7_75t_SL g517 ( .A(n_453), .Y(n_517) );
INVxp67_ASAP7_75t_L g518 ( .A(n_456), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_454), .B(n_41), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_466), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_444), .B(n_46), .Y(n_521) );
OR2x6_ASAP7_75t_L g522 ( .A(n_438), .B(n_320), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_456), .B(n_47), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_454), .B(n_48), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_470), .Y(n_525) );
BUFx3_ASAP7_75t_L g526 ( .A(n_445), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_447), .Y(n_527) );
INVx1_ASAP7_75t_SL g528 ( .A(n_517), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_480), .B(n_479), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_481), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_510), .A2(n_450), .B1(n_431), .B2(n_477), .Y(n_531) );
BUFx2_ASAP7_75t_L g532 ( .A(n_482), .Y(n_532) );
NAND3xp33_ASAP7_75t_L g533 ( .A(n_492), .B(n_471), .C(n_478), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_485), .A2(n_465), .B(n_457), .C(n_478), .Y(n_534) );
INVxp67_ASAP7_75t_L g535 ( .A(n_493), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_520), .B(n_479), .Y(n_536) );
AOI222xp33_ASAP7_75t_L g537 ( .A1(n_482), .A2(n_431), .B1(n_465), .B2(n_477), .C1(n_440), .C2(n_438), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_493), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_497), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_490), .B(n_476), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_499), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_511), .B(n_445), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_488), .A2(n_440), .B1(n_476), .B2(n_432), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_484), .B(n_460), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_486), .B(n_432), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_486), .B(n_432), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_518), .B(n_460), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_525), .B(n_447), .Y(n_548) );
NAND3xp33_ASAP7_75t_L g549 ( .A(n_491), .B(n_474), .C(n_475), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_496), .A2(n_446), .B(n_448), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_501), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_497), .Y(n_552) );
INVxp67_ASAP7_75t_L g553 ( .A(n_483), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_502), .B(n_432), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_495), .B(n_445), .Y(n_555) );
OAI32xp33_ASAP7_75t_L g556 ( .A1(n_489), .A2(n_437), .A3(n_473), .B1(n_475), .B2(n_467), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_483), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_512), .Y(n_558) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_507), .A2(n_448), .B(n_449), .Y(n_559) );
OAI211xp5_ASAP7_75t_L g560 ( .A1(n_498), .A2(n_445), .B(n_473), .C(n_437), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_487), .B(n_459), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_494), .B(n_445), .Y(n_562) );
OAI211xp5_ASAP7_75t_SL g563 ( .A1(n_495), .A2(n_437), .B(n_467), .C(n_462), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_487), .B(n_445), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_512), .Y(n_565) );
INVx1_ASAP7_75t_SL g566 ( .A(n_526), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_527), .Y(n_567) );
OAI21xp33_ASAP7_75t_L g568 ( .A1(n_504), .A2(n_464), .B(n_462), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_527), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_505), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_530), .Y(n_571) );
NOR2xp33_ASAP7_75t_SL g572 ( .A(n_532), .B(n_526), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_540), .B(n_504), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_533), .B(n_515), .Y(n_574) );
OAI211xp5_ASAP7_75t_L g575 ( .A1(n_537), .A2(n_502), .B(n_503), .C(n_506), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_540), .B(n_506), .Y(n_576) );
OAI21xp5_ASAP7_75t_L g577 ( .A1(n_534), .A2(n_503), .B(n_508), .Y(n_577) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_538), .Y(n_578) );
NOR3xp33_ASAP7_75t_SL g579 ( .A(n_560), .B(n_514), .C(n_523), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_541), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_551), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_561), .B(n_521), .Y(n_582) );
AND3x2_ASAP7_75t_L g583 ( .A(n_559), .B(n_509), .C(n_508), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_548), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_528), .B(n_524), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_566), .Y(n_586) );
NOR2x1_ASAP7_75t_L g587 ( .A(n_555), .B(n_519), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_567), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_547), .Y(n_589) );
INVxp67_ASAP7_75t_L g590 ( .A(n_538), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_536), .Y(n_591) );
NOR3xp33_ASAP7_75t_L g592 ( .A(n_549), .B(n_563), .C(n_562), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_570), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_529), .B(n_464), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_545), .B(n_462), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_552), .B(n_500), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_539), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_539), .Y(n_598) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_531), .A2(n_516), .B1(n_513), .B2(n_522), .C(n_164), .Y(n_599) );
NAND2xp33_ASAP7_75t_SL g600 ( .A(n_542), .B(n_500), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_557), .Y(n_601) );
NAND4xp25_ASAP7_75t_SL g602 ( .A(n_543), .B(n_522), .C(n_500), .D(n_318), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_586), .B(n_564), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_575), .A2(n_535), .B1(n_544), .B2(n_550), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_586), .Y(n_605) );
AO22x1_ASAP7_75t_L g606 ( .A1(n_592), .A2(n_535), .B1(n_546), .B2(n_554), .Y(n_606) );
OAI21xp33_ASAP7_75t_L g607 ( .A1(n_574), .A2(n_556), .B(n_568), .Y(n_607) );
XNOR2x1_ASAP7_75t_L g608 ( .A(n_577), .B(n_522), .Y(n_608) );
OAI21xp5_ASAP7_75t_SL g609 ( .A1(n_583), .A2(n_563), .B(n_553), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_571), .Y(n_610) );
NAND4xp75_ASAP7_75t_L g611 ( .A(n_587), .B(n_569), .C(n_565), .D(n_558), .Y(n_611) );
XOR2x2_ASAP7_75t_L g612 ( .A(n_585), .B(n_51), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_584), .B(n_591), .Y(n_613) );
OAI211xp5_ASAP7_75t_L g614 ( .A1(n_600), .A2(n_320), .B(n_280), .C(n_299), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_580), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_602), .A2(n_198), .B1(n_280), .B2(n_201), .Y(n_616) );
INVxp67_ASAP7_75t_L g617 ( .A(n_572), .Y(n_617) );
AOI221xp5_ASAP7_75t_L g618 ( .A1(n_589), .A2(n_201), .B1(n_60), .B2(n_64), .C(n_68), .Y(n_618) );
AOI211xp5_ASAP7_75t_SL g619 ( .A1(n_599), .A2(n_255), .B(n_69), .C(n_57), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_593), .B(n_581), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_604), .A2(n_585), .B1(n_582), .B2(n_573), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_613), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_604), .B(n_579), .Y(n_623) );
NAND2xp33_ASAP7_75t_R g624 ( .A(n_612), .B(n_573), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_607), .A2(n_590), .B1(n_598), .B2(n_597), .C(n_578), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_610), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_617), .Y(n_627) );
INVxp67_ASAP7_75t_L g628 ( .A(n_605), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_606), .A2(n_576), .B1(n_595), .B2(n_594), .C(n_596), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_603), .B(n_595), .Y(n_630) );
AND3x1_ASAP7_75t_L g631 ( .A(n_609), .B(n_601), .C(n_588), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_614), .B(n_588), .Y(n_632) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_608), .B(n_201), .C(n_619), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_620), .B(n_615), .Y(n_634) );
NOR4xp75_ASAP7_75t_L g635 ( .A(n_611), .B(n_616), .C(n_619), .D(n_618), .Y(n_635) );
AND2x4_ASAP7_75t_L g636 ( .A(n_617), .B(n_592), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_613), .Y(n_637) );
AOI21xp33_ASAP7_75t_SL g638 ( .A1(n_606), .A2(n_604), .B(n_617), .Y(n_638) );
INVx1_ASAP7_75t_SL g639 ( .A(n_627), .Y(n_639) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_636), .Y(n_640) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_636), .Y(n_641) );
BUFx2_ASAP7_75t_L g642 ( .A(n_628), .Y(n_642) );
NOR3xp33_ASAP7_75t_SL g643 ( .A(n_624), .B(n_623), .C(n_633), .Y(n_643) );
NOR2x1p5_ASAP7_75t_L g644 ( .A(n_643), .B(n_622), .Y(n_644) );
NAND3xp33_ASAP7_75t_L g645 ( .A(n_640), .B(n_638), .C(n_628), .Y(n_645) );
O2A1O1Ixp33_ASAP7_75t_L g646 ( .A1(n_641), .A2(n_625), .B(n_632), .C(n_637), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_645), .A2(n_639), .B1(n_644), .B2(n_642), .Y(n_647) );
OAI22x1_ASAP7_75t_L g648 ( .A1(n_646), .A2(n_642), .B1(n_621), .B2(n_631), .Y(n_648) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_647), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_648), .Y(n_650) );
AOI222xp33_ASAP7_75t_L g651 ( .A1(n_650), .A2(n_629), .B1(n_626), .B2(n_634), .C1(n_630), .C2(n_635), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_651), .A2(n_649), .B(n_650), .Y(n_652) );
endmodule