module fake_jpeg_30438_n_503 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_503);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_503;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_52),
.B(n_101),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_54),
.B(n_63),
.Y(n_117)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_55),
.Y(n_136)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_65),
.Y(n_154)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_20),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_69),
.B(n_75),
.Y(n_127)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_50),
.B(n_0),
.Y(n_70)
);

NAND2x1_ASAP7_75t_L g164 ( 
.A(n_70),
.B(n_50),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_21),
.B(n_0),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_79),
.Y(n_128)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_81),
.B(n_83),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_41),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_25),
.B(n_23),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_89),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_88),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_21),
.B(n_0),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_91),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_104),
.Y(n_109)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g155 ( 
.A(n_95),
.Y(n_155)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_22),
.B(n_42),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_102),
.Y(n_148)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_103),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_46),
.Y(n_104)
);

AND2x4_ASAP7_75t_SL g105 ( 
.A(n_70),
.B(n_50),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_105),
.B(n_95),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_53),
.A2(n_43),
.B1(n_49),
.B2(n_40),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_111),
.A2(n_98),
.B1(n_57),
.B2(n_25),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_52),
.A2(n_101),
.B1(n_67),
.B2(n_82),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_126),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_60),
.A2(n_49),
.B1(n_43),
.B2(n_40),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_71),
.A2(n_87),
.B1(n_86),
.B2(n_100),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_74),
.A2(n_49),
.B1(n_43),
.B2(n_40),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_58),
.B(n_22),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_132),
.B(n_157),
.Y(n_184)
);

AO22x2_ASAP7_75t_L g140 ( 
.A1(n_94),
.A2(n_27),
.B1(n_50),
.B2(n_38),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g207 ( 
.A1(n_140),
.A2(n_164),
.B1(n_63),
.B2(n_2),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_76),
.B(n_19),
.C(n_27),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_88),
.C(n_55),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_84),
.A2(n_19),
.B1(n_35),
.B2(n_44),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_143),
.A2(n_160),
.B1(n_161),
.B2(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_68),
.B(n_103),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_73),
.B(n_30),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_158),
.B(n_44),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_102),
.A2(n_35),
.B1(n_44),
.B2(n_26),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_93),
.A2(n_35),
.B1(n_44),
.B2(n_26),
.Y(n_161)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_165),
.Y(n_258)
);

INVx4_ASAP7_75t_SL g166 ( 
.A(n_135),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_166),
.B(n_177),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_97),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_167),
.B(n_168),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_138),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_118),
.A2(n_90),
.B1(n_80),
.B2(n_62),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_170),
.A2(n_206),
.B1(n_155),
.B2(n_136),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_110),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_171),
.Y(n_247)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_172),
.Y(n_256)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_78),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_174),
.B(n_180),
.Y(n_241)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_106),
.B(n_96),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_178),
.A2(n_187),
.B1(n_140),
.B2(n_146),
.Y(n_226)
);

INVx3_ASAP7_75t_SL g179 ( 
.A(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_179),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_47),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_117),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_181),
.B(n_185),
.Y(n_234)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_182),
.Y(n_261)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_127),
.B(n_128),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_47),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_186),
.B(n_197),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_105),
.A2(n_99),
.B1(n_91),
.B2(n_66),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_150),
.B(n_30),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_188),
.B(n_190),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_109),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_191),
.Y(n_239)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_105),
.B(n_27),
.CI(n_54),
.CON(n_190),
.SN(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_125),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_72),
.B1(n_56),
.B2(n_64),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_192),
.A2(n_211),
.B1(n_133),
.B2(n_152),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_193),
.B(n_195),
.Y(n_254)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_131),
.Y(n_194)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_196),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_129),
.B(n_37),
.Y(n_197)
);

OR2x2_ASAP7_75t_SL g198 ( 
.A(n_151),
.B(n_27),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_198),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_136),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_199),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_133),
.A2(n_37),
.B1(n_36),
.B2(n_23),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_200),
.A2(n_111),
.B1(n_112),
.B2(n_115),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_208),
.Y(n_240)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_139),
.Y(n_202)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_202),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_203),
.A2(n_141),
.B1(n_146),
.B2(n_7),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_142),
.B(n_44),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_217),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_124),
.B(n_63),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_144),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_125),
.A2(n_35),
.B1(n_45),
.B2(n_54),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g235 ( 
.A(n_207),
.B(n_107),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_148),
.B(n_137),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_107),
.Y(n_209)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_209),
.Y(n_260)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_120),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_212),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_140),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_137),
.B(n_1),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_120),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_139),
.B(n_1),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_215),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_110),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_145),
.B(n_3),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_216),
.B(n_218),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_140),
.B(n_3),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_161),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_143),
.C(n_160),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_221),
.B(n_224),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_145),
.C(n_124),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_225),
.A2(n_179),
.B(n_205),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_226),
.A2(n_250),
.B1(n_198),
.B2(n_179),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_190),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_230),
.B(n_231),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_167),
.B(n_144),
.C(n_121),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_235),
.A2(n_236),
.B1(n_238),
.B2(n_246),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_115),
.B1(n_112),
.B2(n_152),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_180),
.B(n_121),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_186),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_175),
.A2(n_153),
.B1(n_147),
.B2(n_134),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_249),
.A2(n_175),
.B1(n_192),
.B2(n_193),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_263),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_264),
.B(n_266),
.Y(n_320)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_222),
.Y(n_265)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_265),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_174),
.Y(n_266)
);

A2O1A1O1Ixp25_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_190),
.B(n_195),
.C(n_184),
.D(n_207),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_267),
.A2(n_241),
.B(n_254),
.Y(n_302)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_222),
.Y(n_269)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_269),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_239),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_270),
.B(n_271),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_168),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_220),
.B(n_197),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_272),
.B(n_278),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_273),
.A2(n_286),
.B1(n_294),
.B2(n_295),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_234),
.B(n_188),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_274),
.B(n_276),
.Y(n_313)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_223),
.Y(n_275)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_275),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_232),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_232),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_277),
.B(n_283),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_220),
.B(n_169),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_223),
.Y(n_279)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_279),
.Y(n_331)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_280),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_247),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_281),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_245),
.B(n_207),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_282),
.B(n_288),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_234),
.B(n_213),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_236),
.A2(n_218),
.B1(n_207),
.B2(n_211),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_284),
.A2(n_219),
.B1(n_244),
.B2(n_243),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_227),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_285),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_287),
.A2(n_292),
.B(n_250),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_245),
.B(n_183),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_254),
.B(n_241),
.CI(n_224),
.CON(n_289),
.SN(n_289)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_261),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_226),
.A2(n_178),
.B1(n_173),
.B2(n_191),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_290),
.A2(n_296),
.B1(n_297),
.B2(n_251),
.Y(n_323)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

NAND2xp33_ASAP7_75t_SL g305 ( 
.A(n_291),
.B(n_293),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_219),
.A2(n_210),
.B(n_172),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_247),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_256),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_255),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_255),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_235),
.A2(n_196),
.B1(n_194),
.B2(n_182),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_254),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_299),
.B(n_302),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_300),
.A2(n_260),
.B(n_281),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_301),
.A2(n_309),
.B1(n_321),
.B2(n_323),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_262),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_303),
.B(n_308),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_262),
.B(n_231),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_284),
.A2(n_235),
.B1(n_221),
.B2(n_249),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_221),
.C(n_230),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_315),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_266),
.B(n_240),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_240),
.C(n_237),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_317),
.B(n_322),
.Y(n_346)
);

OAI32xp33_ASAP7_75t_L g319 ( 
.A1(n_282),
.A2(n_235),
.A3(n_237),
.B1(n_238),
.B2(n_242),
.Y(n_319)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_268),
.A2(n_242),
.B1(n_246),
.B2(n_251),
.Y(n_321)
);

AOI322xp5_ASAP7_75t_L g324 ( 
.A1(n_276),
.A2(n_253),
.A3(n_176),
.B1(n_228),
.B2(n_258),
.C1(n_215),
.C2(n_233),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_271),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_263),
.A2(n_277),
.B(n_270),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_325),
.A2(n_269),
.B(n_275),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_259),
.C(n_233),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_326),
.B(n_330),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_289),
.B(n_259),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_272),
.Y(n_333)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_333),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_334),
.B(n_345),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_313),
.B(n_274),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_335),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_310),
.A2(n_268),
.B1(n_273),
.B2(n_286),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_336),
.A2(n_318),
.B1(n_330),
.B2(n_322),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_307),
.B(n_285),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_340),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_320),
.B(n_288),
.Y(n_341)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_341),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_320),
.B(n_278),
.Y(n_342)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_342),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_306),
.B(n_264),
.Y(n_343)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_343),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_283),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_325),
.B(n_292),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_347),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_301),
.B(n_293),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_348),
.B(n_351),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_308),
.B(n_267),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_303),
.C(n_299),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_311),
.A2(n_290),
.B1(n_297),
.B2(n_287),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_350),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_258),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_321),
.A2(n_267),
.B1(n_265),
.B2(n_291),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_352),
.A2(n_354),
.B1(n_355),
.B2(n_363),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_353),
.A2(n_361),
.B(n_312),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_309),
.A2(n_279),
.B1(n_280),
.B2(n_296),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_300),
.A2(n_253),
.B1(n_260),
.B2(n_295),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_304),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_356),
.Y(n_393)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_304),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_358),
.B(n_360),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_305),
.Y(n_359)
);

INVx11_ASAP7_75t_L g374 ( 
.A(n_359),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_326),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_311),
.A2(n_199),
.B1(n_209),
.B2(n_281),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_353),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_365),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_368),
.A2(n_377),
.B1(n_382),
.B2(n_383),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_380),
.Y(n_396)
);

NAND2x1_ASAP7_75t_L g372 ( 
.A(n_361),
.B(n_314),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_372),
.Y(n_401)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_344),
.Y(n_373)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_373),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_337),
.A2(n_317),
.B1(n_302),
.B2(n_332),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_375),
.A2(n_388),
.B1(n_389),
.B2(n_391),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_336),
.A2(n_318),
.B1(n_316),
.B2(n_332),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_338),
.B(n_316),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_344),
.A2(n_331),
.B1(n_329),
.B2(n_327),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_347),
.A2(n_331),
.B1(n_329),
.B2(n_327),
.Y(n_383)
);

OAI22x1_ASAP7_75t_SL g384 ( 
.A1(n_350),
.A2(n_312),
.B1(n_166),
.B2(n_171),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_384),
.A2(n_363),
.B1(n_358),
.B2(n_356),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_386),
.B(n_4),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_338),
.B(n_261),
.C(n_257),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_387),
.B(n_339),
.C(n_362),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_337),
.A2(n_312),
.B1(n_257),
.B2(n_202),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_354),
.A2(n_352),
.B1(n_355),
.B2(n_343),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_333),
.A2(n_165),
.B1(n_5),
.B2(n_7),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_402),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_366),
.B(n_335),
.Y(n_397)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_397),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_398),
.A2(n_412),
.B(n_388),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_341),
.Y(n_400)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_400),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_362),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_342),
.Y(n_403)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_403),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_383),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_404),
.B(n_405),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_387),
.B(n_339),
.C(n_349),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_346),
.C(n_357),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_406),
.B(n_381),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_368),
.B(n_357),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_408),
.B(n_416),
.Y(n_423)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_378),
.Y(n_410)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_410),
.Y(n_437)
);

FAx1_ASAP7_75t_SL g411 ( 
.A(n_375),
.B(n_346),
.CI(n_5),
.CON(n_411),
.SN(n_411)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_414),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_369),
.A2(n_17),
.B1(n_5),
.B2(n_7),
.Y(n_413)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_413),
.Y(n_421)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_378),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_367),
.B(n_4),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_415),
.B(n_417),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_377),
.B(n_4),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_385),
.B(n_8),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_373),
.A2(n_367),
.B1(n_390),
.B2(n_369),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_418),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_407),
.A2(n_382),
.B1(n_384),
.B2(n_386),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_422),
.A2(n_364),
.B1(n_399),
.B2(n_389),
.Y(n_439)
);

OA21x2_ASAP7_75t_L g427 ( 
.A1(n_409),
.A2(n_412),
.B(n_410),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_393),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_409),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_430),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_438),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_414),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_399),
.A2(n_401),
.B(n_407),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_431),
.B(n_372),
.Y(n_452)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_435),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_376),
.Y(n_436)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_436),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_396),
.B(n_381),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_441),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_426),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_440),
.B(n_444),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_419),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_434),
.A2(n_371),
.B1(n_376),
.B2(n_411),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_446),
.A2(n_420),
.B(n_434),
.Y(n_456)
);

A2O1A1Ixp33_ASAP7_75t_SL g447 ( 
.A1(n_422),
.A2(n_364),
.B(n_372),
.C(n_401),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_447),
.A2(n_394),
.B1(n_421),
.B2(n_427),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_433),
.B(n_379),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_448),
.B(n_451),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_429),
.B(n_395),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_450),
.B(n_438),
.Y(n_458)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_437),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_452),
.B(n_423),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_425),
.B(n_405),
.C(n_396),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_453),
.B(n_425),
.C(n_402),
.Y(n_457)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_436),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_454),
.B(n_427),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_456),
.B(n_457),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_458),
.B(n_462),
.C(n_465),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_459),
.B(n_466),
.Y(n_473)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_460),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_445),
.A2(n_424),
.B(n_431),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_461),
.B(n_449),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_450),
.B(n_406),
.C(n_423),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_439),
.A2(n_420),
.B1(n_421),
.B2(n_371),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_467),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_453),
.B(n_394),
.C(n_435),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_442),
.A2(n_432),
.B(n_413),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_442),
.B(n_411),
.C(n_408),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_468),
.B(n_8),
.Y(n_481)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_470),
.Y(n_486)
);

AOI221xp5_ASAP7_75t_L g474 ( 
.A1(n_455),
.A2(n_447),
.B1(n_443),
.B2(n_393),
.C(n_432),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_474),
.A2(n_464),
.B1(n_459),
.B2(n_462),
.Y(n_487)
);

AO22x1_ASAP7_75t_L g475 ( 
.A1(n_455),
.A2(n_447),
.B1(n_374),
.B2(n_416),
.Y(n_475)
);

AND2x4_ASAP7_75t_SL g490 ( 
.A(n_475),
.B(n_12),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_SL g477 ( 
.A(n_458),
.B(n_447),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_477),
.A2(n_455),
.B(n_466),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_457),
.B(n_391),
.C(n_374),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_478),
.B(n_479),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_465),
.B(n_8),
.C(n_9),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_481),
.B(n_469),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_483),
.A2(n_484),
.B(n_488),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_480),
.B(n_468),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_485),
.B(n_487),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_472),
.B(n_10),
.C(n_12),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_472),
.B(n_10),
.C(n_12),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_489),
.A2(n_12),
.B(n_13),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_490),
.A2(n_475),
.B1(n_474),
.B2(n_14),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_491),
.B(n_492),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_486),
.A2(n_476),
.B1(n_471),
.B2(n_473),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_495),
.B(n_490),
.C(n_484),
.Y(n_496)
);

AOI31xp33_ASAP7_75t_L g499 ( 
.A1(n_496),
.A2(n_494),
.A3(n_473),
.B(n_15),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_493),
.A2(n_482),
.B(n_490),
.Y(n_497)
);

AOI21x1_ASAP7_75t_L g500 ( 
.A1(n_497),
.A2(n_13),
.B(n_14),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_499),
.A2(n_500),
.B1(n_498),
.B2(n_15),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_501),
.B(n_15),
.Y(n_502)
);

BUFx24_ASAP7_75t_SL g503 ( 
.A(n_502),
.Y(n_503)
);


endmodule