module fake_jpeg_27008_n_294 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_294);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_287;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_11),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_11),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_24),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

AND2x4_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_24),
.Y(n_57)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_32),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_57),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_18),
.B1(n_19),
.B2(n_29),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_54),
.A2(n_19),
.B1(n_39),
.B2(n_44),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_35),
.Y(n_76)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_34),
.Y(n_62)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_61),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_63),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_65),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_43),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_43),
.B1(n_38),
.B2(n_35),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_66),
.A2(n_100),
.B1(n_28),
.B2(n_26),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_41),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_67),
.A2(n_81),
.B(n_103),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_68),
.Y(n_119)
);

OR2x2_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_43),
.Y(n_69)
);

NAND2x1_ASAP7_75t_SL g125 ( 
.A(n_69),
.B(n_74),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_53),
.B(n_33),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_72),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_71),
.Y(n_124)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_37),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_75),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_38),
.B(n_44),
.C(n_18),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_88),
.B1(n_89),
.B2(n_39),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_13),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_79),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_51),
.B(n_13),
.Y(n_80)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_80),
.A2(n_82),
.A3(n_91),
.B1(n_94),
.B2(n_102),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_56),
.B(n_13),
.Y(n_82)
);

AO22x1_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_44),
.B1(n_40),
.B2(n_34),
.Y(n_83)
);

NOR2x1p5_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_99),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_40),
.C(n_36),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_86),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_36),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_49),
.A2(n_39),
.B1(n_45),
.B2(n_19),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_27),
.B1(n_17),
.B2(n_22),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_101),
.B(n_40),
.C(n_31),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_21),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_21),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_97),
.B(n_14),
.Y(n_134)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_59),
.A2(n_27),
.B1(n_22),
.B2(n_28),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_21),
.B1(n_23),
.B2(n_28),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_31),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_55),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_64),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_108),
.B(n_116),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_111),
.A2(n_133),
.B1(n_62),
.B2(n_102),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_134),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_78),
.C(n_65),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_60),
.B1(n_96),
.B2(n_83),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_40),
.C(n_12),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_135),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_77),
.A2(n_42),
.B1(n_14),
.B2(n_20),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_131),
.B1(n_81),
.B2(n_89),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_88),
.A2(n_97),
.B1(n_91),
.B2(n_94),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_78),
.A2(n_23),
.B1(n_26),
.B2(n_31),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_40),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_138),
.A2(n_118),
.B1(n_129),
.B2(n_110),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_67),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_150),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_137),
.A2(n_87),
.B1(n_26),
.B2(n_23),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_145),
.B(n_151),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_146),
.B(n_147),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_124),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_153),
.B1(n_157),
.B2(n_159),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_113),
.B(n_85),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_137),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_154),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_111),
.A2(n_99),
.B1(n_95),
.B2(n_73),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_81),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_122),
.B(n_15),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_125),
.A2(n_83),
.B1(n_42),
.B2(n_15),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_158),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_125),
.A2(n_42),
.B1(n_15),
.B2(n_92),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_132),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_163),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_132),
.B(n_24),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_24),
.Y(n_164)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_20),
.Y(n_165)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_116),
.C(n_108),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_179),
.C(n_180),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_145),
.A2(n_115),
.B1(n_131),
.B2(n_117),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_168),
.A2(n_192),
.B1(n_153),
.B2(n_149),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_174),
.A2(n_175),
.B1(n_20),
.B2(n_16),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_156),
.B1(n_148),
.B2(n_139),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_139),
.A2(n_134),
.B(n_118),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_184),
.B(n_159),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_135),
.C(n_121),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_134),
.C(n_118),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_106),
.B(n_1),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_183),
.A2(n_154),
.B(n_150),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_163),
.A2(n_129),
.B(n_110),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_107),
.C(n_105),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_191),
.C(n_16),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_162),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_16),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_141),
.B(n_8),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_165),
.C(n_9),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_104),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_144),
.A2(n_84),
.B1(n_20),
.B2(n_16),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_176),
.B(n_140),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_195),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_200),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_209),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_155),
.B1(n_161),
.B2(n_147),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_151),
.B1(n_160),
.B2(n_162),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_182),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_204),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_176),
.B(n_84),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_0),
.B(n_1),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_206),
.A2(n_211),
.B1(n_169),
.B2(n_168),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_210),
.C(n_213),
.Y(n_220)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_208),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_12),
.B1(n_10),
.B2(n_9),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_166),
.C(n_179),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_174),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_0),
.C(n_2),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_188),
.B(n_2),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_214),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_3),
.C(n_5),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_187),
.C(n_190),
.Y(n_222)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_173),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_216),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_188),
.B(n_7),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_189),
.Y(n_227)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_232),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_170),
.C(n_181),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_229),
.C(n_207),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_206),
.A2(n_170),
.B1(n_193),
.B2(n_175),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_224),
.A2(n_230),
.B1(n_167),
.B2(n_195),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_227),
.B(n_215),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_181),
.C(n_177),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_196),
.A2(n_167),
.B1(n_172),
.B2(n_183),
.Y(n_230)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_235),
.A2(n_201),
.B(n_211),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_236),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_245),
.C(n_249),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_240),
.A2(n_242),
.B1(n_252),
.B2(n_224),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_198),
.B1(n_216),
.B2(n_197),
.Y(n_242)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_226),
.B(n_203),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_247),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_200),
.C(n_199),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_231),
.Y(n_246)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_213),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_205),
.B(n_177),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_248),
.A2(n_240),
.B1(n_219),
.B2(n_245),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_226),
.B(n_189),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_184),
.C(n_173),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_247),
.C(n_238),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_212),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_242),
.B1(n_236),
.B2(n_249),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_263),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_218),
.B1(n_232),
.B2(n_228),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_260),
.A2(n_248),
.B1(n_252),
.B2(n_237),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_229),
.C(n_221),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_209),
.B(n_244),
.Y(n_272)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_260),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_266),
.Y(n_278)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_269),
.Y(n_280)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_271),
.B(n_273),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_264),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_225),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_258),
.C(n_263),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_277),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_256),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_279),
.A2(n_256),
.B(n_254),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_280),
.A2(n_268),
.B(n_262),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_281),
.A2(n_284),
.B(n_274),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_276),
.A2(n_267),
.B1(n_259),
.B2(n_261),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_277),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_285),
.A2(n_287),
.B(n_278),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_282),
.B(n_275),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_279),
.C(n_259),
.Y(n_290)
);

NAND2x1_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_288),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_291),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_292),
.A2(n_233),
.B(n_222),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_254),
.Y(n_294)
);


endmodule