module fake_jpeg_2359_n_570 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_570);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_570;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_10),
.B(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g114 ( 
.A(n_54),
.Y(n_114)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_9),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_74),
.Y(n_109)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_60),
.Y(n_157)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_65),
.Y(n_164)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_68),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_18),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_69),
.B(n_83),
.Y(n_139)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_21),
.B(n_9),
.Y(n_74)
);

BUFx4f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_76),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_79),
.Y(n_166)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_82),
.Y(n_121)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_18),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_23),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_87),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_42),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_93),
.B(n_100),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_43),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_102),
.Y(n_125)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_95),
.B(n_97),
.Y(n_162)
);

BUFx16f_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_96),
.Y(n_127)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_98),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_99),
.B(n_101),
.Y(n_168)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_19),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_19),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_105),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_104),
.B(n_36),
.Y(n_169)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_19),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_48),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_75),
.A2(n_52),
.B1(n_46),
.B2(n_38),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_108),
.A2(n_147),
.B1(n_150),
.B2(n_28),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_52),
.B1(n_25),
.B2(n_46),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_110),
.A2(n_117),
.B1(n_141),
.B2(n_160),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_52),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_111),
.B(n_29),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_46),
.B1(n_38),
.B2(n_34),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_116),
.A2(n_58),
.B1(n_1),
.B2(n_2),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_30),
.B1(n_29),
.B2(n_25),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_53),
.A2(n_51),
.B1(n_22),
.B2(n_45),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_118),
.B(n_132),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_22),
.C(n_35),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_123),
.B(n_24),
.C(n_36),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_85),
.A2(n_51),
.B1(n_22),
.B2(n_45),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_106),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_62),
.A2(n_48),
.B1(n_31),
.B2(n_25),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_136),
.A2(n_151),
.B1(n_28),
.B2(n_35),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g141 ( 
.A1(n_56),
.A2(n_31),
.B1(n_26),
.B2(n_38),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_24),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_156),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_54),
.B(n_105),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_152),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_55),
.A2(n_31),
.B1(n_26),
.B2(n_27),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_54),
.A2(n_30),
.B1(n_26),
.B2(n_27),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_68),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_67),
.B(n_34),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_100),
.A2(n_51),
.B1(n_45),
.B2(n_36),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_154),
.A2(n_58),
.B1(n_77),
.B2(n_66),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_71),
.B(n_24),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_73),
.A2(n_78),
.B1(n_79),
.B2(n_84),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_98),
.B(n_34),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_104),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_169),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_172),
.Y(n_255)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_121),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_175),
.B(n_178),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_176),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_177),
.B(n_193),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_109),
.B(n_29),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_179),
.B(n_216),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_104),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_181),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_182),
.A2(n_210),
.B1(n_224),
.B2(n_228),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_35),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_183),
.B(n_187),
.Y(n_235)
);

OA22x2_ASAP7_75t_L g244 ( 
.A1(n_184),
.A2(n_122),
.B1(n_137),
.B2(n_118),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_185),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_186),
.B(n_188),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_99),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_139),
.B(n_84),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_189),
.A2(n_198),
.B1(n_114),
.B2(n_122),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_146),
.Y(n_190)
);

BUFx2_ASAP7_75t_SL g257 ( 
.A(n_190),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_124),
.B(n_101),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_191),
.Y(n_271)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_192),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_125),
.B(n_77),
.C(n_66),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_111),
.B(n_10),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_195),
.Y(n_234)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_133),
.Y(n_196)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_196),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_123),
.B(n_0),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_200),
.Y(n_238)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_199),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_131),
.B(n_18),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_201),
.Y(n_263)
);

INVx6_ASAP7_75t_SL g202 ( 
.A(n_127),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_202),
.Y(n_245)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_203),
.Y(n_267)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

AOI32xp33_ASAP7_75t_L g205 ( 
.A1(n_137),
.A2(n_9),
.A3(n_15),
.B1(n_3),
.B2(n_4),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_SL g273 ( 
.A(n_205),
.B(n_144),
.C(n_146),
.Y(n_273)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_144),
.Y(n_206)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_206),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_167),
.A2(n_8),
.B(n_15),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_214),
.B(n_132),
.Y(n_233)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_126),
.B(n_0),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_209),
.B(n_219),
.Y(n_262)
);

INVx11_ASAP7_75t_L g210 ( 
.A(n_133),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_127),
.B(n_8),
.Y(n_211)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_116),
.A2(n_6),
.B1(n_14),
.B2(n_3),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_212),
.A2(n_154),
.B1(n_149),
.B2(n_159),
.Y(n_247)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_107),
.Y(n_213)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_167),
.A2(n_11),
.B(n_14),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_143),
.Y(n_215)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_112),
.B(n_0),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_135),
.B(n_11),
.Y(n_217)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_112),
.B(n_0),
.Y(n_218)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_126),
.B(n_0),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_166),
.Y(n_220)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_220),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_135),
.B(n_4),
.Y(n_221)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_221),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_164),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_222),
.B(n_227),
.Y(n_282)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_160),
.A2(n_4),
.B1(n_5),
.B2(n_11),
.Y(n_224)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_129),
.Y(n_225)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_225),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_112),
.B(n_1),
.Y(n_226)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_226),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_128),
.B(n_141),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g228 ( 
.A(n_140),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_149),
.Y(n_230)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_230),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_158),
.Y(n_231)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_231),
.Y(n_283)
);

BUFx12f_ASAP7_75t_L g232 ( 
.A(n_140),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_232),
.A2(n_114),
.B1(n_115),
.B2(n_133),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_233),
.B(n_273),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_241),
.B(n_244),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_247),
.A2(n_249),
.B1(n_250),
.B2(n_270),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_192),
.A2(n_163),
.B1(n_159),
.B2(n_168),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_163),
.B1(n_165),
.B2(n_170),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_194),
.A2(n_128),
.B1(n_119),
.B2(n_138),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_260),
.A2(n_268),
.B1(n_222),
.B2(n_218),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_194),
.A2(n_119),
.B1(n_138),
.B2(n_165),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_269),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_180),
.A2(n_157),
.B1(n_155),
.B2(n_164),
.Y(n_270)
);

OA22x2_ASAP7_75t_L g275 ( 
.A1(n_229),
.A2(n_107),
.B1(n_157),
.B2(n_155),
.Y(n_275)
);

OA22x2_ASAP7_75t_L g291 ( 
.A1(n_275),
.A2(n_201),
.B1(n_213),
.B2(n_230),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_227),
.A2(n_164),
.B1(n_170),
.B2(n_130),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_279),
.A2(n_281),
.B1(n_210),
.B2(n_120),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_173),
.A2(n_133),
.B1(n_130),
.B2(n_115),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g284 ( 
.A(n_180),
.B(n_113),
.CI(n_120),
.CON(n_284),
.SN(n_284)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_284),
.B(n_183),
.Y(n_292)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_208),
.Y(n_285)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_215),
.Y(n_287)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_287),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_197),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_288),
.B(n_296),
.C(n_297),
.Y(n_354)
);

AND2x2_ASAP7_75t_SL g289 ( 
.A(n_286),
.B(n_179),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_289),
.B(n_291),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_242),
.B(n_175),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g367 ( 
.A(n_290),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_292),
.B(n_304),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_178),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_293),
.B(n_295),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_262),
.B(n_187),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_193),
.C(n_177),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_235),
.B(n_171),
.C(n_179),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_239),
.B(n_209),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_298),
.B(n_299),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_219),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_282),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_301),
.B(n_324),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_262),
.B(n_226),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_302),
.B(n_307),
.Y(n_372)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_258),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_235),
.A2(n_181),
.B1(n_198),
.B2(n_214),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_305),
.A2(n_306),
.B1(n_313),
.B2(n_319),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_236),
.A2(n_181),
.B1(n_207),
.B2(n_218),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_238),
.B(n_236),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_243),
.Y(n_309)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_309),
.Y(n_340)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_237),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_310),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_238),
.B(n_216),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_311),
.B(n_317),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_312),
.A2(n_322),
.B1(n_337),
.B2(n_252),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_282),
.A2(n_216),
.B1(n_226),
.B2(n_185),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_237),
.Y(n_314)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_314),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_233),
.A2(n_202),
.B(n_196),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_315),
.A2(n_316),
.B(n_335),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_271),
.A2(n_206),
.B(n_176),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_234),
.B(n_204),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_243),
.Y(n_318)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_318),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_241),
.A2(n_231),
.B1(n_220),
.B2(n_223),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_248),
.Y(n_320)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_320),
.Y(n_362)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_246),
.Y(n_321)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_321),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_264),
.A2(n_199),
.B1(n_174),
.B2(n_203),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_255),
.B(n_232),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_323),
.B(n_328),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_245),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_277),
.B(n_225),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_325),
.B(n_326),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_277),
.B(n_232),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_248),
.Y(n_327)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_327),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_286),
.B(n_232),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_240),
.B(n_228),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_330),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_280),
.B(n_228),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_331),
.B(n_333),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_254),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_332),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_253),
.B(n_129),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_280),
.B(n_287),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_336),
.A2(n_244),
.B1(n_275),
.B2(n_274),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_268),
.A2(n_260),
.B1(n_270),
.B2(n_284),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_285),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_338),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_341),
.A2(n_344),
.B1(n_350),
.B2(n_358),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_337),
.A2(n_284),
.B1(n_286),
.B2(n_275),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_348),
.A2(n_360),
.B1(n_371),
.B2(n_322),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_315),
.A2(n_244),
.B(n_278),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_349),
.A2(n_359),
.B(n_381),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_301),
.A2(n_275),
.B1(n_278),
.B2(n_253),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_288),
.B(n_244),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_361),
.C(n_363),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_335),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_352),
.B(n_355),
.Y(n_410)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_293),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_353),
.B(n_290),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_331),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_334),
.A2(n_273),
.B1(n_283),
.B2(n_254),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_303),
.A2(n_272),
.B(n_274),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_334),
.A2(n_283),
.B1(n_246),
.B2(n_259),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_296),
.B(n_272),
.C(n_265),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_297),
.B(n_261),
.C(n_259),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_307),
.B(n_261),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_364),
.B(n_369),
.C(n_374),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_295),
.B(n_256),
.C(n_267),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_334),
.A2(n_257),
.B1(n_263),
.B2(n_267),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_303),
.A2(n_228),
.B1(n_263),
.B2(n_256),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_373),
.A2(n_378),
.B1(n_350),
.B2(n_342),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_289),
.B(n_113),
.C(n_1),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_302),
.B(n_4),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_375),
.B(n_306),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_329),
.A2(n_5),
.B(n_12),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_384),
.B(n_387),
.Y(n_441)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_366),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_385),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_299),
.Y(n_386)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_386),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_379),
.B(n_324),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_389),
.B(n_380),
.Y(n_437)
);

XNOR2x1_ASAP7_75t_L g390 ( 
.A(n_351),
.B(n_303),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_390),
.B(n_400),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_369),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_391),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_352),
.B(n_298),
.Y(n_392)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_392),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_366),
.Y(n_394)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_394),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_367),
.B(n_317),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_395),
.B(n_398),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_376),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_396),
.B(n_397),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_339),
.B(n_338),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_345),
.B(n_323),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_345),
.B(n_292),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_399),
.B(n_402),
.Y(n_448)
);

XOR2x2_ASAP7_75t_L g400 ( 
.A(n_354),
.B(n_311),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_339),
.B(n_308),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_401),
.B(n_404),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_365),
.B(n_316),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_354),
.B(n_361),
.C(n_363),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_407),
.C(n_408),
.Y(n_423)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_340),
.Y(n_404)
);

OAI32xp33_ASAP7_75t_L g405 ( 
.A1(n_372),
.A2(n_308),
.A3(n_309),
.B1(n_327),
.B2(n_318),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_405),
.A2(n_409),
.B(n_368),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_356),
.A2(n_294),
.B1(n_289),
.B2(n_305),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_406),
.A2(n_414),
.B1(n_415),
.B2(n_416),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_364),
.B(n_289),
.C(n_328),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_372),
.B(n_313),
.C(n_320),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_378),
.A2(n_312),
.B(n_333),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_373),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_412),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_378),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_413),
.Y(n_433)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_340),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_357),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_383),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_418),
.A2(n_419),
.B1(n_420),
.B2(n_355),
.Y(n_432)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_357),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_300),
.C(n_314),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_421),
.B(n_383),
.C(n_342),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_425),
.B(n_431),
.C(n_421),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_417),
.A2(n_349),
.B(n_359),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_427),
.A2(n_440),
.B(n_449),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_411),
.A2(n_356),
.B1(n_348),
.B2(n_344),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_430),
.B(n_434),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_403),
.B(n_388),
.C(n_400),
.Y(n_431)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_432),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_411),
.A2(n_294),
.B1(n_360),
.B2(n_377),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_415),
.A2(n_347),
.B1(n_358),
.B2(n_371),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_435),
.B(n_443),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_438),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_388),
.B(n_380),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_390),
.B(n_382),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_439),
.B(n_408),
.Y(n_463)
);

OA21x2_ASAP7_75t_L g440 ( 
.A1(n_409),
.A2(n_291),
.B(n_382),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_412),
.A2(n_347),
.B1(n_329),
.B2(n_381),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_413),
.A2(n_368),
.B1(n_362),
.B2(n_343),
.Y(n_444)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_444),
.Y(n_461)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_445),
.Y(n_464)
);

OA21x2_ASAP7_75t_L g449 ( 
.A1(n_410),
.A2(n_291),
.B(n_319),
.Y(n_449)
);

XNOR2x2_ASAP7_75t_L g451 ( 
.A(n_389),
.B(n_375),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_451),
.B(n_407),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_397),
.A2(n_362),
.B1(n_343),
.B2(n_374),
.Y(n_453)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_453),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_410),
.A2(n_346),
.B1(n_300),
.B2(n_291),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_454),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_396),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_456),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_422),
.B(n_386),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_458),
.B(n_459),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_422),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_463),
.B(n_469),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_393),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_465),
.B(n_467),
.C(n_472),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_441),
.B(n_392),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_466),
.B(n_475),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_423),
.B(n_393),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_431),
.B(n_410),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_477),
.C(n_479),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_452),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_474),
.B(n_429),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_446),
.B(n_401),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_450),
.Y(n_476)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_476),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_423),
.B(n_436),
.Y(n_477)
);

AO22x1_ASAP7_75t_SL g478 ( 
.A1(n_426),
.A2(n_406),
.B1(n_405),
.B2(n_417),
.Y(n_478)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_478),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_439),
.B(n_416),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_450),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_480),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_448),
.B(n_321),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_482),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_448),
.B(n_414),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_457),
.A2(n_440),
.B1(n_447),
.B2(n_428),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_485),
.A2(n_486),
.B1(n_501),
.B2(n_503),
.Y(n_507)
);

OAI321xp33_ASAP7_75t_L g486 ( 
.A1(n_464),
.A2(n_440),
.A3(n_428),
.B1(n_424),
.B2(n_447),
.C(n_427),
.Y(n_486)
);

AND3x1_ASAP7_75t_L g489 ( 
.A(n_464),
.B(n_471),
.C(n_470),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_489),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_460),
.A2(n_430),
.B1(n_434),
.B2(n_435),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_491),
.A2(n_496),
.B1(n_468),
.B2(n_404),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_470),
.A2(n_445),
.B(n_424),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_495),
.A2(n_499),
.B(n_505),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_460),
.A2(n_443),
.B1(n_433),
.B2(n_454),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_455),
.A2(n_449),
.B1(n_429),
.B2(n_453),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_497),
.A2(n_468),
.B1(n_457),
.B2(n_478),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_471),
.A2(n_449),
.B(n_425),
.Y(n_499)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_474),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_478),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_455),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_461),
.B(n_444),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_504),
.B(n_13),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_461),
.A2(n_436),
.B(n_437),
.Y(n_505)
);

BUFx12f_ASAP7_75t_SL g506 ( 
.A(n_479),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_506),
.A2(n_463),
.B(n_469),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_488),
.B(n_472),
.C(n_473),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_512),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_510),
.A2(n_520),
.B1(n_496),
.B2(n_498),
.Y(n_527)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_511),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_492),
.B(n_465),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_488),
.B(n_467),
.C(n_477),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_513),
.B(n_517),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_515),
.B(n_499),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_516),
.A2(n_497),
.B1(n_486),
.B2(n_503),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_490),
.B(n_462),
.C(n_451),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_492),
.A2(n_385),
.B1(n_346),
.B2(n_462),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_518),
.B(n_519),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_490),
.B(n_310),
.C(n_332),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_487),
.A2(n_291),
.B1(n_332),
.B2(n_16),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_505),
.B(n_12),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_521),
.B(n_522),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_SL g522 ( 
.A(n_495),
.B(n_13),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_494),
.B(n_13),
.C(n_16),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_523),
.B(n_524),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_494),
.B(n_13),
.C(n_16),
.Y(n_524)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_525),
.Y(n_533)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_527),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_508),
.B(n_484),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_528),
.B(n_513),
.Y(n_551)
);

BUFx24_ASAP7_75t_SL g529 ( 
.A(n_514),
.Y(n_529)
);

BUFx24_ASAP7_75t_SL g549 ( 
.A(n_529),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_531),
.B(n_535),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_534),
.A2(n_511),
.B(n_504),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_519),
.B(n_500),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_507),
.A2(n_498),
.B(n_485),
.Y(n_536)
);

OA21x2_ASAP7_75t_L g546 ( 
.A1(n_536),
.A2(n_487),
.B(n_510),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_509),
.B(n_484),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_540),
.B(n_493),
.Y(n_545)
);

AO21x1_ASAP7_75t_L g541 ( 
.A1(n_536),
.A2(n_509),
.B(n_483),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_541),
.B(n_545),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_532),
.A2(n_514),
.B(n_515),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_543),
.A2(n_521),
.B(n_523),
.Y(n_557)
);

OAI221xp5_ASAP7_75t_L g544 ( 
.A1(n_526),
.A2(n_493),
.B1(n_483),
.B2(n_501),
.C(n_502),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_544),
.A2(n_546),
.B1(n_527),
.B2(n_531),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_547),
.B(n_550),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_533),
.B(n_516),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_551),
.B(n_537),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_552),
.A2(n_553),
.B(n_555),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_550),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_548),
.B(n_530),
.C(n_534),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_556),
.A2(n_557),
.B(n_539),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_555),
.B(n_542),
.C(n_546),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_559),
.B(n_561),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_560),
.A2(n_562),
.B1(n_558),
.B2(n_491),
.Y(n_563)
);

BUFx24_ASAP7_75t_SL g561 ( 
.A(n_554),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_563),
.B(n_517),
.C(n_520),
.Y(n_566)
);

O2A1O1Ixp33_ASAP7_75t_SL g564 ( 
.A1(n_561),
.A2(n_522),
.B(n_489),
.C(n_549),
.Y(n_564)
);

NAND3xp33_ASAP7_75t_L g567 ( 
.A(n_564),
.B(n_524),
.C(n_538),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_566),
.B(n_567),
.C(n_565),
.Y(n_568)
);

FAx1_ASAP7_75t_SL g569 ( 
.A(n_568),
.B(n_506),
.CI(n_538),
.CON(n_569),
.SN(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_569),
.B(n_16),
.Y(n_570)
);


endmodule