module fake_jpeg_26863_n_228 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_29),
.Y(n_47)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_6),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_30),
.B(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_6),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_23),
.B1(n_22),
.B2(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_33),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_25),
.B1(n_13),
.B2(n_22),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_16),
.B1(n_25),
.B2(n_15),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_28),
.B1(n_32),
.B2(n_15),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_33),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_45),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_52),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_28),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_33),
.Y(n_71)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_56),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_32),
.B1(n_28),
.B2(n_25),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_28),
.B1(n_22),
.B2(n_16),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_30),
.B1(n_21),
.B2(n_17),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_34),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_21),
.Y(n_82)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_62),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_74),
.B(n_60),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_38),
.B1(n_37),
.B2(n_36),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_73),
.B1(n_79),
.B2(n_50),
.Y(n_90)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_73)
);

AOI32xp33_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_47),
.A3(n_30),
.B1(n_46),
.B2(n_45),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_49),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_59),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_48),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_50),
.B1(n_53),
.B2(n_61),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_85),
.B(n_94),
.Y(n_109)
);

XOR2x2_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_89),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_56),
.B1(n_52),
.B2(n_54),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_68),
.B1(n_69),
.B2(n_79),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

BUFx8_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

AOI22x1_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_57),
.B1(n_58),
.B2(n_27),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_52),
.B1(n_63),
.B2(n_56),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_69),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_98),
.Y(n_104)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_99),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_107),
.B1(n_94),
.B2(n_83),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_68),
.C(n_65),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_26),
.C(n_39),
.Y(n_122)
);

AOI32xp33_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_69),
.A3(n_78),
.B1(n_72),
.B2(n_79),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_114),
.B(n_116),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_69),
.B1(n_82),
.B2(n_66),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_67),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_80),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_71),
.B(n_70),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_70),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_39),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_SL g116 ( 
.A(n_84),
.B(n_21),
.C(n_14),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_90),
.B1(n_83),
.B2(n_87),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_119),
.B1(n_126),
.B2(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_123),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_117),
.C(n_100),
.Y(n_139)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_13),
.B(n_89),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_125),
.B(n_134),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_41),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_67),
.B1(n_99),
.B2(n_95),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_127),
.Y(n_143)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_129),
.B(n_132),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_27),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_130),
.B(n_112),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_95),
.B(n_1),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

NAND2xp33_ASAP7_75t_SL g136 ( 
.A(n_116),
.B(n_18),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_26),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_144),
.C(n_146),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_117),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_141),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_102),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_145),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_103),
.C(n_102),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_103),
.C(n_114),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_106),
.C(n_116),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_125),
.C(n_123),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_150),
.B1(n_135),
.B2(n_132),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_111),
.B1(n_112),
.B2(n_17),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_121),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_129),
.B(n_112),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_153),
.B(n_131),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_134),
.B(n_125),
.Y(n_162)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_159),
.B(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_163),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_124),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_164),
.C(n_168),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_162),
.A2(n_154),
.B(n_141),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_148),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_155),
.Y(n_178)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_21),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_27),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_42),
.C(n_26),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_170),
.C(n_171),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_42),
.C(n_26),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_42),
.C(n_41),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_173),
.A2(n_9),
.B(n_7),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_171),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_169),
.B1(n_165),
.B2(n_170),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g176 ( 
.A(n_166),
.B(n_137),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_176),
.B(n_182),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_156),
.B(n_140),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_183),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_179),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_159),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_141),
.C(n_145),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_185),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_41),
.C(n_24),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_179),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_10),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_193),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_18),
.C(n_19),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_196),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_10),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_36),
.B1(n_76),
.B2(n_59),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_195),
.Y(n_201)
);

BUFx24_ASAP7_75t_SL g195 ( 
.A(n_178),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_180),
.C(n_182),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_200),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_204),
.B(n_10),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_174),
.C(n_41),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_76),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_205),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_192),
.B(n_8),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_24),
.C(n_33),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_199),
.B(n_8),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_207),
.B(n_1),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_9),
.B1(n_7),
.B2(n_6),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_209),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_198),
.A2(n_12),
.B(n_19),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_210),
.A2(n_211),
.B(n_0),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_12),
.B(n_18),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_202),
.A2(n_12),
.B(n_1),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_213),
.A2(n_1),
.B(n_2),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_215),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_2),
.Y(n_221)
);

AOI21x1_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_212),
.B(n_3),
.Y(n_217)
);

AO21x1_ASAP7_75t_L g222 ( 
.A1(n_217),
.A2(n_219),
.B(n_2),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_222),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_14),
.B1(n_3),
.B2(n_4),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_223),
.A2(n_2),
.B(n_3),
.Y(n_224)
);

AOI321xp33_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_220),
.A3(n_225),
.B1(n_4),
.B2(n_5),
.C(n_24),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_5),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_5),
.B(n_14),
.Y(n_228)
);


endmodule