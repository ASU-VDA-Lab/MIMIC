module fake_jpeg_12318_n_442 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_442);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_442;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_59),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_15),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_60),
.B(n_100),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_65),
.Y(n_171)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_30),
.B(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_71),
.Y(n_118)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_69),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_15),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_70),
.B(n_75),
.Y(n_173)
);

INVx2_ASAP7_75t_R g71 ( 
.A(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_74),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_37),
.B(n_14),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_83),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_79),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_19),
.B(n_0),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_80),
.B(n_95),
.Y(n_149)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_81),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_24),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_28),
.B(n_1),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_84),
.B(n_86),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_28),
.B(n_1),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_29),
.B(n_1),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_88),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_24),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_24),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_90),
.B(n_96),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_92),
.Y(n_175)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_93),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_29),
.Y(n_96)
);

INVx2_ASAP7_75t_R g97 ( 
.A(n_55),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_98),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_42),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_103),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_101),
.B(n_105),
.Y(n_163)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_102),
.B(n_104),
.Y(n_153)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_34),
.B(n_2),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_106),
.B(n_108),
.Y(n_167)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_107),
.B(n_113),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_40),
.Y(n_108)
);

BUFx16f_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_109),
.B(n_110),
.Y(n_168)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_21),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_40),
.B(n_3),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_111),
.B(n_112),
.Y(n_174)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_23),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_45),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_36),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_80),
.A2(n_20),
.B1(n_54),
.B2(n_25),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_115),
.B(n_140),
.C(n_155),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_73),
.B1(n_114),
.B2(n_61),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_SL g188 ( 
.A1(n_116),
.A2(n_152),
.B(n_182),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_33),
.B1(n_22),
.B2(n_26),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_117),
.A2(n_119),
.B1(n_120),
.B2(n_123),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_74),
.A2(n_20),
.B1(n_26),
.B2(n_33),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_59),
.A2(n_22),
.B1(n_25),
.B2(n_47),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_65),
.A2(n_47),
.B1(n_52),
.B2(n_51),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_126),
.B(n_117),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_65),
.A2(n_52),
.B1(n_51),
.B2(n_50),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_134),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_77),
.A2(n_23),
.B1(n_50),
.B2(n_38),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_135),
.A2(n_148),
.B1(n_156),
.B2(n_158),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_58),
.B(n_38),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_138),
.B(n_159),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_103),
.A2(n_53),
.B1(n_46),
.B2(n_39),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_SL g143 ( 
.A(n_67),
.Y(n_143)
);

INVx11_ASAP7_75t_L g240 ( 
.A(n_143),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_66),
.A2(n_53),
.B1(n_46),
.B2(n_39),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_94),
.A2(n_34),
.B1(n_5),
.B2(n_6),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_57),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_81),
.B(n_3),
.C(n_7),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_93),
.A2(n_95),
.B1(n_101),
.B2(n_100),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_63),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_79),
.A2(n_9),
.B1(n_89),
.B2(n_85),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_165),
.B1(n_176),
.B2(n_180),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_107),
.A2(n_9),
.B1(n_71),
.B2(n_97),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_92),
.A2(n_106),
.B1(n_113),
.B2(n_99),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_92),
.A2(n_106),
.B1(n_69),
.B2(n_78),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

OA22x2_ASAP7_75t_L g176 ( 
.A1(n_109),
.A2(n_104),
.B1(n_82),
.B2(n_56),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_91),
.A2(n_24),
.B1(n_29),
.B2(n_20),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_179),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_109),
.A2(n_114),
.B1(n_77),
.B2(n_100),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_74),
.A2(n_24),
.B1(n_29),
.B2(n_20),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g183 ( 
.A1(n_80),
.A2(n_58),
.B1(n_95),
.B2(n_81),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_183),
.A2(n_136),
.B1(n_139),
.B2(n_162),
.Y(n_233)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_131),
.B(n_138),
.C(n_163),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_185),
.B(n_193),
.Y(n_253)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_124),
.Y(n_186)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_186),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_142),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_187),
.B(n_206),
.Y(n_248)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_189),
.B(n_191),
.Y(n_251)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_192),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_130),
.B(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_194),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_197),
.Y(n_266)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_198),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_149),
.B(n_183),
.Y(n_200)
);

NAND2x1_ASAP7_75t_L g268 ( 
.A(n_200),
.B(n_201),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_149),
.B(n_183),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_125),
.Y(n_202)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_202),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_118),
.B(n_174),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_203),
.B(n_208),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_156),
.A2(n_157),
.B1(n_117),
.B2(n_124),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_205),
.A2(n_224),
.B1(n_233),
.B2(n_195),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_141),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_127),
.B(n_151),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_153),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_209),
.B(n_218),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_167),
.B(n_140),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_210),
.B(n_211),
.Y(n_265)
);

NAND2xp33_ASAP7_75t_SL g211 ( 
.A(n_128),
.B(n_172),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_212),
.Y(n_272)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_213),
.Y(n_258)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

INVx13_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

INVx13_ASAP7_75t_L g245 ( 
.A(n_215),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_128),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_217),
.B(n_227),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_155),
.B(n_164),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_164),
.B(n_178),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_219),
.B(n_225),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_117),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_241),
.C(n_234),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_126),
.B(n_115),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_223),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_122),
.Y(n_222)
);

INVx8_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_158),
.B(n_135),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_145),
.A2(n_129),
.B1(n_132),
.B2(n_137),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_177),
.B(n_175),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_129),
.Y(n_226)
);

INVx13_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_133),
.Y(n_228)
);

INVx13_ASAP7_75t_L g285 ( 
.A(n_228),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_145),
.B(n_137),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_236),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_136),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_231),
.B(n_235),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_177),
.B(n_175),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_232),
.B(n_242),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_233),
.A2(n_176),
.B1(n_181),
.B2(n_154),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_139),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_150),
.B(n_176),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_150),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_237),
.Y(n_257)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_162),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_238),
.Y(n_262)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_133),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_239),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_176),
.B(n_133),
.C(n_147),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_147),
.B(n_144),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_244),
.A2(n_262),
.B1(n_250),
.B2(n_269),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_223),
.A2(n_144),
.B1(n_154),
.B2(n_181),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_247),
.A2(n_263),
.B1(n_264),
.B2(n_276),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_191),
.A2(n_147),
.B1(n_220),
.B2(n_184),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_249),
.A2(n_261),
.B1(n_239),
.B2(n_226),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_256),
.A2(n_277),
.B(n_265),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_191),
.A2(n_220),
.B1(n_200),
.B2(n_201),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_190),
.A2(n_221),
.B1(n_195),
.B2(n_199),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_229),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_197),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_189),
.B(n_185),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_275),
.B(n_273),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_190),
.A2(n_230),
.B1(n_236),
.B2(n_201),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_204),
.A2(n_196),
.B1(n_234),
.B2(n_216),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_200),
.B(n_230),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_279),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_186),
.B(n_213),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_212),
.B(n_214),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_262),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_241),
.B(n_188),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_192),
.C(n_207),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_237),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_288),
.B(n_311),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_289),
.B(n_295),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_279),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_290),
.B(n_304),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_246),
.A2(n_204),
.B1(n_196),
.B2(n_216),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_291),
.A2(n_316),
.B1(n_250),
.B2(n_281),
.Y(n_341)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_292),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_293),
.B(n_283),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_268),
.A2(n_228),
.B(n_238),
.Y(n_294)
);

NAND2xp33_ASAP7_75t_SL g332 ( 
.A(n_294),
.B(n_312),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_248),
.B(n_227),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_275),
.B(n_198),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_297),
.B(n_300),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_215),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_298),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_299),
.Y(n_327)
);

INVx8_ASAP7_75t_L g301 ( 
.A(n_255),
.Y(n_301)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_301),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_302),
.Y(n_347)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_282),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_306),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_253),
.B(n_222),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_253),
.B(n_240),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_264),
.A2(n_240),
.B1(n_263),
.B2(n_276),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_307),
.A2(n_320),
.B1(n_322),
.B2(n_272),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_286),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_308),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_252),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_309),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_310),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_270),
.B(n_243),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_259),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_259),
.Y(n_313)
);

OAI21xp33_ASAP7_75t_SL g342 ( 
.A1(n_313),
.A2(n_281),
.B(n_285),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_251),
.B(n_268),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_315),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_251),
.B(n_268),
.C(n_256),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_246),
.A2(n_243),
.B1(n_271),
.B2(n_277),
.Y(n_316)
);

AO21x1_ASAP7_75t_L g317 ( 
.A1(n_271),
.A2(n_280),
.B(n_273),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_317),
.A2(n_260),
.B(n_267),
.Y(n_333)
);

AOI322xp5_ASAP7_75t_L g331 ( 
.A1(n_318),
.A2(n_260),
.A3(n_267),
.B1(n_284),
.B2(n_285),
.C1(n_252),
.C2(n_245),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_258),
.B(n_257),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_321),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_244),
.A2(n_247),
.B1(n_274),
.B2(n_284),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_258),
.B(n_257),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_330),
.B(n_340),
.C(n_293),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_331),
.B(n_289),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_348),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_296),
.A2(n_254),
.B1(n_266),
.B2(n_269),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_336),
.A2(n_344),
.B1(n_309),
.B2(n_301),
.Y(n_353)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_338),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_283),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_341),
.A2(n_307),
.B1(n_322),
.B2(n_290),
.Y(n_361)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_342),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_296),
.A2(n_254),
.B1(n_266),
.B2(n_255),
.Y(n_344)
);

OA21x2_ASAP7_75t_L g346 ( 
.A1(n_320),
.A2(n_285),
.B(n_245),
.Y(n_346)
);

AO22x1_ASAP7_75t_SL g366 ( 
.A1(n_346),
.A2(n_294),
.B1(n_303),
.B2(n_312),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_319),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_298),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_354),
.C(n_355),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_353),
.A2(n_347),
.B1(n_356),
.B2(n_352),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_298),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_340),
.B(n_288),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_308),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_357),
.B(n_326),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_339),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_358),
.B(n_362),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_359),
.B(n_364),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_305),
.C(n_314),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_365),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_361),
.A2(n_367),
.B1(n_370),
.B2(n_338),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_339),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_365),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_305),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_299),
.C(n_311),
.Y(n_365)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_366),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_324),
.A2(n_317),
.B1(n_318),
.B2(n_316),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_325),
.B(n_317),
.C(n_321),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_328),
.Y(n_382)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_337),
.Y(n_369)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_369),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_324),
.A2(n_310),
.B1(n_291),
.B2(n_313),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_337),
.B(n_292),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_355),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_351),
.A2(n_332),
.B(n_333),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_372),
.B(n_387),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_373),
.B(n_385),
.Y(n_390)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_375),
.Y(n_395)
);

NAND2x1_ASAP7_75t_L g376 ( 
.A(n_366),
.B(n_332),
.Y(n_376)
);

BUFx12_ASAP7_75t_L g394 ( 
.A(n_376),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_358),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g401 ( 
.A1(n_378),
.A2(n_356),
.B1(n_323),
.B2(n_343),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_382),
.B(n_360),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_362),
.Y(n_383)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_383),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_384),
.B(n_377),
.C(n_359),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g386 ( 
.A(n_370),
.Y(n_386)
);

INVx11_ASAP7_75t_L g397 ( 
.A(n_386),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_368),
.A2(n_348),
.B(n_334),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_388),
.A2(n_346),
.B1(n_352),
.B2(n_336),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_398),
.C(n_403),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_392),
.B(n_400),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_377),
.C(n_381),
.Y(n_398)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_399),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_381),
.Y(n_400)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_401),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_380),
.A2(n_367),
.B1(n_346),
.B2(n_344),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_402),
.B(n_375),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_350),
.C(n_354),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_395),
.A2(n_380),
.B1(n_387),
.B2(n_389),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_407),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_393),
.A2(n_373),
.B(n_379),
.Y(n_406)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_406),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_400),
.B(n_382),
.C(n_371),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_390),
.B(n_349),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_408),
.B(n_414),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_398),
.B(n_389),
.C(n_364),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_410),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_378),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_392),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_415),
.B(n_417),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_413),
.B(n_383),
.Y(n_417)
);

NOR3xp33_ASAP7_75t_SL g420 ( 
.A(n_412),
.B(n_379),
.C(n_334),
.Y(n_420)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_420),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_391),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_422),
.B(n_405),
.C(n_411),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_424),
.B(n_429),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_419),
.A2(n_372),
.B(n_404),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_425),
.B(n_426),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_420),
.A2(n_395),
.B1(n_402),
.B2(n_399),
.Y(n_426)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_416),
.A2(n_397),
.B(n_345),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_427),
.Y(n_430)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_418),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_428),
.A2(n_421),
.B1(n_397),
.B2(n_327),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_432),
.B(n_425),
.Y(n_435)
);

O2A1O1Ixp33_ASAP7_75t_SL g433 ( 
.A1(n_426),
.A2(n_376),
.B(n_394),
.C(n_366),
.Y(n_433)
);

AOI322xp5_ASAP7_75t_L g437 ( 
.A1(n_433),
.A2(n_394),
.A3(n_376),
.B1(n_369),
.B2(n_346),
.C1(n_341),
.C2(n_396),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_435),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_431),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_436),
.B(n_437),
.C(n_434),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_438),
.B(n_430),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_439),
.C(n_423),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_441),
.B(n_396),
.Y(n_442)
);


endmodule