module fake_jpeg_24404_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_4),
.B(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_22),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_54),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_15),
.B1(n_31),
.B2(n_20),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_53),
.B1(n_61),
.B2(n_22),
.Y(n_72)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_31),
.B1(n_15),
.B2(n_20),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_62),
.B1(n_22),
.B2(n_18),
.Y(n_73)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_55),
.Y(n_89)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_31),
.B1(n_19),
.B2(n_24),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_20),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_28),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_31),
.B1(n_17),
.B2(n_25),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_32),
.A2(n_15),
.B1(n_19),
.B2(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_68),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_63),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

AOI22x1_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_42),
.B1(n_38),
.B2(n_39),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_70),
.A2(n_72),
.B1(n_80),
.B2(n_28),
.Y(n_118)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_78),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_59),
.B1(n_46),
.B2(n_51),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_64),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_74),
.A2(n_86),
.B1(n_88),
.B2(n_59),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_25),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_76),
.A2(n_47),
.B(n_57),
.Y(n_104)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_23),
.B1(n_19),
.B2(n_24),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g107 ( 
.A(n_79),
.B(n_14),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_18),
.B1(n_17),
.B2(n_25),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_84),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_59),
.A2(n_18),
.B1(n_30),
.B2(n_29),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_91),
.Y(n_109)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_40),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_45),
.Y(n_98)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_92),
.B(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_74),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_93),
.A2(n_103),
.B1(n_112),
.B2(n_119),
.Y(n_141)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_100),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_113),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_50),
.B1(n_48),
.B2(n_61),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_111),
.B1(n_74),
.B2(n_77),
.Y(n_134)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_104),
.B(n_116),
.Y(n_135)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_66),
.B1(n_56),
.B2(n_46),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_118),
.B1(n_88),
.B2(n_77),
.Y(n_132)
);

AOI221xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_76),
.B1(n_79),
.B2(n_80),
.C(n_81),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_110),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_76),
.A2(n_66),
.B1(n_29),
.B2(n_30),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_67),
.B(n_23),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_90),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_40),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_89),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_98),
.B1(n_103),
.B2(n_100),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_128),
.B1(n_130),
.B2(n_132),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_121),
.A2(n_28),
.B1(n_101),
.B2(n_16),
.Y(n_163)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_124),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_81),
.C(n_87),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_138),
.C(n_27),
.Y(n_165)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_104),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_131),
.B(n_94),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_72),
.B(n_29),
.C(n_30),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_129),
.B(n_143),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_103),
.B1(n_116),
.B2(n_97),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_27),
.B(n_28),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_134),
.B(n_16),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_69),
.B1(n_71),
.B2(n_91),
.Y(n_137)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_119),
.B(n_36),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_78),
.B1(n_83),
.B2(n_84),
.Y(n_139)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_93),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_144),
.B(n_101),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_83),
.B1(n_84),
.B2(n_27),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_93),
.A2(n_115),
.B1(n_112),
.B2(n_96),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_146),
.A2(n_93),
.B1(n_115),
.B2(n_94),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_125),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_147),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_138),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_161),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_151),
.A2(n_141),
.B(n_144),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_142),
.B(n_128),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_112),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_155),
.B(n_162),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_39),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_163),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_165),
.Y(n_193)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_101),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_166),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_125),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_16),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_17),
.B1(n_25),
.B2(n_108),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_168),
.A2(n_124),
.B1(n_145),
.B2(n_128),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_82),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_171),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_123),
.B(n_108),
.C(n_82),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_130),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_134),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_135),
.B(n_126),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_177),
.A2(n_178),
.B(n_168),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_135),
.B(n_127),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_180),
.A2(n_188),
.B(n_152),
.Y(n_208)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_183),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_149),
.A2(n_163),
.B1(n_158),
.B2(n_153),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_182),
.A2(n_197),
.B1(n_199),
.B2(n_175),
.Y(n_225)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_184),
.A2(n_13),
.B1(n_12),
.B2(n_2),
.Y(n_218)
);

XNOR2x1_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_127),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_200),
.Y(n_201)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_198),
.Y(n_220)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_136),
.Y(n_191)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_131),
.Y(n_194)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_156),
.C(n_170),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_149),
.A2(n_120),
.B1(n_108),
.B2(n_75),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_158),
.A2(n_117),
.B1(n_95),
.B2(n_17),
.Y(n_199)
);

AND2x4_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_167),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_202),
.A2(n_213),
.B(n_178),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_208),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g204 ( 
.A1(n_187),
.A2(n_160),
.B(n_165),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_204),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_153),
.B1(n_168),
.B2(n_160),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_210),
.B(n_211),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_186),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_190),
.A2(n_168),
.B1(n_166),
.B2(n_147),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_214),
.A2(n_216),
.B1(n_219),
.B2(n_183),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_180),
.A2(n_161),
.B1(n_117),
.B2(n_95),
.Y(n_215)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

AOI22x1_ASAP7_75t_L g216 ( 
.A1(n_197),
.A2(n_95),
.B1(n_16),
.B2(n_2),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_184),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_217)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_217),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_221),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_196),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_177),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_223)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_195),
.Y(n_224)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_179),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_244),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_176),
.C(n_193),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_228),
.B(n_229),
.C(n_232),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_176),
.C(n_193),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_200),
.C(n_182),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_220),
.B(n_198),
.Y(n_237)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_240),
.A2(n_247),
.B1(n_214),
.B2(n_225),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_181),
.C(n_179),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_213),
.C(n_222),
.Y(n_252)
);

INVx13_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_202),
.B(n_199),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_241),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_254),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_208),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_255),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_263),
.C(n_265),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_230),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_202),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_258),
.A2(n_239),
.B1(n_217),
.B2(n_223),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_235),
.B1(n_242),
.B2(n_234),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_259),
.A2(n_219),
.B1(n_243),
.B2(n_3),
.Y(n_284)
);

XOR2x2_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_224),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_260),
.A2(n_267),
.B(n_253),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_227),
.B(n_224),
.Y(n_262)
);

MAJx2_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_240),
.C(n_216),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_209),
.C(n_220),
.Y(n_263)
);

BUFx4f_ASAP7_75t_SL g264 ( 
.A(n_236),
.Y(n_264)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_215),
.C(n_207),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_283),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_246),
.C(n_233),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_276),
.C(n_280),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_235),
.B(n_222),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_266),
.A2(n_226),
.B1(n_239),
.B2(n_234),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_277),
.A2(n_281),
.B1(n_284),
.B2(n_282),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_279),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_264),
.B(n_245),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_244),
.C(n_226),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_249),
.A2(n_216),
.B1(n_174),
.B2(n_236),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_282),
.B(n_277),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_249),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_261),
.A2(n_0),
.B(n_1),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_257),
.C(n_264),
.Y(n_288)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_288),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_5),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_283),
.B(n_251),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_293),
.C(n_295),
.Y(n_306)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_292),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_255),
.C(n_256),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_300),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_269),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_295)
);

XNOR2x1_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_3),
.Y(n_297)
);

XNOR2x1_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_6),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_269),
.C(n_270),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_299),
.C(n_7),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_4),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_271),
.Y(n_300)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_302),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_5),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_305),
.A2(n_310),
.B(n_290),
.Y(n_317)
);

FAx1_ASAP7_75t_SL g318 ( 
.A(n_307),
.B(n_9),
.CI(n_10),
.CON(n_318),
.SN(n_318)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_7),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_309),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_7),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_286),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_7),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_8),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_313),
.B(n_8),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_316),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_320),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_318),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_294),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_311),
.A2(n_291),
.B1(n_10),
.B2(n_11),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_305),
.C(n_11),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_304),
.B(n_9),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_322),
.A2(n_307),
.B(n_302),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_317),
.A2(n_301),
.B(n_303),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_323),
.B(n_327),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_324),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_306),
.Y(n_326)
);

MAJx2_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_319),
.C(n_314),
.Y(n_331)
);

NAND4xp25_ASAP7_75t_SL g333 ( 
.A(n_331),
.B(n_329),
.C(n_328),
.D(n_318),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_329),
.B(n_330),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_332),
.C(n_325),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_335),
.B(n_318),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_11),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_11),
.Y(n_339)
);


endmodule