module fake_jpeg_31391_n_485 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_485);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_485;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_17),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_SL g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_53),
.B(n_58),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_55),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_56),
.Y(n_158)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_20),
.B(n_13),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_66),
.B(n_67),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_20),
.B(n_15),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_34),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_80),
.B(n_85),
.Y(n_140)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_34),
.Y(n_85)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

CKINVDCx6p67_ASAP7_75t_R g124 ( 
.A(n_86),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_21),
.B(n_33),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_37),
.Y(n_122)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_97),
.B(n_98),
.Y(n_152)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

BUFx4f_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

BUFx4f_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_58),
.A2(n_21),
.B1(n_32),
.B2(n_33),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_113),
.A2(n_119),
.B1(n_141),
.B2(n_25),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_85),
.B(n_32),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_114),
.B(n_122),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_51),
.A2(n_46),
.B1(n_39),
.B2(n_45),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_115),
.A2(n_64),
.B1(n_71),
.B2(n_94),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_54),
.A2(n_35),
.B1(n_47),
.B2(n_18),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_80),
.A2(n_46),
.B1(n_45),
.B2(n_44),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_132),
.A2(n_156),
.B1(n_140),
.B2(n_37),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_55),
.B(n_18),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_136),
.B(n_25),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_86),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_140),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_56),
.A2(n_44),
.B1(n_43),
.B2(n_41),
.Y(n_141)
);

INVx6_ASAP7_75t_SL g147 ( 
.A(n_87),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_147),
.Y(n_206)
);

BUFx2_ASAP7_75t_R g148 ( 
.A(n_77),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_148),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_74),
.A2(n_43),
.B1(n_41),
.B2(n_39),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_159),
.B(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_160),
.Y(n_228)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_161),
.Y(n_239)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_162),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_63),
.B1(n_68),
.B2(n_62),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_163),
.A2(n_167),
.B1(n_197),
.B2(n_158),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_164),
.Y(n_249)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_108),
.A2(n_36),
.B(n_27),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_166),
.A2(n_208),
.B(n_4),
.Y(n_256)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_124),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_169),
.B(n_171),
.Y(n_234)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_170),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_124),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_172),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_108),
.B(n_27),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_200),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_124),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_176),
.B(n_187),
.Y(n_250)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_177),
.Y(n_254)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_179),
.B(n_189),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_180),
.A2(n_192),
.B(n_1),
.Y(n_252)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_181),
.Y(n_255)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_150),
.A2(n_36),
.B1(n_98),
.B2(n_93),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_185),
.Y(n_235)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_100),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_23),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_193),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_106),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_191),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_109),
.A2(n_23),
.B1(n_13),
.B2(n_22),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_154),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_143),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_194),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_131),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_195),
.Y(n_231)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_135),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_196),
.B(n_198),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_L g197 ( 
.A1(n_120),
.A2(n_127),
.B1(n_104),
.B2(n_116),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_134),
.B(n_83),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

BUFx24_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_128),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_99),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_167),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_133),
.B(n_82),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_203),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_111),
.B(n_75),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_209),
.Y(n_219)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_105),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_SL g245 ( 
.A1(n_205),
.A2(n_130),
.B(n_22),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_110),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_207),
.A2(n_158),
.B1(n_149),
.B2(n_125),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_152),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_116),
.B(n_0),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_117),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_211),
.Y(n_229)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_102),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_115),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_153),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_212),
.A2(n_103),
.B1(n_104),
.B2(n_156),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_216),
.A2(n_245),
.B1(n_252),
.B2(n_175),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_166),
.A2(n_132),
.B(n_145),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_220),
.A2(n_194),
.B(n_211),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_224),
.B(n_236),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_SL g236 ( 
.A(n_208),
.B(n_149),
.C(n_125),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_237),
.A2(n_253),
.B1(n_163),
.B2(n_209),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_238),
.A2(n_207),
.B1(n_164),
.B2(n_204),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_188),
.B(n_121),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_244),
.B(n_251),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_188),
.B(n_1),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_206),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_173),
.B(n_22),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_201),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_4),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_257),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_258),
.A2(n_259),
.B1(n_278),
.B2(n_284),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_201),
.B1(n_197),
.B2(n_159),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_261),
.A2(n_262),
.B1(n_269),
.B2(n_239),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_252),
.A2(n_192),
.B1(n_181),
.B2(n_168),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_234),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_268),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_265),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_266),
.A2(n_273),
.B(n_276),
.Y(n_301)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_267),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_227),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_225),
.A2(n_165),
.B1(n_205),
.B2(n_183),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_220),
.A2(n_161),
.B(n_199),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_270),
.A2(n_6),
.B(n_8),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_222),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_271),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_272),
.B(n_241),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_217),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_274),
.B(n_286),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_232),
.B(n_182),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_279),
.Y(n_300)
);

A2O1A1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_256),
.A2(n_186),
.B(n_191),
.C(n_185),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_277),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_225),
.A2(n_224),
.B1(n_213),
.B2(n_236),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_219),
.B(n_178),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_222),
.Y(n_280)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_280),
.Y(n_318)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_243),
.Y(n_281)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_281),
.Y(n_323)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_223),
.Y(n_282)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_282),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_213),
.A2(n_196),
.B1(n_195),
.B2(n_174),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_226),
.A2(n_235),
.B1(n_231),
.B2(n_254),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_285),
.A2(n_230),
.B(n_223),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_215),
.B(n_5),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_244),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_287),
.A2(n_249),
.B1(n_230),
.B2(n_214),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_240),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_291),
.Y(n_322)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_289),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_250),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_247),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_292),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_215),
.B(n_22),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_221),
.Y(n_311)
);

OA21x2_ASAP7_75t_L g294 ( 
.A1(n_248),
.A2(n_22),
.B(n_7),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_294),
.Y(n_328)
);

O2A1O1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_241),
.A2(n_235),
.B(n_237),
.C(n_218),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_295),
.Y(n_303)
);

OAI32xp33_ASAP7_75t_L g299 ( 
.A1(n_269),
.A2(n_218),
.A3(n_219),
.B1(n_253),
.B2(n_251),
.Y(n_299)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_302),
.B(n_308),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_233),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_306),
.B(n_327),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_266),
.A2(n_239),
.B(n_221),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_307),
.A2(n_276),
.B(n_270),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_275),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_309),
.A2(n_258),
.B1(n_281),
.B2(n_260),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_315),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_261),
.A2(n_246),
.B1(n_242),
.B2(n_228),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_312),
.A2(n_292),
.B1(n_289),
.B2(n_294),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_313),
.A2(n_9),
.B(n_11),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_279),
.B(n_6),
.Y(n_319)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_259),
.A2(n_214),
.B1(n_7),
.B2(n_8),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_321),
.A2(n_286),
.B1(n_265),
.B2(n_280),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_277),
.Y(n_325)
);

BUFx2_ASAP7_75t_SL g351 ( 
.A(n_325),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_283),
.B(n_214),
.C(n_8),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_287),
.C(n_283),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_263),
.B(n_267),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_330),
.A2(n_273),
.B(n_294),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_304),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_331),
.B(n_336),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_332),
.A2(n_359),
.B(n_361),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_333),
.B(n_311),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_290),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_334),
.B(n_340),
.C(n_357),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_304),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_337),
.Y(n_383)
);

BUFx12_ASAP7_75t_L g338 ( 
.A(n_298),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g376 ( 
.A(n_338),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_278),
.C(n_293),
.Y(n_340)
);

NAND3xp33_ASAP7_75t_L g341 ( 
.A(n_322),
.B(n_291),
.C(n_268),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_341),
.B(n_343),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_322),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_300),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_344),
.A2(n_300),
.B(n_302),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_345),
.A2(n_347),
.B1(n_355),
.B2(n_321),
.Y(n_372)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_317),
.Y(n_346)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_346),
.Y(n_367)
);

OAI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_308),
.A2(n_260),
.B1(n_295),
.B2(n_262),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_317),
.Y(n_348)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_348),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_350),
.A2(n_354),
.B1(n_309),
.B2(n_303),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_307),
.A2(n_295),
.B(n_272),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_352),
.A2(n_332),
.B(n_339),
.Y(n_388)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_329),
.Y(n_353)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_353),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_296),
.A2(n_294),
.B1(n_284),
.B2(n_265),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_318),
.Y(n_356)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_356),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_271),
.C(n_282),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_9),
.C(n_10),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_358),
.B(n_330),
.C(n_319),
.Y(n_380)
);

OA21x2_ASAP7_75t_L g361 ( 
.A1(n_303),
.A2(n_9),
.B(n_11),
.Y(n_361)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_362),
.Y(n_389)
);

XOR2x2_ASAP7_75t_L g364 ( 
.A(n_334),
.B(n_299),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_364),
.B(n_369),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_366),
.A2(n_382),
.B1(n_387),
.B2(n_336),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_296),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_370),
.B(n_379),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_351),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_371),
.B(n_372),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_301),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_373),
.B(n_374),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_333),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_335),
.B(n_301),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_381),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_335),
.A2(n_328),
.B1(n_323),
.B2(n_297),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_349),
.A2(n_328),
.B1(n_323),
.B2(n_297),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_343),
.A2(n_305),
.B1(n_315),
.B2(n_320),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_384),
.A2(n_388),
.B(n_337),
.Y(n_395)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_346),
.Y(n_386)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_386),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_355),
.A2(n_305),
.B1(n_312),
.B2(n_316),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_375),
.B(n_370),
.C(n_374),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_390),
.B(n_409),
.C(n_388),
.Y(n_417)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_392),
.Y(n_414)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_377),
.Y(n_394)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_394),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_395),
.B(n_410),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_396),
.A2(n_407),
.B1(n_361),
.B2(n_348),
.Y(n_425)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_367),
.Y(n_398)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_398),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_331),
.Y(n_399)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_399),
.Y(n_429)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_368),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_401),
.Y(n_413)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_378),
.Y(n_401)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_385),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_408),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_373),
.B(n_352),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_406),
.B(n_364),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_383),
.A2(n_344),
.B1(n_342),
.B2(n_354),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_382),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_375),
.B(n_357),
.C(n_342),
.Y(n_409)
);

FAx1_ASAP7_75t_SL g410 ( 
.A(n_379),
.B(n_358),
.CI(n_350),
.CON(n_410),
.SN(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_376),
.Y(n_411)
);

INVxp33_ASAP7_75t_SL g424 ( 
.A(n_411),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_412),
.B(n_425),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_390),
.B(n_369),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_415),
.B(n_402),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_404),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_416),
.B(n_418),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_417),
.B(n_421),
.C(n_422),
.Y(n_431)
);

AOI31xp33_ASAP7_75t_L g418 ( 
.A1(n_410),
.A2(n_383),
.A3(n_314),
.B(n_363),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_372),
.C(n_381),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_397),
.B(n_380),
.C(n_387),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_389),
.A2(n_359),
.B1(n_363),
.B2(n_353),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_395),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_397),
.B(n_318),
.C(n_298),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_427),
.B(n_405),
.C(n_393),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_314),
.Y(n_430)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_430),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_432),
.B(n_433),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_424),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_417),
.B(n_415),
.C(n_422),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_436),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_419),
.A2(n_414),
.B1(n_429),
.B2(n_403),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_428),
.B(n_376),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_440),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_421),
.B(n_405),
.C(n_402),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_413),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_441),
.B(n_442),
.Y(n_453)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_420),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_443),
.B(n_444),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_427),
.B(n_393),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_445),
.B(n_412),
.Y(n_455)
);

XOR2x1_ASAP7_75t_SL g446 ( 
.A(n_438),
.B(n_410),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_446),
.B(n_456),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_435),
.A2(n_407),
.B(n_423),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_447),
.A2(n_454),
.B(n_313),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_437),
.A2(n_411),
.B(n_424),
.Y(n_449)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_449),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_433),
.Y(n_452)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_452),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_431),
.A2(n_411),
.B(n_426),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_455),
.B(n_431),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_438),
.A2(n_396),
.B1(n_391),
.B2(n_406),
.Y(n_456)
);

AOI211xp5_ASAP7_75t_L g458 ( 
.A1(n_440),
.A2(n_361),
.B(n_445),
.C(n_325),
.Y(n_458)
);

OA21x2_ASAP7_75t_L g464 ( 
.A1(n_458),
.A2(n_329),
.B(n_324),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_452),
.Y(n_459)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_459),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_460),
.B(n_462),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_464),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_450),
.B(n_434),
.C(n_432),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_448),
.A2(n_316),
.B(n_324),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_465),
.A2(n_453),
.B(n_447),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_451),
.B(n_310),
.C(n_338),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_467),
.B(n_456),
.C(n_455),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_469),
.B(n_474),
.Y(n_475)
);

AO21x2_ASAP7_75t_L g470 ( 
.A1(n_464),
.A2(n_446),
.B(n_458),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_470),
.A2(n_467),
.B(n_457),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_473),
.A2(n_463),
.B(n_468),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_476),
.A2(n_478),
.B(n_470),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_471),
.B(n_466),
.Y(n_477)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_477),
.Y(n_480)
);

OAI21x1_ASAP7_75t_L g481 ( 
.A1(n_479),
.A2(n_475),
.B(n_472),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_481),
.B(n_480),
.Y(n_482)
);

AO21x1_ASAP7_75t_L g483 ( 
.A1(n_482),
.A2(n_459),
.B(n_338),
.Y(n_483)
);

OAI31xp33_ASAP7_75t_L g484 ( 
.A1(n_483),
.A2(n_310),
.A3(n_11),
.B(n_12),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_484),
.A2(n_12),
.B(n_377),
.Y(n_485)
);


endmodule