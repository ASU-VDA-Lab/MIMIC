module real_aes_9878_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
OAI222xp33_ASAP7_75t_L g602 ( .A1(n_0), .A2(n_39), .B1(n_177), .B2(n_603), .C1(n_605), .C2(n_607), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_0), .A2(n_177), .B1(n_639), .B2(n_641), .C(n_643), .Y(n_638) );
CKINVDCx5p33_ASAP7_75t_R g862 ( .A(n_1), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_2), .A2(n_13), .B1(n_527), .B2(n_662), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_2), .A2(n_13), .B1(n_702), .B2(n_703), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_3), .A2(n_74), .B1(n_1239), .B2(n_1249), .Y(n_1248) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_4), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_4), .B(n_222), .Y(n_406) );
INVx1_ASAP7_75t_L g466 ( .A(n_4), .Y(n_466) );
AND2x2_ASAP7_75t_L g472 ( .A(n_4), .B(n_465), .Y(n_472) );
INVx1_ASAP7_75t_L g1166 ( .A(n_5), .Y(n_1166) );
OAI22xp5_ASAP7_75t_L g1192 ( .A1(n_5), .A2(n_213), .B1(n_337), .B2(n_877), .Y(n_1192) );
INVx1_ASAP7_75t_L g1529 ( .A(n_6), .Y(n_1529) );
AOI22xp33_ASAP7_75t_L g1556 ( .A1(n_6), .A2(n_88), .B1(n_1557), .B2(n_1558), .Y(n_1556) );
AOI22xp33_ASAP7_75t_SL g1184 ( .A1(n_7), .A2(n_53), .B1(n_854), .B2(n_1181), .Y(n_1184) );
INVx1_ASAP7_75t_L g1209 ( .A(n_7), .Y(n_1209) );
OAI221xp5_ASAP7_75t_SL g830 ( .A1(n_8), .A2(n_58), .B1(n_831), .B2(n_833), .C(n_834), .Y(n_830) );
AOI221xp5_ASAP7_75t_L g865 ( .A1(n_8), .A2(n_114), .B1(n_590), .B2(n_866), .C(n_870), .Y(n_865) );
INVx1_ASAP7_75t_L g855 ( .A(n_9), .Y(n_855) );
OAI221xp5_ASAP7_75t_L g1525 ( .A1(n_10), .A2(n_243), .B1(n_719), .B2(n_1035), .C(n_1526), .Y(n_1525) );
OAI22xp33_ASAP7_75t_L g1548 ( .A1(n_10), .A2(n_243), .B1(n_337), .B2(n_877), .Y(n_1548) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_11), .Y(n_794) );
AOI221xp5_ASAP7_75t_L g902 ( .A1(n_12), .A2(n_116), .B1(n_374), .B2(n_556), .C(n_883), .Y(n_902) );
AOI22xp33_ASAP7_75t_SL g920 ( .A1(n_12), .A2(n_170), .B1(n_440), .B2(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g852 ( .A(n_14), .Y(n_852) );
INVx1_ASAP7_75t_L g1064 ( .A(n_15), .Y(n_1064) );
AOI22xp5_ASAP7_75t_L g1242 ( .A1(n_16), .A2(n_79), .B1(n_1235), .B2(n_1239), .Y(n_1242) );
INVxp33_ASAP7_75t_L g492 ( .A(n_17), .Y(n_492) );
AOI221xp5_ASAP7_75t_L g566 ( .A1(n_17), .A2(n_157), .B1(n_567), .B2(n_568), .C(n_569), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_18), .A2(n_117), .B1(n_1019), .B2(n_1020), .Y(n_1018) );
INVxp67_ASAP7_75t_SL g1044 ( .A(n_18), .Y(n_1044) );
INVx1_ASAP7_75t_L g1023 ( .A(n_19), .Y(n_1023) );
INVx1_ASAP7_75t_L g1531 ( .A(n_20), .Y(n_1531) );
AOI221xp5_ASAP7_75t_L g1555 ( .A1(n_20), .A2(n_249), .B1(n_761), .B2(n_968), .C(n_1201), .Y(n_1555) );
OAI221xp5_ASAP7_75t_L g718 ( .A1(n_21), .A2(n_191), .B1(n_719), .B2(n_720), .C(n_721), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_21), .A2(n_191), .B1(n_756), .B2(n_757), .Y(n_755) );
INVx1_ASAP7_75t_L g795 ( .A(n_22), .Y(n_795) );
INVx1_ASAP7_75t_L g1147 ( .A(n_23), .Y(n_1147) );
OR2x2_ASAP7_75t_L g320 ( .A(n_24), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g332 ( .A(n_24), .Y(n_332) );
INVx1_ASAP7_75t_L g578 ( .A(n_25), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g1057 ( .A1(n_26), .A2(n_118), .B1(n_878), .B2(n_1058), .Y(n_1057) );
OAI221xp5_ASAP7_75t_L g1090 ( .A1(n_26), .A2(n_118), .B1(n_495), .B2(n_720), .C(n_721), .Y(n_1090) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_27), .A2(n_47), .B1(n_344), .B2(n_349), .C(n_351), .Y(n_343) );
INVx1_ASAP7_75t_L g468 ( .A(n_27), .Y(n_468) );
OAI221xp5_ASAP7_75t_L g838 ( .A1(n_28), .A2(n_73), .B1(n_503), .B2(n_719), .C(n_839), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_28), .A2(n_73), .B1(n_877), .B2(n_878), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g1241 ( .A1(n_29), .A2(n_141), .B1(n_1223), .B2(n_1231), .Y(n_1241) );
INVx1_ASAP7_75t_L g1021 ( .A(n_30), .Y(n_1021) );
AOI22xp33_ASAP7_75t_SL g1011 ( .A1(n_31), .A2(n_153), .B1(n_563), .B2(n_1012), .Y(n_1011) );
INVxp33_ASAP7_75t_SL g1033 ( .A(n_31), .Y(n_1033) );
BUFx2_ASAP7_75t_L g314 ( .A(n_32), .Y(n_314) );
OR2x2_ASAP7_75t_L g405 ( .A(n_32), .B(n_406), .Y(n_405) );
BUFx2_ASAP7_75t_L g409 ( .A(n_32), .Y(n_409) );
INVx1_ASAP7_75t_L g462 ( .A(n_32), .Y(n_462) );
AOI221xp5_ASAP7_75t_L g779 ( .A1(n_33), .A2(n_43), .B1(n_569), .B2(n_780), .C(n_782), .Y(n_779) );
INVx1_ASAP7_75t_L g804 ( .A(n_33), .Y(n_804) );
INVx1_ASAP7_75t_L g1274 ( .A(n_34), .Y(n_1274) );
INVx1_ASAP7_75t_L g1520 ( .A(n_35), .Y(n_1520) );
AOI221xp5_ASAP7_75t_L g1549 ( .A1(n_35), .A2(n_143), .B1(n_1020), .B2(n_1550), .C(n_1552), .Y(n_1549) );
INVx1_ASAP7_75t_L g1074 ( .A(n_36), .Y(n_1074) );
INVx1_ASAP7_75t_L g736 ( .A(n_37), .Y(n_736) );
AOI22xp33_ASAP7_75t_SL g663 ( .A1(n_38), .A2(n_85), .B1(n_653), .B2(n_655), .Y(n_663) );
INVx1_ASAP7_75t_L g699 ( .A(n_38), .Y(n_699) );
INVx1_ASAP7_75t_L g644 ( .A(n_39), .Y(n_644) );
INVx1_ASAP7_75t_L g1300 ( .A(n_40), .Y(n_1300) );
INVxp67_ASAP7_75t_SL g844 ( .A(n_41), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_41), .A2(n_178), .B1(n_885), .B2(n_886), .Y(n_884) );
AOI22xp33_ASAP7_75t_SL g1475 ( .A1(n_42), .A2(n_115), .B1(n_934), .B2(n_1476), .Y(n_1475) );
AOI221xp5_ASAP7_75t_L g1495 ( .A1(n_42), .A2(n_75), .B1(n_381), .B2(n_1496), .C(n_1498), .Y(n_1495) );
INVx1_ASAP7_75t_L g802 ( .A(n_43), .Y(n_802) );
OAI22xp33_ASAP7_75t_R g961 ( .A1(n_44), .A2(n_259), .B1(n_878), .B2(n_962), .Y(n_961) );
OAI221xp5_ASAP7_75t_L g982 ( .A1(n_44), .A2(n_259), .B1(n_503), .B2(n_719), .C(n_839), .Y(n_982) );
INVx1_ASAP7_75t_L g533 ( .A(n_45), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g652 ( .A1(n_46), .A2(n_230), .B1(n_653), .B2(n_655), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_46), .A2(n_190), .B1(n_562), .B2(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g479 ( .A(n_47), .Y(n_479) );
INVx1_ASAP7_75t_L g401 ( .A(n_48), .Y(n_401) );
INVx1_ASAP7_75t_L g974 ( .A(n_49), .Y(n_974) );
INVx1_ASAP7_75t_L g1024 ( .A(n_50), .Y(n_1024) );
INVxp67_ASAP7_75t_SL g908 ( .A(n_51), .Y(n_908) );
AOI221xp5_ASAP7_75t_L g933 ( .A1(n_51), .A2(n_110), .B1(n_659), .B2(n_934), .C(n_936), .Y(n_933) );
INVxp67_ASAP7_75t_L g713 ( .A(n_52), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g753 ( .A1(n_52), .A2(n_159), .B1(n_359), .B2(n_590), .C(n_700), .Y(n_753) );
INVx1_ASAP7_75t_L g1191 ( .A(n_53), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_54), .A2(n_216), .B1(n_384), .B2(n_387), .Y(n_1072) );
INVxp67_ASAP7_75t_SL g1081 ( .A(n_54), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1222 ( .A1(n_55), .A2(n_106), .B1(n_1223), .B2(n_1231), .Y(n_1222) );
INVxp67_ASAP7_75t_SL g911 ( .A(n_56), .Y(n_911) );
OAI211xp5_ASAP7_75t_SL g925 ( .A1(n_56), .A2(n_537), .B(n_725), .C(n_926), .Y(n_925) );
INVx1_ASAP7_75t_L g913 ( .A(n_57), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_58), .A2(n_133), .B1(n_349), .B2(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g1070 ( .A(n_59), .Y(n_1070) );
XNOR2x2_ASAP7_75t_L g645 ( .A(n_60), .B(n_646), .Y(n_645) );
INVxp33_ASAP7_75t_L g724 ( .A(n_61), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_61), .A2(n_235), .B1(n_567), .B2(n_763), .Y(n_762) );
INVxp33_ASAP7_75t_SL g846 ( .A(n_62), .Y(n_846) );
AOI221xp5_ASAP7_75t_L g881 ( .A1(n_62), .A2(n_238), .B1(n_606), .B2(n_882), .C(n_883), .Y(n_881) );
OAI222xp33_ASAP7_75t_L g609 ( .A1(n_63), .A2(n_150), .B1(n_228), .B2(n_576), .C1(n_610), .C2(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g616 ( .A(n_63), .Y(n_616) );
CKINVDCx5p33_ASAP7_75t_R g1543 ( .A(n_64), .Y(n_1543) );
AOI221xp5_ASAP7_75t_L g953 ( .A1(n_65), .A2(n_149), .B1(n_954), .B2(n_955), .C(n_956), .Y(n_953) );
INVxp33_ASAP7_75t_L g979 ( .A(n_65), .Y(n_979) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_66), .A2(n_190), .B1(n_658), .B2(n_659), .Y(n_657) );
AOI21xp33_ASAP7_75t_L g687 ( .A1(n_66), .A2(n_381), .B(n_688), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g1059 ( .A1(n_67), .A2(n_242), .B1(n_1020), .B2(n_1060), .C(n_1062), .Y(n_1059) );
INVxp33_ASAP7_75t_L g1095 ( .A(n_67), .Y(n_1095) );
INVx1_ASAP7_75t_L g1053 ( .A(n_68), .Y(n_1053) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_69), .A2(n_170), .B1(n_791), .B2(n_900), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_69), .A2(n_116), .B1(n_455), .B2(n_923), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_70), .A2(n_151), .B1(n_563), .B2(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g635 ( .A(n_70), .Y(n_635) );
INVxp33_ASAP7_75t_SL g1104 ( .A(n_71), .Y(n_1104) );
AOI221xp5_ASAP7_75t_L g1138 ( .A1(n_71), .A2(n_267), .B1(n_763), .B2(n_1139), .C(n_1140), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_72), .A2(n_98), .B1(n_387), .B2(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g621 ( .A(n_72), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g1471 ( .A1(n_75), .A2(n_134), .B1(n_1472), .B2(n_1473), .Y(n_1471) );
AOI22xp5_ASAP7_75t_L g1251 ( .A1(n_76), .A2(n_123), .B1(n_1223), .B2(n_1231), .Y(n_1251) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_77), .A2(n_233), .B1(n_457), .B2(n_1179), .Y(n_1185) );
INVx1_ASAP7_75t_L g1199 ( .A(n_77), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_78), .A2(n_104), .B1(n_592), .B2(n_900), .Y(n_903) );
INVxp67_ASAP7_75t_SL g941 ( .A(n_78), .Y(n_941) );
INVx1_ASAP7_75t_L g1175 ( .A(n_80), .Y(n_1175) );
AOI221xp5_ASAP7_75t_L g1193 ( .A1(n_80), .A2(n_111), .B1(n_763), .B2(n_1012), .C(n_1194), .Y(n_1193) );
AOI221xp5_ASAP7_75t_L g904 ( .A1(n_81), .A2(n_171), .B1(n_590), .B2(n_791), .C(n_905), .Y(n_904) );
INVxp33_ASAP7_75t_SL g929 ( .A(n_81), .Y(n_929) );
AOI22xp33_ASAP7_75t_SL g1478 ( .A1(n_82), .A2(n_92), .B1(n_1479), .B2(n_1480), .Y(n_1478) );
INVx1_ASAP7_75t_L g1494 ( .A(n_82), .Y(n_1494) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_83), .A2(n_247), .B1(n_870), .B2(n_972), .Y(n_971) );
INVxp67_ASAP7_75t_SL g992 ( .A(n_83), .Y(n_992) );
CKINVDCx5p33_ASAP7_75t_R g1174 ( .A(n_84), .Y(n_1174) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_85), .B(n_396), .Y(n_678) );
INVx1_ASAP7_75t_L g675 ( .A(n_86), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_86), .A2(n_139), .B1(n_685), .B2(n_688), .Y(n_692) );
INVx1_ASAP7_75t_L g1469 ( .A(n_87), .Y(n_1469) );
AOI221xp5_ASAP7_75t_L g1488 ( .A1(n_87), .A2(n_112), .B1(n_784), .B2(n_1489), .C(n_1491), .Y(n_1488) );
INVx1_ASAP7_75t_L g1537 ( .A(n_88), .Y(n_1537) );
OA22x2_ASAP7_75t_L g944 ( .A1(n_89), .A2(n_945), .B1(n_946), .B2(n_997), .Y(n_944) );
CKINVDCx16_ASAP7_75t_R g997 ( .A(n_89), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g1477 ( .A1(n_90), .A2(n_236), .B1(n_854), .B2(n_934), .Y(n_1477) );
INVx1_ASAP7_75t_L g1504 ( .A(n_90), .Y(n_1504) );
INVx1_ASAP7_75t_L g321 ( .A(n_91), .Y(n_321) );
INVx1_ASAP7_75t_L g364 ( .A(n_91), .Y(n_364) );
INVx1_ASAP7_75t_L g1503 ( .A(n_92), .Y(n_1503) );
INVx1_ASAP7_75t_L g1047 ( .A(n_93), .Y(n_1047) );
CKINVDCx5p33_ASAP7_75t_R g948 ( .A(n_94), .Y(n_948) );
INVx1_ASAP7_75t_L g748 ( .A(n_95), .Y(n_748) );
INVx1_ASAP7_75t_L g667 ( .A(n_96), .Y(n_667) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_96), .A2(n_694), .B(n_695), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_97), .A2(n_277), .B1(n_327), .B2(n_337), .Y(n_326) );
INVx1_ASAP7_75t_L g422 ( .A(n_97), .Y(n_422) );
INVx1_ASAP7_75t_L g618 ( .A(n_98), .Y(n_618) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_99), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g555 ( .A1(n_99), .A2(n_225), .B1(n_553), .B2(n_556), .C(n_557), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g1523 ( .A(n_100), .Y(n_1523) );
AOI22xp5_ASAP7_75t_L g1247 ( .A1(n_101), .A2(n_126), .B1(n_1223), .B2(n_1231), .Y(n_1247) );
INVx1_ASAP7_75t_L g1457 ( .A(n_101), .Y(n_1457) );
AOI22xp33_ASAP7_75t_L g1509 ( .A1(n_101), .A2(n_1510), .B1(n_1514), .B2(n_1564), .Y(n_1509) );
AOI22xp33_ASAP7_75t_L g1264 ( .A1(n_102), .A2(n_229), .B1(n_1223), .B2(n_1231), .Y(n_1264) );
INVxp33_ASAP7_75t_SL g489 ( .A(n_103), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_103), .A2(n_128), .B1(n_571), .B2(n_572), .Y(n_570) );
INVxp33_ASAP7_75t_L g930 ( .A(n_104), .Y(n_930) );
INVxp67_ASAP7_75t_L g717 ( .A(n_105), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_105), .A2(n_205), .B1(n_349), .B2(n_606), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g1234 ( .A1(n_107), .A2(n_144), .B1(n_1235), .B2(n_1239), .Y(n_1234) );
AOI221xp5_ASAP7_75t_L g787 ( .A1(n_108), .A2(n_169), .B1(n_557), .B2(n_568), .C(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g815 ( .A(n_108), .Y(n_815) );
INVx1_ASAP7_75t_L g1257 ( .A(n_109), .Y(n_1257) );
OAI211xp5_ASAP7_75t_SL g897 ( .A1(n_110), .A2(n_319), .B(n_898), .C(n_906), .Y(n_897) );
INVx1_ASAP7_75t_L g1170 ( .A(n_111), .Y(n_1170) );
INVx1_ASAP7_75t_L g1465 ( .A(n_112), .Y(n_1465) );
CKINVDCx5p33_ASAP7_75t_R g1521 ( .A(n_113), .Y(n_1521) );
INVxp33_ASAP7_75t_SL g836 ( .A(n_114), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g1500 ( .A1(n_115), .A2(n_134), .B1(n_384), .B2(n_1501), .Y(n_1500) );
INVxp33_ASAP7_75t_L g1038 ( .A(n_117), .Y(n_1038) );
INVx1_ASAP7_75t_L g1013 ( .A(n_119), .Y(n_1013) );
INVx1_ASAP7_75t_L g768 ( .A(n_120), .Y(n_768) );
INVx1_ASAP7_75t_L g528 ( .A(n_121), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_121), .A2(n_189), .B1(n_560), .B2(n_563), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g778 ( .A(n_122), .Y(n_778) );
OAI22xp33_ASAP7_75t_L g785 ( .A1(n_124), .A2(n_251), .B1(n_576), .B2(n_756), .Y(n_785) );
OAI221xp5_ASAP7_75t_L g807 ( .A1(n_124), .A2(n_251), .B1(n_503), .B2(n_720), .C(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g288 ( .A(n_125), .Y(n_288) );
AO22x1_ASAP7_75t_SL g1254 ( .A1(n_127), .A2(n_237), .B1(n_1223), .B2(n_1231), .Y(n_1254) );
INVxp33_ASAP7_75t_SL g493 ( .A(n_128), .Y(n_493) );
INVx1_ASAP7_75t_L g1121 ( .A(n_129), .Y(n_1121) );
AOI221xp5_ASAP7_75t_L g1132 ( .A1(n_129), .A2(n_224), .B1(n_763), .B2(n_1133), .C(n_1135), .Y(n_1132) );
INVx1_ASAP7_75t_L g1298 ( .A(n_130), .Y(n_1298) );
AO221x2_ASAP7_75t_L g1268 ( .A1(n_131), .A2(n_269), .B1(n_1249), .B2(n_1269), .C(n_1270), .Y(n_1268) );
INVx1_ASAP7_75t_L g372 ( .A(n_132), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_132), .A2(n_180), .B1(n_454), .B2(n_457), .Y(n_453) );
INVxp33_ASAP7_75t_SL g835 ( .A(n_133), .Y(n_835) );
AOI221xp5_ASAP7_75t_L g967 ( .A1(n_135), .A2(n_226), .B1(n_968), .B2(n_969), .C(n_970), .Y(n_967) );
INVxp67_ASAP7_75t_SL g986 ( .A(n_135), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_136), .A2(n_161), .B1(n_1181), .B2(n_1182), .Y(n_1180) );
AOI221xp5_ASAP7_75t_L g1200 ( .A1(n_136), .A2(n_223), .B1(n_381), .B2(n_968), .C(n_1201), .Y(n_1200) );
CKINVDCx5p33_ASAP7_75t_R g1539 ( .A(n_137), .Y(n_1539) );
INVx1_ASAP7_75t_L g1148 ( .A(n_138), .Y(n_1148) );
INVx1_ASAP7_75t_L g671 ( .A(n_139), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_140), .A2(n_200), .B1(n_381), .B2(n_568), .C(n_594), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_140), .A2(n_151), .B1(n_630), .B2(n_632), .C(n_634), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_142), .A2(n_255), .B1(n_384), .B2(n_387), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_142), .A2(n_154), .B1(n_440), .B2(n_445), .Y(n_439) );
INVx1_ASAP7_75t_L g1524 ( .A(n_143), .Y(n_1524) );
INVx1_ASAP7_75t_L g482 ( .A(n_144), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g1515 ( .A1(n_145), .A2(n_1516), .B1(n_1562), .B2(n_1563), .Y(n_1515) );
CKINVDCx5p33_ASAP7_75t_R g1562 ( .A(n_145), .Y(n_1562) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_146), .A2(n_207), .B1(n_327), .B2(n_878), .Y(n_1014) );
OAI221xp5_ASAP7_75t_L g1034 ( .A1(n_146), .A2(n_207), .B1(n_495), .B2(n_721), .C(n_1035), .Y(n_1034) );
CKINVDCx5p33_ASAP7_75t_R g1542 ( .A(n_147), .Y(n_1542) );
AOI221xp5_ASAP7_75t_L g586 ( .A1(n_148), .A2(n_164), .B1(n_587), .B2(n_589), .C(n_590), .Y(n_586) );
INVx1_ASAP7_75t_L g619 ( .A(n_148), .Y(n_619) );
INVxp33_ASAP7_75t_L g981 ( .A(n_149), .Y(n_981) );
INVx1_ASAP7_75t_L g623 ( .A(n_150), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_152), .A2(n_223), .B1(n_655), .B2(n_1179), .Y(n_1178) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_152), .A2(n_161), .B1(n_954), .B2(n_1205), .Y(n_1204) );
INVxp33_ASAP7_75t_L g1029 ( .A(n_153), .Y(n_1029) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_154), .A2(n_163), .B1(n_374), .B2(n_377), .C(n_381), .Y(n_373) );
INVx1_ASAP7_75t_L g1482 ( .A(n_155), .Y(n_1482) );
AOI22xp33_ASAP7_75t_L g1128 ( .A1(n_156), .A2(n_232), .B1(n_478), .B2(n_1129), .Y(n_1128) );
OAI22xp5_ASAP7_75t_L g1150 ( .A1(n_156), .A2(n_250), .B1(n_1151), .B2(n_1153), .Y(n_1150) );
INVxp33_ASAP7_75t_L g490 ( .A(n_157), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g1265 ( .A1(n_158), .A2(n_265), .B1(n_1235), .B2(n_1239), .Y(n_1265) );
INVxp67_ASAP7_75t_L g716 ( .A(n_159), .Y(n_716) );
CKINVDCx5p33_ASAP7_75t_R g1468 ( .A(n_160), .Y(n_1468) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_162), .Y(n_649) );
AOI22xp33_ASAP7_75t_SL g432 ( .A1(n_163), .A2(n_255), .B1(n_433), .B2(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g628 ( .A(n_164), .Y(n_628) );
INVx1_ASAP7_75t_L g398 ( .A(n_165), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_165), .A2(n_199), .B1(n_440), .B2(n_450), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_166), .A2(n_248), .B1(n_572), .B2(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g820 ( .A(n_166), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_167), .A2(n_203), .B1(n_374), .B2(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g800 ( .A(n_167), .Y(n_800) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_168), .Y(n_601) );
INVx1_ASAP7_75t_L g817 ( .A(n_169), .Y(n_817) );
OAI21xp33_ASAP7_75t_SL g917 ( .A1(n_171), .A2(n_918), .B(n_919), .Y(n_917) );
INVx1_ASAP7_75t_L g747 ( .A(n_172), .Y(n_747) );
INVx1_ASAP7_75t_L g1025 ( .A(n_173), .Y(n_1025) );
INVxp67_ASAP7_75t_L g730 ( .A(n_174), .Y(n_730) );
AOI221xp5_ASAP7_75t_L g759 ( .A1(n_174), .A2(n_241), .B1(n_346), .B2(n_760), .C(n_761), .Y(n_759) );
CKINVDCx5p33_ASAP7_75t_R g775 ( .A(n_175), .Y(n_775) );
OAI221xp5_ASAP7_75t_L g494 ( .A1(n_176), .A2(n_278), .B1(n_495), .B2(n_500), .C(n_503), .Y(n_494) );
OAI22xp33_ASAP7_75t_L g573 ( .A1(n_176), .A2(n_278), .B1(n_574), .B2(n_576), .Y(n_573) );
INVxp67_ASAP7_75t_SL g849 ( .A(n_178), .Y(n_849) );
INVx1_ASAP7_75t_L g1112 ( .A(n_179), .Y(n_1112) );
INVx1_ASAP7_75t_L g394 ( .A(n_180), .Y(n_394) );
INVx1_ASAP7_75t_L g959 ( .A(n_181), .Y(n_959) );
INVx1_ASAP7_75t_L g1188 ( .A(n_182), .Y(n_1188) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_183), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g1071 ( .A1(n_184), .A2(n_268), .B1(n_556), .B2(n_557), .C(n_571), .Y(n_1071) );
INVxp33_ASAP7_75t_SL g1084 ( .A(n_184), .Y(n_1084) );
INVx1_ASAP7_75t_L g484 ( .A(n_185), .Y(n_484) );
INVx1_ASAP7_75t_L g1056 ( .A(n_186), .Y(n_1056) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_187), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_187), .B(n_288), .Y(n_1230) );
AND3x2_ASAP7_75t_L g1236 ( .A(n_187), .B(n_288), .C(n_1227), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_188), .A2(n_253), .B1(n_1239), .B2(n_1249), .Y(n_1252) );
INVxp67_ASAP7_75t_SL g514 ( .A(n_189), .Y(n_514) );
INVx1_ASAP7_75t_L g951 ( .A(n_192), .Y(n_951) );
INVx2_ASAP7_75t_L g301 ( .A(n_193), .Y(n_301) );
INVx1_ASAP7_75t_L g907 ( .A(n_194), .Y(n_907) );
XOR2xp5_ASAP7_75t_L g1050 ( .A(n_195), .B(n_1051), .Y(n_1050) );
INVx1_ASAP7_75t_L g1067 ( .A(n_196), .Y(n_1067) );
XNOR2x2_ASAP7_75t_L g1100 ( .A(n_197), .B(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g857 ( .A(n_198), .Y(n_857) );
INVx1_ASAP7_75t_L g317 ( .A(n_199), .Y(n_317) );
INVx1_ASAP7_75t_L g637 ( .A(n_200), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g1172 ( .A(n_201), .Y(n_1172) );
INVxp67_ASAP7_75t_L g707 ( .A(n_202), .Y(n_707) );
INVx1_ASAP7_75t_L g805 ( .A(n_203), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g1545 ( .A(n_204), .Y(n_1545) );
INVxp67_ASAP7_75t_L g712 ( .A(n_205), .Y(n_712) );
INVx1_ASAP7_75t_L g827 ( .A(n_206), .Y(n_827) );
XNOR2xp5_ASAP7_75t_L g769 ( .A(n_208), .B(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g1227 ( .A(n_209), .Y(n_1227) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_210), .A2(n_272), .B1(n_400), .B2(n_557), .C(n_1017), .Y(n_1016) );
INVxp67_ASAP7_75t_SL g1042 ( .A(n_210), .Y(n_1042) );
INVx1_ASAP7_75t_L g1118 ( .A(n_211), .Y(n_1118) );
INVx1_ASAP7_75t_L g1106 ( .A(n_212), .Y(n_1106) );
INVx1_ASAP7_75t_L g1167 ( .A(n_213), .Y(n_1167) );
OAI211xp5_ASAP7_75t_SL g909 ( .A1(n_214), .A2(n_888), .B(n_910), .C(n_915), .Y(n_909) );
INVx1_ASAP7_75t_L g939 ( .A(n_214), .Y(n_939) );
INVx1_ASAP7_75t_L g966 ( .A(n_215), .Y(n_966) );
INVxp33_ASAP7_75t_L g1083 ( .A(n_216), .Y(n_1083) );
INVx1_ASAP7_75t_L g957 ( .A(n_217), .Y(n_957) );
INVx1_ASAP7_75t_L g1075 ( .A(n_218), .Y(n_1075) );
INVx1_ASAP7_75t_L g676 ( .A(n_219), .Y(n_676) );
OAI211xp5_ASAP7_75t_L g697 ( .A1(n_219), .A2(n_610), .B(n_698), .C(n_704), .Y(n_697) );
INVx1_ASAP7_75t_L g536 ( .A(n_220), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g1271 ( .A(n_221), .Y(n_1271) );
INVx1_ASAP7_75t_L g303 ( .A(n_222), .Y(n_303) );
INVx2_ASAP7_75t_L g465 ( .A(n_222), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_224), .A2(n_227), .B1(n_1123), .B2(n_1124), .Y(n_1122) );
INVxp67_ASAP7_75t_SL g525 ( .A(n_225), .Y(n_525) );
INVxp67_ASAP7_75t_SL g990 ( .A(n_226), .Y(n_990) );
INVx1_ASAP7_75t_L g1136 ( .A(n_227), .Y(n_1136) );
INVx1_ASAP7_75t_L g615 ( .A(n_228), .Y(n_615) );
INVx1_ASAP7_75t_L g681 ( .A(n_230), .Y(n_681) );
XOR2x1_ASAP7_75t_L g1162 ( .A(n_231), .B(n_1163), .Y(n_1162) );
AOI221xp5_ASAP7_75t_L g1294 ( .A1(n_231), .A2(n_234), .B1(n_1295), .B2(n_1296), .C(n_1297), .Y(n_1294) );
OAI22xp33_ASAP7_75t_L g1154 ( .A1(n_232), .A2(n_262), .B1(n_345), .B2(n_1155), .Y(n_1154) );
INVx1_ASAP7_75t_L g1208 ( .A(n_233), .Y(n_1208) );
INVxp67_ASAP7_75t_L g733 ( .A(n_235), .Y(n_733) );
INVx1_ASAP7_75t_L g1485 ( .A(n_236), .Y(n_1485) );
INVxp67_ASAP7_75t_SL g848 ( .A(n_238), .Y(n_848) );
INVx1_ASAP7_75t_L g534 ( .A(n_239), .Y(n_534) );
INVx1_ASAP7_75t_L g858 ( .A(n_240), .Y(n_858) );
INVxp33_ASAP7_75t_L g727 ( .A(n_241), .Y(n_727) );
INVxp33_ASAP7_75t_L g1093 ( .A(n_242), .Y(n_1093) );
CKINVDCx5p33_ASAP7_75t_R g1540 ( .A(n_244), .Y(n_1540) );
AOI221xp5_ASAP7_75t_L g1010 ( .A1(n_245), .A2(n_280), .B1(n_590), .B2(n_700), .C(n_791), .Y(n_1010) );
INVxp33_ASAP7_75t_L g1032 ( .A(n_245), .Y(n_1032) );
INVx1_ASAP7_75t_L g1228 ( .A(n_246), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_246), .B(n_1226), .Y(n_1233) );
INVxp67_ASAP7_75t_SL g985 ( .A(n_247), .Y(n_985) );
INVx1_ASAP7_75t_L g812 ( .A(n_248), .Y(n_812) );
INVx1_ASAP7_75t_L g1533 ( .A(n_249), .Y(n_1533) );
INVxp67_ASAP7_75t_SL g1127 ( .A(n_250), .Y(n_1127) );
INVx1_ASAP7_75t_L g914 ( .A(n_252), .Y(n_914) );
INVx1_ASAP7_75t_L g1463 ( .A(n_254), .Y(n_1463) );
OAI22xp5_ASAP7_75t_L g1486 ( .A1(n_254), .A2(n_266), .B1(n_337), .B2(n_1487), .Y(n_1486) );
INVx1_ASAP7_75t_L g739 ( .A(n_256), .Y(n_739) );
CKINVDCx5p33_ASAP7_75t_R g776 ( .A(n_257), .Y(n_776) );
AOI22x1_ASAP7_75t_L g894 ( .A1(n_258), .A2(n_895), .B1(n_942), .B2(n_943), .Y(n_894) );
INVxp67_ASAP7_75t_L g942 ( .A(n_258), .Y(n_942) );
INVx1_ASAP7_75t_L g975 ( .A(n_260), .Y(n_975) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_261), .A2(n_359), .B(n_362), .Y(n_358) );
INVx1_ASAP7_75t_L g476 ( .A(n_261), .Y(n_476) );
INVxp67_ASAP7_75t_SL g1126 ( .A(n_262), .Y(n_1126) );
INVx2_ASAP7_75t_L g300 ( .A(n_263), .Y(n_300) );
XNOR2x1_ASAP7_75t_L g582 ( .A(n_264), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g1462 ( .A(n_266), .Y(n_1462) );
INVxp33_ASAP7_75t_SL g1108 ( .A(n_267), .Y(n_1108) );
INVxp67_ASAP7_75t_L g1079 ( .A(n_268), .Y(n_1079) );
INVx1_ASAP7_75t_L g1110 ( .A(n_270), .Y(n_1110) );
CKINVDCx5p33_ASAP7_75t_R g1466 ( .A(n_271), .Y(n_1466) );
INVxp33_ASAP7_75t_SL g1040 ( .A(n_272), .Y(n_1040) );
INVx1_ASAP7_75t_L g541 ( .A(n_273), .Y(n_541) );
INVx1_ASAP7_75t_L g325 ( .A(n_274), .Y(n_325) );
BUFx3_ASAP7_75t_L g342 ( .A(n_274), .Y(n_342) );
BUFx3_ASAP7_75t_L g324 ( .A(n_275), .Y(n_324) );
INVx1_ASAP7_75t_L g348 ( .A(n_275), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_276), .Y(n_357) );
INVx1_ASAP7_75t_L g417 ( .A(n_277), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g672 ( .A(n_279), .Y(n_672) );
INVxp33_ASAP7_75t_L g1030 ( .A(n_280), .Y(n_1030) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_304), .B(n_1212), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx3_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_291), .Y(n_285) );
AND2x4_ASAP7_75t_L g1508 ( .A(n_286), .B(n_292), .Y(n_1508) );
NOR2xp33_ASAP7_75t_SL g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_SL g1513 ( .A(n_287), .Y(n_1513) );
NAND2xp5_ASAP7_75t_L g1565 ( .A(n_287), .B(n_289), .Y(n_1565) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_289), .B(n_1513), .Y(n_1512) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_293), .B(n_297), .Y(n_292) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g431 ( .A(n_295), .B(n_303), .Y(n_431) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g508 ( .A(n_296), .B(n_509), .Y(n_508) );
OR2x6_ASAP7_75t_L g297 ( .A(n_298), .B(n_302), .Y(n_297) );
OR2x2_ASAP7_75t_L g404 ( .A(n_298), .B(n_405), .Y(n_404) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_298), .Y(n_513) );
BUFx2_ASAP7_75t_L g636 ( .A(n_298), .Y(n_636) );
OAI22xp33_ASAP7_75t_L g643 ( .A1(n_298), .A2(n_539), .B1(n_601), .B2(n_644), .Y(n_643) );
INVx2_ASAP7_75t_SL g746 ( .A(n_298), .Y(n_746) );
INVx2_ASAP7_75t_SL g843 ( .A(n_298), .Y(n_843) );
INVx1_ASAP7_75t_L g938 ( .A(n_298), .Y(n_938) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g421 ( .A(n_300), .Y(n_421) );
INVx1_ASAP7_75t_L g426 ( .A(n_300), .Y(n_426) );
AND2x2_ASAP7_75t_L g435 ( .A(n_300), .B(n_301), .Y(n_435) );
INVx2_ASAP7_75t_L g442 ( .A(n_300), .Y(n_442) );
AND2x4_ASAP7_75t_L g448 ( .A(n_300), .B(n_427), .Y(n_448) );
INVx1_ASAP7_75t_L g415 ( .A(n_301), .Y(n_415) );
INVx2_ASAP7_75t_L g427 ( .A(n_301), .Y(n_427) );
INVx1_ASAP7_75t_L g444 ( .A(n_301), .Y(n_444) );
INVx1_ASAP7_75t_L g518 ( .A(n_301), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_301), .B(n_442), .Y(n_524) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
XNOR2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_1002), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_824), .B1(n_1000), .B2(n_1001), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g1000 ( .A(n_307), .Y(n_1000) );
XNOR2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_580), .Y(n_307) );
XOR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_483), .Y(n_308) );
XNOR2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_482), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_411), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_315), .B1(n_401), .B2(n_402), .Y(n_311) );
INVx2_ASAP7_75t_L g612 ( .A(n_312), .Y(n_612) );
OAI31xp33_ASAP7_75t_L g677 ( .A1(n_312), .A2(n_678), .A3(n_679), .B(n_697), .Y(n_677) );
BUFx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g547 ( .A(n_313), .Y(n_547) );
BUFx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g430 ( .A(n_314), .Y(n_430) );
OR2x6_ASAP7_75t_L g507 ( .A(n_314), .B(n_508), .Y(n_507) );
NAND3xp33_ASAP7_75t_SL g315 ( .A(n_316), .B(n_365), .C(n_393), .Y(n_315) );
AOI211xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B(n_326), .C(n_343), .Y(n_316) );
AOI221xp5_ASAP7_75t_L g565 ( .A1(n_318), .A2(n_534), .B1(n_566), .B2(n_570), .C(n_573), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_318), .A2(n_395), .B1(n_739), .B2(n_747), .Y(n_764) );
AOI221xp5_ASAP7_75t_L g777 ( .A1(n_318), .A2(n_778), .B1(n_779), .B2(n_783), .C(n_785), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_318), .A2(n_395), .B1(n_855), .B2(n_857), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_318), .A2(n_395), .B1(n_974), .B2(n_975), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_318), .A2(n_395), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
AOI22xp33_ASAP7_75t_SL g1073 ( .A1(n_318), .A2(n_395), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_318), .A2(n_395), .B1(n_1208), .B2(n_1209), .Y(n_1207) );
AOI22xp33_ASAP7_75t_L g1502 ( .A1(n_318), .A2(n_395), .B1(n_1503), .B2(n_1504), .Y(n_1502) );
AOI22xp33_ASAP7_75t_L g1560 ( .A1(n_318), .A2(n_395), .B1(n_1539), .B2(n_1542), .Y(n_1560) );
INVx4_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
INVx2_ASAP7_75t_L g371 ( .A(n_320), .Y(n_371) );
OR2x2_ASAP7_75t_L g396 ( .A(n_320), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g330 ( .A(n_321), .Y(n_330) );
INVx1_ASAP7_75t_L g572 ( .A(n_322), .Y(n_572) );
INVx2_ASAP7_75t_L g686 ( .A(n_322), .Y(n_686) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g350 ( .A(n_323), .Y(n_350) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_323), .Y(n_389) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_323), .Y(n_564) );
AND2x4_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx2_ASAP7_75t_L g336 ( .A(n_324), .Y(n_336) );
AND2x2_ASAP7_75t_L g370 ( .A(n_324), .B(n_342), .Y(n_370) );
INVx1_ASAP7_75t_L g355 ( .A(n_325), .Y(n_355) );
INVx2_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g877 ( .A(n_328), .Y(n_877) );
AOI222xp33_ASAP7_75t_L g910 ( .A1(n_328), .A2(n_338), .B1(n_911), .B2(n_912), .C1(n_913), .C2(n_914), .Y(n_910) );
INVx2_ASAP7_75t_SL g962 ( .A(n_328), .Y(n_962) );
INVx1_ASAP7_75t_L g1058 ( .A(n_328), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_328), .A2(n_879), .B1(n_1147), .B2(n_1148), .Y(n_1146) );
INVx2_ASAP7_75t_L g1487 ( .A(n_328), .Y(n_1487) );
AND2x4_ASAP7_75t_L g328 ( .A(n_329), .B(n_333), .Y(n_328) );
AND2x2_ASAP7_75t_L g338 ( .A(n_329), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g392 ( .A(n_329), .Y(n_392) );
AND2x2_ASAP7_75t_L g410 ( .A(n_329), .B(n_361), .Y(n_410) );
AND2x4_ASAP7_75t_L g575 ( .A(n_329), .B(n_333), .Y(n_575) );
AND2x4_ASAP7_75t_L g577 ( .A(n_329), .B(n_339), .Y(n_577) );
BUFx2_ASAP7_75t_L g599 ( .A(n_329), .Y(n_599) );
AND2x2_ASAP7_75t_L g879 ( .A(n_329), .B(n_339), .Y(n_879) );
AND2x4_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
AND2x4_ASAP7_75t_L g363 ( .A(n_331), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g382 ( .A(n_332), .B(n_364), .Y(n_382) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x4_ASAP7_75t_L g361 ( .A(n_336), .B(n_341), .Y(n_361) );
INVx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
BUFx3_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g347 ( .A(n_342), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g592 ( .A(n_346), .Y(n_592) );
INVx1_ASAP7_75t_L g702 ( .A(n_346), .Y(n_702) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_347), .Y(n_376) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_347), .Y(n_400) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_347), .Y(n_553) );
BUFx2_ASAP7_75t_L g571 ( .A(n_347), .Y(n_571) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_347), .Y(n_594) );
BUFx2_ASAP7_75t_L g606 ( .A(n_347), .Y(n_606) );
BUFx3_ASAP7_75t_L g688 ( .A(n_347), .Y(n_688) );
INVx2_ASAP7_75t_SL g789 ( .A(n_347), .Y(n_789) );
INVx1_ASAP7_75t_L g356 ( .A(n_348), .Y(n_356) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g972 ( .A(n_350), .Y(n_972) );
INVx1_ASAP7_75t_L g1020 ( .A(n_350), .Y(n_1020) );
OAI21xp5_ASAP7_75t_SL g351 ( .A1(n_352), .A2(n_357), .B(n_358), .Y(n_351) );
OAI221xp5_ASAP7_75t_L g1135 ( .A1(n_352), .A2(n_375), .B1(n_1118), .B2(n_1136), .C(n_1137), .Y(n_1135) );
INVx2_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g1553 ( .A(n_353), .Y(n_1553) );
BUFx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g604 ( .A(n_354), .Y(n_604) );
BUFx4f_ASAP7_75t_L g683 ( .A(n_354), .Y(n_683) );
INVx2_ASAP7_75t_L g691 ( .A(n_354), .Y(n_691) );
INVx1_ASAP7_75t_L g1063 ( .A(n_354), .Y(n_1063) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
OR2x2_ASAP7_75t_L g397 ( .A(n_355), .B(n_356), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_357), .A2(n_468), .B1(n_469), .B2(n_473), .Y(n_467) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g386 ( .A(n_360), .Y(n_386) );
INVx2_ASAP7_75t_SL g562 ( .A(n_360), .Y(n_562) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_360), .Y(n_597) );
INVx1_ASAP7_75t_L g694 ( .A(n_360), .Y(n_694) );
BUFx6f_ASAP7_75t_L g792 ( .A(n_360), .Y(n_792) );
INVx6_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx2_ASAP7_75t_L g567 ( .A(n_361), .Y(n_567) );
INVx2_ASAP7_75t_L g781 ( .A(n_361), .Y(n_781) );
INVx1_ASAP7_75t_L g960 ( .A(n_362), .Y(n_960) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g569 ( .A(n_363), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_363), .Y(n_590) );
INVx2_ASAP7_75t_SL g695 ( .A(n_363), .Y(n_695) );
HB1xp67_ASAP7_75t_L g1142 ( .A(n_363), .Y(n_1142) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_372), .B1(n_373), .B2(n_383), .C(n_390), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g554 ( .A1(n_366), .A2(n_390), .B1(n_541), .B2(n_555), .C(n_559), .Y(n_554) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g793 ( .A(n_367), .Y(n_793) );
INVx2_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g758 ( .A1(n_368), .A2(n_598), .B1(n_748), .B2(n_759), .C(n_762), .Y(n_758) );
INVx1_ASAP7_75t_L g888 ( .A(n_368), .Y(n_888) );
INVx1_ASAP7_75t_L g965 ( .A(n_368), .Y(n_965) );
AOI221xp5_ASAP7_75t_L g1015 ( .A1(n_368), .A2(n_390), .B1(n_1016), .B2(n_1018), .C(n_1021), .Y(n_1015) );
INVx1_ASAP7_75t_L g1198 ( .A(n_368), .Y(n_1198) );
BUFx6f_ASAP7_75t_L g1493 ( .A(n_368), .Y(n_1493) );
AND2x4_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
BUFx3_ASAP7_75t_L g556 ( .A(n_369), .Y(n_556) );
INVx2_ASAP7_75t_SL g588 ( .A(n_369), .Y(n_588) );
AND2x4_ASAP7_75t_L g598 ( .A(n_369), .B(n_599), .Y(n_598) );
BUFx4f_ASAP7_75t_L g700 ( .A(n_369), .Y(n_700) );
BUFx6f_ASAP7_75t_L g1499 ( .A(n_369), .Y(n_1499) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_370), .Y(n_380) );
AND2x4_ASAP7_75t_L g399 ( .A(n_371), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g552 ( .A(n_371), .B(n_553), .Y(n_552) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_371), .A2(n_395), .B1(n_601), .B2(n_602), .C(n_609), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g698 ( .A1(n_371), .A2(n_699), .B(n_700), .C(n_701), .Y(n_698) );
OAI21xp5_ASAP7_75t_L g1149 ( .A1(n_371), .A2(n_1150), .B(n_1154), .Y(n_1149) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g1061 ( .A(n_376), .Y(n_1061) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g1017 ( .A(n_378), .Y(n_1017) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_L g390 ( .A(n_379), .B(n_391), .Y(n_390) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_379), .Y(n_568) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx6f_ASAP7_75t_L g760 ( .A(n_380), .Y(n_760) );
INVx2_ASAP7_75t_L g869 ( .A(n_380), .Y(n_869) );
BUFx2_ASAP7_75t_L g970 ( .A(n_381), .Y(n_970) );
INVx1_ASAP7_75t_L g1137 ( .A(n_381), .Y(n_1137) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
BUFx3_ASAP7_75t_L g558 ( .A(n_382), .Y(n_558) );
INVx1_ASAP7_75t_L g761 ( .A(n_382), .Y(n_761) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_386), .Y(n_589) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g886 ( .A(n_388), .Y(n_886) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx6f_ASAP7_75t_L g608 ( .A(n_389), .Y(n_608) );
BUFx6f_ASAP7_75t_L g763 ( .A(n_389), .Y(n_763) );
INVx1_ASAP7_75t_L g1559 ( .A(n_389), .Y(n_1559) );
HB1xp67_ASAP7_75t_L g889 ( .A(n_390), .Y(n_889) );
INVx1_ASAP7_75t_L g915 ( .A(n_390), .Y(n_915) );
AOI221xp5_ASAP7_75t_L g963 ( .A1(n_390), .A2(n_964), .B1(n_966), .B2(n_967), .C(n_971), .Y(n_963) );
AOI221xp5_ASAP7_75t_L g1069 ( .A1(n_390), .A2(n_964), .B1(n_1070), .B2(n_1071), .C(n_1072), .Y(n_1069) );
AOI221xp5_ASAP7_75t_L g1196 ( .A1(n_390), .A2(n_1197), .B1(n_1199), .B2(n_1200), .C(n_1204), .Y(n_1196) );
AOI221xp5_ASAP7_75t_L g1492 ( .A1(n_390), .A2(n_1493), .B1(n_1494), .B2(n_1495), .C(n_1500), .Y(n_1492) );
AOI221xp5_ASAP7_75t_L g1554 ( .A1(n_390), .A2(n_1197), .B1(n_1543), .B2(n_1555), .C(n_1556), .Y(n_1554) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B1(n_398), .B2(n_399), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_395), .A2(n_533), .B1(n_536), .B2(n_550), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_395), .A2(n_552), .B1(n_775), .B2(n_776), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_395), .A2(n_399), .B1(n_907), .B2(n_908), .Y(n_906) );
INVx6_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx2_ASAP7_75t_L g958 ( .A(n_397), .Y(n_958) );
INVx1_ASAP7_75t_L g1066 ( .A(n_397), .Y(n_1066) );
INVx2_ASAP7_75t_L g1152 ( .A(n_397), .Y(n_1152) );
INVx1_ASAP7_75t_L g875 ( .A(n_399), .Y(n_875) );
HB1xp67_ASAP7_75t_L g952 ( .A(n_399), .Y(n_952) );
AOI221xp5_ASAP7_75t_L g1009 ( .A1(n_399), .A2(n_1010), .B1(n_1011), .B2(n_1013), .C(n_1014), .Y(n_1009) );
AOI211xp5_ASAP7_75t_L g1055 ( .A1(n_399), .A2(n_1056), .B(n_1057), .C(n_1059), .Y(n_1055) );
AOI211xp5_ASAP7_75t_L g1190 ( .A1(n_399), .A2(n_1191), .B(n_1192), .C(n_1193), .Y(n_1190) );
AOI211xp5_ASAP7_75t_SL g1484 ( .A1(n_399), .A2(n_1485), .B(n_1486), .C(n_1488), .Y(n_1484) );
AOI211xp5_ASAP7_75t_L g1547 ( .A1(n_399), .A2(n_1540), .B(n_1548), .C(n_1549), .Y(n_1547) );
BUFx3_ASAP7_75t_L g1012 ( .A(n_400), .Y(n_1012) );
INVx1_ASAP7_75t_L g1551 ( .A(n_400), .Y(n_1551) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_402), .A2(n_772), .B1(n_1008), .B2(n_1025), .Y(n_1007) );
AOI21xp33_ASAP7_75t_L g1052 ( .A1(n_402), .A2(n_1053), .B(n_1054), .Y(n_1052) );
AOI21xp5_ASAP7_75t_L g1481 ( .A1(n_402), .A2(n_1482), .B(n_1483), .Y(n_1481) );
INVx5_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g579 ( .A(n_403), .Y(n_579) );
INVx2_ASAP7_75t_SL g767 ( .A(n_403), .Y(n_767) );
INVx2_ASAP7_75t_L g796 ( .A(n_403), .Y(n_796) );
INVx1_ASAP7_75t_L g1187 ( .A(n_403), .Y(n_1187) );
AND2x4_ASAP7_75t_L g403 ( .A(n_404), .B(n_407), .Y(n_403) );
INVx2_ASAP7_75t_L g624 ( .A(n_404), .Y(n_624) );
INVx3_ASAP7_75t_L g416 ( .A(n_405), .Y(n_416) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx2_ASAP7_75t_L g610 ( .A(n_410), .Y(n_610) );
AND4x1_ASAP7_75t_L g411 ( .A(n_412), .B(n_428), .C(n_467), .D(n_475), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_417), .B1(n_418), .B2(n_422), .C(n_423), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_413), .A2(n_418), .B1(n_423), .B2(n_615), .C(n_616), .Y(n_614) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_413), .A2(n_418), .B1(n_423), .B2(n_649), .C(n_650), .Y(n_648) );
INVx1_ASAP7_75t_L g1160 ( .A(n_413), .Y(n_1160) );
AOI221xp5_ASAP7_75t_L g1165 ( .A1(n_413), .A2(n_1157), .B1(n_1166), .B2(n_1167), .C(n_1168), .Y(n_1165) );
AND2x4_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g499 ( .A(n_415), .Y(n_499) );
AND2x4_ASAP7_75t_L g418 ( .A(n_416), .B(n_419), .Y(n_418) );
AND2x4_ASAP7_75t_L g423 ( .A(n_416), .B(n_424), .Y(n_423) );
NAND2x1_ASAP7_75t_SL g497 ( .A(n_416), .B(n_498), .Y(n_497) );
NAND2x1p5_ASAP7_75t_L g500 ( .A(n_416), .B(n_501), .Y(n_500) );
NAND2x1p5_ASAP7_75t_L g504 ( .A(n_416), .B(n_474), .Y(n_504) );
AOI32xp33_ASAP7_75t_L g919 ( .A1(n_416), .A2(n_920), .A3(n_922), .B1(n_924), .B2(n_925), .Y(n_919) );
INVx1_ASAP7_75t_L g1158 ( .A(n_418), .Y(n_1158) );
HB1xp67_ASAP7_75t_L g1461 ( .A(n_418), .Y(n_1461) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g517 ( .A(n_421), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_421), .B(n_518), .Y(n_540) );
AOI221xp5_ASAP7_75t_L g1156 ( .A1(n_423), .A2(n_1147), .B1(n_1148), .B2(n_1157), .C(n_1159), .Y(n_1156) );
HB1xp67_ASAP7_75t_L g1168 ( .A(n_423), .Y(n_1168) );
AOI221xp5_ASAP7_75t_L g1460 ( .A1(n_423), .A2(n_1159), .B1(n_1461), .B2(n_1462), .C(n_1463), .Y(n_1460) );
BUFx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_425), .Y(n_438) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_425), .Y(n_458) );
BUFx3_ASAP7_75t_L g474 ( .A(n_425), .Y(n_474) );
INVx1_ASAP7_75t_L g656 ( .A(n_425), .Y(n_656) );
BUFx3_ASAP7_75t_L g1130 ( .A(n_425), .Y(n_1130) );
AND2x4_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
AOI33xp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_432), .A3(n_439), .B1(n_449), .B2(n_453), .B3(n_459), .Y(n_428) );
AOI222xp33_ASAP7_75t_L g625 ( .A1(n_429), .A2(n_459), .B1(n_626), .B2(n_628), .C1(n_629), .C2(n_638), .Y(n_625) );
AOI33xp33_ASAP7_75t_L g651 ( .A1(n_429), .A2(n_652), .A3(n_657), .B1(n_661), .B2(n_663), .B3(n_664), .Y(n_651) );
AND2x4_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
AND2x2_ASAP7_75t_L g664 ( .A(n_430), .B(n_665), .Y(n_664) );
BUFx2_ASAP7_75t_L g766 ( .A(n_430), .Y(n_766) );
AND2x4_ASAP7_75t_L g924 ( .A(n_430), .B(n_431), .Y(n_924) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx3_ASAP7_75t_L g654 ( .A(n_434), .Y(n_654) );
BUFx2_ASAP7_75t_L g1179 ( .A(n_434), .Y(n_1179) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx3_ASAP7_75t_L g456 ( .A(n_435), .Y(n_456) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g1124 ( .A(n_437), .Y(n_1124) );
INVx2_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
BUFx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_441), .Y(n_481) );
INVx1_ASAP7_75t_L g631 ( .A(n_441), .Y(n_631) );
INVx1_ASAP7_75t_L g640 ( .A(n_441), .Y(n_640) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_441), .Y(n_658) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_441), .Y(n_662) );
AND2x4_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
INVx1_ASAP7_75t_L g502 ( .A(n_442), .Y(n_502) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_445), .Y(n_850) );
BUFx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x4_ASAP7_75t_L g470 ( .A(n_446), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g1088 ( .A(n_446), .Y(n_1088) );
INVx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx3_ASAP7_75t_L g452 ( .A(n_447), .Y(n_452) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_447), .Y(n_660) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_448), .Y(n_527) );
INVx1_ASAP7_75t_L g743 ( .A(n_448), .Y(n_743) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_451), .A2(n_776), .B1(n_778), .B2(n_818), .Y(n_822) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g633 ( .A(n_452), .Y(n_633) );
INVx2_ASAP7_75t_L g642 ( .A(n_452), .Y(n_642) );
AND2x2_ASAP7_75t_L g674 ( .A(n_452), .B(n_471), .Y(n_674) );
INVx1_ASAP7_75t_L g1536 ( .A(n_452), .Y(n_1536) );
BUFx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_SL g478 ( .A(n_456), .Y(n_478) );
INVx2_ASAP7_75t_SL g627 ( .A(n_456), .Y(n_627) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g714 ( .A(n_458), .B(n_471), .Y(n_714) );
INVx2_ASAP7_75t_SL g1474 ( .A(n_458), .Y(n_1474) );
INVx1_ASAP7_75t_L g749 ( .A(n_459), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g932 ( .A1(n_459), .A2(n_469), .B1(n_933), .B2(n_941), .Y(n_932) );
AOI33xp33_ASAP7_75t_L g1176 ( .A1(n_459), .A2(n_1177), .A3(n_1178), .B1(n_1180), .B2(n_1184), .B3(n_1185), .Y(n_1176) );
AOI33xp33_ASAP7_75t_L g1470 ( .A1(n_459), .A2(n_1177), .A3(n_1471), .B1(n_1475), .B2(n_1477), .B3(n_1478), .Y(n_1470) );
INVx6_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx5_ASAP7_75t_L g543 ( .A(n_460), .Y(n_543) );
OR2x6_ASAP7_75t_L g460 ( .A(n_461), .B(n_463), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x4_ASAP7_75t_L g471 ( .A(n_462), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g665 ( .A(n_463), .Y(n_665) );
NAND2x1p5_ASAP7_75t_L g463 ( .A(n_464), .B(n_466), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g509 ( .A(n_465), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_469), .A2(n_473), .B1(n_489), .B2(n_490), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_469), .A2(n_473), .B1(n_1029), .B2(n_1030), .Y(n_1028) );
BUFx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g622 ( .A(n_470), .Y(n_622) );
BUFx2_ASAP7_75t_L g801 ( .A(n_470), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_470), .A2(n_835), .B1(n_836), .B2(n_837), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_470), .A2(n_837), .B1(n_957), .B2(n_981), .Y(n_980) );
BUFx2_ASAP7_75t_L g1105 ( .A(n_470), .Y(n_1105) );
BUFx2_ASAP7_75t_L g1171 ( .A(n_470), .Y(n_1171) );
AND2x6_ASAP7_75t_L g473 ( .A(n_471), .B(n_474), .Y(n_473) );
AND2x4_ASAP7_75t_L g477 ( .A(n_471), .B(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g480 ( .A(n_471), .B(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g626 ( .A(n_471), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g670 ( .A(n_471), .B(n_481), .Y(n_670) );
AND2x2_ASAP7_75t_L g806 ( .A(n_471), .B(n_481), .Y(n_806) );
AND2x2_ASAP7_75t_L g931 ( .A(n_471), .B(n_481), .Y(n_931) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_471), .B(n_481), .Y(n_1109) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_473), .A2(n_480), .B1(n_618), .B2(n_619), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_473), .A2(n_670), .B1(n_671), .B2(n_672), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_473), .A2(n_800), .B1(n_801), .B2(n_802), .Y(n_799) );
BUFx2_ASAP7_75t_L g837 ( .A(n_473), .Y(n_837) );
INVx1_ASAP7_75t_SL g918 ( .A(n_473), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_473), .A2(n_801), .B1(n_1064), .B2(n_1093), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_473), .A2(n_1104), .B1(n_1105), .B2(n_1106), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_473), .A2(n_1170), .B1(n_1171), .B2(n_1172), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g1464 ( .A1(n_473), .A2(n_1105), .B1(n_1465), .B2(n_1466), .Y(n_1464) );
AOI22xp33_ASAP7_75t_L g1519 ( .A1(n_473), .A2(n_622), .B1(n_1520), .B2(n_1521), .Y(n_1519) );
BUFx2_ASAP7_75t_L g923 ( .A(n_474), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B1(n_479), .B2(n_480), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_477), .A2(n_480), .B1(n_492), .B2(n_493), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_477), .B(n_667), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_477), .A2(n_804), .B1(n_805), .B2(n_806), .Y(n_803) );
BUFx2_ASAP7_75t_L g832 ( .A(n_477), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_477), .A2(n_929), .B1(n_930), .B2(n_931), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_477), .A2(n_931), .B1(n_1032), .B2(n_1033), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_477), .A2(n_480), .B1(n_1067), .B2(n_1095), .Y(n_1094) );
AOI21xp5_ASAP7_75t_L g1111 ( .A1(n_477), .A2(n_1112), .B(n_1113), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1173 ( .A1(n_477), .A2(n_931), .B1(n_1174), .B2(n_1175), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1467 ( .A1(n_477), .A2(n_931), .B1(n_1468), .B2(n_1469), .Y(n_1467) );
AOI22xp33_ASAP7_75t_L g1522 ( .A1(n_477), .A2(n_1109), .B1(n_1523), .B2(n_1524), .Y(n_1522) );
BUFx3_ASAP7_75t_L g1479 ( .A(n_478), .Y(n_1479) );
INVx2_ASAP7_75t_SL g935 ( .A(n_481), .Y(n_935) );
XNOR2x1_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_544), .Y(n_485) );
NOR3xp33_ASAP7_75t_L g486 ( .A(n_487), .B(n_494), .C(n_505), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_491), .Y(n_487) );
INVx2_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g719 ( .A(n_496), .Y(n_719) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_497), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_498), .A2(n_501), .B1(n_913), .B2(n_914), .Y(n_926) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx4f_ASAP7_75t_L g720 ( .A(n_500), .Y(n_720) );
BUFx4f_ASAP7_75t_L g1035 ( .A(n_500), .Y(n_1035) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx3_ASAP7_75t_L g721 ( .A(n_504), .Y(n_721) );
BUFx2_ASAP7_75t_L g1526 ( .A(n_504), .Y(n_1526) );
OAI33xp33_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_510), .A3(n_520), .B1(n_529), .B2(n_535), .B3(n_542), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OAI33xp33_ASAP7_75t_L g722 ( .A1(n_507), .A2(n_723), .A3(n_729), .B1(n_735), .B2(n_744), .B3(n_749), .Y(n_722) );
OAI33xp33_ASAP7_75t_L g809 ( .A1(n_507), .A2(n_542), .A3(n_810), .B1(n_816), .B2(n_822), .B3(n_823), .Y(n_809) );
OAI33xp33_ASAP7_75t_L g840 ( .A1(n_507), .A2(n_841), .A3(n_847), .B1(n_851), .B2(n_856), .B3(n_859), .Y(n_840) );
OAI33xp33_ASAP7_75t_L g983 ( .A1(n_507), .A2(n_749), .A3(n_984), .B1(n_987), .B2(n_993), .B3(n_996), .Y(n_983) );
OAI33xp33_ASAP7_75t_L g1036 ( .A1(n_507), .A2(n_542), .A3(n_1037), .B1(n_1041), .B2(n_1045), .B3(n_1046), .Y(n_1036) );
OAI33xp33_ASAP7_75t_L g1077 ( .A1(n_507), .A2(n_542), .A3(n_1078), .B1(n_1082), .B2(n_1087), .B3(n_1089), .Y(n_1077) );
OAI22xp5_ASAP7_75t_L g1113 ( .A1(n_507), .A2(n_542), .B1(n_1114), .B2(n_1125), .Y(n_1113) );
OAI33xp33_ASAP7_75t_L g1527 ( .A1(n_507), .A2(n_542), .A3(n_1528), .B1(n_1532), .B2(n_1538), .B3(n_1541), .Y(n_1527) );
OAI22xp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_514), .B1(n_515), .B2(n_519), .Y(n_510) );
OAI22xp33_ASAP7_75t_L g535 ( .A1(n_511), .A2(n_536), .B1(n_537), .B2(n_541), .Y(n_535) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx2_ASAP7_75t_L g1039 ( .A(n_513), .Y(n_1039) );
OAI22xp33_ASAP7_75t_L g1538 ( .A1(n_513), .A2(n_530), .B1(n_1539), .B2(n_1540), .Y(n_1538) );
OAI22xp33_ASAP7_75t_L g1089 ( .A1(n_515), .A2(n_842), .B1(n_1070), .B2(n_1074), .Y(n_1089) );
BUFx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g1086 ( .A(n_516), .Y(n_1086) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g728 ( .A(n_517), .Y(n_728) );
BUFx2_ASAP7_75t_L g814 ( .A(n_517), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_525), .B1(n_526), .B2(n_528), .Y(n_520) );
BUFx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g732 ( .A(n_523), .Y(n_732) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_523), .Y(n_989) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g532 ( .A(n_524), .Y(n_532) );
BUFx2_ASAP7_75t_L g1117 ( .A(n_524), .Y(n_1117) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_526), .A2(n_530), .B1(n_533), .B2(n_534), .Y(n_529) );
INVx2_ASAP7_75t_L g921 ( .A(n_526), .Y(n_921) );
INVx2_ASAP7_75t_SL g1472 ( .A(n_526), .Y(n_1472) );
INVx4_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g854 ( .A(n_527), .Y(n_854) );
INVx2_ASAP7_75t_SL g991 ( .A(n_527), .Y(n_991) );
INVx2_ASAP7_75t_SL g1183 ( .A(n_527), .Y(n_1183) );
OAI22xp5_ASAP7_75t_L g847 ( .A1(n_530), .A2(n_848), .B1(n_849), .B2(n_850), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_530), .A2(n_852), .B1(n_853), .B2(n_855), .Y(n_851) );
BUFx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g819 ( .A(n_531), .Y(n_819) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx3_ASAP7_75t_L g738 ( .A(n_532), .Y(n_738) );
OAI22xp5_ASAP7_75t_SL g744 ( .A1(n_537), .A2(n_745), .B1(n_747), .B2(n_748), .Y(n_744) );
OAI22xp33_ASAP7_75t_L g823 ( .A1(n_537), .A2(n_775), .B1(n_794), .B2(n_811), .Y(n_823) );
OAI22xp33_ASAP7_75t_L g984 ( .A1(n_537), .A2(n_745), .B1(n_985), .B2(n_986), .Y(n_984) );
OAI22xp33_ASAP7_75t_L g996 ( .A1(n_537), .A2(n_966), .B1(n_975), .B2(n_991), .Y(n_996) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g940 ( .A(n_538), .Y(n_940) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_539), .A2(n_635), .B1(n_636), .B2(n_637), .Y(n_634) );
BUFx3_ASAP7_75t_L g845 ( .A(n_539), .Y(n_845) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g860 ( .A(n_542), .Y(n_860) );
CKINVDCx8_ASAP7_75t_R g542 ( .A(n_543), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_548), .B1(n_578), .B2(n_579), .Y(n_544) );
INVx1_ASAP7_75t_SL g891 ( .A(n_545), .Y(n_891) );
OAI21xp33_ASAP7_75t_L g896 ( .A1(n_545), .A2(n_897), .B(n_909), .Y(n_896) );
INVx5_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AOI31xp33_ASAP7_75t_L g1054 ( .A1(n_546), .A2(n_1055), .A3(n_1069), .B(n_1073), .Y(n_1054) );
BUFx8_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g772 ( .A(n_547), .Y(n_772) );
AOI31xp33_ASAP7_75t_L g949 ( .A1(n_547), .A2(n_950), .A3(n_963), .B(n_973), .Y(n_949) );
NAND3xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_554), .C(n_565), .Y(n_548) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g752 ( .A1(n_552), .A2(n_736), .B1(n_753), .B2(n_754), .C(n_755), .Y(n_752) );
BUFx2_ASAP7_75t_L g873 ( .A(n_553), .Y(n_873) );
INVx1_ASAP7_75t_L g1490 ( .A(n_553), .Y(n_1490) );
INVx1_ASAP7_75t_L g1497 ( .A(n_553), .Y(n_1497) );
INVx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g883 ( .A(n_558), .Y(n_883) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx3_ASAP7_75t_L g784 ( .A(n_564), .Y(n_784) );
INVx1_ASAP7_75t_L g901 ( .A(n_564), .Y(n_901) );
A2O1A1Ixp33_ASAP7_75t_L g1144 ( .A1(n_567), .A2(n_568), .B(n_1110), .C(n_1145), .Y(n_1144) );
HB1xp67_ASAP7_75t_L g882 ( .A(n_568), .Y(n_882) );
INVx1_ASAP7_75t_L g1153 ( .A(n_572), .Y(n_1153) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_SL g611 ( .A(n_575), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_575), .A2(n_577), .B1(n_649), .B2(n_650), .Y(n_704) );
INVx4_ASAP7_75t_L g756 ( .A(n_575), .Y(n_756) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_SL g757 ( .A(n_577), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g861 ( .A1(n_579), .A2(n_862), .B(n_863), .Y(n_861) );
XOR2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_705), .Y(n_580) );
XNOR2x1_ASAP7_75t_L g581 ( .A(n_582), .B(n_645), .Y(n_581) );
NOR2x1_ASAP7_75t_L g583 ( .A(n_584), .B(n_613), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_600), .B(n_612), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_591), .B1(n_593), .B2(n_595), .C(n_598), .Y(n_585) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g782 ( .A(n_588), .Y(n_782) );
INVx1_ASAP7_75t_L g905 ( .A(n_588), .Y(n_905) );
HB1xp67_ASAP7_75t_L g885 ( .A(n_589), .Y(n_885) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g696 ( .A(n_598), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g786 ( .A1(n_598), .A2(n_787), .B1(n_790), .B2(n_793), .C(n_794), .Y(n_786) );
BUFx3_ASAP7_75t_L g1145 ( .A(n_599), .Y(n_1145) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g912 ( .A(n_610), .Y(n_912) );
AOI31xp33_ASAP7_75t_L g1483 ( .A1(n_612), .A2(n_1484), .A3(n_1492), .B(n_1502), .Y(n_1483) );
NAND4xp25_ASAP7_75t_L g613 ( .A(n_614), .B(n_617), .C(n_620), .D(n_625), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B1(n_623), .B2(n_624), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_624), .A2(n_674), .B1(n_675), .B2(n_676), .Y(n_673) );
AOI22xp33_ASAP7_75t_SL g1107 ( .A1(n_624), .A2(n_1108), .B1(n_1109), .B2(n_1110), .Y(n_1107) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_626), .A2(n_670), .B1(n_716), .B2(n_717), .Y(n_715) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g821 ( .A(n_632), .Y(n_821) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_SL g726 ( .A(n_636), .Y(n_726) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g734 ( .A(n_641), .Y(n_734) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_668), .C(n_677), .Y(n_646) );
AND3x1_ASAP7_75t_L g647 ( .A(n_648), .B(n_651), .C(n_666), .Y(n_647) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g1123 ( .A(n_654), .Y(n_1123) );
INVx2_ASAP7_75t_SL g1476 ( .A(n_654), .Y(n_1476) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g1120 ( .A(n_660), .Y(n_1120) );
BUFx3_ASAP7_75t_L g1181 ( .A(n_662), .Y(n_1181) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_673), .Y(n_668) );
OAI211xp5_ASAP7_75t_L g689 ( .A1(n_672), .A2(n_690), .B(n_692), .C(n_693), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_674), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_711) );
NAND3xp33_ASAP7_75t_L g679 ( .A(n_680), .B(n_689), .C(n_696), .Y(n_679) );
OAI211xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_682), .B(n_684), .C(n_687), .Y(n_680) );
OAI221xp5_ASAP7_75t_L g956 ( .A1(n_682), .A2(n_957), .B1(n_958), .B2(n_959), .C(n_960), .Y(n_956) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g1141 ( .A(n_683), .Y(n_1141) );
INVx2_ASAP7_75t_SL g1155 ( .A(n_683), .Y(n_1155) );
INVx1_ASAP7_75t_L g1195 ( .A(n_683), .Y(n_1195) );
BUFx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g703 ( .A(n_686), .Y(n_703) );
BUFx3_ASAP7_75t_L g955 ( .A(n_688), .Y(n_955) );
BUFx3_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g1134 ( .A(n_694), .Y(n_1134) );
HB1xp67_ASAP7_75t_L g1557 ( .A(n_694), .Y(n_1557) );
INVx1_ASAP7_75t_L g1068 ( .A(n_695), .Y(n_1068) );
BUFx2_ASAP7_75t_L g969 ( .A(n_700), .Y(n_969) );
INVx1_ASAP7_75t_L g1139 ( .A(n_702), .Y(n_1139) );
INVx1_ASAP7_75t_L g954 ( .A(n_703), .Y(n_954) );
XNOR2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_769), .Y(n_705) );
XNOR2x1_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
AND2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_750), .Y(n_708) );
NOR3xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_718), .C(n_722), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_711), .B(n_715), .Y(n_710) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_720), .Y(n_839) );
OAI22xp33_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .B1(n_727), .B2(n_728), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_SL g811 ( .A(n_726), .Y(n_811) );
OAI22xp33_ASAP7_75t_L g1037 ( .A1(n_728), .A2(n_1038), .B1(n_1039), .B2(n_1040), .Y(n_1037) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B1(n_733), .B2(n_734), .Y(n_729) );
BUFx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI22xp5_ASAP7_75t_SL g735 ( .A1(n_736), .A2(n_737), .B1(n_739), .B2(n_740), .Y(n_735) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_SL g995 ( .A(n_738), .Y(n_995) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OAI22xp33_ASAP7_75t_L g993 ( .A1(n_745), .A2(n_951), .B1(n_974), .B2(n_994), .Y(n_993) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_765), .B1(n_767), .B2(n_768), .Y(n_750) );
NAND3xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_758), .C(n_764), .Y(n_751) );
HB1xp67_ASAP7_75t_L g1501 ( .A(n_763), .Y(n_1501) );
OAI31xp33_ASAP7_75t_SL g1131 ( .A1(n_765), .A2(n_1132), .A3(n_1138), .B(n_1143), .Y(n_1131) );
INVx2_ASAP7_75t_L g1561 ( .A(n_765), .Y(n_1561) );
CKINVDCx8_ASAP7_75t_R g765 ( .A(n_766), .Y(n_765) );
AOI31xp33_ASAP7_75t_L g1189 ( .A1(n_766), .A2(n_1190), .A3(n_1196), .B(n_1207), .Y(n_1189) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_797), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_773), .B1(n_795), .B2(n_796), .Y(n_771) );
NAND3xp33_ASAP7_75t_SL g773 ( .A(n_774), .B(n_777), .C(n_786), .Y(n_773) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g1019 ( .A(n_781), .Y(n_1019) );
INVx2_ASAP7_75t_SL g1206 ( .A(n_781), .Y(n_1206) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx2_ASAP7_75t_SL g968 ( .A(n_789), .Y(n_968) );
INVx4_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g871 ( .A(n_792), .Y(n_871) );
AOI21xp5_ASAP7_75t_L g947 ( .A1(n_796), .A2(n_948), .B(n_949), .Y(n_947) );
NOR3xp33_ASAP7_75t_L g797 ( .A(n_798), .B(n_807), .C(n_809), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_803), .Y(n_798) );
INVx1_ASAP7_75t_L g833 ( .A(n_806), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_806), .A2(n_832), .B1(n_959), .B2(n_979), .Y(n_978) );
OAI22xp33_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_812), .B1(n_813), .B2(n_815), .Y(n_810) );
OAI22xp33_ASAP7_75t_L g1046 ( .A1(n_813), .A2(n_1021), .B1(n_1023), .B2(n_1039), .Y(n_1046) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_818), .B1(n_820), .B2(n_821), .Y(n_816) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx2_ASAP7_75t_L g1043 ( .A(n_819), .Y(n_1043) );
INVx2_ASAP7_75t_L g1080 ( .A(n_819), .Y(n_1080) );
INVx1_ASAP7_75t_L g1001 ( .A(n_824), .Y(n_1001) );
XNOR2xp5_ASAP7_75t_L g824 ( .A(n_825), .B(n_892), .Y(n_824) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
XNOR2xp5_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
OAI22xp5_ASAP7_75t_SL g1255 ( .A1(n_827), .A2(n_1256), .B1(n_1257), .B2(n_1258), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_829), .B(n_861), .Y(n_828) );
NOR3xp33_ASAP7_75t_SL g829 ( .A(n_830), .B(n_838), .C(n_840), .Y(n_829) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
OAI22xp33_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_844), .B1(n_845), .B2(n_846), .Y(n_841) );
OAI22xp33_ASAP7_75t_L g856 ( .A1(n_842), .A2(n_845), .B1(n_857), .B2(n_858), .Y(n_856) );
OAI22xp33_ASAP7_75t_L g1528 ( .A1(n_842), .A2(n_1529), .B1(n_1530), .B2(n_1531), .Y(n_1528) );
INVx3_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
OAI22xp5_ASAP7_75t_L g1045 ( .A1(n_850), .A2(n_1013), .B1(n_1024), .B2(n_1043), .Y(n_1045) );
OAI22xp5_ASAP7_75t_L g1078 ( .A1(n_850), .A2(n_1079), .B1(n_1080), .B2(n_1081), .Y(n_1078) );
OAI22xp33_ASAP7_75t_L g1541 ( .A1(n_850), .A2(n_1530), .B1(n_1542), .B2(n_1543), .Y(n_1541) );
AOI221xp5_ASAP7_75t_SL g864 ( .A1(n_852), .A2(n_865), .B1(n_872), .B2(n_874), .C(n_876), .Y(n_864) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
AOI221xp5_ASAP7_75t_L g880 ( .A1(n_858), .A2(n_881), .B1(n_884), .B2(n_887), .C(n_889), .Y(n_880) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
AOI31xp33_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_880), .A3(n_890), .B(n_891), .Y(n_863) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx3_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx2_ASAP7_75t_L g1203 ( .A(n_869), .Y(n_1203) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx3_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
CKINVDCx5p33_ASAP7_75t_R g887 ( .A(n_888), .Y(n_887) );
AOI22xp5_ASAP7_75t_L g892 ( .A1(n_893), .A2(n_944), .B1(n_998), .B2(n_999), .Y(n_892) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g999 ( .A(n_894), .Y(n_999) );
INVx2_ASAP7_75t_SL g943 ( .A(n_895), .Y(n_943) );
AND2x2_ASAP7_75t_L g895 ( .A(n_896), .B(n_916), .Y(n_895) );
AOI22xp5_ASAP7_75t_L g898 ( .A1(n_899), .A2(n_902), .B1(n_903), .B2(n_904), .Y(n_898) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
OAI22xp33_ASAP7_75t_L g936 ( .A1(n_907), .A2(n_937), .B1(n_939), .B2(n_940), .Y(n_936) );
NOR2xp33_ASAP7_75t_L g916 ( .A(n_917), .B(n_927), .Y(n_916) );
BUFx3_ASAP7_75t_L g1177 ( .A(n_924), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_928), .B(n_932), .Y(n_927) );
INVx3_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVx2_ASAP7_75t_SL g998 ( .A(n_944), .Y(n_998) );
INVx1_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_947), .B(n_976), .Y(n_946) );
AOI211xp5_ASAP7_75t_L g950 ( .A1(n_951), .A2(n_952), .B(n_953), .C(n_961), .Y(n_950) );
OAI221xp5_ASAP7_75t_L g1194 ( .A1(n_960), .A2(n_1065), .B1(n_1172), .B2(n_1174), .C(n_1195), .Y(n_1194) );
OAI221xp5_ASAP7_75t_L g1552 ( .A1(n_960), .A2(n_1065), .B1(n_1521), .B2(n_1523), .C(n_1553), .Y(n_1552) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
NOR3xp33_ASAP7_75t_L g976 ( .A(n_977), .B(n_982), .C(n_983), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_978), .B(n_980), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_988), .A2(n_990), .B1(n_991), .B2(n_992), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
OAI22xp5_ASAP7_75t_SL g1041 ( .A1(n_991), .A2(n_1042), .B1(n_1043), .B2(n_1044), .Y(n_1041) );
OAI221xp5_ASAP7_75t_L g1125 ( .A1(n_991), .A2(n_995), .B1(n_1126), .B2(n_1127), .C(n_1128), .Y(n_1125) );
BUFx2_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_1003), .A2(n_1097), .B1(n_1098), .B2(n_1211), .Y(n_1002) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1003), .Y(n_1211) );
AO22x1_ASAP7_75t_L g1003 ( .A1(n_1004), .A2(n_1048), .B1(n_1049), .B2(n_1096), .Y(n_1003) );
BUFx2_ASAP7_75t_SL g1004 ( .A(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1005), .Y(n_1096) );
XOR2x2_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1047), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1026), .Y(n_1006) );
NAND3xp33_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1015), .C(n_1022), .Y(n_1008) );
NOR3xp33_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1034), .C(n_1036), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1031), .Y(n_1027) );
OAI22xp33_ASAP7_75t_L g1082 ( .A1(n_1039), .A2(n_1083), .B1(n_1084), .B2(n_1085), .Y(n_1082) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_1043), .A2(n_1056), .B1(n_1075), .B2(n_1088), .Y(n_1087) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1076), .Y(n_1051) );
INVx2_ASAP7_75t_SL g1060 ( .A(n_1061), .Y(n_1060) );
OAI221xp5_ASAP7_75t_L g1062 ( .A1(n_1063), .A2(n_1064), .B1(n_1065), .B2(n_1067), .C(n_1068), .Y(n_1062) );
OAI221xp5_ASAP7_75t_L g1491 ( .A1(n_1063), .A2(n_1065), .B1(n_1142), .B2(n_1466), .C(n_1468), .Y(n_1491) );
OAI221xp5_ASAP7_75t_L g1140 ( .A1(n_1065), .A2(n_1106), .B1(n_1112), .B2(n_1141), .C(n_1142), .Y(n_1140) );
INVx2_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
NOR3xp33_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1090), .C(n_1091), .Y(n_1076) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1086), .Y(n_1530) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_1092), .B(n_1094), .Y(n_1091) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
AO22x2_ASAP7_75t_L g1098 ( .A1(n_1099), .A2(n_1161), .B1(n_1162), .B2(n_1210), .Y(n_1098) );
HB1xp67_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1100), .Y(n_1210) );
NAND4xp25_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1111), .C(n_1131), .D(n_1156), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1107), .Y(n_1102) );
OAI221xp5_ASAP7_75t_L g1114 ( .A1(n_1115), .A2(n_1118), .B1(n_1119), .B2(n_1121), .C(n_1122), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g1532 ( .A1(n_1115), .A2(n_1533), .B1(n_1534), .B2(n_1537), .Y(n_1532) );
INVx2_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
INVx2_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
BUFx6f_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
NAND3xp33_ASAP7_75t_L g1143 ( .A(n_1144), .B(n_1146), .C(n_1149), .Y(n_1143) );
INVx2_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_SL g1161 ( .A(n_1162), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1186), .Y(n_1163) );
AND4x1_ASAP7_75t_L g1164 ( .A(n_1165), .B(n_1169), .C(n_1173), .D(n_1176), .Y(n_1164) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
AOI21xp33_ASAP7_75t_L g1186 ( .A1(n_1187), .A2(n_1188), .B(n_1189), .Y(n_1186) );
AOI21xp5_ASAP7_75t_L g1544 ( .A1(n_1187), .A2(n_1545), .B(n_1546), .Y(n_1544) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
BUFx2_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
OAI221xp5_ASAP7_75t_L g1212 ( .A1(n_1213), .A2(n_1453), .B1(n_1455), .B2(n_1505), .C(n_1509), .Y(n_1212) );
NOR2xp33_ASAP7_75t_L g1213 ( .A(n_1214), .B(n_1385), .Y(n_1213) );
OAI211xp5_ASAP7_75t_L g1214 ( .A1(n_1215), .A2(n_1329), .B(n_1356), .C(n_1372), .Y(n_1214) );
AOI21xp33_ASAP7_75t_L g1215 ( .A1(n_1216), .A2(n_1304), .B(n_1305), .Y(n_1215) );
AOI21xp5_ASAP7_75t_L g1329 ( .A1(n_1216), .A2(n_1330), .B(n_1355), .Y(n_1329) );
OAI211xp5_ASAP7_75t_L g1216 ( .A1(n_1217), .A2(n_1243), .B(n_1259), .C(n_1284), .Y(n_1216) );
NOR2xp33_ASAP7_75t_L g1414 ( .A(n_1217), .B(n_1415), .Y(n_1414) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1219), .B(n_1240), .Y(n_1218) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1219), .Y(n_1312) );
NOR2xp33_ASAP7_75t_L g1348 ( .A(n_1219), .B(n_1240), .Y(n_1348) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1220), .B(n_1262), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1220), .B(n_1263), .Y(n_1289) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1221), .B(n_1281), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1221), .B(n_1263), .Y(n_1337) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1234), .Y(n_1221) );
AND2x4_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1229), .Y(n_1223) );
OAI21xp33_ASAP7_75t_SL g1564 ( .A1(n_1224), .A2(n_1513), .B(n_1565), .Y(n_1564) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1273 ( .A(n_1225), .B(n_1230), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1228), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1228), .Y(n_1238) );
AND2x4_ASAP7_75t_L g1231 ( .A(n_1229), .B(n_1232), .Y(n_1231) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
OR2x2_ASAP7_75t_L g1276 ( .A(n_1230), .B(n_1233), .Y(n_1276) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1236), .B(n_1237), .Y(n_1235) );
AND2x4_ASAP7_75t_L g1239 ( .A(n_1236), .B(n_1238), .Y(n_1239) );
AND2x4_ASAP7_75t_L g1249 ( .A(n_1236), .B(n_1237), .Y(n_1249) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
INVx2_ASAP7_75t_L g1258 ( .A(n_1239), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1240), .B(n_1267), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1240), .B(n_1280), .Y(n_1279) );
CKINVDCx5p33_ASAP7_75t_R g1291 ( .A(n_1240), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1240), .B(n_1312), .Y(n_1311) );
OR2x2_ASAP7_75t_L g1321 ( .A(n_1240), .B(n_1312), .Y(n_1321) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1240), .B(n_1263), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1240), .B(n_1289), .Y(n_1327) );
OR2x2_ASAP7_75t_L g1366 ( .A(n_1240), .B(n_1346), .Y(n_1366) );
NOR2xp33_ASAP7_75t_L g1375 ( .A(n_1240), .B(n_1345), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1420 ( .A(n_1240), .B(n_1261), .Y(n_1420) );
AND2x4_ASAP7_75t_SL g1240 ( .A(n_1241), .B(n_1242), .Y(n_1240) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1243), .Y(n_1359) );
NOR2xp33_ASAP7_75t_L g1383 ( .A(n_1243), .B(n_1384), .Y(n_1383) );
OR2x2_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1253), .Y(n_1243) );
INVx2_ASAP7_75t_L g1389 ( .A(n_1244), .Y(n_1389) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1244), .Y(n_1416) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1245), .B(n_1250), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1245), .B(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1246), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1246), .B(n_1287), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_1246), .B(n_1250), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1354 ( .A(n_1246), .B(n_1253), .Y(n_1354) );
BUFx6f_ASAP7_75t_L g1362 ( .A(n_1246), .Y(n_1362) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1247), .B(n_1248), .Y(n_1246) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1249), .Y(n_1256) );
BUFx3_ASAP7_75t_L g1295 ( .A(n_1249), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1250), .B(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1250), .Y(n_1287) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1250), .Y(n_1328) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1250), .Y(n_1352) );
AOI321xp33_ASAP7_75t_L g1372 ( .A1(n_1250), .A2(n_1373), .A3(n_1376), .B1(n_1378), .B2(n_1380), .C(n_1383), .Y(n_1372) );
NAND2xp5_ASAP7_75t_SL g1378 ( .A(n_1250), .B(n_1379), .Y(n_1378) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1251), .B(n_1252), .Y(n_1250) );
CKINVDCx6p67_ASAP7_75t_R g1278 ( .A(n_1253), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1303 ( .A(n_1253), .B(n_1293), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1253), .B(n_1283), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_1253), .B(n_1351), .Y(n_1350) );
CKINVDCx5p33_ASAP7_75t_R g1355 ( .A(n_1253), .Y(n_1355) );
OR2x2_ASAP7_75t_L g1430 ( .A(n_1253), .B(n_1283), .Y(n_1430) );
OR2x6_ASAP7_75t_L g1253 ( .A(n_1254), .B(n_1255), .Y(n_1253) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_1254), .B(n_1255), .Y(n_1435) );
INVx2_ASAP7_75t_L g1269 ( .A(n_1258), .Y(n_1269) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1258), .Y(n_1296) );
AOI22xp5_ASAP7_75t_L g1259 ( .A1(n_1260), .A2(n_1277), .B1(n_1279), .B2(n_1282), .Y(n_1259) );
O2A1O1Ixp33_ASAP7_75t_L g1313 ( .A1(n_1260), .A2(n_1314), .B(n_1318), .C(n_1319), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1261), .B(n_1266), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1261), .B(n_1391), .Y(n_1390) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1261), .B(n_1291), .Y(n_1411) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
INVxp67_ASAP7_75t_SL g1281 ( .A(n_1263), .Y(n_1281) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1263), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1264), .B(n_1265), .Y(n_1263) );
AOI211xp5_ASAP7_75t_L g1333 ( .A1(n_1266), .A2(n_1320), .B(n_1334), .C(n_1338), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1266), .B(n_1280), .Y(n_1405) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1266), .B(n_1289), .Y(n_1418) );
INVx2_ASAP7_75t_SL g1310 ( .A(n_1267), .Y(n_1310) );
BUFx2_ASAP7_75t_L g1316 ( .A(n_1267), .Y(n_1316) );
NOR2xp33_ASAP7_75t_L g1336 ( .A(n_1267), .B(n_1287), .Y(n_1336) );
BUFx3_ASAP7_75t_L g1343 ( .A(n_1267), .Y(n_1343) );
INVx2_ASAP7_75t_SL g1267 ( .A(n_1268), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1268), .B(n_1291), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1434 ( .A(n_1268), .B(n_1287), .Y(n_1434) );
OAI22xp33_ASAP7_75t_L g1270 ( .A1(n_1271), .A2(n_1272), .B1(n_1274), .B2(n_1275), .Y(n_1270) );
BUFx3_ASAP7_75t_L g1299 ( .A(n_1272), .Y(n_1299) );
BUFx6f_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
HB1xp67_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1276), .Y(n_1302) );
AOI22xp33_ASAP7_75t_L g1426 ( .A1(n_1277), .A2(n_1324), .B1(n_1427), .B2(n_1429), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1278), .B(n_1283), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1278), .B(n_1292), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1438 ( .A(n_1278), .B(n_1307), .Y(n_1438) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1279), .Y(n_1384) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1280), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1280), .B(n_1291), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_1280), .B(n_1290), .Y(n_1450) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1282), .Y(n_1379) );
AOI21xp33_ASAP7_75t_SL g1431 ( .A1(n_1282), .A2(n_1327), .B(n_1432), .Y(n_1431) );
NAND2xp5_ASAP7_75t_L g1377 ( .A(n_1283), .B(n_1292), .Y(n_1377) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1283), .Y(n_1445) );
A2O1A1Ixp33_ASAP7_75t_SL g1284 ( .A1(n_1285), .A2(n_1288), .B(n_1292), .C(n_1303), .Y(n_1284) );
NOR2xp33_ASAP7_75t_L g1451 ( .A(n_1285), .B(n_1452), .Y(n_1451) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_1286), .B(n_1310), .Y(n_1394) );
OAI21xp33_ASAP7_75t_L g1419 ( .A1(n_1286), .A2(n_1357), .B(n_1420), .Y(n_1419) );
OAI21xp5_ASAP7_75t_L g1423 ( .A1(n_1286), .A2(n_1408), .B(n_1424), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1289), .B(n_1290), .Y(n_1288) );
INVx2_ASAP7_75t_L g1320 ( .A(n_1289), .Y(n_1320) );
OAI21xp5_ASAP7_75t_SL g1367 ( .A1(n_1289), .A2(n_1368), .B(n_1369), .Y(n_1367) );
NAND2xp5_ASAP7_75t_L g1382 ( .A(n_1289), .B(n_1310), .Y(n_1382) );
OR2x2_ASAP7_75t_L g1339 ( .A(n_1291), .B(n_1315), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1291), .B(n_1358), .Y(n_1357) );
OR2x2_ASAP7_75t_L g1381 ( .A(n_1291), .B(n_1382), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1291), .B(n_1337), .Y(n_1397) );
INVx2_ASAP7_75t_L g1371 ( .A(n_1292), .Y(n_1371) );
A2O1A1Ixp33_ASAP7_75t_L g1395 ( .A1(n_1292), .A2(n_1361), .B(n_1396), .C(n_1398), .Y(n_1395) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
OAI22xp33_ASAP7_75t_L g1297 ( .A1(n_1298), .A2(n_1299), .B1(n_1300), .B2(n_1301), .Y(n_1297) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1299), .Y(n_1454) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1303), .Y(n_1439) );
OAI211xp5_ASAP7_75t_SL g1305 ( .A1(n_1306), .A2(n_1308), .B(n_1313), .C(n_1323), .Y(n_1305) );
A2O1A1Ixp33_ASAP7_75t_L g1387 ( .A1(n_1306), .A2(n_1308), .B(n_1325), .C(n_1388), .Y(n_1387) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
NAND2xp5_ASAP7_75t_L g1322 ( .A(n_1307), .B(n_1316), .Y(n_1322) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1309), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1309 ( .A(n_1310), .B(n_1311), .Y(n_1309) );
NOR2xp33_ASAP7_75t_L g1338 ( .A(n_1310), .B(n_1317), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1310), .B(n_1348), .Y(n_1347) );
NOR2x1p5_ASAP7_75t_L g1358 ( .A(n_1310), .B(n_1320), .Y(n_1358) );
HB1xp67_ASAP7_75t_L g1410 ( .A(n_1310), .Y(n_1410) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1311), .B(n_1343), .Y(n_1425) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
OR2x2_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1317), .Y(n_1315) );
OR2x2_ASAP7_75t_L g1325 ( .A(n_1316), .B(n_1326), .Y(n_1325) );
NOR2xp33_ASAP7_75t_L g1365 ( .A(n_1316), .B(n_1366), .Y(n_1365) );
NAND2xp5_ASAP7_75t_L g1374 ( .A(n_1316), .B(n_1375), .Y(n_1374) );
INVx2_ASAP7_75t_L g1400 ( .A(n_1316), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_1316), .B(n_1445), .Y(n_1444) );
NOR2xp33_ASAP7_75t_L g1392 ( .A(n_1317), .B(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1318), .Y(n_1342) );
AOI21xp33_ASAP7_75t_SL g1319 ( .A1(n_1320), .A2(n_1321), .B(n_1322), .Y(n_1319) );
OAI21xp33_ASAP7_75t_L g1427 ( .A1(n_1321), .A2(n_1400), .B(n_1428), .Y(n_1427) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1322), .Y(n_1369) );
OAI21xp5_ASAP7_75t_L g1323 ( .A1(n_1324), .A2(n_1327), .B(n_1328), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1326), .Y(n_1442) );
NAND2xp67_ASAP7_75t_L g1404 ( .A(n_1328), .B(n_1405), .Y(n_1404) );
NAND2xp5_ASAP7_75t_L g1449 ( .A(n_1328), .B(n_1450), .Y(n_1449) );
OAI211xp5_ASAP7_75t_L g1330 ( .A1(n_1331), .A2(n_1333), .B(n_1339), .C(n_1340), .Y(n_1330) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1336), .B(n_1337), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1413 ( .A(n_1336), .B(n_1411), .Y(n_1413) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1337), .Y(n_1436) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_1337), .B(n_1438), .Y(n_1437) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1339), .Y(n_1360) );
A2O1A1Ixp33_ASAP7_75t_L g1340 ( .A1(n_1341), .A2(n_1344), .B(n_1347), .C(n_1349), .Y(n_1340) );
NOR2xp33_ASAP7_75t_L g1341 ( .A(n_1342), .B(n_1343), .Y(n_1341) );
O2A1O1Ixp33_ASAP7_75t_SL g1363 ( .A1(n_1342), .A2(n_1364), .B(n_1367), .C(n_1370), .Y(n_1363) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1343), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1396 ( .A(n_1343), .B(n_1397), .Y(n_1396) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1350), .B(n_1353), .Y(n_1349) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1351), .Y(n_1402) );
INVx3_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
AOI31xp33_ASAP7_75t_L g1406 ( .A1(n_1355), .A2(n_1407), .A3(n_1417), .B(n_1419), .Y(n_1406) );
AOI221xp5_ASAP7_75t_L g1356 ( .A1(n_1357), .A2(n_1359), .B1(n_1360), .B2(n_1361), .C(n_1363), .Y(n_1356) );
AOI211xp5_ASAP7_75t_L g1407 ( .A1(n_1361), .A2(n_1408), .B(n_1412), .C(n_1414), .Y(n_1407) );
CKINVDCx14_ASAP7_75t_R g1361 ( .A(n_1362), .Y(n_1361) );
OAI21xp33_ASAP7_75t_L g1417 ( .A1(n_1362), .A2(n_1403), .B(n_1418), .Y(n_1417) );
OAI221xp5_ASAP7_75t_L g1440 ( .A1(n_1362), .A2(n_1396), .B1(n_1441), .B2(n_1443), .C(n_1446), .Y(n_1440) );
INVxp67_ASAP7_75t_SL g1364 ( .A(n_1365), .Y(n_1364) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1368), .Y(n_1428) );
AOI21xp5_ASAP7_75t_L g1388 ( .A1(n_1370), .A2(n_1389), .B(n_1390), .Y(n_1388) );
AOI22xp5_ASAP7_75t_L g1421 ( .A1(n_1370), .A2(n_1422), .B1(n_1439), .B2(n_1440), .Y(n_1421) );
INVx3_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1375), .B(n_1400), .Y(n_1399) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
INVx2_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
NAND2xp5_ASAP7_75t_L g1385 ( .A(n_1386), .B(n_1421), .Y(n_1385) );
O2A1O1Ixp33_ASAP7_75t_L g1386 ( .A1(n_1387), .A2(n_1392), .B(n_1395), .C(n_1406), .Y(n_1386) );
NAND2xp5_ASAP7_75t_L g1415 ( .A(n_1391), .B(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1397), .Y(n_1452) );
AOI21xp5_ASAP7_75t_L g1398 ( .A1(n_1399), .A2(n_1401), .B(n_1403), .Y(n_1398) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1402), .Y(n_1447) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1404), .Y(n_1403) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
NAND2xp5_ASAP7_75t_L g1409 ( .A(n_1410), .B(n_1411), .Y(n_1409) );
NOR2xp33_ASAP7_75t_L g1441 ( .A(n_1411), .B(n_1442), .Y(n_1441) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
AOI211xp5_ASAP7_75t_SL g1446 ( .A1(n_1418), .A2(n_1447), .B(n_1448), .C(n_1451), .Y(n_1446) );
NAND4xp25_ASAP7_75t_L g1422 ( .A(n_1423), .B(n_1426), .C(n_1431), .D(n_1437), .Y(n_1422) );
INVxp67_ASAP7_75t_SL g1424 ( .A(n_1425), .Y(n_1424) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
NOR3xp33_ASAP7_75t_L g1432 ( .A(n_1433), .B(n_1435), .C(n_1436), .Y(n_1432) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
XNOR2x1_ASAP7_75t_L g1456 ( .A(n_1457), .B(n_1458), .Y(n_1456) );
AND2x4_ASAP7_75t_L g1458 ( .A(n_1459), .B(n_1481), .Y(n_1458) );
AND4x1_ASAP7_75t_L g1459 ( .A(n_1460), .B(n_1464), .C(n_1467), .D(n_1470), .Y(n_1459) );
INVx2_ASAP7_75t_SL g1473 ( .A(n_1474), .Y(n_1473) );
INVx2_ASAP7_75t_L g1480 ( .A(n_1474), .Y(n_1480) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
BUFx2_ASAP7_75t_SL g1498 ( .A(n_1499), .Y(n_1498) );
INVx4_ASAP7_75t_SL g1505 ( .A(n_1506), .Y(n_1505) );
BUFx3_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
BUFx2_ASAP7_75t_L g1507 ( .A(n_1508), .Y(n_1507) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
CKINVDCx5p33_ASAP7_75t_R g1511 ( .A(n_1512), .Y(n_1511) );
INVxp33_ASAP7_75t_SL g1514 ( .A(n_1515), .Y(n_1514) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1516), .Y(n_1563) );
AND2x2_ASAP7_75t_L g1516 ( .A(n_1517), .B(n_1544), .Y(n_1516) );
NOR3xp33_ASAP7_75t_L g1517 ( .A(n_1518), .B(n_1525), .C(n_1527), .Y(n_1517) );
NAND2xp5_ASAP7_75t_L g1518 ( .A(n_1519), .B(n_1522), .Y(n_1518) );
INVx2_ASAP7_75t_SL g1534 ( .A(n_1535), .Y(n_1534) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
AOI31xp33_ASAP7_75t_L g1546 ( .A1(n_1547), .A2(n_1554), .A3(n_1560), .B(n_1561), .Y(n_1546) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
endmodule