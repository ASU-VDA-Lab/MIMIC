module real_aes_7113_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_532;
wire n_284;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_735;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_283;
wire n_252;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g271 ( .A1(n_0), .A2(n_272), .B(n_273), .C(n_276), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_1), .B(n_260), .Y(n_277) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_2), .B(n_109), .C(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g123 ( .A(n_2), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_3), .B(n_188), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_4), .A2(n_149), .B(n_152), .C(n_532), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_5), .A2(n_144), .B(n_556), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_6), .A2(n_144), .B(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_7), .B(n_260), .Y(n_562) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_8), .A2(n_179), .B(n_216), .Y(n_215) );
AND2x6_ASAP7_75t_L g149 ( .A(n_9), .B(n_150), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_10), .A2(n_149), .B(n_152), .C(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g500 ( .A(n_11), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_12), .B(n_40), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_12), .B(n_40), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_13), .B(n_236), .Y(n_534) );
INVx1_ASAP7_75t_L g170 ( .A(n_14), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_15), .B(n_188), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_16), .A2(n_189), .B(n_518), .C(n_520), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_17), .B(n_260), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_18), .B(n_164), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g151 ( .A1(n_19), .A2(n_152), .B(n_155), .C(n_163), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_20), .A2(n_224), .B(n_275), .C(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_21), .B(n_236), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_22), .A2(n_54), .B1(n_754), .B2(n_755), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_22), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_23), .B(n_236), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_24), .Y(n_547) );
INVx1_ASAP7_75t_L g472 ( .A(n_25), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_26), .A2(n_152), .B(n_163), .C(n_219), .Y(n_218) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_27), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_28), .Y(n_530) );
INVx1_ASAP7_75t_L g488 ( .A(n_29), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_30), .A2(n_144), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g147 ( .A(n_31), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_32), .A2(n_192), .B(n_201), .C(n_203), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_33), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_34), .A2(n_275), .B(n_559), .C(n_561), .Y(n_558) );
INVxp67_ASAP7_75t_L g489 ( .A(n_35), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_36), .B(n_221), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_37), .A2(n_152), .B(n_163), .C(n_471), .Y(n_470) );
CKINVDCx14_ASAP7_75t_R g557 ( .A(n_38), .Y(n_557) );
AOI222xp33_ASAP7_75t_SL g126 ( .A1(n_39), .A2(n_127), .B1(n_133), .B2(n_738), .C1(n_739), .C2(n_743), .Y(n_126) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_41), .A2(n_276), .B(n_498), .C(n_499), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_42), .B(n_143), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_43), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_44), .B(n_188), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_45), .B(n_144), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_46), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_47), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_48), .A2(n_192), .B(n_201), .C(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g274 ( .A(n_49), .Y(n_274) );
OAI22xp5_ASAP7_75t_SL g751 ( .A1(n_50), .A2(n_752), .B1(n_753), .B2(n_756), .Y(n_751) );
CKINVDCx16_ASAP7_75t_R g756 ( .A(n_50), .Y(n_756) );
INVx1_ASAP7_75t_L g246 ( .A(n_51), .Y(n_246) );
INVx1_ASAP7_75t_L g506 ( .A(n_52), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_53), .B(n_144), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_54), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_55), .Y(n_172) );
CKINVDCx14_ASAP7_75t_R g496 ( .A(n_56), .Y(n_496) );
INVx1_ASAP7_75t_L g150 ( .A(n_57), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_58), .B(n_144), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_59), .B(n_260), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_60), .A2(n_162), .B(n_185), .C(n_257), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_61), .Y(n_125) );
INVx1_ASAP7_75t_L g169 ( .A(n_62), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g128 ( .A1(n_63), .A2(n_102), .B1(n_129), .B2(n_130), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_63), .Y(n_130) );
INVx1_ASAP7_75t_SL g560 ( .A(n_64), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_65), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_66), .B(n_188), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_67), .B(n_260), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_68), .B(n_189), .Y(n_234) );
INVx1_ASAP7_75t_L g550 ( .A(n_69), .Y(n_550) );
CKINVDCx16_ASAP7_75t_R g270 ( .A(n_70), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_71), .B(n_157), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g182 ( .A1(n_72), .A2(n_152), .B(n_183), .C(n_192), .Y(n_182) );
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_73), .Y(n_255) );
INVx1_ASAP7_75t_L g112 ( .A(n_74), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_75), .A2(n_144), .B(n_495), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_76), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_77), .A2(n_144), .B(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_78), .A2(n_104), .B1(n_113), .B2(n_758), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_79), .A2(n_143), .B(n_484), .Y(n_483) );
CKINVDCx16_ASAP7_75t_R g469 ( .A(n_80), .Y(n_469) );
INVx1_ASAP7_75t_L g516 ( .A(n_81), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_82), .B(n_160), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_83), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_84), .A2(n_144), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g519 ( .A(n_85), .Y(n_519) );
INVx2_ASAP7_75t_L g167 ( .A(n_86), .Y(n_167) );
INVx1_ASAP7_75t_L g533 ( .A(n_87), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_88), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_89), .B(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g109 ( .A(n_90), .Y(n_109) );
OR2x2_ASAP7_75t_L g120 ( .A(n_90), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g461 ( .A(n_90), .B(n_122), .Y(n_461) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_91), .A2(n_128), .B1(n_131), .B2(n_132), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_91), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_92), .A2(n_152), .B(n_192), .C(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_93), .B(n_144), .Y(n_199) );
INVx1_ASAP7_75t_L g204 ( .A(n_94), .Y(n_204) );
INVxp67_ASAP7_75t_L g258 ( .A(n_95), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_96), .B(n_179), .Y(n_501) );
INVx2_ASAP7_75t_L g509 ( .A(n_97), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g184 ( .A(n_99), .Y(n_184) );
INVx1_ASAP7_75t_L g230 ( .A(n_100), .Y(n_230) );
AND2x2_ASAP7_75t_L g248 ( .A(n_101), .B(n_166), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_102), .Y(n_129) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g758 ( .A(n_106), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
OR2x2_ASAP7_75t_L g737 ( .A(n_109), .B(n_122), .Y(n_737) );
NOR2x2_ASAP7_75t_L g745 ( .A(n_109), .B(n_121), .Y(n_745) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AOI22x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_126), .B1(n_746), .B2(n_748), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g747 ( .A(n_117), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_118), .A2(n_749), .B(n_757), .Y(n_748) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_125), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g757 ( .A(n_120), .Y(n_757) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g738 ( .A(n_127), .Y(n_738) );
INVx1_ASAP7_75t_L g131 ( .A(n_128), .Y(n_131) );
OAI22xp5_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_459), .B1(n_462), .B2(n_735), .Y(n_133) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_134), .A2(n_741), .B1(n_750), .B2(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx2_ASAP7_75t_L g741 ( .A(n_135), .Y(n_741) );
AND3x1_ASAP7_75t_L g135 ( .A(n_136), .B(n_363), .C(n_420), .Y(n_135) );
NOR3xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_308), .C(n_344), .Y(n_136) );
OAI211xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_210), .B(n_262), .C(n_295), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_174), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x4_ASAP7_75t_L g265 ( .A(n_140), .B(n_266), .Y(n_265) );
INVx5_ASAP7_75t_L g294 ( .A(n_140), .Y(n_294) );
AND2x2_ASAP7_75t_L g367 ( .A(n_140), .B(n_283), .Y(n_367) );
AND2x2_ASAP7_75t_L g405 ( .A(n_140), .B(n_311), .Y(n_405) );
AND2x2_ASAP7_75t_L g425 ( .A(n_140), .B(n_267), .Y(n_425) );
OR2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_171), .Y(n_140) );
AOI21xp5_ASAP7_75t_SL g141 ( .A1(n_142), .A2(n_151), .B(n_164), .Y(n_141) );
BUFx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_149), .Y(n_144) );
NAND2x1p5_ASAP7_75t_L g231 ( .A(n_145), .B(n_149), .Y(n_231) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
INVx1_ASAP7_75t_L g162 ( .A(n_146), .Y(n_162) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx1_ASAP7_75t_L g225 ( .A(n_147), .Y(n_225) );
INVx1_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_148), .Y(n_158) );
INVx3_ASAP7_75t_L g189 ( .A(n_148), .Y(n_189) );
INVx1_ASAP7_75t_L g221 ( .A(n_148), .Y(n_221) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_148), .Y(n_236) );
BUFx3_ASAP7_75t_L g163 ( .A(n_149), .Y(n_163) );
INVx4_ASAP7_75t_SL g193 ( .A(n_149), .Y(n_193) );
INVx5_ASAP7_75t_L g202 ( .A(n_152), .Y(n_202) );
AND2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_153), .Y(n_191) );
BUFx3_ASAP7_75t_L g207 ( .A(n_153), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_159), .B(n_161), .Y(n_155) );
INVx2_ASAP7_75t_L g160 ( .A(n_157), .Y(n_160) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx4_ASAP7_75t_L g186 ( .A(n_158), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_160), .A2(n_204), .B(n_205), .C(n_206), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_160), .A2(n_206), .B(n_246), .C(n_247), .Y(n_245) );
O2A1O1Ixp5_ASAP7_75t_L g532 ( .A1(n_160), .A2(n_533), .B(n_534), .C(n_535), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_L g549 ( .A1(n_160), .A2(n_535), .B(n_550), .C(n_551), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_161), .A2(n_188), .B(n_472), .C(n_473), .Y(n_471) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_162), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_165), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g173 ( .A(n_166), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_166), .A2(n_199), .B(n_200), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_166), .A2(n_243), .B(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_166), .A2(n_231), .B(n_469), .C(n_470), .Y(n_468) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_166), .A2(n_494), .B(n_501), .Y(n_493) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_167), .B(n_168), .Y(n_166) );
AND2x2_ASAP7_75t_L g180 ( .A(n_167), .B(n_168), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_173), .A2(n_529), .B(n_536), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_174), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_197), .Y(n_174) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_175), .Y(n_306) );
AND2x2_ASAP7_75t_L g320 ( .A(n_175), .B(n_266), .Y(n_320) );
INVx1_ASAP7_75t_L g343 ( .A(n_175), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_175), .B(n_294), .Y(n_382) );
OR2x2_ASAP7_75t_L g419 ( .A(n_175), .B(n_264), .Y(n_419) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_176), .Y(n_355) );
AND2x2_ASAP7_75t_L g362 ( .A(n_176), .B(n_267), .Y(n_362) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g283 ( .A(n_177), .B(n_267), .Y(n_283) );
BUFx2_ASAP7_75t_L g311 ( .A(n_177), .Y(n_311) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_181), .B(n_195), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_178), .B(n_196), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_178), .B(n_209), .Y(n_208) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_178), .A2(n_229), .B(n_237), .Y(n_228) );
INVx3_ASAP7_75t_L g260 ( .A(n_178), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_178), .B(n_475), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_178), .B(n_537), .Y(n_536) );
AO21x2_ASAP7_75t_L g545 ( .A1(n_178), .A2(n_546), .B(n_552), .Y(n_545) );
INVx4_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_179), .A2(n_217), .B(n_218), .Y(n_216) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_179), .Y(n_252) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g239 ( .A(n_180), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_194), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_187), .C(n_190), .Y(n_183) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_186), .A2(n_188), .B1(n_488), .B2(n_489), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_186), .B(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_186), .B(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_188), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g272 ( .A(n_188), .Y(n_272) );
INVx5_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_189), .B(n_500), .Y(n_499) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx3_ASAP7_75t_L g561 ( .A(n_191), .Y(n_561) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_193), .A2(n_202), .B(n_255), .C(n_256), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_SL g269 ( .A1(n_193), .A2(n_202), .B(n_270), .C(n_271), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_SL g484 ( .A1(n_193), .A2(n_202), .B(n_485), .C(n_486), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_SL g495 ( .A1(n_193), .A2(n_202), .B(n_496), .C(n_497), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_SL g505 ( .A1(n_193), .A2(n_202), .B(n_506), .C(n_507), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_SL g515 ( .A1(n_193), .A2(n_202), .B(n_516), .C(n_517), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_L g556 ( .A1(n_193), .A2(n_202), .B(n_557), .C(n_558), .Y(n_556) );
INVx5_ASAP7_75t_L g264 ( .A(n_197), .Y(n_264) );
BUFx2_ASAP7_75t_L g287 ( .A(n_197), .Y(n_287) );
AND2x2_ASAP7_75t_L g444 ( .A(n_197), .B(n_298), .Y(n_444) );
OR2x6_ASAP7_75t_L g197 ( .A(n_198), .B(n_208), .Y(n_197) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g276 ( .A(n_207), .Y(n_276) );
INVx1_ASAP7_75t_L g520 ( .A(n_207), .Y(n_520) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp33_ASAP7_75t_L g211 ( .A(n_212), .B(n_249), .Y(n_211) );
OAI221xp5_ASAP7_75t_L g344 ( .A1(n_212), .A2(n_345), .B1(n_352), .B2(n_353), .C(n_356), .Y(n_344) );
OR2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_226), .Y(n_212) );
AND2x2_ASAP7_75t_L g250 ( .A(n_213), .B(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_213), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g279 ( .A(n_214), .B(n_227), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_214), .B(n_228), .Y(n_289) );
OR2x2_ASAP7_75t_L g300 ( .A(n_214), .B(n_251), .Y(n_300) );
AND2x2_ASAP7_75t_L g303 ( .A(n_214), .B(n_291), .Y(n_303) );
AND2x2_ASAP7_75t_L g319 ( .A(n_214), .B(n_240), .Y(n_319) );
OR2x2_ASAP7_75t_L g335 ( .A(n_214), .B(n_228), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_214), .B(n_251), .Y(n_397) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_215), .B(n_240), .Y(n_389) );
AND2x2_ASAP7_75t_L g392 ( .A(n_215), .B(n_228), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_222), .B(n_223), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_223), .A2(n_234), .B(n_235), .Y(n_233) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
OR2x2_ASAP7_75t_L g313 ( .A(n_226), .B(n_300), .Y(n_313) );
INVx2_ASAP7_75t_L g339 ( .A(n_226), .Y(n_339) );
OR2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_240), .Y(n_226) );
AND2x2_ASAP7_75t_L g261 ( .A(n_227), .B(n_241), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_227), .B(n_251), .Y(n_318) );
OR2x2_ASAP7_75t_L g329 ( .A(n_227), .B(n_241), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_227), .B(n_291), .Y(n_388) );
OAI221xp5_ASAP7_75t_L g421 ( .A1(n_227), .A2(n_422), .B1(n_424), .B2(n_426), .C(n_429), .Y(n_421) );
INVx5_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_228), .B(n_251), .Y(n_360) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_232), .Y(n_229) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_231), .A2(n_530), .B(n_531), .Y(n_529) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_231), .A2(n_547), .B(n_548), .Y(n_546) );
INVx4_ASAP7_75t_L g275 ( .A(n_236), .Y(n_275) );
INVx2_ASAP7_75t_L g498 ( .A(n_236), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx2_ASAP7_75t_L g481 ( .A(n_239), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_240), .B(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_240), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g307 ( .A(n_240), .B(n_279), .Y(n_307) );
OR2x2_ASAP7_75t_L g351 ( .A(n_240), .B(n_251), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_240), .B(n_303), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_240), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g416 ( .A(n_240), .B(n_417), .Y(n_416) );
INVx5_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_SL g280 ( .A(n_241), .B(n_250), .Y(n_280) );
O2A1O1Ixp33_ASAP7_75t_SL g284 ( .A1(n_241), .A2(n_285), .B(n_288), .C(n_292), .Y(n_284) );
OR2x2_ASAP7_75t_L g322 ( .A(n_241), .B(n_318), .Y(n_322) );
OR2x2_ASAP7_75t_L g358 ( .A(n_241), .B(n_300), .Y(n_358) );
OAI311xp33_ASAP7_75t_L g364 ( .A1(n_241), .A2(n_303), .A3(n_365), .B1(n_368), .C1(n_375), .Y(n_364) );
AND2x2_ASAP7_75t_L g415 ( .A(n_241), .B(n_251), .Y(n_415) );
AND2x2_ASAP7_75t_L g423 ( .A(n_241), .B(n_278), .Y(n_423) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_241), .Y(n_441) );
AND2x2_ASAP7_75t_L g458 ( .A(n_241), .B(n_279), .Y(n_458) );
OR2x6_ASAP7_75t_L g241 ( .A(n_242), .B(n_248), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_261), .Y(n_249) );
AND2x2_ASAP7_75t_L g286 ( .A(n_250), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g442 ( .A(n_250), .Y(n_442) );
AND2x2_ASAP7_75t_L g278 ( .A(n_251), .B(n_279), .Y(n_278) );
INVx3_ASAP7_75t_L g291 ( .A(n_251), .Y(n_291) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_251), .Y(n_334) );
INVxp67_ASAP7_75t_L g373 ( .A(n_251), .Y(n_373) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_253), .B(n_259), .Y(n_251) );
OA21x2_ASAP7_75t_L g503 ( .A1(n_252), .A2(n_504), .B(n_510), .Y(n_503) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_252), .A2(n_514), .B(n_521), .Y(n_513) );
OA21x2_ASAP7_75t_L g554 ( .A1(n_252), .A2(n_555), .B(n_562), .Y(n_554) );
OA21x2_ASAP7_75t_L g267 ( .A1(n_260), .A2(n_268), .B(n_277), .Y(n_267) );
AND2x2_ASAP7_75t_L g451 ( .A(n_261), .B(n_299), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_278), .B1(n_280), .B2(n_281), .C(n_284), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_264), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g304 ( .A(n_264), .B(n_294), .Y(n_304) );
AND2x2_ASAP7_75t_L g312 ( .A(n_264), .B(n_266), .Y(n_312) );
OR2x2_ASAP7_75t_L g324 ( .A(n_264), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g342 ( .A(n_264), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g366 ( .A(n_264), .B(n_367), .Y(n_366) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_264), .Y(n_386) );
AND2x2_ASAP7_75t_L g438 ( .A(n_264), .B(n_362), .Y(n_438) );
OAI31xp33_ASAP7_75t_L g446 ( .A1(n_264), .A2(n_315), .A3(n_414), .B(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_265), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_SL g410 ( .A(n_265), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_265), .B(n_419), .Y(n_418) );
AND2x4_ASAP7_75t_L g298 ( .A(n_266), .B(n_294), .Y(n_298) );
INVx1_ASAP7_75t_L g385 ( .A(n_266), .Y(n_385) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g435 ( .A(n_267), .B(n_294), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_275), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g535 ( .A(n_276), .Y(n_535) );
INVx1_ASAP7_75t_SL g445 ( .A(n_278), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_279), .B(n_350), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_280), .A2(n_392), .B1(n_430), .B2(n_433), .Y(n_429) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g293 ( .A(n_283), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g352 ( .A(n_283), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_283), .B(n_304), .Y(n_457) );
INVx1_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g427 ( .A(n_286), .B(n_428), .Y(n_427) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_287), .A2(n_346), .B(n_348), .Y(n_345) );
OR2x2_ASAP7_75t_L g353 ( .A(n_287), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g374 ( .A(n_287), .B(n_362), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_287), .B(n_385), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_287), .B(n_425), .Y(n_424) );
OAI221xp5_ASAP7_75t_SL g401 ( .A1(n_288), .A2(n_402), .B1(n_407), .B2(n_410), .C(n_411), .Y(n_401) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
OR2x2_ASAP7_75t_L g378 ( .A(n_289), .B(n_351), .Y(n_378) );
INVx1_ASAP7_75t_L g417 ( .A(n_289), .Y(n_417) );
INVx2_ASAP7_75t_L g393 ( .A(n_290), .Y(n_393) );
INVx1_ASAP7_75t_L g327 ( .A(n_291), .Y(n_327) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g332 ( .A(n_294), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_294), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g361 ( .A(n_294), .B(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g449 ( .A(n_294), .B(n_419), .Y(n_449) );
AOI222xp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_299), .B1(n_301), .B2(n_304), .C1(n_305), .C2(n_307), .Y(n_295) );
INVxp67_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g305 ( .A(n_298), .B(n_306), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_298), .A2(n_348), .B1(n_376), .B2(n_377), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_298), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OAI21xp33_ASAP7_75t_SL g336 ( .A1(n_307), .A2(n_337), .B(n_340), .Y(n_336) );
OAI211xp5_ASAP7_75t_SL g308 ( .A1(n_309), .A2(n_313), .B(n_314), .C(n_336), .Y(n_308) );
INVxp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
AOI221xp5_ASAP7_75t_L g314 ( .A1(n_312), .A2(n_315), .B1(n_320), .B2(n_321), .C(n_323), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_312), .B(n_400), .Y(n_399) );
INVxp67_ASAP7_75t_L g406 ( .A(n_312), .Y(n_406) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
AND2x2_ASAP7_75t_L g408 ( .A(n_317), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g325 ( .A(n_320), .Y(n_325) );
AND2x2_ASAP7_75t_L g331 ( .A(n_320), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_326), .B1(n_330), .B2(n_333), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_327), .B(n_339), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_328), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g428 ( .A(n_332), .Y(n_428) );
AND2x2_ASAP7_75t_L g447 ( .A(n_332), .B(n_362), .Y(n_447) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_339), .B(n_396), .Y(n_455) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_342), .B(n_410), .Y(n_453) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g376 ( .A(n_354), .Y(n_376) );
BUFx2_ASAP7_75t_L g400 ( .A(n_355), .Y(n_400) );
OAI21xp5_ASAP7_75t_SL g356 ( .A1(n_357), .A2(n_359), .B(n_361), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NOR3xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_379), .C(n_401), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI21xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_371), .B(n_374), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
A2O1A1Ixp33_ASAP7_75t_SL g379 ( .A1(n_380), .A2(n_383), .B(n_387), .C(n_390), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_380), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp67_ASAP7_75t_SL g384 ( .A(n_385), .B(n_386), .Y(n_384) );
OR2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_SL g409 ( .A(n_389), .Y(n_409) );
OAI21xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_394), .B(n_398), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
AND2x2_ASAP7_75t_L g414 ( .A(n_392), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_414), .B1(n_416), .B2(n_418), .Y(n_411) );
INVx2_ASAP7_75t_SL g432 ( .A(n_419), .Y(n_432) );
NOR3xp33_ASAP7_75t_L g420 ( .A(n_421), .B(n_436), .C(n_448), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_432), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI221xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_439), .B1(n_443), .B2(n_445), .C(n_446), .Y(n_436) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_437), .A2(n_449), .B(n_450), .C(n_452), .Y(n_448) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVxp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B1(n_456), .B2(n_458), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g740 ( .A(n_460), .Y(n_740) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_SL g742 ( .A(n_462), .Y(n_742) );
OR5x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_629), .C(n_693), .D(n_709), .E(n_724), .Y(n_462) );
NAND4xp25_ASAP7_75t_L g463 ( .A(n_464), .B(n_563), .C(n_590), .D(n_613), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_511), .B(n_522), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_476), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx3_ASAP7_75t_SL g542 ( .A(n_467), .Y(n_542) );
AND2x4_ASAP7_75t_L g576 ( .A(n_467), .B(n_565), .Y(n_576) );
OR2x2_ASAP7_75t_L g586 ( .A(n_467), .B(n_544), .Y(n_586) );
OR2x2_ASAP7_75t_L g632 ( .A(n_467), .B(n_479), .Y(n_632) );
AND2x2_ASAP7_75t_L g646 ( .A(n_467), .B(n_543), .Y(n_646) );
AND2x2_ASAP7_75t_L g689 ( .A(n_467), .B(n_579), .Y(n_689) );
AND2x2_ASAP7_75t_L g696 ( .A(n_467), .B(n_554), .Y(n_696) );
AND2x2_ASAP7_75t_L g715 ( .A(n_467), .B(n_605), .Y(n_715) );
AND2x2_ASAP7_75t_L g733 ( .A(n_467), .B(n_575), .Y(n_733) );
OR2x6_ASAP7_75t_L g467 ( .A(n_468), .B(n_474), .Y(n_467) );
INVx1_ASAP7_75t_L g698 ( .A(n_476), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_492), .Y(n_476) );
AND2x2_ASAP7_75t_L g608 ( .A(n_477), .B(n_543), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_477), .B(n_628), .Y(n_627) );
AOI32xp33_ASAP7_75t_L g641 ( .A1(n_477), .A2(n_642), .A3(n_645), .B1(n_647), .B2(n_651), .Y(n_641) );
AND2x2_ASAP7_75t_L g711 ( .A(n_477), .B(n_605), .Y(n_711) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g575 ( .A(n_479), .B(n_544), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_479), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g617 ( .A(n_479), .B(n_564), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_479), .B(n_696), .Y(n_695) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_482), .B(n_490), .Y(n_479) );
INVx1_ASAP7_75t_L g580 ( .A(n_480), .Y(n_580) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OA21x2_ASAP7_75t_L g579 ( .A1(n_483), .A2(n_491), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g582 ( .A(n_492), .B(n_526), .Y(n_582) );
AND2x2_ASAP7_75t_L g658 ( .A(n_492), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g730 ( .A(n_492), .Y(n_730) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_502), .Y(n_492) );
OR2x2_ASAP7_75t_L g525 ( .A(n_493), .B(n_503), .Y(n_525) );
AND2x2_ASAP7_75t_L g539 ( .A(n_493), .B(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_493), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g589 ( .A(n_493), .Y(n_589) );
AND2x2_ASAP7_75t_L g616 ( .A(n_493), .B(n_503), .Y(n_616) );
BUFx3_ASAP7_75t_L g619 ( .A(n_493), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_493), .B(n_594), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_493), .B(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g570 ( .A(n_502), .Y(n_570) );
AND2x2_ASAP7_75t_L g588 ( .A(n_502), .B(n_568), .Y(n_588) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g599 ( .A(n_503), .B(n_513), .Y(n_599) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_503), .Y(n_612) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_512), .B(n_619), .Y(n_669) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_SL g540 ( .A(n_513), .Y(n_540) );
NAND3xp33_ASAP7_75t_L g587 ( .A(n_513), .B(n_588), .C(n_589), .Y(n_587) );
OR2x2_ASAP7_75t_L g595 ( .A(n_513), .B(n_568), .Y(n_595) );
AND2x2_ASAP7_75t_L g615 ( .A(n_513), .B(n_568), .Y(n_615) );
AND2x2_ASAP7_75t_L g659 ( .A(n_513), .B(n_528), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_538), .B(n_541), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_524), .B(n_526), .Y(n_523) );
AND2x2_ASAP7_75t_L g734 ( .A(n_524), .B(n_659), .Y(n_734) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_525), .A2(n_632), .B1(n_674), .B2(n_676), .Y(n_673) );
OR2x2_ASAP7_75t_L g680 ( .A(n_525), .B(n_595), .Y(n_680) );
OR2x2_ASAP7_75t_L g704 ( .A(n_525), .B(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_525), .B(n_624), .Y(n_717) );
AND2x2_ASAP7_75t_L g610 ( .A(n_526), .B(n_611), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_526), .A2(n_683), .B(n_698), .Y(n_697) );
AOI32xp33_ASAP7_75t_L g718 ( .A1(n_526), .A2(n_608), .A3(n_719), .B1(n_721), .B2(n_722), .Y(n_718) );
OR2x2_ASAP7_75t_L g729 ( .A(n_526), .B(n_730), .Y(n_729) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g597 ( .A(n_527), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_527), .B(n_611), .Y(n_676) );
BUFx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx4_ASAP7_75t_L g568 ( .A(n_528), .Y(n_568) );
AND2x2_ASAP7_75t_L g634 ( .A(n_528), .B(n_599), .Y(n_634) );
AND3x2_ASAP7_75t_L g643 ( .A(n_528), .B(n_539), .C(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g569 ( .A(n_540), .B(n_570), .Y(n_569) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_540), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_540), .B(n_568), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
AND2x2_ASAP7_75t_L g564 ( .A(n_542), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g604 ( .A(n_542), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g622 ( .A(n_542), .B(n_554), .Y(n_622) );
AND2x2_ASAP7_75t_L g640 ( .A(n_542), .B(n_544), .Y(n_640) );
OR2x2_ASAP7_75t_L g654 ( .A(n_542), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g700 ( .A(n_542), .B(n_628), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_543), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_554), .Y(n_543) );
AND2x2_ASAP7_75t_L g601 ( .A(n_544), .B(n_579), .Y(n_601) );
OR2x2_ASAP7_75t_L g655 ( .A(n_544), .B(n_579), .Y(n_655) );
AND2x2_ASAP7_75t_L g708 ( .A(n_544), .B(n_565), .Y(n_708) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
BUFx2_ASAP7_75t_L g606 ( .A(n_545), .Y(n_606) );
AND2x2_ASAP7_75t_L g628 ( .A(n_545), .B(n_554), .Y(n_628) );
INVx2_ASAP7_75t_L g565 ( .A(n_554), .Y(n_565) );
INVx1_ASAP7_75t_L g585 ( .A(n_554), .Y(n_585) );
AOI211xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_566), .B(n_571), .C(n_583), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_564), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g727 ( .A(n_564), .Y(n_727) );
AND2x2_ASAP7_75t_L g605 ( .A(n_565), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_568), .B(n_569), .Y(n_577) );
INVx1_ASAP7_75t_L g662 ( .A(n_568), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_568), .B(n_589), .Y(n_686) );
AND2x2_ASAP7_75t_L g702 ( .A(n_568), .B(n_616), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_569), .B(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g593 ( .A(n_570), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_577), .B1(n_578), .B2(n_581), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_574), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_575), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g600 ( .A(n_576), .B(n_601), .Y(n_600) );
AOI221xp5_ASAP7_75t_SL g665 ( .A1(n_576), .A2(n_618), .B1(n_666), .B2(n_671), .C(n_673), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_576), .B(n_639), .Y(n_672) );
INVx1_ASAP7_75t_L g732 ( .A(n_578), .Y(n_732) );
BUFx3_ASAP7_75t_L g639 ( .A(n_579), .Y(n_639) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AOI21xp33_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_586), .B(n_587), .Y(n_583) );
INVx1_ASAP7_75t_L g648 ( .A(n_585), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_585), .B(n_639), .Y(n_692) );
INVx1_ASAP7_75t_L g649 ( .A(n_586), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_586), .B(n_639), .Y(n_650) );
INVxp67_ASAP7_75t_L g670 ( .A(n_588), .Y(n_670) );
AND2x2_ASAP7_75t_L g611 ( .A(n_589), .B(n_612), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_596), .B(n_600), .C(n_602), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_SL g625 ( .A(n_593), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_594), .B(n_625), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_594), .B(n_616), .Y(n_667) );
INVx2_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_597), .A2(n_603), .B1(n_607), .B2(n_609), .Y(n_602) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g618 ( .A(n_599), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g663 ( .A(n_599), .B(n_664), .Y(n_663) );
OAI21xp33_ASAP7_75t_L g666 ( .A1(n_601), .A2(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_605), .A2(n_614), .B1(n_617), .B2(n_618), .C(n_620), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_605), .B(n_639), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_605), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g721 ( .A(n_611), .Y(n_721) );
INVxp67_ASAP7_75t_L g644 ( .A(n_612), .Y(n_644) );
INVx1_ASAP7_75t_L g651 ( .A(n_614), .Y(n_651) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
AND2x2_ASAP7_75t_L g690 ( .A(n_615), .B(n_619), .Y(n_690) );
INVx1_ASAP7_75t_L g664 ( .A(n_619), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_619), .B(n_634), .Y(n_694) );
OAI32xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_623), .A3(n_625), .B1(n_626), .B2(n_627), .Y(n_620) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_SL g633 ( .A(n_628), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_628), .B(n_660), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_628), .B(n_689), .Y(n_720) );
NAND2x1p5_ASAP7_75t_L g728 ( .A(n_628), .B(n_639), .Y(n_728) );
NAND5xp2_ASAP7_75t_L g629 ( .A(n_630), .B(n_652), .C(n_665), .D(n_677), .E(n_678), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_634), .B1(n_635), .B2(n_637), .C(n_641), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND2xp33_ASAP7_75t_SL g656 ( .A(n_636), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_639), .B(n_708), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_640), .A2(n_653), .B1(n_656), .B2(n_660), .Y(n_652) );
INVx2_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
OAI211xp5_ASAP7_75t_SL g647 ( .A1(n_643), .A2(n_648), .B(n_649), .C(n_650), .Y(n_647) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g675 ( .A(n_655), .Y(n_675) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_664), .B(n_713), .Y(n_723) );
OR2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI222xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_681), .B1(n_683), .B2(n_687), .C1(n_690), .C2(n_691), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B1(n_697), .B2(n_699), .C(n_701), .Y(n_693) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
OAI21xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B(n_706), .Y(n_701) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g713 ( .A(n_705), .Y(n_713) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_712), .B1(n_714), .B2(n_716), .C(n_718), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_728), .B(n_729), .C(n_731), .Y(n_724) );
INVxp67_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OAI21xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B(n_734), .Y(n_731) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_737), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
endmodule