module fake_jpeg_30328_n_68 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_68);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_68;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_18),
.C(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_27),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_30),
.Y(n_34)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_21),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_22),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_31),
.B1(n_25),
.B2(n_22),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_4),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_25),
.B1(n_2),
.B2(n_3),
.Y(n_37)
);

NOR2x1_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_1),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_24),
.B(n_6),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_48),
.B(n_5),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_45)
);

AO22x1_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_49),
.B1(n_43),
.B2(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_47),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_24),
.C(n_5),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_15),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_34),
.C(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_55),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_57),
.B(n_7),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_39),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_56),
.Y(n_60)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_58),
.B(n_14),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_51),
.B(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_63),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_59),
.C(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_50),
.Y(n_66)
);

MAJx2_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_53),
.C(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_53),
.Y(n_68)
);


endmodule