module fake_jpeg_29353_n_118 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_118);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_2),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_30),
.Y(n_47)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_38),
.Y(n_54)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_0),
.C(n_1),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_16),
.C(n_21),
.Y(n_59)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_1),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_12),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_32),
.B(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_12),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_29),
.B(n_17),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_57),
.A2(n_21),
.B1(n_35),
.B2(n_33),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_39),
.B1(n_41),
.B2(n_40),
.Y(n_60)
);

NAND2x1_ASAP7_75t_SL g81 ( 
.A(n_60),
.B(n_56),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_66),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_58),
.A2(n_49),
.B1(n_43),
.B2(n_57),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_52),
.B(n_54),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_68),
.Y(n_78)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_70),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_74),
.Y(n_86)
);

AOI32xp33_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_71),
.B(n_47),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_82),
.Y(n_89)
);

AO21x1_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_81),
.B(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_59),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_54),
.C(n_45),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_87),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_56),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_45),
.B(n_60),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_95),
.B(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_92),
.Y(n_98)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_66),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_94),
.B(n_86),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_67),
.B(n_61),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_76),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_96),
.B(n_99),
.Y(n_105)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_102),
.Y(n_106)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_104),
.B(n_107),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_91),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_105),
.B(n_6),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_110),
.B(n_106),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_106),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_SL g114 ( 
.A1(n_111),
.A2(n_100),
.B(n_68),
.C(n_70),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_100),
.C(n_84),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_93),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_114),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_84),
.B(n_43),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_70),
.C(n_56),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_73),
.Y(n_118)
);


endmodule