module fake_jpeg_8213_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_16),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_42),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_48),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx5_ASAP7_75t_SL g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_53),
.B(n_56),
.Y(n_84)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_34),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_25),
.Y(n_72)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_21),
.B1(n_29),
.B2(n_32),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_21),
.B1(n_29),
.B2(n_36),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_67),
.B(n_68),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_69),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_72),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_21),
.B1(n_29),
.B2(n_25),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_76),
.B(n_20),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_25),
.B1(n_30),
.B2(n_28),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_77),
.Y(n_106)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_42),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_81),
.Y(n_104)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_36),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_89),
.Y(n_107)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_49),
.A2(n_30),
.B1(n_24),
.B2(n_17),
.Y(n_94)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

NAND2x1_ASAP7_75t_SL g95 ( 
.A(n_58),
.B(n_46),
.Y(n_95)
);

MAJx3_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_45),
.C(n_61),
.Y(n_121)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_98),
.Y(n_108)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_71),
.B(n_18),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_101),
.B(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_125),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_58),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_115),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_79),
.B(n_18),
.Y(n_110)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_47),
.C(n_55),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_113),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_46),
.C(n_38),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_59),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_59),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_95),
.B(n_91),
.Y(n_138)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_126),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_97),
.B1(n_90),
.B2(n_96),
.Y(n_140)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_69),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_30),
.Y(n_127)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_129),
.B(n_134),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_72),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_141),
.Y(n_164)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_135),
.B(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_78),
.B1(n_82),
.B2(n_90),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_152),
.B1(n_123),
.B2(n_116),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_139),
.B(n_150),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_97),
.B(n_83),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_98),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_89),
.B1(n_87),
.B2(n_74),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_143),
.A2(n_145),
.B1(n_155),
.B2(n_140),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_106),
.A2(n_85),
.B1(n_63),
.B2(n_88),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_120),
.B1(n_122),
.B2(n_118),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_63),
.B1(n_92),
.B2(n_31),
.Y(n_145)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_149),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_109),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_103),
.A2(n_28),
.B1(n_23),
.B2(n_24),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_35),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_106),
.A2(n_22),
.B1(n_31),
.B2(n_36),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_156),
.A2(n_22),
.B(n_31),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_117),
.C(n_115),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_165),
.C(n_186),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_134),
.B(n_110),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_159),
.B(n_185),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_160),
.A2(n_163),
.B1(n_176),
.B2(n_35),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_154),
.A2(n_125),
.B1(n_99),
.B2(n_124),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_111),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_131),
.B1(n_155),
.B2(n_151),
.Y(n_196)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_179),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_99),
.B1(n_105),
.B2(n_116),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_171),
.A2(n_178),
.B1(n_20),
.B2(n_1),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_172),
.A2(n_114),
.B1(n_129),
.B2(n_136),
.Y(n_191)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_177),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_175),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_145),
.A2(n_149),
.B1(n_142),
.B2(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_99),
.B1(n_120),
.B2(n_118),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_139),
.A2(n_22),
.B(n_33),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_180),
.A2(n_182),
.B(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_181),
.A2(n_187),
.B1(n_0),
.B2(n_1),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_128),
.A2(n_33),
.B(n_23),
.Y(n_182)
);

OA21x2_ASAP7_75t_L g183 ( 
.A1(n_135),
.A2(n_33),
.B(n_122),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_184),
.B(n_152),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_128),
.A2(n_45),
.B(n_93),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_150),
.B(n_17),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_132),
.B(n_114),
.C(n_24),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_197),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_191),
.A2(n_202),
.B1(n_216),
.B2(n_183),
.Y(n_237)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_194),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_162),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_131),
.C(n_130),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_205),
.C(n_213),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_196),
.Y(n_242)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_199),
.Y(n_230)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_200),
.A2(n_203),
.B(n_204),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_130),
.B1(n_28),
.B2(n_27),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_183),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_35),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_206),
.A2(n_208),
.B1(n_167),
.B2(n_182),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_0),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_207),
.A2(n_210),
.B(n_214),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_163),
.A2(n_27),
.B1(n_23),
.B2(n_17),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_209),
.A2(n_215),
.B(n_217),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_161),
.A2(n_27),
.B(n_35),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_211),
.A2(n_203),
.B1(n_190),
.B2(n_160),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_157),
.B(n_16),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_161),
.A2(n_168),
.B(n_180),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

OA21x2_ASAP7_75t_L g217 ( 
.A1(n_187),
.A2(n_0),
.B(n_1),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_218),
.B(n_222),
.Y(n_262)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_237),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_189),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_168),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_233),
.C(n_240),
.Y(n_248)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_212),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_231),
.B(n_235),
.Y(n_263)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_173),
.C(n_186),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_192),
.B(n_159),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_236),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_215),
.A2(n_173),
.B1(n_177),
.B2(n_172),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_239),
.A2(n_200),
.B1(n_208),
.B2(n_199),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_169),
.C(n_175),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_214),
.B(n_185),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_188),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_217),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_1),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_207),
.Y(n_244)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_246),
.A2(n_254),
.B1(n_235),
.B2(n_243),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_220),
.A2(n_204),
.B1(n_211),
.B2(n_194),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_249),
.A2(n_256),
.B1(n_228),
.B2(n_239),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_251),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_205),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_253),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_228),
.A2(n_217),
.B1(n_169),
.B2(n_207),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_232),
.A2(n_179),
.B1(n_170),
.B2(n_210),
.Y(n_256)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_259),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_213),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_SL g268 ( 
.A(n_261),
.B(n_227),
.C(n_240),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_2),
.C(n_3),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_259),
.C(n_266),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_221),
.B(n_2),
.Y(n_266)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_266),
.Y(n_277)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_267),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_261),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_260),
.A2(n_230),
.B1(n_242),
.B2(n_241),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_272),
.A2(n_276),
.B1(n_282),
.B2(n_284),
.Y(n_288)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_226),
.C(n_219),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_280),
.C(n_281),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_246),
.A2(n_219),
.B1(n_229),
.B2(n_225),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_278),
.A2(n_283),
.B1(n_257),
.B2(n_255),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_258),
.A2(n_229),
.B1(n_238),
.B2(n_9),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_279),
.B(n_247),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_238),
.C(n_3),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_8),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_254),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_257),
.A2(n_8),
.B(n_15),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_245),
.A2(n_16),
.B1(n_13),
.B2(n_12),
.Y(n_284)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_256),
.Y(n_286)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_271),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_251),
.Y(n_289)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_245),
.Y(n_290)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_290),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_249),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_292),
.B(n_296),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_253),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_271),
.C(n_272),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_258),
.C(n_265),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_290),
.C(n_291),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_263),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_299),
.B(n_288),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_284),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_312),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_307),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_305),
.C(n_311),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_276),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_293),
.A2(n_267),
.B(n_283),
.Y(n_309)
);

OAI22x1_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_281),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_304),
.A2(n_291),
.B(n_298),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_314),
.B(n_322),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_297),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_303),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_250),
.B1(n_295),
.B2(n_264),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_317),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_309),
.A2(n_11),
.B(n_8),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_318),
.A2(n_4),
.B(n_5),
.Y(n_327)
);

A2O1A1Ixp33_ASAP7_75t_SL g328 ( 
.A1(n_319),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_2),
.C(n_3),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_319),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_302),
.A2(n_11),
.B1(n_5),
.B2(n_6),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_325),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_313),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_326),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_328),
.A2(n_318),
.B(n_7),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_329),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_320),
.C(n_313),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_335),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_315),
.C(n_321),
.Y(n_337)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_337),
.Y(n_338)
);

NAND3xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_331),
.C(n_323),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_330),
.B(n_328),
.Y(n_340)
);


endmodule