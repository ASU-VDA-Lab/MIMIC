module real_aes_11766_n_267 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_267);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_267;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_602;
wire n_733;
wire n_402;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1482;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_578;
wire n_372;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_559;
wire n_466;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_269;
wire n_430;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
CKINVDCx5p33_ASAP7_75t_R g910 ( .A(n_0), .Y(n_910) );
XNOR2xp5_ASAP7_75t_L g720 ( .A(n_1), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g1264 ( .A(n_2), .Y(n_1264) );
CKINVDCx5p33_ASAP7_75t_R g737 ( .A(n_3), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_4), .A2(n_82), .B1(n_1000), .B2(n_1003), .Y(n_1174) );
INVx1_ASAP7_75t_L g1205 ( .A(n_4), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_5), .A2(n_257), .B1(n_876), .B2(n_877), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_5), .A2(n_257), .B1(n_885), .B2(n_886), .Y(n_884) );
AO22x2_ASAP7_75t_L g660 ( .A1(n_6), .A2(n_661), .B1(n_715), .B2(n_716), .Y(n_660) );
INVxp67_ASAP7_75t_L g715 ( .A(n_6), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_7), .A2(n_229), .B1(n_301), .B2(n_309), .Y(n_300) );
INVx1_ASAP7_75t_L g423 ( .A(n_7), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_8), .A2(n_239), .B1(n_705), .B2(n_1005), .Y(n_1036) );
INVx1_ASAP7_75t_L g1044 ( .A(n_8), .Y(n_1044) );
CKINVDCx5p33_ASAP7_75t_R g927 ( .A(n_9), .Y(n_927) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_10), .Y(n_280) );
INVx1_ASAP7_75t_L g467 ( .A(n_10), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_10), .B(n_208), .Y(n_509) );
AND2x2_ASAP7_75t_L g513 ( .A(n_10), .B(n_305), .Y(n_513) );
INVx1_ASAP7_75t_L g1245 ( .A(n_11), .Y(n_1245) );
CKINVDCx5p33_ASAP7_75t_R g852 ( .A(n_12), .Y(n_852) );
OAI22xp33_ASAP7_75t_L g750 ( .A1(n_13), .A2(n_196), .B1(n_551), .B2(n_560), .Y(n_750) );
INVx1_ASAP7_75t_L g777 ( .A(n_13), .Y(n_777) );
INVx1_ASAP7_75t_L g610 ( .A(n_14), .Y(n_610) );
OAI22xp33_ASAP7_75t_L g645 ( .A1(n_14), .A2(n_154), .B1(n_646), .B2(n_649), .Y(n_645) );
INVx1_ASAP7_75t_L g807 ( .A(n_15), .Y(n_807) );
OAI221xp5_ASAP7_75t_L g819 ( .A1(n_15), .A2(n_522), .B1(n_767), .B2(n_820), .C(n_823), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_16), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g926 ( .A(n_17), .Y(n_926) );
INVx1_ASAP7_75t_L g1017 ( .A(n_18), .Y(n_1017) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_18), .A2(n_89), .B1(n_965), .B2(n_1042), .Y(n_1041) );
INVx1_ASAP7_75t_L g1310 ( .A(n_19), .Y(n_1310) );
CKINVDCx16_ASAP7_75t_R g1324 ( .A(n_20), .Y(n_1324) );
XNOR2x2_ASAP7_75t_L g470 ( .A(n_21), .B(n_471), .Y(n_470) );
AOI21xp33_ASAP7_75t_L g494 ( .A1(n_22), .A2(n_495), .B(n_496), .Y(n_494) );
INVx1_ASAP7_75t_L g574 ( .A(n_22), .Y(n_574) );
INVxp67_ASAP7_75t_SL g595 ( .A(n_23), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_23), .A2(n_247), .B1(n_630), .B2(n_640), .Y(n_639) );
AOI221xp5_ASAP7_75t_L g774 ( .A1(n_24), .A2(n_228), .B1(n_495), .B2(n_496), .C(n_775), .Y(n_774) );
OAI22xp33_ASAP7_75t_L g788 ( .A1(n_24), .A2(n_102), .B1(n_789), .B2(n_791), .Y(n_788) );
INVx1_ASAP7_75t_L g829 ( .A(n_25), .Y(n_829) );
OAI22xp33_ASAP7_75t_L g838 ( .A1(n_25), .A2(n_34), .B1(n_789), .B2(n_791), .Y(n_838) );
INVx1_ASAP7_75t_L g968 ( .A(n_26), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_26), .A2(n_206), .B1(n_1005), .B2(n_1006), .Y(n_1004) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_27), .A2(n_54), .B1(n_354), .B2(n_362), .Y(n_353) );
INVx1_ASAP7_75t_L g455 ( .A(n_27), .Y(n_455) );
AO22x2_ASAP7_75t_L g1107 ( .A1(n_28), .A2(n_1108), .B1(n_1109), .B2(n_1159), .Y(n_1107) );
INVxp67_ASAP7_75t_SL g1108 ( .A(n_28), .Y(n_1108) );
INVx2_ASAP7_75t_L g348 ( .A(n_29), .Y(n_348) );
OR2x2_ASAP7_75t_L g573 ( .A(n_29), .B(n_558), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_30), .A2(n_173), .B1(n_511), .B2(n_517), .Y(n_510) );
INVx1_ASAP7_75t_L g549 ( .A(n_30), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_31), .Y(n_498) );
AOI22xp33_ASAP7_75t_SL g622 ( .A1(n_32), .A2(n_95), .B1(n_619), .B2(n_623), .Y(n_622) );
INVxp33_ASAP7_75t_L g656 ( .A(n_32), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_33), .A2(n_152), .B1(n_581), .B2(n_584), .Y(n_1065) );
INVx1_ASAP7_75t_L g1088 ( .A(n_33), .Y(n_1088) );
AOI221xp5_ASAP7_75t_L g832 ( .A1(n_34), .A2(n_144), .B1(n_495), .B2(n_496), .C(n_606), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_35), .A2(n_118), .B1(n_977), .B2(n_978), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_35), .A2(n_118), .B1(n_998), .B2(n_1031), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1176 ( .A1(n_36), .A2(n_225), .B1(n_1005), .B2(n_1006), .Y(n_1176) );
OAI22xp5_ASAP7_75t_L g1212 ( .A1(n_36), .A2(n_225), .B1(n_517), .B2(n_1092), .Y(n_1212) );
BUFx2_ASAP7_75t_L g296 ( .A(n_37), .Y(n_296) );
BUFx2_ASAP7_75t_L g394 ( .A(n_37), .Y(n_394) );
INVx1_ASAP7_75t_L g465 ( .A(n_37), .Y(n_465) );
INVx1_ASAP7_75t_L g1257 ( .A(n_38), .Y(n_1257) );
INVx1_ASAP7_75t_L g1308 ( .A(n_39), .Y(n_1308) );
INVx1_ASAP7_75t_L g603 ( .A(n_40), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_40), .A2(n_74), .B1(n_636), .B2(n_637), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g670 ( .A1(n_41), .A2(n_236), .B1(n_649), .B2(n_671), .C(n_672), .Y(n_670) );
INVx1_ASAP7_75t_L g682 ( .A(n_41), .Y(n_682) );
INVx1_ASAP7_75t_L g745 ( .A(n_42), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_42), .A2(n_87), .B1(n_511), .B2(n_517), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_43), .A2(n_120), .B1(n_633), .B2(n_902), .Y(n_901) );
AOI221xp5_ASAP7_75t_L g921 ( .A1(n_43), .A2(n_120), .B1(n_433), .B2(n_499), .C(n_775), .Y(n_921) );
AOI221xp5_ASAP7_75t_L g1485 ( .A1(n_44), .A2(n_69), .B1(n_433), .B2(n_604), .C(n_1486), .Y(n_1485) );
AOI22xp33_ASAP7_75t_L g1511 ( .A1(n_44), .A2(n_69), .B1(n_1000), .B2(n_1512), .Y(n_1511) );
OAI22xp33_ASAP7_75t_L g521 ( .A1(n_45), .A2(n_52), .B1(n_522), .B2(n_524), .Y(n_521) );
AOI221xp5_ASAP7_75t_L g542 ( .A1(n_45), .A2(n_52), .B1(n_531), .B2(n_543), .C(n_545), .Y(n_542) );
OAI22xp33_ASAP7_75t_L g814 ( .A1(n_46), .A2(n_67), .B1(n_551), .B2(n_560), .Y(n_814) );
INVx1_ASAP7_75t_L g835 ( .A(n_46), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_47), .A2(n_81), .B1(n_1144), .B2(n_1147), .Y(n_1146) );
INVxp67_ASAP7_75t_SL g1152 ( .A(n_47), .Y(n_1152) );
CKINVDCx16_ASAP7_75t_R g1235 ( .A(n_48), .Y(n_1235) );
INVx1_ASAP7_75t_L g773 ( .A(n_49), .Y(n_773) );
OAI22xp33_ASAP7_75t_L g786 ( .A1(n_49), .A2(n_228), .B1(n_584), .B2(n_787), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g912 ( .A(n_50), .Y(n_912) );
XNOR2xp5_ASAP7_75t_L g1164 ( .A(n_51), .B(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g1304 ( .A(n_51), .Y(n_1304) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_53), .Y(n_477) );
INVx1_ASAP7_75t_L g333 ( .A(n_54), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_55), .A2(n_96), .B1(n_619), .B2(n_621), .Y(n_618) );
AOI22xp33_ASAP7_75t_SL g629 ( .A1(n_55), .A2(n_96), .B1(n_630), .B2(n_631), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_56), .A2(n_262), .B1(n_980), .B2(n_981), .Y(n_979) );
AOI22xp33_ASAP7_75t_SL g992 ( .A1(n_56), .A2(n_262), .B1(n_993), .B2(n_995), .Y(n_992) );
AOI22xp33_ASAP7_75t_SL g907 ( .A1(n_57), .A2(n_263), .B1(n_576), .B2(n_631), .Y(n_907) );
INVx1_ASAP7_75t_L g916 ( .A(n_57), .Y(n_916) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_58), .Y(n_402) );
INVx1_ASAP7_75t_L g1022 ( .A(n_59), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_59), .A2(n_248), .B1(n_983), .B2(n_986), .Y(n_1027) );
INVx1_ASAP7_75t_L g949 ( .A(n_60), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_60), .A2(n_161), .B1(n_983), .B2(n_986), .Y(n_982) );
AOI221xp5_ASAP7_75t_L g1476 ( .A1(n_61), .A2(n_219), .B1(n_978), .B2(n_1081), .C(n_1196), .Y(n_1476) );
INVx1_ASAP7_75t_L g1494 ( .A(n_61), .Y(n_1494) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_62), .A2(n_172), .B1(n_1092), .B2(n_1093), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_62), .A2(n_172), .B1(n_1104), .B2(n_1105), .Y(n_1103) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_63), .Y(n_480) );
INVx1_ASAP7_75t_L g1060 ( .A(n_64), .Y(n_1060) );
INVx1_ASAP7_75t_L g752 ( .A(n_65), .Y(n_752) );
INVx1_ASAP7_75t_L g810 ( .A(n_66), .Y(n_810) );
OAI211xp5_ASAP7_75t_L g827 ( .A1(n_66), .A2(n_524), .B(n_828), .C(n_833), .Y(n_827) );
INVx1_ASAP7_75t_L g834 ( .A(n_67), .Y(n_834) );
AO221x2_ASAP7_75t_L g1255 ( .A1(n_68), .A2(n_84), .B1(n_1232), .B2(n_1234), .C(n_1256), .Y(n_1255) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_70), .A2(n_107), .B1(n_616), .B2(n_625), .Y(n_624) );
INVxp67_ASAP7_75t_SL g644 ( .A(n_70), .Y(n_644) );
INVx1_ASAP7_75t_L g954 ( .A(n_71), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_71), .A2(n_136), .B1(n_604), .B2(n_988), .Y(n_987) );
AOI22xp33_ASAP7_75t_SL g1131 ( .A1(n_72), .A2(n_132), .B1(n_606), .B2(n_1132), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_72), .A2(n_132), .B1(n_1144), .B2(n_1145), .Y(n_1143) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_73), .Y(n_488) );
INVxp33_ASAP7_75t_L g598 ( .A(n_74), .Y(n_598) );
AO22x2_ASAP7_75t_L g1008 ( .A1(n_75), .A2(n_1009), .B1(n_1048), .B2(n_1049), .Y(n_1008) );
INVxp67_ASAP7_75t_SL g1048 ( .A(n_75), .Y(n_1048) );
INVx1_ASAP7_75t_L g1319 ( .A(n_76), .Y(n_1319) );
CKINVDCx16_ASAP7_75t_R g1322 ( .A(n_77), .Y(n_1322) );
AOI222xp33_ASAP7_75t_L g1467 ( .A1(n_77), .A2(n_1468), .B1(n_1519), .B2(n_1523), .C1(n_1528), .C2(n_1532), .Y(n_1467) );
AO221x1_ASAP7_75t_L g924 ( .A1(n_78), .A2(n_103), .B1(n_495), .B2(n_496), .C(n_626), .Y(n_924) );
INVx1_ASAP7_75t_L g935 ( .A(n_78), .Y(n_935) );
OAI221xp5_ASAP7_75t_L g1069 ( .A1(n_79), .A2(n_522), .B1(n_767), .B2(n_1070), .C(n_1074), .Y(n_1069) );
AOI22xp33_ASAP7_75t_SL g1101 ( .A1(n_79), .A2(n_212), .B1(n_1003), .B2(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g859 ( .A(n_80), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_80), .A2(n_148), .B1(n_630), .B2(n_886), .Y(n_889) );
INVxp33_ASAP7_75t_L g1158 ( .A(n_81), .Y(n_1158) );
INVx1_ASAP7_75t_L g1203 ( .A(n_82), .Y(n_1203) );
CKINVDCx5p33_ASAP7_75t_R g1183 ( .A(n_83), .Y(n_1183) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_85), .A2(n_241), .B1(n_569), .B2(n_1102), .Y(n_1175) );
OAI211xp5_ASAP7_75t_SL g1187 ( .A1(n_85), .A2(n_524), .B(n_1188), .C(n_1199), .Y(n_1187) );
INVx1_ASAP7_75t_L g680 ( .A(n_86), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_86), .A2(n_217), .B1(n_576), .B2(n_705), .Y(n_714) );
INVx1_ASAP7_75t_L g748 ( .A(n_87), .Y(n_748) );
INVxp67_ASAP7_75t_SL g1118 ( .A(n_88), .Y(n_1118) );
AOI22xp33_ASAP7_75t_SL g1137 ( .A1(n_88), .A2(n_127), .B1(n_978), .B2(n_1132), .Y(n_1137) );
INVx1_ASAP7_75t_L g1019 ( .A(n_89), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_90), .A2(n_226), .B1(n_619), .B2(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_90), .A2(n_226), .B1(n_630), .B2(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g861 ( .A(n_91), .Y(n_861) );
AOI22xp33_ASAP7_75t_SL g888 ( .A1(n_91), .A2(n_210), .B1(n_531), .B2(n_713), .Y(n_888) );
INVx1_ASAP7_75t_L g1073 ( .A(n_92), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_92), .A2(n_213), .B1(n_1098), .B2(n_1099), .Y(n_1097) );
INVx1_ASAP7_75t_L g1265 ( .A(n_93), .Y(n_1265) );
OAI22xp5_ASAP7_75t_L g1478 ( .A1(n_94), .A2(n_140), .B1(n_782), .B2(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g1506 ( .A(n_94), .Y(n_1506) );
INVxp67_ASAP7_75t_SL g657 ( .A(n_95), .Y(n_657) );
INVx1_ASAP7_75t_L g855 ( .A(n_97), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_97), .A2(n_143), .B1(n_619), .B2(n_872), .Y(n_871) );
XNOR2x2_ASAP7_75t_L g944 ( .A(n_98), .B(n_945), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g1149 ( .A1(n_99), .A2(n_135), .B1(n_1005), .B2(n_1006), .Y(n_1149) );
INVxp33_ASAP7_75t_SL g1155 ( .A(n_99), .Y(n_1155) );
INVx1_ASAP7_75t_L g1180 ( .A(n_100), .Y(n_1180) );
AOI221xp5_ASAP7_75t_L g1195 ( .A1(n_100), .A2(n_191), .B1(n_626), .B2(n_1196), .C(n_1198), .Y(n_1195) );
INVx1_ASAP7_75t_L g813 ( .A(n_101), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_101), .A2(n_160), .B1(n_511), .B2(n_517), .Y(n_818) );
INVx1_ASAP7_75t_L g771 ( .A(n_102), .Y(n_771) );
INVx1_ASAP7_75t_L g937 ( .A(n_103), .Y(n_937) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_104), .Y(n_414) );
AO22x2_ASAP7_75t_L g841 ( .A1(n_105), .A2(n_842), .B1(n_843), .B2(n_892), .Y(n_841) );
INVxp67_ASAP7_75t_SL g842 ( .A(n_105), .Y(n_842) );
OAI222xp33_ASAP7_75t_L g846 ( .A1(n_106), .A2(n_188), .B1(n_224), .B2(n_646), .C1(n_649), .C2(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g862 ( .A(n_106), .Y(n_862) );
INVxp33_ASAP7_75t_L g651 ( .A(n_107), .Y(n_651) );
INVx1_ASAP7_75t_L g392 ( .A(n_108), .Y(n_392) );
INVx1_ASAP7_75t_L g558 ( .A(n_108), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_109), .A2(n_125), .B1(n_695), .B2(n_880), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_109), .A2(n_125), .B1(n_531), .B2(n_633), .Y(n_883) );
CKINVDCx5p33_ASAP7_75t_R g929 ( .A(n_110), .Y(n_929) );
AOI22xp5_ASAP7_75t_L g1248 ( .A1(n_111), .A2(n_157), .B1(n_1249), .B2(n_1252), .Y(n_1248) );
INVx1_ASAP7_75t_L g1482 ( .A(n_112), .Y(n_1482) );
AOI22xp33_ASAP7_75t_SL g1517 ( .A1(n_112), .A2(n_113), .B1(n_1034), .B2(n_1518), .Y(n_1517) );
INVx1_ASAP7_75t_L g1483 ( .A(n_113), .Y(n_1483) );
AOI22xp33_ASAP7_75t_L g1475 ( .A1(n_114), .A2(n_235), .B1(n_876), .B2(n_1135), .Y(n_1475) );
INVx1_ASAP7_75t_L g1497 ( .A(n_114), .Y(n_1497) );
AOI22x1_ASAP7_75t_L g894 ( .A1(n_115), .A2(n_895), .B1(n_896), .B2(n_938), .Y(n_894) );
INVxp67_ASAP7_75t_SL g938 ( .A(n_115), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_116), .Y(n_411) );
INVx1_ASAP7_75t_L g851 ( .A(n_117), .Y(n_851) );
AOI22xp33_ASAP7_75t_SL g869 ( .A1(n_117), .A2(n_224), .B1(n_695), .B2(n_870), .Y(n_869) );
XNOR2xp5_ASAP7_75t_L g794 ( .A(n_119), .B(n_795), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g1170 ( .A(n_121), .Y(n_1170) );
INVx1_ASAP7_75t_L g1242 ( .A(n_122), .Y(n_1242) );
CKINVDCx5p33_ASAP7_75t_R g1169 ( .A(n_123), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_124), .A2(n_185), .B1(n_995), .B2(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1207 ( .A(n_124), .Y(n_1207) );
INVx1_ASAP7_75t_L g1477 ( .A(n_126), .Y(n_1477) );
AOI22xp33_ASAP7_75t_L g1515 ( .A1(n_126), .A2(n_253), .B1(n_1512), .B2(n_1516), .Y(n_1515) );
INVxp33_ASAP7_75t_SL g1112 ( .A(n_127), .Y(n_1112) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_128), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g453 ( .A(n_128), .Y(n_453) );
AO221x2_ASAP7_75t_L g1262 ( .A1(n_129), .A2(n_192), .B1(n_1218), .B2(n_1234), .C(n_1263), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_130), .A2(n_259), .B1(n_616), .B2(n_617), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_130), .A2(n_259), .B1(n_373), .B2(n_633), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_131), .A2(n_190), .B1(n_531), .B2(n_904), .Y(n_903) );
OAI221xp5_ASAP7_75t_L g923 ( .A1(n_131), .A2(n_524), .B1(n_924), .B2(n_925), .C(n_928), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_133), .A2(n_220), .B1(n_886), .B2(n_900), .Y(n_899) );
AOI22xp33_ASAP7_75t_SL g919 ( .A1(n_133), .A2(n_220), .B1(n_762), .B2(n_920), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_134), .A2(n_246), .B1(n_980), .B2(n_981), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_134), .A2(n_246), .B1(n_705), .B2(n_1034), .Y(n_1033) );
INVxp67_ASAP7_75t_SL g1156 ( .A(n_135), .Y(n_1156) );
INVx1_ASAP7_75t_L g948 ( .A(n_136), .Y(n_948) );
INVx1_ASAP7_75t_L g272 ( .A(n_137), .Y(n_272) );
OA22x2_ASAP7_75t_L g293 ( .A1(n_138), .A2(n_294), .B1(n_468), .B2(n_469), .Y(n_293) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_138), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g1524 ( .A1(n_139), .A2(n_1525), .B1(n_1526), .B2(n_1527), .Y(n_1524) );
CKINVDCx5p33_ASAP7_75t_R g1525 ( .A(n_139), .Y(n_1525) );
INVx1_ASAP7_75t_L g1507 ( .A(n_140), .Y(n_1507) );
CKINVDCx5p33_ASAP7_75t_R g1012 ( .A(n_141), .Y(n_1012) );
INVx1_ASAP7_75t_L g673 ( .A(n_142), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_142), .A2(n_156), .B1(n_616), .B2(n_696), .Y(n_701) );
INVx1_ASAP7_75t_L g854 ( .A(n_143), .Y(n_854) );
OAI22xp33_ASAP7_75t_L g837 ( .A1(n_144), .A2(n_168), .B1(n_584), .B2(n_787), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g1254 ( .A1(n_145), .A2(n_183), .B1(n_1232), .B2(n_1234), .Y(n_1254) );
INVx1_ASAP7_75t_L g963 ( .A(n_146), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_146), .A2(n_209), .B1(n_1000), .B2(n_1003), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_147), .A2(n_249), .B1(n_1003), .B2(n_1031), .Y(n_1035) );
INVx1_ASAP7_75t_L g1047 ( .A(n_147), .Y(n_1047) );
INVx1_ASAP7_75t_L g858 ( .A(n_148), .Y(n_858) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_149), .Y(n_503) );
OAI221xp5_ASAP7_75t_L g550 ( .A1(n_149), .A2(n_551), .B1(n_559), .B2(n_560), .C(n_563), .Y(n_550) );
XOR2xp5_ASAP7_75t_L g1055 ( .A(n_150), .B(n_1056), .Y(n_1055) );
CKINVDCx5p33_ASAP7_75t_R g800 ( .A(n_151), .Y(n_800) );
INVx1_ASAP7_75t_L g1079 ( .A(n_152), .Y(n_1079) );
INVx1_ASAP7_75t_L g1258 ( .A(n_153), .Y(n_1258) );
INVxp67_ASAP7_75t_SL g607 ( .A(n_154), .Y(n_607) );
INVx1_ASAP7_75t_L g689 ( .A(n_155), .Y(n_689) );
AOI22xp33_ASAP7_75t_SL g712 ( .A1(n_155), .A2(n_159), .B1(n_531), .B2(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g665 ( .A(n_156), .Y(n_665) );
INVx1_ASAP7_75t_L g1064 ( .A(n_158), .Y(n_1064) );
INVx1_ASAP7_75t_L g684 ( .A(n_159), .Y(n_684) );
INVx1_ASAP7_75t_L g812 ( .A(n_160), .Y(n_812) );
INVx1_ASAP7_75t_L g952 ( .A(n_161), .Y(n_952) );
INVx1_ASAP7_75t_L g1063 ( .A(n_162), .Y(n_1063) );
CKINVDCx5p33_ASAP7_75t_R g951 ( .A(n_163), .Y(n_951) );
INVx1_ASAP7_75t_L g1061 ( .A(n_164), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_165), .A2(n_195), .B1(n_695), .B2(n_696), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_165), .A2(n_195), .B1(n_531), .B2(n_633), .Y(n_707) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_166), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_167), .A2(n_189), .B1(n_977), .B2(n_978), .Y(n_976) );
AOI22xp33_ASAP7_75t_SL g997 ( .A1(n_167), .A2(n_189), .B1(n_998), .B2(n_1000), .Y(n_997) );
INVx1_ASAP7_75t_L g831 ( .A(n_168), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g1270 ( .A1(n_169), .A2(n_177), .B1(n_1249), .B2(n_1252), .Y(n_1270) );
CKINVDCx5p33_ASAP7_75t_R g801 ( .A(n_170), .Y(n_801) );
INVx1_ASAP7_75t_L g1075 ( .A(n_171), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_171), .A2(n_199), .B1(n_902), .B2(n_998), .Y(n_1096) );
INVx1_ASAP7_75t_L g546 ( .A(n_173), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g730 ( .A(n_174), .Y(n_730) );
INVxp33_ASAP7_75t_SL g1113 ( .A(n_175), .Y(n_1113) );
AOI22xp33_ASAP7_75t_SL g1134 ( .A1(n_175), .A2(n_207), .B1(n_1128), .B2(n_1135), .Y(n_1134) );
INVx1_ASAP7_75t_L g1185 ( .A(n_176), .Y(n_1185) );
AOI22xp5_ASAP7_75t_L g1271 ( .A1(n_178), .A2(n_215), .B1(n_1218), .B2(n_1272), .Y(n_1271) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_179), .Y(n_274) );
AND3x2_ASAP7_75t_L g1222 ( .A(n_179), .B(n_272), .C(n_1223), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_179), .B(n_272), .Y(n_1239) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_180), .Y(n_334) );
INVx2_ASAP7_75t_L g285 ( .A(n_181), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g668 ( .A(n_182), .Y(n_668) );
CKINVDCx5p33_ASAP7_75t_R g732 ( .A(n_184), .Y(n_732) );
INVx1_ASAP7_75t_L g1209 ( .A(n_185), .Y(n_1209) );
INVx1_ASAP7_75t_L g803 ( .A(n_186), .Y(n_803) );
AOI21xp33_ASAP7_75t_L g825 ( .A1(n_186), .A2(n_433), .B(n_826), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g1487 ( .A1(n_187), .A2(n_205), .B1(n_980), .B2(n_981), .Y(n_1487) );
AOI22xp33_ASAP7_75t_L g1509 ( .A1(n_187), .A2(n_205), .B1(n_705), .B2(n_1510), .Y(n_1509) );
INVx1_ASAP7_75t_L g863 ( .A(n_188), .Y(n_863) );
INVx1_ASAP7_75t_L g922 ( .A(n_190), .Y(n_922) );
INVx1_ASAP7_75t_L g1182 ( .A(n_191), .Y(n_1182) );
AOI22xp5_ASAP7_75t_L g1289 ( .A1(n_193), .A2(n_200), .B1(n_1232), .B2(n_1234), .Y(n_1289) );
AOI22xp33_ASAP7_75t_L g1127 ( .A1(n_194), .A2(n_211), .B1(n_1128), .B2(n_1129), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_194), .A2(n_211), .B1(n_1140), .B2(n_1141), .Y(n_1139) );
INVx1_ASAP7_75t_L g780 ( .A(n_196), .Y(n_780) );
INVx1_ASAP7_75t_L g1223 ( .A(n_197), .Y(n_1223) );
INVx1_ASAP7_75t_L g955 ( .A(n_198), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_198), .A2(n_222), .B1(n_965), .B2(n_966), .Y(n_964) );
INVx1_ASAP7_75t_L g1076 ( .A(n_199), .Y(n_1076) );
INVx1_ASAP7_75t_L g816 ( .A(n_201), .Y(n_816) );
CKINVDCx16_ASAP7_75t_R g587 ( .A(n_202), .Y(n_587) );
INVx1_ASAP7_75t_L g1306 ( .A(n_203), .Y(n_1306) );
INVx1_ASAP7_75t_L g739 ( .A(n_204), .Y(n_739) );
OAI221xp5_ASAP7_75t_L g759 ( .A1(n_204), .A2(n_522), .B1(n_760), .B2(n_763), .C(n_767), .Y(n_759) );
INVx1_ASAP7_75t_L g969 ( .A(n_206), .Y(n_969) );
INVxp33_ASAP7_75t_L g1116 ( .A(n_207), .Y(n_1116) );
INVx1_ASAP7_75t_L g287 ( .A(n_208), .Y(n_287) );
INVx2_ASAP7_75t_L g305 ( .A(n_208), .Y(n_305) );
INVx1_ASAP7_75t_L g971 ( .A(n_209), .Y(n_971) );
INVx1_ASAP7_75t_L g865 ( .A(n_210), .Y(n_865) );
OAI221xp5_ASAP7_75t_L g1077 ( .A1(n_212), .A2(n_524), .B1(n_1078), .B2(n_1083), .C(n_1089), .Y(n_1077) );
INVx1_ASAP7_75t_L g1071 ( .A(n_213), .Y(n_1071) );
AOI22xp5_ASAP7_75t_L g1288 ( .A1(n_214), .A2(n_242), .B1(n_1249), .B2(n_1252), .Y(n_1288) );
INVx1_ASAP7_75t_L g482 ( .A(n_216), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g530 ( .A1(n_216), .A2(n_237), .B1(n_531), .B2(n_533), .C(n_536), .Y(n_530) );
INVx1_ASAP7_75t_L g679 ( .A(n_217), .Y(n_679) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_218), .Y(n_299) );
INVx1_ASAP7_75t_L g1498 ( .A(n_219), .Y(n_1498) );
CKINVDCx5p33_ASAP7_75t_R g734 ( .A(n_221), .Y(n_734) );
INVx1_ASAP7_75t_L g959 ( .A(n_222), .Y(n_959) );
INVx1_ASAP7_75t_L g1021 ( .A(n_223), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_223), .A2(n_230), .B1(n_977), .B2(n_978), .Y(n_1028) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_227), .Y(n_492) );
INVx1_ASAP7_75t_L g425 ( .A(n_229), .Y(n_425) );
INVx1_ASAP7_75t_L g1015 ( .A(n_230), .Y(n_1015) );
INVx1_ASAP7_75t_L g502 ( .A(n_231), .Y(n_502) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_231), .Y(n_559) );
OAI211xp5_ASAP7_75t_L g370 ( .A1(n_232), .A2(n_371), .B(n_376), .C(n_387), .Y(n_370) );
INVx1_ASAP7_75t_L g460 ( .A(n_232), .Y(n_460) );
INVx1_ASAP7_75t_L g599 ( .A(n_233), .Y(n_599) );
INVx1_ASAP7_75t_L g1320 ( .A(n_234), .Y(n_1320) );
INVx1_ASAP7_75t_L g1495 ( .A(n_235), .Y(n_1495) );
INVx1_ASAP7_75t_L g683 ( .A(n_236), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g484 ( .A1(n_237), .A2(n_433), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g1221 ( .A(n_238), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_238), .B(n_1241), .Y(n_1244) );
INVx1_ASAP7_75t_L g1045 ( .A(n_239), .Y(n_1045) );
INVx1_ASAP7_75t_L g1119 ( .A(n_240), .Y(n_1119) );
OAI22xp5_ASAP7_75t_L g1153 ( .A1(n_240), .A2(n_254), .B1(n_609), .B2(n_1042), .Y(n_1153) );
OAI221xp5_ASAP7_75t_L g1200 ( .A1(n_241), .A2(n_522), .B1(n_1201), .B2(n_1206), .C(n_1211), .Y(n_1200) );
INVx1_ASAP7_75t_L g1067 ( .A(n_243), .Y(n_1067) );
INVx1_ASAP7_75t_L g1115 ( .A(n_244), .Y(n_1115) );
OAI211xp5_ASAP7_75t_L g315 ( .A1(n_245), .A2(n_316), .B(n_321), .C(n_328), .Y(n_315) );
INVx1_ASAP7_75t_L g421 ( .A(n_245), .Y(n_421) );
INVx1_ASAP7_75t_L g593 ( .A(n_247), .Y(n_593) );
INVx1_ASAP7_75t_L g1013 ( .A(n_248), .Y(n_1013) );
INVx1_ASAP7_75t_L g1039 ( .A(n_249), .Y(n_1039) );
INVx2_ASAP7_75t_L g284 ( .A(n_250), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g1499 ( .A(n_251), .B(n_1500), .Y(n_1499) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_252), .Y(n_804) );
INVx1_ASAP7_75t_L g1488 ( .A(n_253), .Y(n_1488) );
INVx1_ASAP7_75t_L g1120 ( .A(n_254), .Y(n_1120) );
INVx1_ASAP7_75t_L g669 ( .A(n_255), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_255), .A2(n_256), .B1(n_619), .B2(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g666 ( .A(n_256), .Y(n_666) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_258), .Y(n_406) );
INVx1_ASAP7_75t_L g352 ( .A(n_260), .Y(n_352) );
BUFx3_ASAP7_75t_L g368 ( .A(n_260), .Y(n_368) );
BUFx3_ASAP7_75t_L g351 ( .A(n_261), .Y(n_351) );
INVx1_ASAP7_75t_L g361 ( .A(n_261), .Y(n_361) );
INVx1_ASAP7_75t_L g917 ( .A(n_263), .Y(n_917) );
CKINVDCx5p33_ASAP7_75t_R g1179 ( .A(n_264), .Y(n_1179) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_265), .Y(n_380) );
INVx1_ASAP7_75t_L g742 ( .A(n_266), .Y(n_742) );
OAI211xp5_ASAP7_75t_L g768 ( .A1(n_266), .A2(n_524), .B(n_769), .C(n_776), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_288), .B(n_1215), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_275), .Y(n_269) );
AND2x4_ASAP7_75t_L g1522 ( .A(n_270), .B(n_276), .Y(n_1522) );
NOR2xp33_ASAP7_75t_SL g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_SL g1531 ( .A(n_271), .Y(n_1531) );
NAND2xp5_ASAP7_75t_L g1536 ( .A(n_271), .B(n_273), .Y(n_1536) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g1530 ( .A(n_273), .B(n_1531), .Y(n_1530) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_281), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g295 ( .A(n_278), .B(n_296), .Y(n_295) );
OR2x6_ASAP7_75t_L g590 ( .A(n_278), .B(n_296), .Y(n_590) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g614 ( .A(n_279), .B(n_287), .Y(n_614) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g433 ( .A(n_280), .B(n_304), .Y(n_433) );
INVx8_ASAP7_75t_L g298 ( .A(n_281), .Y(n_298) );
OR2x6_ASAP7_75t_L g281 ( .A(n_282), .B(n_286), .Y(n_281) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_282), .Y(n_435) );
OR2x6_ASAP7_75t_L g601 ( .A(n_282), .B(n_303), .Y(n_601) );
INVx1_ASAP7_75t_L g765 ( .A(n_282), .Y(n_765) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx2_ASAP7_75t_L g308 ( .A(n_284), .Y(n_308) );
AND2x4_ASAP7_75t_L g313 ( .A(n_284), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g320 ( .A(n_284), .Y(n_320) );
INVx1_ASAP7_75t_L g327 ( .A(n_284), .Y(n_327) );
AND2x2_ASAP7_75t_L g332 ( .A(n_284), .B(n_285), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_285), .B(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g314 ( .A(n_285), .Y(n_314) );
INVx1_ASAP7_75t_L g319 ( .A(n_285), .Y(n_319) );
INVx1_ASAP7_75t_L g336 ( .A(n_285), .Y(n_336) );
INVx1_ASAP7_75t_L g516 ( .A(n_285), .Y(n_516) );
AND2x4_ASAP7_75t_L g335 ( .A(n_286), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g966 ( .A(n_287), .B(n_339), .Y(n_966) );
OR2x2_ASAP7_75t_L g1042 ( .A(n_287), .B(n_339), .Y(n_1042) );
OAI22xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_939), .B1(n_940), .B2(n_1214), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g1214 ( .A(n_290), .Y(n_1214) );
XNOR2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_718), .Y(n_290) );
XNOR2x1_ASAP7_75t_L g291 ( .A(n_292), .B(n_585), .Y(n_291) );
XNOR2x1_ASAP7_75t_L g292 ( .A(n_293), .B(n_470), .Y(n_292) );
INVx1_ASAP7_75t_L g468 ( .A(n_294), .Y(n_468) );
OAI211xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_297), .B(n_342), .C(n_395), .Y(n_294) );
AOI31xp33_ASAP7_75t_L g1037 ( .A1(n_295), .A2(n_1038), .A3(n_1043), .B(n_1046), .Y(n_1037) );
AOI31xp33_ASAP7_75t_L g1150 ( .A1(n_295), .A2(n_1151), .A3(n_1154), .B(n_1157), .Y(n_1150) );
AND2x4_ASAP7_75t_L g428 ( .A(n_296), .B(n_429), .Y(n_428) );
AND2x4_ASAP7_75t_L g577 ( .A(n_296), .B(n_578), .Y(n_577) );
AND2x4_ASAP7_75t_L g641 ( .A(n_296), .B(n_429), .Y(n_641) );
AOI211xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B(n_300), .C(n_315), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_298), .A2(n_598), .B1(n_599), .B2(n_600), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_298), .A2(n_600), .B1(n_668), .B2(n_689), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_298), .A2(n_852), .B1(n_865), .B2(n_866), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_298), .A2(n_600), .B1(n_951), .B2(n_971), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_298), .A2(n_866), .B1(n_1012), .B2(n_1047), .Y(n_1046) );
AOI22xp33_ASAP7_75t_SL g1157 ( .A1(n_298), .A2(n_866), .B1(n_1115), .B2(n_1158), .Y(n_1157) );
OAI22xp33_ASAP7_75t_L g418 ( .A1(n_299), .A2(n_412), .B1(n_419), .B2(n_421), .Y(n_418) );
OR2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_306), .Y(n_301) );
AOI322xp5_ASAP7_75t_L g328 ( .A1(n_302), .A2(n_329), .A3(n_333), .B1(n_334), .B2(n_335), .C1(n_337), .C2(n_341), .Y(n_328) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x4_ASAP7_75t_L g310 ( .A(n_303), .B(n_311), .Y(n_310) );
AND2x4_ASAP7_75t_L g594 ( .A(n_303), .B(n_514), .Y(n_594) );
AND2x4_ASAP7_75t_L g596 ( .A(n_303), .B(n_311), .Y(n_596) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g325 ( .A(n_305), .Y(n_325) );
INVx2_ASAP7_75t_L g441 ( .A(n_306), .Y(n_441) );
BUFx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g448 ( .A(n_307), .Y(n_448) );
INVx1_ASAP7_75t_L g476 ( .A(n_307), .Y(n_476) );
INVx1_ASAP7_75t_L g505 ( .A(n_308), .Y(n_505) );
AND2x4_ASAP7_75t_L g514 ( .A(n_308), .B(n_515), .Y(n_514) );
INVx5_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_310), .A2(n_594), .B1(n_1044), .B2(n_1045), .Y(n_1043) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g444 ( .A(n_313), .Y(n_444) );
INVx3_ASAP7_75t_L g452 ( .A(n_313), .Y(n_452) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_313), .Y(n_762) );
AND2x4_ASAP7_75t_L g326 ( .A(n_314), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g438 ( .A(n_318), .Y(n_438) );
INVx3_ASAP7_75t_L g483 ( .A(n_318), .Y(n_483) );
INVx2_ASAP7_75t_L g493 ( .A(n_318), .Y(n_493) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_319), .B(n_320), .Y(n_459) );
INVx1_ASAP7_75t_L g339 ( .A(n_320), .Y(n_339) );
NAND4xp25_ASAP7_75t_SL g591 ( .A(n_321), .B(n_592), .C(n_597), .D(n_602), .Y(n_591) );
NAND4xp25_ASAP7_75t_SL g677 ( .A(n_321), .B(n_678), .C(n_681), .D(n_688), .Y(n_677) );
NAND4xp25_ASAP7_75t_SL g856 ( .A(n_321), .B(n_857), .C(n_860), .D(n_864), .Y(n_856) );
CKINVDCx11_ASAP7_75t_R g321 ( .A(n_322), .Y(n_321) );
AOI211xp5_ASAP7_75t_L g962 ( .A1(n_322), .A2(n_696), .B(n_963), .C(n_964), .Y(n_962) );
AOI211xp5_ASAP7_75t_L g1038 ( .A1(n_322), .A2(n_1039), .B(n_1040), .C(n_1041), .Y(n_1038) );
AOI211xp5_ASAP7_75t_L g1151 ( .A1(n_322), .A2(n_1040), .B(n_1152), .C(n_1153), .Y(n_1151) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_326), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVxp67_ASAP7_75t_L g340 ( .A(n_324), .Y(n_340) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2x1p5_ASAP7_75t_L g466 ( .A(n_325), .B(n_467), .Y(n_466) );
BUFx3_ASAP7_75t_L g526 ( .A(n_326), .Y(n_526) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_326), .Y(n_606) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_326), .Y(n_626) );
BUFx2_ASAP7_75t_L g687 ( .A(n_326), .Y(n_687) );
BUFx3_ASAP7_75t_L g775 ( .A(n_326), .Y(n_775) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g695 ( .A(n_330), .Y(n_695) );
INVx2_ASAP7_75t_SL g826 ( .A(n_330), .Y(n_826) );
INVx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_331), .Y(n_499) );
AND2x4_ASAP7_75t_L g523 ( .A(n_331), .B(n_513), .Y(n_523) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx3_ASAP7_75t_L g486 ( .A(n_332), .Y(n_486) );
AOI322xp5_ASAP7_75t_L g376 ( .A1(n_334), .A2(n_341), .A3(n_377), .B1(n_379), .B2(n_380), .C1(n_381), .C2(n_385), .Y(n_376) );
INVx2_ASAP7_75t_L g609 ( .A(n_335), .Y(n_609) );
AOI222xp33_ASAP7_75t_L g681 ( .A1(n_335), .A2(n_337), .B1(n_682), .B2(n_683), .C1(n_684), .C2(n_685), .Y(n_681) );
INVx2_ASAP7_75t_L g965 ( .A(n_335), .Y(n_965) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_336), .A2(n_502), .B1(n_503), .B2(n_504), .Y(n_501) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_336), .Y(n_779) );
INVx1_ASAP7_75t_L g933 ( .A(n_336), .Y(n_933) );
AOI222xp33_ASAP7_75t_L g602 ( .A1(n_337), .A2(n_603), .B1(n_604), .B2(n_607), .C1(n_608), .C2(n_610), .Y(n_602) );
AOI222xp33_ASAP7_75t_L g860 ( .A1(n_337), .A2(n_604), .B1(n_608), .B2(n_861), .C1(n_862), .C2(n_863), .Y(n_860) );
AND2x4_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g931 ( .A1(n_338), .A2(n_910), .B1(n_912), .B2(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI31xp33_ASAP7_75t_SL g342 ( .A1(n_343), .A2(n_353), .A3(n_370), .B(n_390), .Y(n_342) );
INVx4_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_345), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_345), .A2(n_664), .B1(n_665), .B2(n_666), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_345), .A2(n_655), .B1(n_854), .B2(n_855), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_345), .A2(n_363), .B1(n_951), .B2(n_952), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_345), .A2(n_363), .B1(n_1012), .B2(n_1013), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_345), .A2(n_363), .B1(n_1115), .B2(n_1116), .Y(n_1114) );
AND2x6_ASAP7_75t_L g345 ( .A(n_346), .B(n_349), .Y(n_345) );
AND2x4_ASAP7_75t_L g652 ( .A(n_346), .B(n_653), .Y(n_652) );
AND2x4_ASAP7_75t_L g664 ( .A(n_346), .B(n_653), .Y(n_664) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g647 ( .A(n_347), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g357 ( .A(n_348), .Y(n_357) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_348), .Y(n_365) );
AND2x2_ASAP7_75t_L g399 ( .A(n_348), .B(n_392), .Y(n_399) );
INVx2_ASAP7_75t_L g430 ( .A(n_348), .Y(n_430) );
INVx1_ASAP7_75t_L g426 ( .A(n_349), .Y(n_426) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_349), .Y(n_631) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_349), .Y(n_640) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_349), .Y(n_747) );
INVx2_ASAP7_75t_L g996 ( .A(n_349), .Y(n_996) );
INVx1_ASAP7_75t_L g1142 ( .A(n_349), .Y(n_1142) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g409 ( .A(n_350), .Y(n_409) );
INVx1_ASAP7_75t_L g539 ( .A(n_350), .Y(n_539) );
INVx1_ASAP7_75t_L g582 ( .A(n_350), .Y(n_582) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_350), .Y(n_706) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx2_ASAP7_75t_L g369 ( .A(n_351), .Y(n_369) );
AND2x2_ASAP7_75t_L g375 ( .A(n_351), .B(n_368), .Y(n_375) );
INVx1_ASAP7_75t_L g359 ( .A(n_352), .Y(n_359) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_358), .Y(n_354) );
INVx1_ASAP7_75t_L g379 ( .A(n_355), .Y(n_379) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g372 ( .A(n_356), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g389 ( .A(n_356), .Y(n_389) );
AND2x6_ASAP7_75t_L g655 ( .A(n_356), .B(n_378), .Y(n_655) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x6_ASAP7_75t_L g385 ( .A(n_357), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g413 ( .A(n_358), .Y(n_413) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
AND2x2_ASAP7_75t_L g417 ( .A(n_359), .B(n_360), .Y(n_417) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g378 ( .A(n_361), .B(n_368), .Y(n_378) );
INVx4_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_363), .A2(n_599), .B1(n_651), .B2(n_652), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g667 ( .A1(n_363), .A2(n_655), .B1(n_668), .B2(n_669), .C(n_670), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_363), .A2(n_664), .B1(n_851), .B2(n_852), .Y(n_850) );
AND2x4_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
AND2x2_ASAP7_75t_SL g381 ( .A(n_364), .B(n_382), .Y(n_381) );
AND2x4_ASAP7_75t_L g958 ( .A(n_364), .B(n_382), .Y(n_958) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx6_ASAP7_75t_L g535 ( .A(n_366), .Y(n_535) );
INVx2_ASAP7_75t_L g570 ( .A(n_366), .Y(n_570) );
AND2x2_ASAP7_75t_L g578 ( .A(n_366), .B(n_556), .Y(n_578) );
BUFx2_ASAP7_75t_L g636 ( .A(n_366), .Y(n_636) );
AND2x4_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
INVx1_ASAP7_75t_L g386 ( .A(n_367), .Y(n_386) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g384 ( .A(n_369), .Y(n_384) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI211xp5_ASAP7_75t_L g643 ( .A1(n_372), .A2(n_388), .B(n_644), .C(n_645), .Y(n_643) );
HB1xp67_ASAP7_75t_L g1016 ( .A(n_373), .Y(n_1016) );
HB1xp67_ASAP7_75t_L g1145 ( .A(n_373), .Y(n_1145) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_L g388 ( .A(n_374), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g532 ( .A(n_374), .Y(n_532) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_374), .Y(n_674) );
INVx1_ASAP7_75t_L g725 ( .A(n_374), .Y(n_725) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_375), .Y(n_565) );
INVx2_ASAP7_75t_L g405 ( .A(n_377), .Y(n_405) );
INVx1_ASAP7_75t_L g744 ( .A(n_377), .Y(n_744) );
INVx2_ASAP7_75t_SL g799 ( .A(n_377), .Y(n_799) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_SL g424 ( .A(n_378), .Y(n_424) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_378), .Y(n_538) );
BUFx2_ASAP7_75t_L g630 ( .A(n_378), .Y(n_630) );
BUFx3_ASAP7_75t_L g729 ( .A(n_378), .Y(n_729) );
BUFx6f_ASAP7_75t_L g793 ( .A(n_378), .Y(n_793) );
BUFx2_ASAP7_75t_L g885 ( .A(n_378), .Y(n_885) );
BUFx6f_ASAP7_75t_L g994 ( .A(n_378), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_380), .A2(n_446), .B1(n_449), .B2(n_453), .Y(n_445) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g648 ( .A(n_383), .Y(n_648) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g553 ( .A(n_384), .Y(n_553) );
INVx3_ASAP7_75t_L g649 ( .A(n_385), .Y(n_649) );
AOI222xp33_ASAP7_75t_L g953 ( .A1(n_385), .A2(n_902), .B1(n_954), .B2(n_955), .C1(n_956), .C2(n_959), .Y(n_953) );
AOI222xp33_ASAP7_75t_L g1014 ( .A1(n_385), .A2(n_1015), .B1(n_1016), .B2(n_1017), .C1(n_1018), .C2(n_1019), .Y(n_1014) );
AOI222xp33_ASAP7_75t_L g1117 ( .A1(n_385), .A2(n_958), .B1(n_1102), .B2(n_1118), .C1(n_1119), .C2(n_1120), .Y(n_1117) );
BUFx3_ASAP7_75t_L g562 ( .A(n_386), .Y(n_562) );
CKINVDCx8_ASAP7_75t_R g387 ( .A(n_388), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g845 ( .A(n_388), .B(n_846), .Y(n_845) );
INVx5_ASAP7_75t_L g960 ( .A(n_388), .Y(n_960) );
OAI21xp33_ASAP7_75t_L g672 ( .A1(n_389), .A2(n_673), .B(n_674), .Y(n_672) );
INVx1_ASAP7_75t_SL g658 ( .A(n_390), .Y(n_658) );
AND2x4_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
AND2x4_ASAP7_75t_L g676 ( .A(n_391), .B(n_393), .Y(n_676) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x4_ASAP7_75t_L g429 ( .A(n_392), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g784 ( .A(n_393), .Y(n_784) );
BUFx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g400 ( .A(n_394), .Y(n_400) );
OR2x6_ASAP7_75t_L g432 ( .A(n_394), .B(n_433), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_431), .Y(n_395) );
OAI33xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_401), .A3(n_410), .B1(n_418), .B2(n_422), .B3(n_427), .Y(n_396) );
INVx1_ASAP7_75t_SL g628 ( .A(n_397), .Y(n_628) );
OAI33xp33_ASAP7_75t_L g726 ( .A1(n_397), .A2(n_727), .A3(n_733), .B1(n_738), .B2(n_743), .B3(n_749), .Y(n_726) );
OAI33xp33_ASAP7_75t_L g797 ( .A1(n_397), .A2(n_749), .A3(n_798), .B1(n_802), .B2(n_805), .B3(n_811), .Y(n_797) );
OR2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_400), .Y(n_397) );
OR2x6_ASAP7_75t_L g541 ( .A(n_398), .B(n_400), .Y(n_541) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g710 ( .A(n_399), .Y(n_710) );
INVx2_ASAP7_75t_L g528 ( .A(n_400), .Y(n_528) );
AND2x4_ASAP7_75t_L g613 ( .A(n_400), .B(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g709 ( .A(n_400), .B(n_710), .Y(n_709) );
AND2x4_ASAP7_75t_L g975 ( .A(n_400), .B(n_614), .Y(n_975) );
BUFx2_ASAP7_75t_L g1491 ( .A(n_400), .Y(n_1491) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_406), .B2(n_407), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_402), .A2(n_406), .B1(n_440), .B2(n_442), .Y(n_439) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_405), .A2(n_546), .B1(n_547), .B2(n_549), .Y(n_545) );
INVx2_ASAP7_75t_SL g1104 ( .A(n_405), .Y(n_1104) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g548 ( .A(n_409), .Y(n_548) );
OAI22xp33_ASAP7_75t_SL g410 ( .A1(n_411), .A2(n_412), .B1(n_414), .B2(n_415), .Y(n_410) );
OAI22xp33_ASAP7_75t_L g434 ( .A1(n_411), .A2(n_414), .B1(n_435), .B2(n_436), .Y(n_434) );
OAI22xp33_ASAP7_75t_L g733 ( .A1(n_412), .A2(n_734), .B1(n_735), .B2(n_737), .Y(n_733) );
OAI22xp33_ASAP7_75t_L g738 ( .A1(n_412), .A2(n_739), .B1(n_740), .B2(n_742), .Y(n_738) );
OAI22xp33_ASAP7_75t_L g802 ( .A1(n_412), .A2(n_735), .B1(n_803), .B2(n_804), .Y(n_802) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g790 ( .A(n_413), .Y(n_790) );
INVx2_ASAP7_75t_L g806 ( .A(n_413), .Y(n_806) );
BUFx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g809 ( .A(n_416), .Y(n_809) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g420 ( .A(n_417), .Y(n_420) );
BUFx2_ASAP7_75t_L g736 ( .A(n_417), .Y(n_736) );
BUFx4f_ASAP7_75t_L g741 ( .A(n_417), .Y(n_741) );
INVx1_ASAP7_75t_L g849 ( .A(n_417), .Y(n_849) );
BUFx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OR2x6_ASAP7_75t_L g584 ( .A(n_420), .B(n_572), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B1(n_425), .B2(n_426), .Y(n_422) );
INVx2_ASAP7_75t_L g576 ( .A(n_424), .Y(n_576) );
INVx1_ASAP7_75t_L g900 ( .A(n_424), .Y(n_900) );
INVx4_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g529 ( .A1(n_428), .A2(n_530), .B1(n_540), .B2(n_542), .C(n_550), .Y(n_529) );
BUFx4f_ASAP7_75t_L g1007 ( .A(n_428), .Y(n_1007) );
AOI33xp33_ASAP7_75t_L g1029 ( .A1(n_428), .A2(n_991), .A3(n_1030), .B1(n_1033), .B2(n_1035), .B3(n_1036), .Y(n_1029) );
BUFx4f_ASAP7_75t_L g1106 ( .A(n_428), .Y(n_1106) );
AOI33xp33_ASAP7_75t_L g1138 ( .A1(n_428), .A2(n_991), .A3(n_1139), .B1(n_1143), .B2(n_1146), .B3(n_1149), .Y(n_1138) );
AND2x4_ASAP7_75t_L g556 ( .A(n_430), .B(n_557), .Y(n_556) );
OAI33xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_434), .A3(n_439), .B1(n_445), .B2(n_454), .B3(n_461), .Y(n_431) );
OAI22xp33_ASAP7_75t_L g454 ( .A1(n_435), .A2(n_455), .B1(n_456), .B2(n_460), .Y(n_454) );
OAI221xp5_ASAP7_75t_L g1074 ( .A1(n_435), .A2(n_458), .B1(n_766), .B2(n_1075), .C(n_1076), .Y(n_1074) );
OAI221xp5_ASAP7_75t_L g1078 ( .A1(n_435), .A2(n_483), .B1(n_1064), .B2(n_1079), .C(n_1080), .Y(n_1078) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_438), .B(n_501), .Y(n_500) );
OR2x6_ASAP7_75t_L g767 ( .A(n_438), .B(n_507), .Y(n_767) );
OR2x2_ASAP7_75t_L g1211 ( .A(n_438), .B(n_507), .Y(n_1211) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_440), .A2(n_800), .B1(n_801), .B2(n_821), .Y(n_820) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x4_ASAP7_75t_L g518 ( .A(n_443), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g1194 ( .A(n_444), .Y(n_1194) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_446), .A2(n_730), .B1(n_732), .B2(n_761), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g1070 ( .A1(n_446), .A2(n_1071), .B1(n_1072), .B2(n_1073), .Y(n_1070) );
INVx2_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g1208 ( .A(n_447), .Y(n_1208) );
BUFx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g1190 ( .A(n_448), .Y(n_1190) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g700 ( .A(n_451), .Y(n_700) );
INVx3_ASAP7_75t_L g1087 ( .A(n_451), .Y(n_1087) );
INVx2_ASAP7_75t_L g1130 ( .A(n_451), .Y(n_1130) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx3_ASAP7_75t_L g479 ( .A(n_452), .Y(n_479) );
INVx3_ASAP7_75t_L g822 ( .A(n_452), .Y(n_822) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI221xp5_ASAP7_75t_L g763 ( .A1(n_458), .A2(n_734), .B1(n_737), .B2(n_764), .C(n_766), .Y(n_763) );
BUFx3_ASAP7_75t_L g824 ( .A(n_458), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_458), .B(n_931), .Y(n_930) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AOI33xp33_ASAP7_75t_L g612 ( .A1(n_462), .A2(n_613), .A3(n_615), .B1(n_618), .B2(n_622), .B3(n_624), .Y(n_612) );
AOI33xp33_ASAP7_75t_L g973 ( .A1(n_462), .A2(n_974), .A3(n_976), .B1(n_979), .B2(n_982), .B3(n_987), .Y(n_973) );
AOI33xp33_ASAP7_75t_L g1024 ( .A1(n_462), .A2(n_974), .A3(n_1025), .B1(n_1026), .B2(n_1027), .B3(n_1028), .Y(n_1024) );
INVx6_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx5_ASAP7_75t_L g702 ( .A(n_463), .Y(n_702) );
OR2x6_ASAP7_75t_L g463 ( .A(n_464), .B(n_466), .Y(n_463) );
NAND2x1p5_ASAP7_75t_L g555 ( .A(n_464), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g572 ( .A(n_465), .B(n_573), .Y(n_572) );
BUFx2_ASAP7_75t_L g496 ( .A(n_466), .Y(n_496) );
INVx2_ASAP7_75t_L g1082 ( .A(n_466), .Y(n_1082) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_472), .B(n_529), .C(n_567), .D(n_579), .Y(n_471) );
OAI31xp33_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_510), .A3(n_521), .B(n_527), .Y(n_472) );
OAI221xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_481), .B1(n_487), .B2(n_491), .C(n_497), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_477), .B1(n_478), .B2(n_480), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_475), .A2(n_488), .B1(n_489), .B2(n_490), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_475), .A2(n_489), .B1(n_926), .B2(n_927), .Y(n_925) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g770 ( .A(n_476), .Y(n_770) );
INVx1_ASAP7_75t_L g1085 ( .A(n_476), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_477), .A2(n_480), .B1(n_537), .B2(n_539), .Y(n_536) );
INVx2_ASAP7_75t_L g623 ( .A(n_478), .Y(n_623) );
INVx2_ASAP7_75t_SL g693 ( .A(n_478), .Y(n_693) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g489 ( .A(n_479), .Y(n_489) );
INVx2_ASAP7_75t_L g873 ( .A(n_479), .Y(n_873) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B(n_484), .Y(n_481) );
BUFx2_ASAP7_75t_L g1202 ( .A(n_483), .Y(n_1202) );
BUFx2_ASAP7_75t_L g616 ( .A(n_485), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_485), .B(n_756), .Y(n_755) );
INVx2_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g495 ( .A(n_486), .Y(n_495) );
INVx2_ASAP7_75t_SL g1133 ( .A(n_486), .Y(n_1133) );
AOI222xp33_ASAP7_75t_L g567 ( .A1(n_488), .A2(n_498), .B1(n_568), .B2(n_574), .C1(n_575), .C2(n_577), .Y(n_567) );
INVx1_ASAP7_75t_L g621 ( .A(n_489), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_490), .A2(n_492), .B1(n_580), .B2(n_583), .Y(n_579) );
OAI21xp33_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .B(n_494), .Y(n_491) );
BUFx3_ASAP7_75t_L g977 ( .A(n_495), .Y(n_977) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B(n_500), .C(n_506), .Y(n_497) );
INVx1_ASAP7_75t_L g989 ( .A(n_499), .Y(n_989) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OR2x6_ASAP7_75t_L g782 ( .A(n_505), .B(n_507), .Y(n_782) );
A2O1A1Ixp33_ASAP7_75t_L g928 ( .A1(n_506), .A2(n_695), .B(n_929), .C(n_930), .Y(n_928) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g756 ( .A(n_507), .Y(n_756) );
INVx1_ASAP7_75t_L g1480 ( .A(n_507), .Y(n_1480) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_512), .A2(n_518), .B1(n_916), .B2(n_917), .Y(n_915) );
INVx3_ASAP7_75t_L g1092 ( .A(n_512), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g1481 ( .A1(n_512), .A2(n_518), .B1(n_1482), .B2(n_1483), .Y(n_1481) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
INVx2_ASAP7_75t_L g520 ( .A(n_513), .Y(n_520) );
INVx1_ASAP7_75t_L g620 ( .A(n_514), .Y(n_620) );
BUFx2_ASAP7_75t_L g876 ( .A(n_514), .Y(n_876) );
BUFx6f_ASAP7_75t_L g920 ( .A(n_514), .Y(n_920) );
BUFx2_ASAP7_75t_L g980 ( .A(n_514), .Y(n_980) );
BUFx6f_ASAP7_75t_L g985 ( .A(n_514), .Y(n_985) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx3_ASAP7_75t_L g1093 ( .A(n_518), .Y(n_1093) );
AND2x4_ASAP7_75t_L g525 ( .A(n_519), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
CKINVDCx6p67_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g918 ( .A1(n_523), .A2(n_919), .B1(n_921), .B2(n_922), .Y(n_918) );
AOI221xp5_ASAP7_75t_L g1484 ( .A1(n_523), .A2(n_1485), .B1(n_1487), .B2(n_1488), .C(n_1489), .Y(n_1484) );
INVx8_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AOI221xp5_ASAP7_75t_L g1474 ( .A1(n_525), .A2(n_1475), .B1(n_1476), .B2(n_1477), .C(n_1478), .Y(n_1474) );
INVx1_ASAP7_75t_L g881 ( .A(n_526), .Y(n_881) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NOR2xp67_ASAP7_75t_L g754 ( .A(n_528), .B(n_755), .Y(n_754) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_535), .Y(n_544) );
INVx2_ASAP7_75t_L g634 ( .A(n_535), .Y(n_634) );
INVx2_ASAP7_75t_L g653 ( .A(n_535), .Y(n_653) );
INVx1_ASAP7_75t_L g713 ( .A(n_535), .Y(n_713) );
INVx2_ASAP7_75t_SL g906 ( .A(n_535), .Y(n_906) );
INVx2_ASAP7_75t_L g999 ( .A(n_535), .Y(n_999) );
INVx1_ASAP7_75t_L g1514 ( .A(n_535), .Y(n_1514) );
INVx1_ASAP7_75t_L g1098 ( .A(n_537), .Y(n_1098) );
INVx1_ASAP7_75t_L g1173 ( .A(n_537), .Y(n_1173) );
INVx2_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
BUFx3_ASAP7_75t_L g1034 ( .A(n_538), .Y(n_1034) );
OAI22xp33_ASAP7_75t_L g798 ( .A1(n_539), .A2(n_799), .B1(n_800), .B2(n_801), .Y(n_798) );
INVx1_ASAP7_75t_L g1006 ( .A(n_539), .Y(n_1006) );
INVx1_ASAP7_75t_L g1518 ( .A(n_539), .Y(n_1518) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g991 ( .A(n_541), .Y(n_991) );
CKINVDCx5p33_ASAP7_75t_R g1095 ( .A(n_541), .Y(n_1095) );
INVx4_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g886 ( .A(n_547), .Y(n_886) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g909 ( .A(n_551), .Y(n_909) );
INVx1_ASAP7_75t_L g1059 ( .A(n_551), .Y(n_1059) );
INVx2_ASAP7_75t_L g1505 ( .A(n_551), .Y(n_1505) );
NAND2x1p5_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
OR2x6_ASAP7_75t_L g560 ( .A(n_555), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g566 ( .A(n_555), .Y(n_566) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g911 ( .A(n_560), .Y(n_911) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND3xp33_ASAP7_75t_SL g1167 ( .A(n_563), .B(n_1168), .C(n_1171), .Y(n_1167) );
INVx1_ASAP7_75t_L g1503 ( .A(n_563), .Y(n_1503) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
INVx1_ASAP7_75t_L g1148 ( .A(n_564), .Y(n_1148) );
HB1xp67_ASAP7_75t_L g1516 ( .A(n_564), .Y(n_1516) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g638 ( .A(n_565), .Y(n_638) );
BUFx4f_ASAP7_75t_L g902 ( .A(n_565), .Y(n_902) );
INVx2_ASAP7_75t_SL g1001 ( .A(n_565), .Y(n_1001) );
BUFx3_ASAP7_75t_L g1102 ( .A(n_565), .Y(n_1102) );
AND2x2_ASAP7_75t_L g723 ( .A(n_566), .B(n_724), .Y(n_723) );
AOI222xp33_ASAP7_75t_L g934 ( .A1(n_568), .A2(n_577), .B1(n_580), .B2(n_926), .C1(n_929), .C2(n_935), .Y(n_934) );
AOI221xp5_ASAP7_75t_L g1062 ( .A1(n_568), .A2(n_575), .B1(n_1063), .B2(n_1064), .C(n_1065), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1181 ( .A1(n_568), .A2(n_575), .B1(n_1182), .B2(n_1183), .Y(n_1181) );
AOI22xp33_ASAP7_75t_L g1493 ( .A1(n_568), .A2(n_575), .B1(n_1494), .B2(n_1495), .Y(n_1493) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
BUFx2_ASAP7_75t_L g1144 ( .A(n_569), .Y(n_1144) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g1003 ( .A(n_570), .Y(n_1003) );
AND2x2_ASAP7_75t_L g575 ( .A(n_571), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x6_ASAP7_75t_L g581 ( .A(n_572), .B(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g787 ( .A(n_572), .B(n_582), .Y(n_787) );
OR2x2_ASAP7_75t_L g789 ( .A(n_572), .B(n_790), .Y(n_789) );
OR2x2_ASAP7_75t_L g791 ( .A(n_572), .B(n_792), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g936 ( .A1(n_575), .A2(n_583), .B1(n_927), .B2(n_937), .Y(n_936) );
OR2x6_ASAP7_75t_L g753 ( .A(n_577), .B(n_754), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_580), .A2(n_583), .B1(n_1179), .B2(n_1180), .Y(n_1178) );
AOI22xp33_ASAP7_75t_L g1496 ( .A1(n_580), .A2(n_583), .B1(n_1497), .B2(n_1498), .Y(n_1496) );
CKINVDCx6p67_ASAP7_75t_R g580 ( .A(n_581), .Y(n_580) );
CKINVDCx6p67_ASAP7_75t_R g583 ( .A(n_584), .Y(n_583) );
OA22x2_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_659), .B1(n_660), .B2(n_717), .Y(n_585) );
INVx1_ASAP7_75t_L g717 ( .A(n_586), .Y(n_717) );
XNOR2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g1230 ( .A1(n_587), .A2(n_1231), .B1(n_1233), .B2(n_1235), .Y(n_1230) );
AOI211xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_591), .B(n_611), .C(n_642), .Y(n_588) );
AOI221x1_ASAP7_75t_L g661 ( .A1(n_589), .A2(n_662), .B1(n_675), .B2(n_677), .C(n_690), .Y(n_661) );
AOI221x1_ASAP7_75t_L g843 ( .A1(n_589), .A2(n_675), .B1(n_844), .B2(n_856), .C(n_867), .Y(n_843) );
CKINVDCx16_ASAP7_75t_R g589 ( .A(n_590), .Y(n_589) );
AOI31xp33_ASAP7_75t_L g961 ( .A1(n_590), .A2(n_962), .A3(n_967), .B(n_970), .Y(n_961) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B1(n_595), .B2(n_596), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_594), .A2(n_596), .B1(n_679), .B2(n_680), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_594), .A2(n_596), .B1(n_858), .B2(n_859), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_594), .A2(n_596), .B1(n_968), .B2(n_969), .Y(n_967) );
AOI22xp33_ASAP7_75t_SL g1154 ( .A1(n_594), .A2(n_596), .B1(n_1155), .B2(n_1156), .Y(n_1154) );
INVx4_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx5_ASAP7_75t_L g866 ( .A(n_601), .Y(n_866) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_SL g978 ( .A(n_605), .Y(n_978) );
INVx2_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_606), .Y(n_617) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_612), .B(n_627), .Y(n_611) );
NAND3xp33_ASAP7_75t_L g691 ( .A(n_613), .B(n_692), .C(n_694), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g874 ( .A(n_613), .B(n_875), .C(n_879), .Y(n_874) );
BUFx2_ASAP7_75t_SL g766 ( .A(n_614), .Y(n_766) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
BUFx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_SL g697 ( .A(n_626), .Y(n_697) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_626), .Y(n_870) );
AOI33xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .A3(n_632), .B1(n_635), .B2(n_639), .B3(n_641), .Y(n_627) );
AOI33xp33_ASAP7_75t_L g898 ( .A1(n_628), .A2(n_641), .A3(n_899), .B1(n_901), .B2(n_903), .B3(n_907), .Y(n_898) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g711 ( .A(n_641), .B(n_712), .C(n_714), .Y(n_711) );
INVx1_ASAP7_75t_L g749 ( .A(n_641), .Y(n_749) );
INVx1_ASAP7_75t_L g891 ( .A(n_641), .Y(n_891) );
AOI31xp33_ASAP7_75t_SL g642 ( .A1(n_643), .A2(n_650), .A3(n_654), .B(n_658), .Y(n_642) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g671 ( .A(n_647), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_652), .A2(n_655), .B1(n_1112), .B2(n_1113), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_655), .A2(n_664), .B1(n_948), .B2(n_949), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_655), .A2(n_664), .B1(n_1021), .B2(n_1022), .Y(n_1020) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g716 ( .A(n_661), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_667), .Y(n_662) );
INVx1_ASAP7_75t_L g1032 ( .A(n_674), .Y(n_1032) );
AOI211x1_ASAP7_75t_L g945 ( .A1(n_675), .A2(n_946), .B(n_961), .C(n_972), .Y(n_945) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI211x1_ASAP7_75t_SL g1009 ( .A1(n_676), .A2(n_1010), .B(n_1023), .C(n_1037), .Y(n_1009) );
INVx1_ASAP7_75t_L g1122 ( .A(n_676), .Y(n_1122) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND4xp25_ASAP7_75t_L g690 ( .A(n_691), .B(n_698), .C(n_703), .D(n_711), .Y(n_690) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_701), .C(n_702), .Y(n_698) );
NAND3xp33_ASAP7_75t_L g868 ( .A(n_702), .B(n_869), .C(n_871), .Y(n_868) );
AOI33xp33_ASAP7_75t_L g1124 ( .A1(n_702), .A2(n_1125), .A3(n_1127), .B1(n_1131), .B2(n_1134), .B3(n_1137), .Y(n_1124) );
NAND3xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_707), .C(n_708), .Y(n_703) );
BUFx6f_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g731 ( .A(n_706), .Y(n_731) );
INVx1_ASAP7_75t_L g1100 ( .A(n_706), .Y(n_1100) );
NAND3xp33_ASAP7_75t_L g882 ( .A(n_708), .B(n_883), .C(n_884), .Y(n_882) );
INVx3_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
XNOR2xp5_ASAP7_75t_L g718 ( .A(n_719), .B(n_839), .Y(n_718) );
XOR2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_794), .Y(n_719) );
AND4x1_ASAP7_75t_L g721 ( .A(n_722), .B(n_751), .C(n_757), .D(n_785), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_726), .C(n_750), .Y(n_722) );
NOR3xp33_ASAP7_75t_L g796 ( .A(n_723), .B(n_797), .C(n_814), .Y(n_796) );
AOI221xp5_ASAP7_75t_L g908 ( .A1(n_723), .A2(n_909), .B1(n_910), .B2(n_911), .C(n_912), .Y(n_908) );
AOI221xp5_ASAP7_75t_L g1058 ( .A1(n_723), .A2(n_911), .B1(n_1059), .B2(n_1060), .C(n_1061), .Y(n_1058) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OAI22xp33_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_727) );
INVx2_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
BUFx3_ASAP7_75t_L g1140 ( .A(n_729), .Y(n_1140) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_731), .A2(n_744), .B1(n_812), .B2(n_813), .Y(n_811) );
INVx2_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B1(n_746), .B2(n_748), .Y(n_743) );
INVx2_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_753), .B(n_816), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_753), .B(n_1067), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1184 ( .A(n_753), .B(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1500 ( .A(n_753), .Y(n_1500) );
AND2x2_ASAP7_75t_L g778 ( .A(n_756), .B(n_779), .Y(n_778) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_756), .B(n_779), .Y(n_1090) );
OAI31xp33_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_759), .A3(n_768), .B(n_783), .Y(n_757) );
INVx2_ASAP7_75t_SL g981 ( .A(n_761), .Y(n_981) );
INVx4_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_SL g772 ( .A(n_762), .Y(n_772) );
INVx2_ASAP7_75t_SL g830 ( .A(n_762), .Y(n_830) );
BUFx3_ASAP7_75t_L g986 ( .A(n_762), .Y(n_986) );
INVx2_ASAP7_75t_SL g1072 ( .A(n_762), .Y(n_1072) );
INVx2_ASAP7_75t_SL g1136 ( .A(n_762), .Y(n_1136) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g1204 ( .A(n_765), .Y(n_1204) );
OAI221xp5_ASAP7_75t_L g1201 ( .A1(n_766), .A2(n_1202), .B1(n_1203), .B2(n_1204), .C(n_1205), .Y(n_1201) );
INVx2_ASAP7_75t_L g1489 ( .A(n_767), .Y(n_1489) );
OAI221xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_771), .B1(n_772), .B2(n_773), .C(n_774), .Y(n_769) );
OAI221xp5_ASAP7_75t_L g828 ( .A1(n_770), .A2(n_829), .B1(n_830), .B2(n_831), .C(n_832), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_778), .B1(n_780), .B2(n_781), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_778), .A2(n_781), .B1(n_834), .B2(n_835), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_778), .A2(n_781), .B1(n_1169), .B2(n_1170), .Y(n_1199) );
AOI22xp5_ASAP7_75t_L g1089 ( .A1(n_781), .A2(n_1060), .B1(n_1061), .B2(n_1090), .Y(n_1089) );
CKINVDCx11_ASAP7_75t_R g781 ( .A(n_782), .Y(n_781) );
OAI31xp33_ASAP7_75t_L g817 ( .A1(n_783), .A2(n_818), .A3(n_819), .B(n_827), .Y(n_817) );
OAI21xp5_ASAP7_75t_L g913 ( .A1(n_783), .A2(n_914), .B(n_923), .Y(n_913) );
OAI31xp33_ASAP7_75t_L g1068 ( .A1(n_783), .A2(n_1069), .A3(n_1077), .B(n_1091), .Y(n_1068) );
OAI31xp33_ASAP7_75t_L g1186 ( .A1(n_783), .A2(n_1187), .A3(n_1200), .B(n_1212), .Y(n_1186) );
BUFx8_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_786), .B(n_788), .Y(n_785) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
BUFx2_ASAP7_75t_L g1005 ( .A(n_793), .Y(n_1005) );
AND4x1_ASAP7_75t_L g795 ( .A(n_796), .B(n_815), .C(n_817), .D(n_836), .Y(n_795) );
OAI21xp33_ASAP7_75t_SL g823 ( .A1(n_804), .A2(n_824), .B(n_825), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_807), .B1(n_808), .B2(n_810), .Y(n_805) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g878 ( .A(n_822), .Y(n_878) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
OAI22x1_ASAP7_75t_L g839 ( .A1(n_840), .A2(n_841), .B1(n_893), .B2(n_894), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g892 ( .A(n_843), .Y(n_892) );
NAND3xp33_ASAP7_75t_L g844 ( .A(n_845), .B(n_850), .C(n_853), .Y(n_844) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
NAND4xp25_ASAP7_75t_L g867 ( .A(n_868), .B(n_874), .C(n_882), .D(n_887), .Y(n_867) );
INVx2_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g1040 ( .A(n_881), .Y(n_1040) );
NAND3xp33_ASAP7_75t_L g887 ( .A(n_888), .B(n_889), .C(n_890), .Y(n_887) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx2_ASAP7_75t_SL g893 ( .A(n_894), .Y(n_893) );
INVx2_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
NAND4xp75_ASAP7_75t_L g896 ( .A(n_897), .B(n_913), .C(n_934), .D(n_936), .Y(n_896) );
AND2x2_ASAP7_75t_L g897 ( .A(n_898), .B(n_908), .Y(n_897) );
INVx2_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g1168 ( .A1(n_911), .A2(n_1059), .B1(n_1169), .B2(n_1170), .Y(n_1168) );
AOI22xp5_ASAP7_75t_L g1504 ( .A1(n_911), .A2(n_1505), .B1(n_1506), .B2(n_1507), .Y(n_1504) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_915), .B(n_918), .Y(n_914) );
BUFx3_ASAP7_75t_L g1128 ( .A(n_920), .Y(n_1128) );
NAND2x1p5_ASAP7_75t_L g1479 ( .A(n_932), .B(n_1480), .Y(n_1479) );
INVx2_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
XNOR2xp5_ASAP7_75t_L g940 ( .A(n_941), .B(n_1051), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_943), .A2(n_944), .B1(n_1008), .B2(n_1050), .Y(n_942) );
INVx2_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
NAND4xp25_ASAP7_75t_SL g946 ( .A(n_947), .B(n_950), .C(n_953), .D(n_960), .Y(n_946) );
INVx1_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
BUFx4f_ASAP7_75t_L g1018 ( .A(n_958), .Y(n_1018) );
NAND4xp25_ASAP7_75t_L g1010 ( .A(n_960), .B(n_1011), .C(n_1014), .D(n_1020), .Y(n_1010) );
NAND4xp25_ASAP7_75t_L g1110 ( .A(n_960), .B(n_1111), .C(n_1114), .D(n_1117), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_973), .B(n_990), .Y(n_972) );
BUFx3_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
INVx2_ASAP7_75t_L g1126 ( .A(n_975), .Y(n_1126) );
INVx3_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
INVx2_ASAP7_75t_SL g984 ( .A(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g1210 ( .A(n_986), .Y(n_1210) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
AOI33xp33_ASAP7_75t_L g990 ( .A1(n_991), .A2(n_992), .A3(n_997), .B1(n_1002), .B2(n_1004), .B3(n_1007), .Y(n_990) );
AOI33xp33_ASAP7_75t_L g1171 ( .A1(n_991), .A2(n_1007), .A3(n_1172), .B1(n_1174), .B2(n_1175), .B3(n_1176), .Y(n_1171) );
AOI33xp33_ASAP7_75t_L g1508 ( .A1(n_991), .A2(n_1007), .A3(n_1509), .B1(n_1511), .B2(n_1515), .B3(n_1517), .Y(n_1508) );
BUFx3_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
BUFx2_ASAP7_75t_L g1510 ( .A(n_994), .Y(n_1510) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g1105 ( .A(n_996), .Y(n_1105) );
BUFx3_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx2_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
INVx2_ASAP7_75t_L g1050 ( .A(n_1008), .Y(n_1050) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1009), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1029), .Y(n_1023) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
AOI22xp5_ASAP7_75t_L g1051 ( .A1(n_1052), .A2(n_1053), .B1(n_1162), .B2(n_1213), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
AO22x1_ASAP7_75t_L g1053 ( .A1(n_1054), .A2(n_1107), .B1(n_1160), .B2(n_1161), .Y(n_1053) );
HB1xp67_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1055), .Y(n_1161) );
NAND4xp75_ASAP7_75t_SL g1056 ( .A(n_1057), .B(n_1066), .C(n_1068), .D(n_1094), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1062), .Y(n_1057) );
OAI22xp5_ASAP7_75t_L g1083 ( .A1(n_1063), .A2(n_1084), .B1(n_1086), .B2(n_1088), .Y(n_1083) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
INVx2_ASAP7_75t_SL g1081 ( .A(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1082), .Y(n_1198) );
BUFx2_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
AOI33xp33_ASAP7_75t_L g1094 ( .A1(n_1095), .A2(n_1096), .A3(n_1097), .B1(n_1101), .B2(n_1103), .B3(n_1106), .Y(n_1094) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
INVx2_ASAP7_75t_L g1160 ( .A(n_1107), .Y(n_1160) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1109), .Y(n_1159) );
AOI211x1_ASAP7_75t_L g1109 ( .A1(n_1110), .A2(n_1121), .B(n_1123), .C(n_1150), .Y(n_1109) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1138), .Y(n_1123) );
INVx2_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
HB1xp67_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
BUFx3_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1133), .Y(n_1197) );
BUFx2_ASAP7_75t_L g1486 ( .A(n_1133), .Y(n_1486) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1162), .Y(n_1213) );
HB1xp67_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
AND3x1_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1184), .C(n_1186), .Y(n_1165) );
NOR2xp33_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1177), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1181), .Y(n_1177) );
OAI221xp5_ASAP7_75t_L g1188 ( .A1(n_1179), .A2(n_1183), .B1(n_1189), .B2(n_1191), .C(n_1195), .Y(n_1188) );
BUFx2_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
OAI22xp5_ASAP7_75t_L g1206 ( .A1(n_1207), .A2(n_1208), .B1(n_1209), .B2(n_1210), .Y(n_1206) );
OAI21xp5_ASAP7_75t_L g1215 ( .A1(n_1216), .A2(n_1224), .B(n_1467), .Y(n_1215) );
CKINVDCx5p33_ASAP7_75t_R g1216 ( .A(n_1217), .Y(n_1216) );
BUFx3_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1218), .Y(n_1305) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1218), .Y(n_1323) );
AND2x4_ASAP7_75t_L g1218 ( .A(n_1219), .B(n_1222), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1219), .B(n_1222), .Y(n_1232) );
HB1xp67_ASAP7_75t_L g1535 ( .A(n_1219), .Y(n_1535) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
AND2x4_ASAP7_75t_L g1234 ( .A(n_1220), .B(n_1222), .Y(n_1234) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1221), .B(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1223), .Y(n_1241) );
NOR2x1_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1404), .Y(n_1224) );
NAND3xp33_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1325), .C(n_1364), .Y(n_1225) );
OAI21xp5_ASAP7_75t_L g1226 ( .A1(n_1227), .A2(n_1281), .B(n_1299), .Y(n_1226) );
AOI22xp5_ASAP7_75t_L g1227 ( .A1(n_1228), .A2(n_1259), .B1(n_1275), .B2(n_1277), .Y(n_1227) );
NOR2xp33_ASAP7_75t_L g1390 ( .A(n_1228), .B(n_1285), .Y(n_1390) );
OR2x2_ASAP7_75t_L g1228 ( .A(n_1229), .B(n_1246), .Y(n_1228) );
CKINVDCx6p67_ASAP7_75t_R g1274 ( .A(n_1229), .Y(n_1274) );
OAI222xp33_ASAP7_75t_L g1281 ( .A1(n_1229), .A2(n_1282), .B1(n_1285), .B2(n_1290), .C1(n_1294), .C2(n_1298), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1229), .B(n_1247), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1229), .B(n_1297), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_1229), .B(n_1279), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1229), .B(n_1296), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1229), .B(n_1344), .Y(n_1368) );
OR2x2_ASAP7_75t_L g1388 ( .A(n_1229), .B(n_1297), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1229), .B(n_1267), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1229), .B(n_1403), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1229), .B(n_1371), .Y(n_1410) );
OR2x6_ASAP7_75t_SL g1229 ( .A(n_1230), .B(n_1236), .Y(n_1229) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
OAI22xp5_ASAP7_75t_L g1321 ( .A1(n_1233), .A2(n_1322), .B1(n_1323), .B2(n_1324), .Y(n_1321) );
INVx1_ASAP7_75t_SL g1233 ( .A(n_1234), .Y(n_1233) );
INVx2_ASAP7_75t_L g1273 ( .A(n_1234), .Y(n_1273) );
OAI22xp5_ASAP7_75t_L g1236 ( .A1(n_1237), .A2(n_1242), .B1(n_1243), .B2(n_1245), .Y(n_1236) );
OAI22xp33_ASAP7_75t_L g1263 ( .A1(n_1237), .A2(n_1243), .B1(n_1264), .B2(n_1265), .Y(n_1263) );
BUFx3_ASAP7_75t_L g1309 ( .A(n_1237), .Y(n_1309) );
OAI22xp33_ASAP7_75t_L g1318 ( .A1(n_1237), .A2(n_1312), .B1(n_1319), .B2(n_1320), .Y(n_1318) );
BUFx6f_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
OAI22xp5_ASAP7_75t_L g1256 ( .A1(n_1238), .A2(n_1243), .B1(n_1257), .B2(n_1258), .Y(n_1256) );
OR2x2_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1240), .Y(n_1238) );
OR2x2_ASAP7_75t_L g1243 ( .A(n_1239), .B(n_1244), .Y(n_1243) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1239), .Y(n_1251) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1240), .Y(n_1250) );
HB1xp67_ASAP7_75t_L g1534 ( .A(n_1241), .Y(n_1534) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1243), .Y(n_1313) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1244), .Y(n_1253) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1246), .Y(n_1344) );
OAI221xp5_ASAP7_75t_L g1365 ( .A1(n_1246), .A2(n_1366), .B1(n_1372), .B2(n_1375), .C(n_1377), .Y(n_1365) );
NOR2xp33_ASAP7_75t_L g1403 ( .A(n_1246), .B(n_1280), .Y(n_1403) );
OR2x2_ASAP7_75t_L g1246 ( .A(n_1247), .B(n_1255), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1247), .B(n_1255), .Y(n_1267) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1247), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1247), .B(n_1328), .Y(n_1371) );
NOR2xp33_ASAP7_75t_SL g1442 ( .A(n_1247), .B(n_1443), .Y(n_1442) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1248), .B(n_1254), .Y(n_1247) );
AND2x4_ASAP7_75t_L g1249 ( .A(n_1250), .B(n_1251), .Y(n_1249) );
AND2x4_ASAP7_75t_L g1252 ( .A(n_1251), .B(n_1253), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1255), .B(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1255), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1422 ( .A(n_1255), .B(n_1274), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1260), .B(n_1266), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1453 ( .A(n_1260), .B(n_1408), .Y(n_1453) );
NAND2xp5_ASAP7_75t_L g1459 ( .A(n_1260), .B(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1261), .Y(n_1260) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1261), .Y(n_1276) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1261), .Y(n_1341) );
NAND2xp5_ASAP7_75t_L g1381 ( .A(n_1261), .B(n_1382), .Y(n_1381) );
NAND2xp5_ASAP7_75t_L g1418 ( .A(n_1261), .B(n_1368), .Y(n_1418) );
HB1xp67_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1262), .B(n_1287), .Y(n_1286) );
INVx2_ASAP7_75t_SL g1293 ( .A(n_1262), .Y(n_1293) );
OR2x2_ASAP7_75t_L g1348 ( .A(n_1262), .B(n_1287), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1267), .B(n_1268), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1267), .B(n_1280), .Y(n_1279) );
AOI322xp5_ASAP7_75t_L g1454 ( .A1(n_1267), .A2(n_1315), .A3(n_1328), .B1(n_1354), .B2(n_1431), .C1(n_1455), .C2(n_1456), .Y(n_1454) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1268), .B(n_1296), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1461 ( .A(n_1268), .B(n_1344), .Y(n_1461) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1274), .Y(n_1268) );
INVx4_ASAP7_75t_L g1280 ( .A(n_1269), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1269), .B(n_1292), .Y(n_1291) );
NOR2xp33_ASAP7_75t_L g1345 ( .A(n_1269), .B(n_1274), .Y(n_1345) );
INVx2_ASAP7_75t_L g1361 ( .A(n_1269), .Y(n_1361) );
NAND2xp5_ASAP7_75t_L g1389 ( .A(n_1269), .B(n_1293), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1412 ( .A(n_1269), .B(n_1410), .Y(n_1412) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_1269), .B(n_1317), .Y(n_1431) );
A2O1A1Ixp33_ASAP7_75t_SL g1438 ( .A1(n_1269), .A2(n_1439), .B(n_1440), .C(n_1447), .Y(n_1438) );
NAND2xp5_ASAP7_75t_L g1443 ( .A(n_1269), .B(n_1354), .Y(n_1443) );
OR2x2_ASAP7_75t_L g1446 ( .A(n_1269), .B(n_1362), .Y(n_1446) );
AND2x6_ASAP7_75t_L g1269 ( .A(n_1270), .B(n_1271), .Y(n_1269) );
INVx2_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
OAI22xp5_ASAP7_75t_L g1303 ( .A1(n_1273), .A2(n_1304), .B1(n_1305), .B2(n_1306), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1274), .B(n_1279), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1274), .B(n_1296), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1370 ( .A(n_1274), .B(n_1371), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1274), .B(n_1328), .Y(n_1382) );
NOR3xp33_ASAP7_75t_SL g1423 ( .A(n_1274), .B(n_1280), .C(n_1424), .Y(n_1423) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_1274), .B(n_1328), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1452 ( .A(n_1274), .B(n_1297), .Y(n_1452) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1280), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1330 ( .A(n_1280), .B(n_1292), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1280), .B(n_1332), .Y(n_1331) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_1280), .B(n_1295), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1280), .B(n_1370), .Y(n_1408) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1280), .B(n_1437), .Y(n_1436) );
NAND2xp5_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1284), .Y(n_1282) );
OAI211xp5_ASAP7_75t_L g1391 ( .A1(n_1285), .A2(n_1392), .B(n_1395), .C(n_1399), .Y(n_1391) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1287), .B(n_1293), .Y(n_1292) );
OR2x2_ASAP7_75t_L g1298 ( .A(n_1287), .B(n_1293), .Y(n_1298) );
AOI22xp5_ASAP7_75t_L g1327 ( .A1(n_1287), .A2(n_1328), .B1(n_1329), .B2(n_1331), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1287), .B(n_1317), .Y(n_1339) );
OR2x2_ASAP7_75t_L g1350 ( .A(n_1287), .B(n_1316), .Y(n_1350) );
INVx2_ASAP7_75t_L g1374 ( .A(n_1287), .Y(n_1374) );
NAND2xp5_ASAP7_75t_L g1386 ( .A(n_1287), .B(n_1387), .Y(n_1386) );
OAI21xp5_ASAP7_75t_L g1406 ( .A1(n_1287), .A2(n_1407), .B(n_1409), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1287), .B(n_1316), .Y(n_1417) );
O2A1O1Ixp33_ASAP7_75t_L g1457 ( .A1(n_1287), .A2(n_1401), .B(n_1458), .C(n_1459), .Y(n_1457) );
AND2x4_ASAP7_75t_L g1287 ( .A(n_1288), .B(n_1289), .Y(n_1287) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1292), .B(n_1335), .Y(n_1334) );
NAND2xp5_ASAP7_75t_L g1409 ( .A(n_1292), .B(n_1410), .Y(n_1409) );
INVx2_ASAP7_75t_SL g1354 ( .A(n_1293), .Y(n_1354) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1293), .B(n_1316), .Y(n_1463) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1295), .B(n_1353), .Y(n_1379) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1296), .Y(n_1428) );
INVx2_ASAP7_75t_L g1376 ( .A(n_1298), .Y(n_1376) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_1301), .B(n_1314), .Y(n_1300) );
OAI21xp5_ASAP7_75t_L g1364 ( .A1(n_1301), .A2(n_1365), .B(n_1391), .Y(n_1364) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_1301), .B(n_1374), .Y(n_1414) );
CKINVDCx5p33_ASAP7_75t_R g1301 ( .A(n_1302), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1337 ( .A(n_1302), .B(n_1315), .Y(n_1337) );
AOI221xp5_ASAP7_75t_L g1405 ( .A1(n_1302), .A2(n_1406), .B1(n_1411), .B2(n_1413), .C(n_1415), .Y(n_1405) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1302), .Y(n_1448) );
OR2x6_ASAP7_75t_SL g1302 ( .A(n_1303), .B(n_1307), .Y(n_1302) );
OAI22xp5_ASAP7_75t_L g1307 ( .A1(n_1308), .A2(n_1309), .B1(n_1310), .B2(n_1311), .Y(n_1307) );
HB1xp67_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1357 ( .A(n_1314), .B(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_SL g1314 ( .A(n_1315), .Y(n_1314) );
NOR3xp33_ASAP7_75t_L g1445 ( .A(n_1315), .B(n_1393), .C(n_1446), .Y(n_1445) );
INVx3_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1316), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1425 ( .A(n_1316), .B(n_1374), .Y(n_1425) );
INVx3_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
OR2x2_ASAP7_75t_L g1347 ( .A(n_1317), .B(n_1348), .Y(n_1347) );
OR2x2_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1321), .Y(n_1317) );
XNOR2xp5_ASAP7_75t_L g1471 ( .A(n_1322), .B(n_1472), .Y(n_1471) );
NOR2xp33_ASAP7_75t_L g1325 ( .A(n_1326), .B(n_1349), .Y(n_1325) );
A2O1A1Ixp33_ASAP7_75t_L g1326 ( .A1(n_1327), .A2(n_1333), .B(n_1337), .C(n_1338), .Y(n_1326) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
AOI22xp5_ASAP7_75t_L g1338 ( .A1(n_1331), .A2(n_1339), .B1(n_1340), .B2(n_1346), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1383 ( .A(n_1332), .B(n_1384), .Y(n_1383) );
INVxp67_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1339), .Y(n_1385) );
AND2x2_ASAP7_75t_L g1420 ( .A(n_1339), .B(n_1354), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1341), .B(n_1342), .Y(n_1340) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1342), .Y(n_1464) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1344), .B(n_1345), .Y(n_1343) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1345), .Y(n_1394) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
NOR2xp33_ASAP7_75t_L g1439 ( .A(n_1347), .B(n_1428), .Y(n_1439) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1348), .Y(n_1437) );
A2O1A1Ixp33_ASAP7_75t_L g1349 ( .A1(n_1350), .A2(n_1351), .B(n_1356), .C(n_1357), .Y(n_1349) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1350), .Y(n_1378) );
INVxp67_ASAP7_75t_SL g1351 ( .A(n_1352), .Y(n_1351) );
OAI21xp5_ASAP7_75t_L g1395 ( .A1(n_1352), .A2(n_1396), .B(n_1398), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1353), .B(n_1355), .Y(n_1352) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1354), .Y(n_1362) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1354), .Y(n_1401) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1355), .B(n_1376), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1456 ( .A(n_1355), .B(n_1437), .Y(n_1456) );
OAI22xp5_ASAP7_75t_L g1462 ( .A1(n_1356), .A2(n_1463), .B1(n_1464), .B2(n_1465), .Y(n_1462) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1359), .B(n_1363), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
NOR2xp33_ASAP7_75t_L g1455 ( .A(n_1360), .B(n_1393), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1361), .B(n_1362), .Y(n_1360) );
NOR2xp33_ASAP7_75t_L g1373 ( .A(n_1361), .B(n_1374), .Y(n_1373) );
INVx2_ASAP7_75t_L g1384 ( .A(n_1361), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1421 ( .A(n_1361), .B(n_1422), .Y(n_1421) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1367), .B(n_1369), .Y(n_1366) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1368), .Y(n_1367) );
OAI221xp5_ASAP7_75t_L g1440 ( .A1(n_1369), .A2(n_1416), .B1(n_1424), .B2(n_1441), .C(n_1444), .Y(n_1440) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
OAI21xp5_ASAP7_75t_SL g1433 ( .A1(n_1370), .A2(n_1434), .B(n_1436), .Y(n_1433) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1371), .Y(n_1393) );
INVxp67_ASAP7_75t_SL g1372 ( .A(n_1373), .Y(n_1372) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1374), .Y(n_1466) );
OAI211xp5_ASAP7_75t_L g1450 ( .A1(n_1375), .A2(n_1451), .B(n_1453), .C(n_1454), .Y(n_1450) );
NAND3xp33_ASAP7_75t_L g1430 ( .A(n_1376), .B(n_1431), .C(n_1432), .Y(n_1430) );
AOI211xp5_ASAP7_75t_L g1377 ( .A1(n_1378), .A2(n_1379), .B(n_1380), .C(n_1390), .Y(n_1377) );
A2O1A1Ixp33_ASAP7_75t_L g1380 ( .A1(n_1381), .A2(n_1383), .B(n_1385), .C(n_1386), .Y(n_1380) );
NOR2xp33_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1389), .Y(n_1387) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1388), .Y(n_1432) );
OR2x2_ASAP7_75t_L g1392 ( .A(n_1393), .B(n_1394), .Y(n_1392) );
AND2x2_ASAP7_75t_L g1427 ( .A(n_1393), .B(n_1428), .Y(n_1427) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1398), .Y(n_1458) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
NOR2xp33_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1402), .Y(n_1400) );
NAND3xp33_ASAP7_75t_L g1404 ( .A(n_1405), .B(n_1438), .C(n_1449), .Y(n_1404) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
OAI211xp5_ASAP7_75t_L g1415 ( .A1(n_1416), .A2(n_1418), .B(n_1419), .C(n_1433), .Y(n_1415) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
AOI221xp5_ASAP7_75t_L g1419 ( .A1(n_1420), .A2(n_1421), .B1(n_1423), .B2(n_1426), .C(n_1429), .Y(n_1419) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
INVx1_ASAP7_75t_SL g1429 ( .A(n_1430), .Y(n_1429) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
INVxp67_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1445), .Y(n_1444) );
OAI31xp33_ASAP7_75t_SL g1449 ( .A1(n_1447), .A2(n_1450), .A3(n_1457), .B(n_1462), .Y(n_1449) );
CKINVDCx14_ASAP7_75t_R g1447 ( .A(n_1448), .Y(n_1447) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1469), .Y(n_1468) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
HB1xp67_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
HB1xp67_ASAP7_75t_L g1526 ( .A(n_1472), .Y(n_1526) );
NOR4xp75_ASAP7_75t_L g1472 ( .A(n_1473), .B(n_1492), .C(n_1499), .D(n_1501), .Y(n_1472) );
AOI31xp33_ASAP7_75t_SL g1473 ( .A1(n_1474), .A2(n_1481), .A3(n_1484), .B(n_1490), .Y(n_1473) );
CKINVDCx8_ASAP7_75t_R g1490 ( .A(n_1491), .Y(n_1490) );
NAND2xp5_ASAP7_75t_L g1492 ( .A(n_1493), .B(n_1496), .Y(n_1492) );
NAND3xp33_ASAP7_75t_SL g1501 ( .A(n_1502), .B(n_1504), .C(n_1508), .Y(n_1501) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1503), .Y(n_1502) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1514), .Y(n_1513) );
BUFx2_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
INVxp67_ASAP7_75t_L g1527 ( .A(n_1526), .Y(n_1527) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
CKINVDCx5p33_ASAP7_75t_R g1529 ( .A(n_1530), .Y(n_1529) );
A2O1A1Ixp33_ASAP7_75t_L g1532 ( .A1(n_1531), .A2(n_1533), .B(n_1535), .C(n_1536), .Y(n_1532) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
endmodule