module real_jpeg_4781_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_1),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_1),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_1),
.Y(n_162)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_1),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_1),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_3),
.B(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_3),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_3),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_3),
.B(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_3),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_3),
.B(n_52),
.Y(n_396)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_5),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_5),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_6),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_6),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_6),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_6),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_6),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_6),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_6),
.B(n_377),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_7),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_7),
.B(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_7),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_7),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_7),
.B(n_410),
.Y(n_409)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_8),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_8),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_8),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_8),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_8),
.B(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_8),
.Y(n_250)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_10),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_10),
.Y(n_136)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_10),
.Y(n_173)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_10),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_11),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_11),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_11),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_11),
.B(n_91),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_11),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_11),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_11),
.B(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_12),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_12),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_12),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_12),
.B(n_91),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_12),
.B(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_12),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_12),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_12),
.B(n_356),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_13),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_13),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_13),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_13),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_13),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_13),
.B(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_13),
.Y(n_190)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_14),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_14),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_15),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_15),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_15),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_15),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_15),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_203),
.B1(n_452),
.B2(n_453),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g452 ( 
.A(n_18),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_202),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_164),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_21),
.B(n_164),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_101),
.C(n_138),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_22),
.B(n_335),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_68),
.C(n_81),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_23),
.B(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.C(n_55),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_24),
.B(n_290),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_35),
.B2(n_36),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_27),
.A2(n_28),
.B1(n_106),
.B2(n_107),
.Y(n_307)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_28),
.B(n_31),
.C(n_36),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_28),
.B(n_107),
.C(n_221),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_29),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g348 ( 
.A(n_30),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_31),
.A2(n_34),
.B1(n_110),
.B2(n_114),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_31),
.B(n_110),
.C(n_149),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_31),
.A2(n_34),
.B1(n_362),
.B2(n_363),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

OR2x2_ASAP7_75t_SL g57 ( 
.A(n_32),
.B(n_58),
.Y(n_57)
);

OR2x2_ASAP7_75t_SL g89 ( 
.A(n_32),
.B(n_90),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_32),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_34),
.B(n_362),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_35),
.A2(n_36),
.B1(n_193),
.B2(n_197),
.Y(n_192)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_38),
.Y(n_130)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_38),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_39),
.B(n_55),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_51),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_40),
.B(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_44),
.Y(n_270)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_45),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_45),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_46),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_46),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_46),
.B(n_51),
.Y(n_284)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_49),
.Y(n_123)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_50),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_50),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g382 ( 
.A(n_50),
.Y(n_382)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_60),
.B2(n_67),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_79),
.C(n_80),
.Y(n_78)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_59),
.Y(n_279)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_65),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_68),
.B(n_81),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_78),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_74),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_74),
.B(n_76),
.C(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_74),
.A2(n_77),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_77),
.B(n_158),
.C(n_161),
.Y(n_186)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_95),
.C(n_97),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_83),
.B(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_89),
.C(n_93),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_84),
.A2(n_93),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_84),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_84),
.A2(n_239),
.B1(n_267),
.B2(n_268),
.Y(n_371)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_88),
.Y(n_215)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_88),
.Y(n_228)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_88),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_89),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_89),
.Y(n_235)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_93),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_95),
.B(n_97),
.Y(n_296)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_101),
.B(n_138),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_115),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_102),
.B(n_116),
.C(n_124),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_103),
.B(n_107),
.C(n_110),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_110),
.B2(n_114),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_106),
.A2(n_107),
.B1(n_175),
.B2(n_179),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_109),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_110),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_110),
.B(n_309),
.C(n_313),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_110),
.A2(n_114),
.B1(n_358),
.B2(n_359),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_111),
.Y(n_252)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_111),
.Y(n_412)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_112),
.Y(n_389)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_112),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_124),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.C(n_121),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_117),
.A2(n_143),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_117),
.B(n_175),
.C(n_258),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_121),
.Y(n_144)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_133),
.B2(n_137),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_127),
.B(n_132),
.C(n_133),
.Y(n_183)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g364 ( 
.A(n_129),
.Y(n_364)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_130),
.Y(n_275)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_136),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_154),
.B2(n_163),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_155),
.C(n_157),
.Y(n_165)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_146),
.C(n_147),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_141),
.A2(n_142),
.B1(n_146),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_146),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_147),
.B(n_327),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_152),
.B2(n_153),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_151),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g456 ( 
.A(n_164),
.Y(n_456)
);

FAx1_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_166),
.CI(n_184),
.CON(n_164),
.SN(n_164)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_180),
.B2(n_181),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_174),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_175),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_175),
.A2(n_179),
.B1(n_257),
.B2(n_261),
.Y(n_256)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_178),
.Y(n_353)
);

INVx5_ASAP7_75t_L g370 ( 
.A(n_178),
.Y(n_370)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_191),
.B1(n_192),
.B2(n_198),
.Y(n_187)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_199),
.Y(n_201)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_203),
.Y(n_453)
);

AO21x1_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_333),
.B(n_336),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_322),
.B(n_332),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_299),
.B(n_321),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_206),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_286),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_207),
.B(n_286),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_255),
.C(n_280),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_208),
.B(n_320),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_233),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_209),
.B(n_234),
.C(n_240),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_220),
.C(n_224),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_210),
.B(n_317),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g454 ( 
.A(n_210),
.Y(n_454)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_213),
.CI(n_216),
.CON(n_210),
.SN(n_210)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_211),
.B(n_213),
.C(n_216),
.Y(n_285)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_220),
.A2(n_224),
.B1(n_225),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_220),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_221),
.B(n_307),
.Y(n_306)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_226),
.A2(n_227),
.B1(n_229),
.B2(n_230),
.Y(n_315)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_240),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_248),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_242),
.B(n_244),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_241),
.B(n_249),
.C(n_253),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_247),
.B(n_389),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_254),
.B(n_355),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_254),
.B(n_367),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_254),
.B(n_403),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_255),
.B(n_280),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_262),
.C(n_264),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_256),
.A2(n_262),
.B1(n_263),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_256),
.Y(n_304)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_257),
.Y(n_261)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_258),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_264),
.B(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_271),
.C(n_276),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_265),
.A2(n_266),
.B1(n_439),
.B2(n_440),
.Y(n_438)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_271),
.A2(n_272),
.B1(n_276),
.B2(n_277),
.Y(n_440)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx4_ASAP7_75t_SL g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_285),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_283),
.C(n_285),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_287),
.B(n_289),
.C(n_298),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_291),
.B1(n_297),
.B2(n_298),
.Y(n_288)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_289),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_292),
.B(n_294),
.C(n_295),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_319),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_300),
.B(n_319),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_305),
.C(n_316),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_301),
.A2(n_302),
.B1(n_445),
.B2(n_446),
.Y(n_444)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_305),
.B(n_316),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.C(n_315),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_306),
.B(n_432),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_308),
.B(n_315),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_309),
.A2(n_310),
.B1(n_313),
.B2(n_314),
.Y(n_359)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_312),
.Y(n_356)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_323),
.B(n_333),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_325),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_334),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_325),
.B(n_334),
.Y(n_451)
);

FAx1_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_329),
.CI(n_331),
.CON(n_325),
.SN(n_325)
);

OAI31xp33_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_448),
.A3(n_449),
.B(n_451),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_442),
.B(n_447),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_339),
.A2(n_427),
.B(n_441),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_384),
.B(n_426),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_372),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_341),
.B(n_372),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_360),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_357),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_343),
.B(n_357),
.C(n_360),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_349),
.C(n_354),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_344),
.A2(n_345),
.B1(n_349),
.B2(n_350),
.Y(n_374)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx8_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_354),
.B(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_361),
.B(n_365),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_361),
.B(n_436),
.C(n_437),
.Y(n_435)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_371),
.Y(n_365)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_366),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx5_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_371),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_375),
.C(n_383),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_373),
.B(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_375),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_375),
.A2(n_383),
.B1(n_418),
.B2(n_424),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_380),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_376),
.Y(n_416)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_379),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_380),
.Y(n_417)
);

INVx5_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_383),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_420),
.B(n_425),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_405),
.B(n_419),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_387),
.A2(n_394),
.B(n_404),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_390),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_402),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_402),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_397),
.B(n_401),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_396),
.B(n_397),
.Y(n_401)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_401),
.A2(n_407),
.B1(n_413),
.B2(n_414),
.Y(n_406)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_401),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_415),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_406),
.B(n_415),
.Y(n_419)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_407),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_408),
.A2(n_409),
.B(n_413),
.Y(n_421)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_416),
.A2(n_417),
.B(n_418),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_422),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_421),
.B(n_422),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_428),
.B(n_429),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_431),
.B1(n_433),
.B2(n_434),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_430),
.B(n_435),
.C(n_438),
.Y(n_443)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_438),
.Y(n_434)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_444),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_443),
.B(n_444),
.Y(n_447)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_445),
.Y(n_446)
);


endmodule