module fake_jpeg_31354_n_446 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_446);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_446;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_6),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_9),
.B(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_44),
.B(n_46),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_48),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_47),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_24),
.B(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_49),
.B(n_54),
.Y(n_106)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_50),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_21),
.B(n_18),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_55),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_56),
.B(n_59),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_21),
.B(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_69),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_17),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_27),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_61),
.B(n_66),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_22),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_0),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_42),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_85),
.B(n_25),
.Y(n_96)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_86),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_88),
.Y(n_118)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_25),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_90),
.B(n_94),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_47),
.A2(n_25),
.B1(n_41),
.B2(n_36),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_93),
.A2(n_100),
.B1(n_62),
.B2(n_36),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_45),
.B(n_38),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_73),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_55),
.A2(n_23),
.B1(n_41),
.B2(n_27),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_98),
.A2(n_72),
.B1(n_71),
.B2(n_74),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_50),
.A2(n_41),
.B1(n_36),
.B2(n_23),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

OR2x2_ASAP7_75t_SL g110 ( 
.A(n_69),
.B(n_23),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_52),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_70),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_111),
.B(n_82),
.Y(n_163)
);

NAND2x1_ASAP7_75t_L g121 ( 
.A(n_53),
.B(n_36),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_121),
.B(n_73),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_136),
.B(n_145),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_146),
.Y(n_177)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_139),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_64),
.B1(n_87),
.B2(n_58),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_140),
.A2(n_157),
.B1(n_160),
.B2(n_165),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_92),
.A2(n_51),
.B1(n_78),
.B2(n_65),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_141),
.A2(n_148),
.B1(n_134),
.B2(n_119),
.Y(n_178)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_90),
.A2(n_63),
.B1(n_31),
.B2(n_38),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_115),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_77),
.B1(n_88),
.B2(n_86),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_46),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_150),
.B(n_151),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_34),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_75),
.C(n_76),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_156),
.C(n_101),
.Y(n_190)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_81),
.B1(n_79),
.B2(n_68),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_158),
.A2(n_164),
.B1(n_170),
.B2(n_171),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_84),
.B1(n_67),
.B2(n_34),
.Y(n_160)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_168),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_60),
.B1(n_62),
.B2(n_83),
.Y(n_165)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_167),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_106),
.B(n_129),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_109),
.Y(n_169)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_100),
.A2(n_35),
.B1(n_17),
.B2(n_16),
.Y(n_170)
);

AOI32xp33_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_171),
.A3(n_159),
.B1(n_156),
.B2(n_149),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_93),
.A2(n_35),
.B1(n_15),
.B2(n_14),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_91),
.B(n_80),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_118),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_174),
.B(n_190),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_178),
.A2(n_194),
.B1(n_95),
.B2(n_167),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_114),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_193),
.Y(n_222)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_191),
.Y(n_206)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_136),
.A2(n_148),
.A3(n_159),
.B1(n_141),
.B2(n_145),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_126),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_158),
.A2(n_99),
.B1(n_95),
.B2(n_131),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_196),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_202),
.Y(n_213)
);

INVx3_ASAP7_75t_SL g203 ( 
.A(n_198),
.Y(n_203)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_199),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_204),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_205),
.A2(n_192),
.B1(n_178),
.B2(n_175),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_163),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_208),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_162),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_209),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_161),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_216),
.Y(n_234)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_212),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_174),
.B(n_146),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_215),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_173),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_153),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_120),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_221),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_180),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_224),
.Y(n_251)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_219),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_122),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_180),
.A2(n_154),
.B1(n_143),
.B2(n_195),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_223),
.A2(n_175),
.B(n_176),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_193),
.B(n_121),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_184),
.Y(n_225)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_190),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_230),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_233),
.A2(n_238),
.B1(n_243),
.B2(n_249),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_197),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_222),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_213),
.A2(n_217),
.B1(n_205),
.B2(n_206),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_197),
.B1(n_192),
.B2(n_175),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_239),
.A2(n_215),
.B1(n_216),
.B2(n_227),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_206),
.A2(n_224),
.B(n_214),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_241),
.A2(n_245),
.B(n_223),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_196),
.C(n_187),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_242),
.B(n_250),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_205),
.A2(n_186),
.B1(n_138),
.B2(n_176),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_210),
.A2(n_183),
.B(n_182),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_211),
.A2(n_186),
.B1(n_155),
.B2(n_154),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_208),
.C(n_207),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_251),
.Y(n_252)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_251),
.Y(n_253)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_253),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_231),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_255),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_256),
.B(n_262),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_258),
.A2(n_268),
.B1(n_269),
.B2(n_273),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_227),
.Y(n_259)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_227),
.Y(n_260)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_260),
.Y(n_291)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

AO22x1_ASAP7_75t_SL g263 ( 
.A1(n_238),
.A2(n_248),
.B1(n_228),
.B2(n_241),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_263),
.B(n_266),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_231),
.B(n_220),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_264),
.B(n_248),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_230),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_265),
.B(n_267),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_233),
.A2(n_203),
.B1(n_209),
.B2(n_220),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_230),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_239),
.A2(n_203),
.B1(n_209),
.B2(n_225),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_230),
.A2(n_203),
.B1(n_209),
.B2(n_225),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_234),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_271),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_272),
.B(n_274),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_236),
.A2(n_218),
.B1(n_212),
.B2(n_219),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_218),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_229),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_229),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_279),
.Y(n_281)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_240),
.Y(n_279)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_257),
.A2(n_235),
.B(n_242),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_286),
.A2(n_293),
.B(n_295),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_255),
.B(n_232),
.Y(n_287)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_287),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_254),
.A2(n_261),
.B1(n_277),
.B2(n_270),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_290),
.A2(n_299),
.B1(n_266),
.B2(n_218),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_262),
.A2(n_236),
.B(n_228),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_259),
.A2(n_242),
.B(n_247),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g296 ( 
.A(n_260),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_296),
.B(n_308),
.Y(n_326)
);

NAND2x1_ASAP7_75t_SL g297 ( 
.A(n_263),
.B(n_246),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_298),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_254),
.A2(n_246),
.B1(n_247),
.B2(n_240),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_264),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_300),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_232),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_301),
.B(n_302),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_183),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_243),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_273),
.Y(n_313)
);

OAI32xp33_ASAP7_75t_L g306 ( 
.A1(n_252),
.A2(n_244),
.A3(n_181),
.B1(n_189),
.B2(n_201),
.Y(n_306)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_306),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_274),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_283),
.B(n_275),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_311),
.B(n_313),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_277),
.C(n_256),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_316),
.C(n_318),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_292),
.B(n_253),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_300),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_258),
.C(n_268),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_279),
.Y(n_317)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_317),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_278),
.C(n_276),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_298),
.A2(n_247),
.B1(n_244),
.B2(n_212),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_320),
.A2(n_284),
.B1(n_281),
.B2(n_291),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_322),
.A2(n_307),
.B1(n_297),
.B2(n_289),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_181),
.C(n_189),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_323),
.B(n_288),
.C(n_280),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_294),
.B(n_219),
.Y(n_324)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_324),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_293),
.A2(n_226),
.B(n_130),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_286),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_283),
.B(n_103),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_318),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_201),
.Y(n_329)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_329),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_303),
.A2(n_179),
.B1(n_144),
.B2(n_155),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_331),
.A2(n_285),
.B1(n_307),
.B2(n_289),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_285),
.A2(n_144),
.B1(n_143),
.B2(n_139),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_334),
.A2(n_299),
.B1(n_290),
.B2(n_291),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_335),
.B(n_351),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_340),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_341),
.A2(n_343),
.B1(n_348),
.B2(n_327),
.Y(n_363)
);

OAI31xp33_ASAP7_75t_L g342 ( 
.A1(n_319),
.A2(n_303),
.A3(n_297),
.B(n_304),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_342),
.B(n_344),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_321),
.B(n_282),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_345),
.B(n_352),
.Y(n_365)
);

XNOR2x1_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_349),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_333),
.A2(n_288),
.B1(n_280),
.B2(n_304),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_350),
.B(n_357),
.C(n_358),
.Y(n_362)
);

XNOR2x1_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_306),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_312),
.A2(n_226),
.B(n_123),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_332),
.A2(n_169),
.B1(n_124),
.B2(n_133),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_355),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_310),
.B(n_166),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_354),
.B(n_324),
.Y(n_374)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_317),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_333),
.A2(n_124),
.B1(n_133),
.B2(n_131),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_356),
.B(n_357),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_323),
.B(n_115),
.C(n_101),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_313),
.B(n_226),
.C(n_108),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_338),
.B(n_326),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_359),
.B(n_363),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_348),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_361),
.B(n_378),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_366),
.A2(n_337),
.B1(n_339),
.B2(n_343),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_338),
.B(n_316),
.Y(n_367)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_350),
.B(n_314),
.Y(n_368)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_368),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_336),
.B(n_330),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_369),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_310),
.C(n_311),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_372),
.B(n_376),
.C(n_347),
.Y(n_380)
);

OAI32xp33_ASAP7_75t_L g373 ( 
.A1(n_342),
.A2(n_312),
.A3(n_327),
.B1(n_322),
.B2(n_325),
.Y(n_373)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_373),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_374),
.B(n_375),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_347),
.B(n_334),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_329),
.C(n_331),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_344),
.B(n_14),
.Y(n_377)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_377),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_341),
.A2(n_130),
.B1(n_127),
.B2(n_108),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_380),
.B(n_383),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_362),
.B(n_335),
.C(n_354),
.Y(n_383)
);

BUFx4f_ASAP7_75t_SL g385 ( 
.A(n_373),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_385),
.B(n_379),
.Y(n_397)
);

NOR2xp67_ASAP7_75t_SL g387 ( 
.A(n_364),
.B(n_351),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_387),
.A2(n_392),
.B(n_389),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_390),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_362),
.B(n_352),
.C(n_166),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_364),
.B(n_166),
.C(n_127),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_395),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_370),
.B(n_372),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_125),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_396),
.B(n_374),
.Y(n_401)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_397),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_379),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_401),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_384),
.A2(n_360),
.B1(n_365),
.B2(n_375),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_399),
.B(n_402),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_381),
.B(n_376),
.C(n_370),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_405),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_166),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_116),
.C(n_97),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_386),
.A2(n_125),
.B(n_116),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_385),
.B(n_97),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_407),
.B(n_408),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_383),
.B(n_390),
.C(n_391),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_393),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_410),
.B(n_415),
.C(n_1),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_398),
.B(n_394),
.Y(n_411)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_411),
.Y(n_425)
);

BUFx24_ASAP7_75t_SL g414 ( 
.A(n_400),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_414),
.B(n_417),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_385),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_397),
.A2(n_396),
.B1(n_14),
.B2(n_11),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_420),
.B(n_35),
.Y(n_423)
);

AOI321xp33_ASAP7_75t_L g421 ( 
.A1(n_406),
.A2(n_104),
.A3(n_97),
.B1(n_35),
.B2(n_4),
.C(n_5),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_421),
.A2(n_2),
.B(n_3),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_412),
.A2(n_104),
.B(n_2),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_422),
.A2(n_3),
.B(n_4),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_423),
.B(n_429),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_416),
.B(n_1),
.Y(n_424)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_424),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_418),
.B(n_1),
.Y(n_426)
);

AO21x1_ASAP7_75t_L g431 ( 
.A1(n_426),
.A2(n_427),
.B(n_3),
.Y(n_431)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_413),
.A2(n_1),
.B(n_2),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_430),
.B(n_415),
.Y(n_435)
);

NAND3xp33_ASAP7_75t_L g439 ( 
.A(n_431),
.B(n_435),
.C(n_4),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_425),
.B(n_410),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_434),
.A2(n_432),
.B(n_5),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_436),
.A2(n_424),
.B(n_5),
.Y(n_438)
);

NOR3xp33_ASAP7_75t_SL g437 ( 
.A(n_433),
.B(n_419),
.C(n_428),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_437),
.A2(n_4),
.B(n_6),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_438),
.A2(n_439),
.B(n_440),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_441),
.B(n_8),
.C(n_6),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_443),
.A2(n_442),
.B1(n_7),
.B2(n_8),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_444),
.B(n_7),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_445),
.A2(n_8),
.B(n_412),
.Y(n_446)
);


endmodule