module fake_jpeg_544_n_219 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_219);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_24),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_25),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_30),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_10),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

BUFx4f_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_84),
.B(n_87),
.Y(n_88)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_54),
.B1(n_65),
.B2(n_62),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_94),
.B1(n_75),
.B2(n_77),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_58),
.B1(n_68),
.B2(n_62),
.Y(n_93)
);

BUFx4f_ASAP7_75t_SL g107 ( 
.A(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_68),
.B1(n_59),
.B2(n_74),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_55),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_61),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_80),
.Y(n_101)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_109),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_73),
.B1(n_74),
.B2(n_59),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_104),
.B1(n_108),
.B2(n_111),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_82),
.B1(n_81),
.B2(n_78),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_105),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_70),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_84),
.B1(n_67),
.B2(n_73),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_75),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NOR2x1_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_100),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_115),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_117),
.Y(n_137)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_56),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_60),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_21),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_109),
.A2(n_99),
.B1(n_89),
.B2(n_86),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_89),
.C(n_71),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_125),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_141),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_76),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_77),
.B1(n_66),
.B2(n_69),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_126),
.A2(n_107),
.B1(n_72),
.B2(n_2),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_136),
.B(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_113),
.B(n_0),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_152),
.B1(n_164),
.B2(n_143),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_137),
.B(n_0),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_144),
.B(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_134),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_1),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_150),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_SL g150 ( 
.A(n_131),
.B(n_107),
.C(n_22),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_128),
.A2(n_107),
.B1(n_2),
.B2(n_3),
.Y(n_152)
);

AOI32xp33_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_1),
.A3(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_12),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_4),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_160),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_157),
.B1(n_13),
.B2(n_14),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_28),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_163),
.C(n_33),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_129),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_165),
.Y(n_180)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_32),
.C(n_50),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_29),
.B(n_49),
.Y(n_164)
);

NOR2x1_ASAP7_75t_SL g183 ( 
.A(n_164),
.B(n_35),
.Y(n_183)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_159),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_171),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_139),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_169),
.B(n_173),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_149),
.B1(n_150),
.B2(n_18),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_26),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_174),
.A2(n_175),
.B1(n_181),
.B2(n_184),
.Y(n_190)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_176),
.B(n_16),
.CI(n_17),
.CON(n_192),
.SN(n_192)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_23),
.C(n_48),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_179),
.B(n_46),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_148),
.B(n_15),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_182),
.A2(n_183),
.B(n_40),
.Y(n_191)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_188),
.B1(n_193),
.B2(n_179),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_175),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_192),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_170),
.A2(n_19),
.B1(n_34),
.B2(n_43),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_176),
.Y(n_199)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_185),
.B(n_169),
.CI(n_168),
.CON(n_196),
.SN(n_196)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_199),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_202),
.B1(n_190),
.B2(n_187),
.Y(n_205)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g200 ( 
.A(n_195),
.B(n_180),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_201),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_178),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_202),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_205),
.A2(n_196),
.B1(n_186),
.B2(n_203),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_201),
.C(n_200),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_209),
.B(n_210),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_208),
.A2(n_177),
.B1(n_172),
.B2(n_183),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_204),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_209),
.C(n_207),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_206),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_216),
.A2(n_212),
.B(n_166),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_194),
.C(n_51),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_192),
.Y(n_219)
);


endmodule