module fake_jpeg_13491_n_645 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_645);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_645;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_519;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_378;
wire n_133;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx8_ASAP7_75t_SL g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_8),
.B(n_0),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_13),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_61),
.Y(n_152)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g171 ( 
.A(n_62),
.Y(n_171)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_64),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_69),
.B(n_72),
.Y(n_132)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_71),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_31),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_73),
.Y(n_172)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_75),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_76),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_37),
.B(n_9),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_78),
.B(n_79),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_22),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_80),
.Y(n_181)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_9),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_82),
.B(n_83),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_9),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_84),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_21),
.B(n_8),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_85),
.B(n_91),
.Y(n_155)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_87),
.Y(n_207)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_88),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_89),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_21),
.B(n_8),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_95),
.Y(n_188)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_96),
.Y(n_190)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_100),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_19),
.Y(n_101)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_102),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_19),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_103),
.B(n_105),
.Y(n_160)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_47),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_106),
.B(n_107),
.Y(n_170)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_28),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_19),
.Y(n_116)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_117),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_19),
.Y(n_118)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_19),
.Y(n_119)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_119),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_34),
.B(n_8),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_120),
.B(n_56),
.Y(n_196)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_41),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g186 ( 
.A(n_121),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_18),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_18),
.Y(n_123)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_18),
.Y(n_124)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_26),
.Y(n_125)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_125),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_90),
.A2(n_44),
.B1(n_35),
.B2(n_26),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_129),
.A2(n_149),
.B1(n_51),
.B2(n_49),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_115),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_130),
.B(n_131),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_62),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_65),
.A2(n_35),
.B1(n_29),
.B2(n_20),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_142),
.A2(n_145),
.B1(n_49),
.B2(n_55),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_71),
.A2(n_34),
.B1(n_45),
.B2(n_56),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_78),
.B(n_124),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_148),
.B(n_193),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_67),
.A2(n_27),
.B1(n_58),
.B2(n_38),
.Y(n_149)
);

BUFx10_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

INVxp67_ASAP7_75t_SL g226 ( 
.A(n_154),
.Y(n_226)
);

INVx5_ASAP7_75t_SL g158 ( 
.A(n_66),
.Y(n_158)
);

BUFx2_ASAP7_75t_R g238 ( 
.A(n_158),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_64),
.B(n_57),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_166),
.B(n_169),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_93),
.B(n_57),
.Y(n_169)
);

BUFx8_ASAP7_75t_L g177 ( 
.A(n_101),
.Y(n_177)
);

INVx13_ASAP7_75t_L g264 ( 
.A(n_177),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_123),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_196),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_61),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_182),
.B(n_189),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_77),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_187),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_121),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_122),
.B(n_26),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_75),
.B(n_45),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_194),
.B(n_27),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_89),
.Y(n_195)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_195),
.Y(n_259)
);

INVx4_ASAP7_75t_SL g197 ( 
.A(n_116),
.Y(n_197)
);

INVx11_ASAP7_75t_L g250 ( 
.A(n_197),
.Y(n_250)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_118),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_119),
.Y(n_202)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_209),
.Y(n_288)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_152),
.Y(n_211)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_211),
.Y(n_285)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_156),
.Y(n_213)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_213),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_148),
.B(n_51),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_214),
.B(n_223),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_215),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_186),
.A2(n_39),
.B1(n_52),
.B2(n_36),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_216),
.A2(n_224),
.B1(n_233),
.B2(n_253),
.Y(n_322)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_149),
.A2(n_87),
.B1(n_112),
.B2(n_98),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_217),
.A2(n_234),
.B1(n_241),
.B2(n_246),
.Y(n_298)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_136),
.Y(n_218)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_218),
.Y(n_286)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_127),
.Y(n_221)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_221),
.Y(n_287)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_126),
.Y(n_222)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_222),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_138),
.B(n_38),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_186),
.A2(n_36),
.B1(n_52),
.B2(n_39),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_143),
.Y(n_225)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_225),
.Y(n_309)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_128),
.Y(n_227)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_227),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_138),
.A2(n_32),
.B(n_20),
.C(n_29),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_228),
.B(n_230),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_229),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_170),
.B(n_58),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_146),
.Y(n_231)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_231),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_160),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_162),
.A2(n_76),
.B1(n_84),
.B2(n_94),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_142),
.A2(n_32),
.B1(n_55),
.B2(n_46),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_163),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_235),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_236),
.B(n_249),
.Y(n_307)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_162),
.Y(n_237)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_206),
.Y(n_240)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_240),
.Y(n_320)
);

OR2x2_ASAP7_75t_SL g242 ( 
.A(n_150),
.B(n_40),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_242),
.B(n_267),
.Y(n_295)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_147),
.Y(n_243)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_243),
.Y(n_297)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_150),
.A2(n_104),
.B1(n_92),
.B2(n_117),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_175),
.Y(n_247)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_247),
.Y(n_313)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_188),
.Y(n_248)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_248),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_170),
.B(n_132),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_251),
.A2(n_185),
.B1(n_161),
.B2(n_176),
.Y(n_291)
);

CKINVDCx12_ASAP7_75t_R g252 ( 
.A(n_171),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_252),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_190),
.A2(n_46),
.B1(n_26),
.B2(n_40),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_155),
.B(n_26),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_254),
.B(n_261),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_132),
.B(n_155),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_256),
.B(n_257),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_160),
.B(n_178),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_159),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_258),
.B(n_268),
.Y(n_319)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_167),
.Y(n_260)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_260),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_192),
.B(n_0),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_140),
.A2(n_40),
.B1(n_43),
.B2(n_5),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_262),
.A2(n_263),
.B1(n_280),
.B2(n_195),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_144),
.A2(n_204),
.B1(n_135),
.B2(n_134),
.Y(n_263)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_159),
.Y(n_265)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_265),
.Y(n_327)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_168),
.Y(n_266)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_266),
.Y(n_330)
);

OR2x6_ASAP7_75t_SL g267 ( 
.A(n_187),
.B(n_43),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_137),
.B(n_3),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_157),
.Y(n_269)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_269),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_207),
.Y(n_270)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_270),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_193),
.B(n_3),
.Y(n_271)
);

XNOR2x1_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_180),
.Y(n_292)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_191),
.Y(n_272)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_272),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_141),
.B(n_4),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_273),
.B(n_276),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_L g274 ( 
.A1(n_129),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_274),
.A2(n_165),
.B1(n_205),
.B2(n_179),
.Y(n_341)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_136),
.Y(n_275)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_275),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_173),
.Y(n_276)
);

INVx11_ASAP7_75t_L g277 ( 
.A(n_154),
.Y(n_277)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_277),
.Y(n_303)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_207),
.Y(n_278)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_278),
.Y(n_337)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_173),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_279),
.B(n_281),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_151),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_280)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_161),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_187),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_282),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_251),
.A2(n_174),
.B1(n_164),
.B2(n_176),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_289),
.A2(n_291),
.B1(n_299),
.B2(n_314),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_212),
.B(n_172),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_290),
.B(n_304),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_292),
.B(n_264),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_214),
.A2(n_254),
.B1(n_232),
.B2(n_271),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_261),
.B(n_199),
.Y(n_304)
);

BUFx8_ASAP7_75t_L g305 ( 
.A(n_250),
.Y(n_305)
);

INVx6_ASAP7_75t_SL g370 ( 
.A(n_305),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_219),
.B(n_181),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_311),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_223),
.A2(n_185),
.B1(n_200),
.B2(n_184),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_222),
.B(n_153),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_316),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_225),
.B(n_197),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_323),
.B(n_335),
.C(n_338),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_250),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_328),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_267),
.Y(n_328)
);

NAND2xp33_ASAP7_75t_SL g333 ( 
.A(n_246),
.B(n_267),
.Y(n_333)
);

NAND2xp33_ASAP7_75t_SL g347 ( 
.A(n_333),
.B(n_341),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_242),
.B(n_230),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_231),
.B(n_235),
.Y(n_338)
);

AO21x2_ASAP7_75t_L g340 ( 
.A1(n_274),
.A2(n_154),
.B(n_139),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_340),
.A2(n_259),
.B1(n_277),
.B2(n_239),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_342),
.A2(n_226),
.B1(n_278),
.B2(n_240),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_312),
.B(n_208),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_344),
.B(n_346),
.Y(n_412)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_313),
.Y(n_345)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_345),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_307),
.B(n_255),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_283),
.B(n_220),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_348),
.B(n_354),
.Y(n_413)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_320),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_350),
.Y(n_418)
);

OR2x2_ASAP7_75t_SL g351 ( 
.A(n_335),
.B(n_228),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_351),
.Y(n_393)
);

INVx8_ASAP7_75t_L g352 ( 
.A(n_303),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_352),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_334),
.B(n_247),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_353),
.B(n_366),
.C(n_325),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_321),
.B(n_237),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_338),
.Y(n_356)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_356),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_357),
.Y(n_401)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_296),
.Y(n_358)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_358),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_334),
.B(n_245),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_359),
.B(n_365),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_302),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_361),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_299),
.B(n_213),
.Y(n_361)
);

AND2x2_ASAP7_75t_SL g362 ( 
.A(n_295),
.B(n_238),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_362),
.B(n_376),
.Y(n_396)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_338),
.Y(n_363)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_363),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_310),
.B(n_265),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_292),
.B(n_238),
.C(n_244),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_304),
.B(n_260),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_371),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_319),
.B(n_211),
.Y(n_368)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_368),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_304),
.B(n_210),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_311),
.B(n_266),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_372),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_295),
.A2(n_272),
.B(n_239),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_373),
.A2(n_389),
.B(n_326),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_331),
.B(n_210),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_374),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_375),
.A2(n_340),
.B1(n_303),
.B2(n_323),
.Y(n_403)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_320),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_289),
.A2(n_281),
.B1(n_275),
.B2(n_218),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_378),
.A2(n_385),
.B1(n_340),
.B2(n_337),
.Y(n_416)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_327),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_379),
.B(n_388),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_298),
.A2(n_270),
.B1(n_215),
.B2(n_229),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_380),
.A2(n_383),
.B1(n_386),
.B2(n_375),
.Y(n_414)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_300),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_381),
.B(n_384),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_290),
.A2(n_239),
.B1(n_259),
.B2(n_269),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_382),
.A2(n_341),
.B(n_316),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_298),
.A2(n_209),
.B1(n_183),
.B2(n_165),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_339),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_333),
.A2(n_239),
.B1(n_177),
.B2(n_157),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_331),
.A2(n_264),
.B1(n_171),
.B2(n_133),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_387),
.B(n_323),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_316),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_290),
.A2(n_5),
.B(n_11),
.Y(n_389)
);

OAI21xp33_ASAP7_75t_SL g391 ( 
.A1(n_362),
.A2(n_294),
.B(n_322),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_391),
.A2(n_416),
.B1(n_362),
.B2(n_369),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_353),
.B(n_311),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_392),
.B(n_400),
.C(n_402),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_297),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_349),
.B(n_293),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_403),
.A2(n_426),
.B1(n_382),
.B2(n_385),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_406),
.B(n_409),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_407),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_370),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_408),
.B(n_427),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_347),
.A2(n_340),
.B(n_326),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_410),
.A2(n_411),
.B(n_347),
.Y(n_441)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_414),
.Y(n_430)
);

OAI32xp33_ASAP7_75t_L g417 ( 
.A1(n_361),
.A2(n_340),
.A3(n_287),
.B1(n_318),
.B2(n_330),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_417),
.B(n_419),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_359),
.B(n_365),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_368),
.B(n_308),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_360),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_364),
.A2(n_336),
.B1(n_286),
.B2(n_329),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_421),
.A2(n_425),
.B1(n_383),
.B2(n_352),
.Y(n_442)
);

AND2x2_ASAP7_75t_SL g424 ( 
.A(n_366),
.B(n_305),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_424),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_364),
.A2(n_336),
.B1(n_286),
.B2(n_329),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_380),
.A2(n_288),
.B1(n_315),
.B2(n_306),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_370),
.Y(n_427)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_415),
.Y(n_432)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_432),
.Y(n_470)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_429),
.Y(n_433)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_433),
.Y(n_474)
);

AND2x6_ASAP7_75t_L g435 ( 
.A(n_393),
.B(n_351),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_435),
.A2(n_441),
.B(n_448),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_412),
.B(n_346),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_436),
.B(n_437),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_405),
.B(n_374),
.Y(n_437)
);

INVx13_ASAP7_75t_L g438 ( 
.A(n_418),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_438),
.Y(n_469)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_440),
.Y(n_487)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_442),
.Y(n_496)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_429),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_443),
.Y(n_492)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_429),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_444),
.B(n_446),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_394),
.B(n_420),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_445),
.B(n_447),
.Y(n_483)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_404),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_394),
.B(n_384),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_451),
.B(n_454),
.Y(n_491)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_404),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_452),
.B(n_456),
.Y(n_489)
);

AND2x6_ASAP7_75t_L g454 ( 
.A(n_393),
.B(n_362),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_386),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_455),
.B(n_457),
.Y(n_486)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_398),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_423),
.B(n_369),
.Y(n_457)
);

INVx6_ASAP7_75t_SL g458 ( 
.A(n_395),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_458),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_SL g459 ( 
.A(n_396),
.B(n_377),
.C(n_349),
.Y(n_459)
);

AOI322xp5_ASAP7_75t_SL g479 ( 
.A1(n_459),
.A2(n_343),
.A3(n_371),
.B1(n_367),
.B2(n_396),
.C1(n_406),
.C2(n_392),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_403),
.A2(n_373),
.B1(n_343),
.B2(n_388),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_460),
.B(n_463),
.Y(n_497)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_398),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_461),
.B(n_462),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_397),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_397),
.B(n_345),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_428),
.B(n_284),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_464),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_419),
.B(n_363),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_465),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_399),
.B(n_356),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_466),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_434),
.B(n_402),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_467),
.B(n_472),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_434),
.B(n_409),
.C(n_424),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_468),
.B(n_481),
.C(n_482),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_441),
.A2(n_411),
.B(n_396),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_471),
.A2(n_449),
.B(n_460),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_450),
.B(n_400),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_430),
.A2(n_414),
.B1(n_410),
.B2(n_401),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_475),
.B(n_494),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_450),
.B(n_424),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_476),
.B(n_466),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_479),
.B(n_480),
.Y(n_526)
);

HAxp5_ASAP7_75t_SL g480 ( 
.A(n_458),
.B(n_401),
.CON(n_480),
.SN(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_422),
.C(n_399),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_422),
.C(n_377),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_433),
.B(n_377),
.C(n_423),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_490),
.B(n_443),
.C(n_444),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_430),
.A2(n_426),
.B1(n_417),
.B2(n_416),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_437),
.B(n_436),
.Y(n_495)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_495),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_462),
.B(n_418),
.Y(n_498)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_498),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_439),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_486),
.Y(n_515)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_473),
.Y(n_502)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_502),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_477),
.Y(n_505)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_505),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_SL g506 ( 
.A(n_476),
.B(n_465),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_506),
.B(n_508),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_SL g508 ( 
.A(n_467),
.B(n_435),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_509),
.B(n_513),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_510),
.A2(n_524),
.B(n_527),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_495),
.A2(n_431),
.B1(n_447),
.B2(n_442),
.Y(n_512)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_512),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_472),
.B(n_448),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_473),
.Y(n_514)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_514),
.Y(n_541)
);

AOI31xp33_ASAP7_75t_L g542 ( 
.A1(n_515),
.A2(n_531),
.A3(n_483),
.B(n_474),
.Y(n_542)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_493),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_516),
.B(n_517),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_471),
.A2(n_449),
.B(n_431),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_518),
.B(n_519),
.C(n_481),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_468),
.B(n_461),
.C(n_456),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_493),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_520),
.B(n_521),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_491),
.A2(n_457),
.B(n_445),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_498),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_522),
.B(n_523),
.Y(n_555)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_489),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_491),
.A2(n_454),
.B(n_440),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_478),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_525),
.B(n_529),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_497),
.A2(n_463),
.B(n_451),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_489),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_528),
.Y(n_550)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_470),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_470),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_530),
.A2(n_469),
.B1(n_478),
.B2(n_446),
.Y(n_556)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_487),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_533),
.B(n_538),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_507),
.B(n_490),
.C(n_492),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_534),
.B(n_546),
.C(n_510),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_504),
.A2(n_497),
.B1(n_496),
.B2(n_488),
.Y(n_537)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_537),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_507),
.B(n_499),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_518),
.B(n_499),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_540),
.B(n_557),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_542),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_524),
.A2(n_474),
.B(n_492),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g569 ( 
.A1(n_545),
.A2(n_527),
.B(n_517),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_519),
.B(n_492),
.C(n_482),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_504),
.A2(n_496),
.B1(n_494),
.B2(n_475),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_548),
.A2(n_554),
.B1(n_541),
.B2(n_553),
.Y(n_575)
);

CKINVDCx14_ASAP7_75t_R g549 ( 
.A(n_526),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_549),
.B(n_503),
.Y(n_579)
);

AOI21xp33_ASAP7_75t_L g552 ( 
.A1(n_521),
.A2(n_484),
.B(n_486),
.Y(n_552)
);

OA21x2_ASAP7_75t_SL g566 ( 
.A1(n_552),
.A2(n_501),
.B(n_483),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_516),
.A2(n_488),
.B1(n_485),
.B2(n_487),
.Y(n_554)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_556),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_509),
.B(n_506),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_559),
.B(n_567),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_550),
.B(n_484),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_560),
.B(n_563),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_547),
.Y(n_562)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_562),
.Y(n_585)
);

OAI32xp33_ASAP7_75t_L g563 ( 
.A1(n_551),
.A2(n_511),
.A3(n_520),
.B1(n_531),
.B2(n_502),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_566),
.A2(n_577),
.B1(n_579),
.B2(n_555),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_534),
.B(n_503),
.C(n_513),
.Y(n_567)
);

CKINVDCx16_ASAP7_75t_R g568 ( 
.A(n_544),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_568),
.B(n_576),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_569),
.A2(n_573),
.B(n_355),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_533),
.B(n_546),
.C(n_557),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_570),
.B(n_532),
.C(n_540),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_SL g572 ( 
.A(n_536),
.B(n_508),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_572),
.B(n_532),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_543),
.A2(n_485),
.B(n_514),
.Y(n_573)
);

BUFx12_ASAP7_75t_L g574 ( 
.A(n_556),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_574),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_575),
.A2(n_578),
.B1(n_537),
.B2(n_541),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_548),
.A2(n_500),
.B1(n_525),
.B2(n_530),
.Y(n_576)
);

INVx13_ASAP7_75t_L g577 ( 
.A(n_545),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_554),
.A2(n_530),
.B1(n_469),
.B2(n_432),
.Y(n_578)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_581),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_571),
.A2(n_543),
.B1(n_535),
.B2(n_539),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_582),
.B(n_583),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_559),
.B(n_538),
.Y(n_583)
);

OAI22xp33_ASAP7_75t_SL g604 ( 
.A1(n_586),
.A2(n_574),
.B1(n_563),
.B2(n_378),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_564),
.A2(n_558),
.B1(n_579),
.B2(n_571),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_587),
.A2(n_591),
.B1(n_352),
.B2(n_379),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_588),
.B(n_593),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_589),
.B(n_592),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_558),
.A2(n_544),
.B1(n_536),
.B2(n_425),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_573),
.A2(n_452),
.B1(n_390),
.B2(n_421),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_561),
.B(n_390),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_561),
.B(n_407),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_595),
.B(n_596),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_570),
.B(n_418),
.C(n_376),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_597),
.B(n_389),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_583),
.B(n_565),
.C(n_567),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_598),
.B(n_601),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_SL g599 ( 
.A(n_580),
.B(n_565),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_SL g623 ( 
.A(n_599),
.B(n_610),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_589),
.B(n_564),
.C(n_569),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_596),
.B(n_572),
.C(n_577),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_602),
.B(n_603),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_586),
.B(n_574),
.C(n_562),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_604),
.A2(n_611),
.B1(n_591),
.B2(n_595),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_593),
.B(n_350),
.C(n_438),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_606),
.B(n_585),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_SL g610 ( 
.A(n_582),
.B(n_381),
.Y(n_610)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_612),
.Y(n_621)
);

AOI21xp33_ASAP7_75t_L g613 ( 
.A1(n_609),
.A2(n_594),
.B(n_584),
.Y(n_613)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_613),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_615),
.B(n_617),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_SL g616 ( 
.A1(n_601),
.A2(n_587),
.B1(n_597),
.B2(n_590),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g625 ( 
.A(n_616),
.B(n_602),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_607),
.B(n_588),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_618),
.B(n_317),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_600),
.A2(n_358),
.B1(n_315),
.B2(n_288),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_619),
.B(n_620),
.Y(n_631)
);

A2O1A1Ixp33_ASAP7_75t_SL g620 ( 
.A1(n_604),
.A2(n_306),
.B(n_305),
.C(n_332),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_L g624 ( 
.A1(n_614),
.A2(n_598),
.B(n_603),
.Y(n_624)
);

AO21x1_ASAP7_75t_L g632 ( 
.A1(n_624),
.A2(n_626),
.B(n_622),
.Y(n_632)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_625),
.Y(n_634)
);

AOI322xp5_ASAP7_75t_L g626 ( 
.A1(n_623),
.A2(n_608),
.A3(n_605),
.B1(n_606),
.B2(n_285),
.C1(n_308),
.C2(n_309),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_627),
.B(n_628),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_SL g628 ( 
.A(n_621),
.B(n_317),
.Y(n_628)
);

A2O1A1Ixp33_ASAP7_75t_SL g637 ( 
.A1(n_632),
.A2(n_633),
.B(n_629),
.C(n_631),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g633 ( 
.A1(n_630),
.A2(n_613),
.B(n_620),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_629),
.Y(n_635)
);

AOI322xp5_ASAP7_75t_L g639 ( 
.A1(n_635),
.A2(n_285),
.A3(n_301),
.B1(n_15),
.B2(n_16),
.C1(n_12),
.C2(n_13),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_SL g641 ( 
.A1(n_637),
.A2(n_639),
.B(n_15),
.Y(n_641)
);

AOI31xp33_ASAP7_75t_SL g638 ( 
.A1(n_634),
.A2(n_620),
.A3(n_309),
.B(n_301),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_638),
.A2(n_636),
.B(n_15),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_SL g642 ( 
.A(n_640),
.B(n_641),
.Y(n_642)
);

XNOR2xp5_ASAP7_75t_L g643 ( 
.A(n_642),
.B(n_15),
.Y(n_643)
);

INVxp33_ASAP7_75t_L g644 ( 
.A(n_643),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_L g645 ( 
.A(n_644),
.B(n_16),
.Y(n_645)
);


endmodule