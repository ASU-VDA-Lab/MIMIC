module real_jpeg_18105_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_22),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_1),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_1),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_1),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_1),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_1),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_1),
.B(n_256),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_1),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_1),
.B(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_2),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_2),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_3),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_3),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_4),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_4),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_4),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_4),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_4),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_4),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_4),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_4),
.B(n_89),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_5),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_5),
.B(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_5),
.A2(n_13),
.B1(n_120),
.B2(n_123),
.Y(n_119)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_5),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_5),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_5),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_5),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_6),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_6),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_6),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_6),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_6),
.B(n_362),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_6),
.B(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_6),
.B(n_414),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_7),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_7),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_7),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_7),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_7),
.B(n_122),
.Y(n_181)
);

NAND2x1p5_ASAP7_75t_L g193 ( 
.A(n_7),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_7),
.B(n_264),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_7),
.B(n_106),
.Y(n_297)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_8),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_8),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_8),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_8),
.Y(n_144)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_9),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_9),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_9),
.Y(n_226)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_9),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_10),
.A2(n_19),
.B(n_21),
.Y(n_18)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_11),
.Y(n_266)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_11),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_12),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_12),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_12),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_12),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_12),
.B(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_12),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_13),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_13),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_13),
.B(n_102),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_13),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_13),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_13),
.B(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_13),
.B(n_477),
.Y(n_476)
);

NAND2x1_ASAP7_75t_SL g502 ( 
.A(n_13),
.B(n_503),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_14),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_15),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_15),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_15),
.B(n_152),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_15),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_15),
.B(n_361),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_15),
.B(n_66),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_15),
.B(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_15),
.B(n_400),
.Y(n_418)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_16),
.Y(n_112)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g106 ( 
.A(n_17),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g449 ( 
.A(n_17),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

A2O1A1O1Ixp25_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_430),
.B(n_522),
.C(n_529),
.D(n_531),
.Y(n_22)
);

NAND2x1_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_321),
.Y(n_23)
);

A2O1A1O1Ixp25_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_234),
.B(n_283),
.C(n_284),
.D(n_320),
.Y(n_24)
);

OAI21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_205),
.B(n_233),
.Y(n_25)
);

NOR2x1_ASAP7_75t_L g322 ( 
.A(n_26),
.B(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_157),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_27),
.B(n_157),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_103),
.C(n_128),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_28),
.B(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_68),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_46),
.Y(n_29)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_30),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_42),
.B2(n_43),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_36),
.B1(n_40),
.B2(n_41),
.Y(n_32)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_33),
.B(n_41),
.C(n_42),
.Y(n_183)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_35),
.Y(n_171)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_35),
.Y(n_459)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_36),
.A2(n_41),
.B1(n_58),
.B2(n_131),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_36),
.A2(n_41),
.B1(n_193),
.B2(n_198),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_36),
.B(n_131),
.C(n_505),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_39),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_41),
.B(n_198),
.C(n_313),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_42),
.A2(n_43),
.B1(n_316),
.B2(n_319),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_43),
.B(n_313),
.C(n_319),
.Y(n_460)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_46),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_57),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B1(n_52),
.B2(n_56),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_48),
.A2(n_52),
.B(n_57),
.C(n_202),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_50),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_50),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_50),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_51),
.B(n_56),
.Y(n_202)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.C(n_65),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_58),
.A2(n_65),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_58),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_58),
.A2(n_101),
.B1(n_131),
.B2(n_217),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_58),
.B(n_217),
.C(n_457),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_61),
.B(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g253 ( 
.A(n_63),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_65),
.B(n_272),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_68),
.B(n_159),
.C(n_160),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_84),
.C(n_94),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_69),
.B(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_75),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_76),
.C(n_80),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_78),
.Y(n_398)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_79),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_79),
.Y(n_344)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_79),
.Y(n_370)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_84),
.A2(n_85),
.B1(n_94),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_91),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_86),
.A2(n_87),
.B1(n_91),
.B2(n_180),
.Y(n_218)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_90),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_91),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_91),
.Y(n_180)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_94),
.Y(n_212)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.C(n_101),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_95),
.A2(n_101),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_95),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_97),
.B(n_215),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_100),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_101),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_101),
.A2(n_147),
.B1(n_217),
.B2(n_268),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_101),
.B(n_268),
.C(n_305),
.Y(n_461)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_102),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_102),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_103),
.B(n_128),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_116),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_104),
.B(n_118),
.C(n_127),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_105),
.B(n_109),
.C(n_113),
.Y(n_199)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g469 ( 
.A(n_106),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_113),
.B2(n_115),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_111),
.Y(n_417)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_113),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_115),
.B(n_147),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_127),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_134),
.B(n_140),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.C(n_145),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_129),
.B(n_133),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_132),
.B(n_273),
.C(n_280),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_135),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_135),
.B(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_145),
.B(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.C(n_153),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_146),
.B(n_334),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_147),
.A2(n_181),
.B1(n_182),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_147),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_147),
.B(n_182),
.C(n_263),
.Y(n_298)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_334)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_158),
.B(n_186),
.C(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_186),
.B2(n_187),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_163),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_175),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_164),
.B(n_183),
.C(n_184),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g258 ( 
.A(n_165),
.B(n_170),
.C(n_172),
.Y(n_258)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_172),
.A2(n_440),
.B1(n_441),
.B2(n_442),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_172),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_172),
.B(n_441),
.C(n_446),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_174),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_175)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

XNOR2x1_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_177),
.B(n_180),
.C(n_182),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_181),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_181),
.B(n_343),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_182),
.B(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_188),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_189)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_199),
.B2(n_200),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_192)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_193),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_193),
.A2(n_198),
.B1(n_263),
.B2(n_518),
.Y(n_517)
);

NAND3xp33_ASAP7_75t_L g530 ( 
.A(n_193),
.B(n_446),
.C(n_518),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_195),
.Y(n_257)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_195),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_196),
.B(n_198),
.C(n_200),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_199),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_231),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_206),
.B(n_231),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.C(n_213),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_207),
.B(n_327),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_209),
.A2(n_210),
.B1(n_213),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_213),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.C(n_219),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_214),
.B(n_332),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_218),
.B(n_219),
.Y(n_332)
);

MAJx2_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.C(n_227),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_220),
.B(n_227),
.Y(n_377)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_224),
.B(n_377),
.Y(n_376)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NAND4xp25_ASAP7_75t_SL g321 ( 
.A(n_234),
.B(n_284),
.C(n_322),
.D(n_324),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_235),
.B(n_237),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_242),
.Y(n_237)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_238),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.C(n_241),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_261),
.B1(n_281),
.B2(n_282),
.Y(n_242)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_243),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_260),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_244),
.B(n_247),
.C(n_259),
.Y(n_288)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_259),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_249),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_258),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_252),
.B(n_254),
.C(n_258),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_254),
.A2(n_255),
.B1(n_475),
.B2(n_476),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_254),
.B(n_473),
.C(n_476),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_255),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_255),
.B(n_300),
.C(n_452),
.Y(n_451)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_281),
.C(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_269),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_270),
.C(n_271),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_267),
.Y(n_262)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_263),
.Y(n_518)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_266),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_276),
.B2(n_280),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_275),
.Y(n_318)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_276),
.Y(n_280)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_287),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_288),
.B(n_290),
.C(n_302),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_302),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_301),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_291),
.B(n_294),
.C(n_295),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

AO22x1_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_295)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_296),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g452 ( 
.A(n_297),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_298),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_310),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_303),
.B(n_311),
.C(n_312),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_306),
.B(n_458),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_306),
.B(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_SL g499 ( 
.A(n_313),
.B(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_316),
.Y(n_319)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

OAI21x1_ASAP7_75t_SL g324 ( 
.A1(n_325),
.A2(n_345),
.B(n_429),
.Y(n_324)
);

NOR2xp67_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_329),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_326),
.B(n_329),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_333),
.C(n_335),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_330),
.A2(n_331),
.B1(n_426),
.B2(n_427),
.Y(n_425)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_333),
.B(n_335),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.C(n_342),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_336),
.A2(n_337),
.B1(n_338),
.B2(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_336),
.Y(n_380)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_342),
.B(n_379),
.Y(n_378)
);

AOI21x1_ASAP7_75t_SL g345 ( 
.A1(n_346),
.A2(n_423),
.B(n_428),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_381),
.B(n_422),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_373),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_348),
.B(n_373),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_364),
.C(n_371),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_349),
.A2(n_350),
.B1(n_389),
.B2(n_391),
.Y(n_388)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_360),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_357),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_357),
.C(n_360),
.Y(n_375)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_364),
.A2(n_371),
.B1(n_372),
.B2(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_364),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_365),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.Y(n_384)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_378),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_375),
.B(n_376),
.C(n_378),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_392),
.B(n_421),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_388),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_383),
.B(n_388),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_385),
.C(n_387),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_404),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_385),
.A2(n_386),
.B1(n_387),
.B2(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_387),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_389),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_393),
.A2(n_406),
.B(n_420),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_403),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_394),
.B(n_403),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_399),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_395),
.B(n_399),
.Y(n_411)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_412),
.B(n_419),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_411),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_408),
.B(n_411),
.Y(n_419)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_418),
.Y(n_412)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_424),
.B(n_425),
.Y(n_428)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

NOR3xp33_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_492),
.C(n_511),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_488),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_433),
.A2(n_525),
.B(n_526),
.Y(n_524)
);

NOR2xp67_ASAP7_75t_SL g433 ( 
.A(n_434),
.B(n_482),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_434),
.B(n_482),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_453),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_435),
.B(n_454),
.C(n_462),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.C(n_451),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_436),
.B(n_484),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_437),
.B(n_451),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_438),
.A2(n_439),
.B1(n_446),
.B2(n_450),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_446),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_446),
.A2(n_450),
.B1(n_517),
.B2(n_519),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_448),
.Y(n_503)
);

INVx8_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_452),
.A2(n_515),
.B(n_530),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_462),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_460),
.C(n_461),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_455),
.B(n_486),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

INVx6_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_460),
.B(n_461),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_463),
.A2(n_464),
.B1(n_471),
.B2(n_472),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_465),
.B(n_466),
.C(n_471),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_470),
.Y(n_466)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_467),
.Y(n_505)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_473),
.B(n_474),
.Y(n_472)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_485),
.C(n_487),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_483),
.B(n_485),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_487),
.B(n_490),
.Y(n_489)
);

OR2x6_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_491),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_489),
.B(n_491),
.Y(n_525)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

A2O1A1O1Ixp25_ASAP7_75t_L g523 ( 
.A1(n_493),
.A2(n_512),
.B(n_524),
.C(n_527),
.D(n_528),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_494),
.B(n_510),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_494),
.B(n_510),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_495),
.B(n_497),
.C(n_509),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_497),
.A2(n_498),
.B1(n_508),
.B2(n_509),
.Y(n_496)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_497),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_498),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_501),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_499),
.B(n_504),
.C(n_506),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_504),
.B1(n_506),
.B2(n_507),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_502),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_504),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_521),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_513),
.B(n_521),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_520),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_516),
.Y(n_514)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_517),
.Y(n_519)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_530),
.Y(n_529)
);


endmodule