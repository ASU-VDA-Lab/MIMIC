module fake_jpeg_17014_n_375 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_375);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_375;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_SL g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_13),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_38),
.B(n_41),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_12),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_50),
.Y(n_66)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_23),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_10),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_26),
.B(n_9),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_1),
.Y(n_107)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_29),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_57),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_29),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_63),
.Y(n_77)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_24),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_33),
.B1(n_35),
.B2(n_14),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_65),
.A2(n_78),
.B1(n_101),
.B2(n_109),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_37),
.A2(n_33),
.B1(n_36),
.B2(n_28),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_68),
.A2(n_72),
.B1(n_82),
.B2(n_84),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_30),
.B1(n_27),
.B2(n_25),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_35),
.B1(n_18),
.B2(n_22),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_21),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_79),
.B(n_81),
.Y(n_120)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_21),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_37),
.A2(n_36),
.B1(n_28),
.B2(n_30),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_27),
.B1(n_25),
.B2(n_34),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_38),
.B(n_16),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_95),
.Y(n_118)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_16),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_54),
.A2(n_35),
.B1(n_22),
.B2(n_24),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_43),
.B(n_16),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_105),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_45),
.B(n_1),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_110),
.Y(n_151)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_42),
.Y(n_108)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_47),
.A2(n_22),
.B1(n_15),
.B2(n_34),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_59),
.Y(n_111)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_7),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_49),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_75),
.A2(n_63),
.B1(n_64),
.B2(n_61),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_115),
.A2(n_137),
.B1(n_139),
.B2(n_157),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_61),
.B1(n_34),
.B2(n_64),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_117),
.A2(n_119),
.B1(n_132),
.B2(n_127),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_73),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_122),
.B(n_123),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_100),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_41),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_124),
.B(n_116),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_69),
.B(n_2),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_125),
.B(n_140),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_114),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_143),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_34),
.C(n_3),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_129),
.B(n_140),
.C(n_139),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_2),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_132),
.A2(n_145),
.B(n_125),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_134),
.B(n_135),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_114),
.Y(n_135)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_136),
.B(n_149),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_75),
.A2(n_34),
.B1(n_4),
.B2(n_5),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_77),
.B(n_6),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_82),
.B(n_6),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_85),
.B(n_7),
.Y(n_145)
);

NAND2xp33_ASAP7_75t_SL g148 ( 
.A(n_65),
.B(n_7),
.Y(n_148)
);

XNOR2x1_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_112),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_150),
.B(n_162),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_76),
.A2(n_86),
.B1(n_78),
.B2(n_96),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_152),
.A2(n_128),
.B1(n_134),
.B2(n_143),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_153),
.Y(n_172)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_97),
.A2(n_8),
.B1(n_110),
.B2(n_67),
.Y(n_157)
);

AOI32xp33_ASAP7_75t_L g158 ( 
.A1(n_66),
.A2(n_101),
.A3(n_68),
.B1(n_109),
.B2(n_87),
.Y(n_158)
);

A2O1A1O1Ixp25_ASAP7_75t_L g203 ( 
.A1(n_158),
.A2(n_164),
.B(n_130),
.C(n_153),
.D(n_147),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_90),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_163),
.Y(n_174)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_74),
.B(n_111),
.Y(n_161)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_88),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_67),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_165),
.B(n_87),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_166),
.B(n_167),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_168),
.B(n_184),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_169),
.A2(n_189),
.B1(n_200),
.B2(n_183),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_118),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_173),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_121),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_175),
.B(n_193),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_117),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_177),
.A2(n_192),
.B(n_197),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_141),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_178),
.B(n_198),
.Y(n_229)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_181),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_182),
.B(n_183),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_117),
.Y(n_183)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_128),
.A2(n_152),
.B1(n_119),
.B2(n_132),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_203),
.B1(n_177),
.B2(n_170),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_117),
.B(n_121),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_133),
.A2(n_138),
.B1(n_131),
.B2(n_127),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_194),
.A2(n_189),
.B1(n_200),
.B2(n_176),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_120),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g219 ( 
.A(n_196),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_133),
.B(n_138),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_131),
.B(n_154),
.Y(n_198)
);

NAND2xp33_ASAP7_75t_SL g199 ( 
.A(n_150),
.B(n_165),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_199),
.A2(n_192),
.B(n_208),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_144),
.A2(n_159),
.B1(n_163),
.B2(n_145),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_144),
.B(n_155),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_201),
.B(n_204),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_116),
.B(n_147),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_206),
.Y(n_232)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_126),
.Y(n_207)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

AND2x6_ASAP7_75t_L g209 ( 
.A(n_134),
.B(n_158),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_171),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_212),
.B(n_214),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_166),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_184),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_215),
.B(n_236),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_217),
.B(n_227),
.Y(n_262)
);

OA21x2_ASAP7_75t_L g222 ( 
.A1(n_168),
.A2(n_191),
.B(n_203),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_222),
.B(n_223),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_174),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_225),
.A2(n_213),
.B1(n_241),
.B2(n_237),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_250),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_169),
.A2(n_209),
.B1(n_178),
.B2(n_173),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_228),
.A2(n_233),
.B1(n_238),
.B2(n_246),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_185),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_230),
.B(n_231),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_210),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_232),
.B(n_247),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_186),
.B1(n_199),
.B2(n_207),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_234),
.A2(n_213),
.B(n_221),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_197),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_197),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_237),
.B(n_239),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_179),
.A2(n_198),
.B1(n_201),
.B2(n_181),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_201),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_187),
.Y(n_245)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_195),
.A2(n_172),
.B1(n_193),
.B2(n_182),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_187),
.B(n_195),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_187),
.B(n_180),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_174),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_207),
.Y(n_251)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_214),
.B(n_248),
.C(n_222),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_252),
.B(n_273),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_247),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_254),
.B(n_258),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_235),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_229),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_240),
.A2(n_222),
.B1(n_250),
.B2(n_235),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_256),
.A2(n_274),
.B1(n_283),
.B2(n_262),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_224),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_220),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_265),
.B(n_266),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_218),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_271),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_227),
.B1(n_244),
.B2(n_226),
.Y(n_288)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_220),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_216),
.Y(n_272)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_239),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_245),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_271),
.Y(n_305)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_279),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_243),
.A2(n_235),
.B(n_244),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_279),
.A2(n_282),
.B(n_277),
.Y(n_307)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_216),
.Y(n_280)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_234),
.A2(n_212),
.B(n_225),
.Y(n_282)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_229),
.C(n_248),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_285),
.B(n_303),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_289),
.C(n_269),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_276),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_287),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_288),
.A2(n_300),
.B1(n_263),
.B2(n_278),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_256),
.Y(n_289)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_297),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_254),
.B(n_232),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_298),
.Y(n_313)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_259),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_299),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_262),
.A2(n_219),
.B1(n_249),
.B2(n_267),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_264),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_301),
.Y(n_326)
);

INVx13_ASAP7_75t_L g304 ( 
.A(n_264),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_304),
.A2(n_306),
.B1(n_309),
.B2(n_280),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_305),
.B(n_308),
.Y(n_321)
);

INVx13_ASAP7_75t_L g306 ( 
.A(n_272),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_307),
.A2(n_311),
.B(n_273),
.Y(n_330)
);

BUFx12_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_258),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_267),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_252),
.A2(n_253),
.B(n_283),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_312),
.B(n_322),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_281),
.C(n_263),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_327),
.C(n_294),
.Y(n_339)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_315),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_281),
.Y(n_318)
);

AOI221xp5_ASAP7_75t_L g335 ( 
.A1(n_319),
.A2(n_310),
.B1(n_300),
.B2(n_292),
.C(n_296),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g323 ( 
.A1(n_291),
.A2(n_290),
.B(n_298),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_308),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_257),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_288),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_291),
.A2(n_253),
.B1(n_261),
.B2(n_278),
.Y(n_328)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_328),
.Y(n_334)
);

AOI21xp33_ASAP7_75t_L g329 ( 
.A1(n_285),
.A2(n_257),
.B(n_261),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_329),
.A2(n_330),
.B(n_302),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_311),
.A2(n_273),
.B1(n_260),
.B2(n_275),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_331),
.A2(n_301),
.B1(n_304),
.B2(n_306),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_321),
.B(n_309),
.Y(n_332)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_332),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_335),
.A2(n_322),
.B1(n_323),
.B2(n_319),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_336),
.A2(n_345),
.B(n_317),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_337),
.A2(n_313),
.B(n_315),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_326),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_338),
.B(n_342),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_339),
.B(n_341),
.Y(n_347)
);

OAI32xp33_ASAP7_75t_L g340 ( 
.A1(n_323),
.A2(n_260),
.A3(n_293),
.B1(n_270),
.B2(n_259),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_328),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_325),
.B(n_308),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_316),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_343),
.A2(n_320),
.B1(n_314),
.B2(n_318),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_324),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_295),
.C(n_287),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_346),
.B(n_317),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_333),
.A2(n_331),
.B(n_343),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_348),
.A2(n_357),
.B(n_346),
.Y(n_358)
);

AO21x1_ASAP7_75t_L g363 ( 
.A1(n_349),
.A2(n_356),
.B(n_351),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_350),
.B(n_354),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_355),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_339),
.B(n_327),
.Y(n_354)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_358),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_353),
.B(n_334),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_360),
.B(n_361),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_350),
.B(n_341),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_363),
.B(n_340),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_365),
.A2(n_363),
.B(n_355),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_359),
.A2(n_352),
.B1(n_349),
.B2(n_348),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_366),
.B(n_362),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_368),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_369),
.A2(n_367),
.B1(n_364),
.B2(n_354),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_371),
.B(n_347),
.C(n_344),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_372),
.Y(n_373)
);

AO21x1_ASAP7_75t_L g374 ( 
.A1(n_373),
.A2(n_370),
.B(n_365),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_374),
.B(n_347),
.Y(n_375)
);


endmodule