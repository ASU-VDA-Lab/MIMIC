module fake_jpeg_48_n_63 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_26),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_0),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_23),
.Y(n_30)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_25),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_22),
.C(n_24),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_23),
.B(n_19),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

AOI22x1_ASAP7_75t_SL g38 ( 
.A1(n_31),
.A2(n_26),
.B1(n_24),
.B2(n_21),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_22),
.B1(n_20),
.B2(n_31),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_SL g40 ( 
.A(n_34),
.B(n_24),
.C(n_23),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_1),
.C(n_2),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_22),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_20),
.B1(n_21),
.B2(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_49),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_21),
.C(n_20),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_50),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_1),
.C(n_2),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_5),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_41),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_6),
.C(n_7),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_47),
.B1(n_7),
.B2(n_8),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_57),
.C(n_58),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_9),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

OAI321xp33_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_53),
.C(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_11),
.Y(n_63)
);


endmodule