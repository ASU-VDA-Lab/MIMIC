module real_jpeg_9843_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_300, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_300;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_249;
wire n_292;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_271;
wire n_281;
wire n_131;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_293;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_160;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_202;
wire n_213;
wire n_167;
wire n_179;
wire n_216;
wire n_133;
wire n_295;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx24_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_1),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_1),
.A2(n_35),
.B1(n_63),
.B2(n_66),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_1),
.A2(n_35),
.B1(n_47),
.B2(n_48),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_2),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

AOI21xp33_ASAP7_75t_L g222 ( 
.A1(n_2),
.A2(n_3),
.B(n_32),
.Y(n_222)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_3),
.A2(n_48),
.B(n_58),
.C(n_127),
.D(n_128),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_3),
.B(n_48),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_3),
.B(n_46),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_3),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_3),
.A2(n_83),
.B(n_146),
.Y(n_166)
);

A2O1A1O1Ixp25_ASAP7_75t_L g179 ( 
.A1(n_3),
.A2(n_31),
.B(n_42),
.C(n_180),
.D(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_3),
.B(n_31),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_3),
.B(n_115),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_3),
.A2(n_27),
.B1(n_34),
.B2(n_161),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_4),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_4),
.B(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_4),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_4),
.A2(n_164),
.B(n_190),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx6f_ASAP7_75t_SL g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_9),
.A2(n_51),
.B1(n_63),
.B2(n_66),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_54),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_10),
.A2(n_54),
.B1(n_63),
.B2(n_66),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_11),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_11),
.A2(n_63),
.B1(n_66),
.B2(n_141),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_141),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_11),
.A2(n_27),
.B1(n_34),
.B2(n_141),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_12),
.A2(n_27),
.B1(n_34),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_12),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_12),
.A2(n_47),
.B1(n_48),
.B2(n_92),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_12),
.A2(n_63),
.B1(n_66),
.B2(n_92),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_92),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_14),
.A2(n_27),
.B1(n_34),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_14),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_14),
.A2(n_37),
.B1(n_63),
.B2(n_66),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_15),
.A2(n_27),
.B1(n_34),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_15),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_15),
.A2(n_63),
.B1(n_66),
.B2(n_113),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_15),
.A2(n_47),
.B1(n_48),
.B2(n_113),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_113),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_16),
.A2(n_47),
.B1(n_48),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_16),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_16),
.A2(n_63),
.B1(n_66),
.B2(n_69),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_118),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_116),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_94),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_20),
.B(n_94),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_79),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_71),
.B2(n_72),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_38),
.B2(n_39),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_25)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_26),
.A2(n_112),
.B(n_114),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_26),
.A2(n_30),
.B1(n_112),
.B2(n_251),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_28),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_27),
.A2(n_28),
.B(n_161),
.C(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_30),
.A2(n_33),
.B(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_30),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_30),
.A2(n_90),
.B(n_251),
.Y(n_250)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_43),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_55),
.B1(n_56),
.B2(n_70),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_40),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_41),
.A2(n_52),
.B1(n_200),
.B2(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_41),
.A2(n_235),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_46),
.B1(n_50),
.B2(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_42),
.A2(n_46),
.B1(n_74),
.B2(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_42),
.B(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_44),
.B(n_47),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_45),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_46),
.Y(n_52)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_59),
.B(n_61),
.C(n_62),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_59),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_48),
.A2(n_180),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_52),
.B(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_52),
.A2(n_200),
.B(n_201),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_52),
.A2(n_201),
.B(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_67),
.B(n_68),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_67),
.B1(n_77),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_57),
.A2(n_67),
.B1(n_87),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_57),
.A2(n_67),
.B1(n_140),
.B2(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_57),
.A2(n_178),
.B(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_57),
.A2(n_67),
.B1(n_107),
.B2(n_232),
.Y(n_246)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_62),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_58),
.B(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_66),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_59),
.B(n_66),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_61),
.A2(n_63),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_62),
.Y(n_67)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_84),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_66),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_67),
.B(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_67),
.A2(n_140),
.B(n_142),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_67),
.B(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_67),
.A2(n_142),
.B(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_72),
.A2(n_73),
.B(n_75),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_88),
.B(n_89),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_81),
.B1(n_96),
.B2(n_98),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_82),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_88),
.B1(n_89),
.B2(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_82),
.A2(n_86),
.B1(n_88),
.B2(n_281),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B(n_85),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_83),
.A2(n_145),
.B(n_146),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_83),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_83),
.B(n_148),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_83),
.A2(n_84),
.B1(n_191),
.B2(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_83),
.A2(n_84),
.B1(n_205),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_83),
.A2(n_84),
.B1(n_105),
.B2(n_225),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_84),
.A2(n_153),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_84),
.B(n_161),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_86),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_93),
.A2(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.C(n_101),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_95),
.A2(n_99),
.B1(n_100),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_95),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_96),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_101),
.A2(n_102),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.C(n_110),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_103),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_104),
.B(n_106),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_108),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_109),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_114),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI321xp33_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_274),
.A3(n_287),
.B1(n_293),
.B2(n_298),
.C(n_300),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_241),
.C(n_271),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_215),
.B(n_240),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_194),
.B(n_214),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_172),
.B(n_193),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_149),
.B(n_171),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_134),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_125),
.B(n_134),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_126),
.A2(n_130),
.B1(n_131),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_127),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_128),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_129),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_144),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_139),
.C(n_144),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_145),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_158),
.B(n_170),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_151),
.B(n_156),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_165),
.B(n_169),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_160),
.B(n_162),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_173),
.B(n_174),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_185),
.B2(n_192),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_179),
.B1(n_183),
.B2(n_184),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_177),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_179),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_184),
.C(n_192),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_181),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_182),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_185),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_189),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_195),
.B(n_196),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_210),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_211),
.C(n_212),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_203),
.B2(n_209),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_206),
.C(n_207),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_204),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_206),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_216),
.B(n_217),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_229),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_219),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_219),
.B(n_228),
.C(n_229),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_224),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_226),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_237),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_233),
.B1(n_234),
.B2(n_236),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_231),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_236),
.C(n_237),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

AOI21xp33_ASAP7_75t_L g294 ( 
.A1(n_242),
.A2(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_257),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_243),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_243),
.B(n_257),
.Y(n_296)
);

FAx1_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_247),
.CI(n_248),
.CON(n_243),
.SN(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_246),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_256),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_252),
.B1(n_253),
.B2(n_255),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_250),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_255),
.C(n_256),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_269),
.B2(n_270),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_261),
.C(n_270),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_266),
.C(n_268),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_264),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_269),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_273),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_283),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_275),
.B(n_283),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_280),
.C(n_282),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_276),
.A2(n_277),
.B1(n_280),
.B2(n_292),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_288),
.A2(n_294),
.B(n_297),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_289),
.B(n_290),
.Y(n_297)
);


endmodule