module fake_jpeg_10389_n_207 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_207);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_207;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_6),
.B(n_5),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_2),
.B(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp67_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_36),
.B(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_24),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_0),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_29),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_63),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_67),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_20),
.B1(n_26),
.B2(n_22),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_61),
.B1(n_64),
.B2(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_59),
.B(n_62),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_26),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_65),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_20),
.B1(n_22),
.B2(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_33),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_35),
.A2(n_20),
.B1(n_31),
.B2(n_23),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_30),
.C(n_31),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_35),
.A2(n_17),
.B1(n_18),
.B2(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_77),
.Y(n_103)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_52),
.B(n_21),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_78),
.B(n_79),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_21),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_48),
.A2(n_28),
.B1(n_24),
.B2(n_30),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_94),
.B1(n_4),
.B2(n_5),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_82),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_29),
.B1(n_27),
.B2(n_33),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_83),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_116)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_91),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_1),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_16),
.B(n_38),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_51),
.B(n_1),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_29),
.B(n_38),
.C(n_27),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_98),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_40),
.B1(n_1),
.B2(n_2),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_97),
.Y(n_106)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_49),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_123),
.B1(n_94),
.B2(n_82),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_74),
.B(n_0),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_88),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_3),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_113),
.B(n_95),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_3),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_4),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_119),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_117),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_7),
.C(n_11),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_73),
.B(n_7),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_122),
.B(n_7),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_80),
.B1(n_91),
.B2(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_125),
.B(n_126),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_134),
.B1(n_104),
.B2(n_102),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_75),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_133),
.Y(n_153)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_100),
.B1(n_94),
.B2(n_99),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_135),
.B(n_110),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_75),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_143),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_103),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_103),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_72),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_144),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_145),
.B(n_147),
.Y(n_167)
);

FAx1_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_115),
.CI(n_114),
.CON(n_147),
.SN(n_147)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_149),
.A2(n_152),
.B(n_157),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_150),
.B(n_125),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_108),
.C(n_109),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_159),
.C(n_124),
.Y(n_165)
);

NAND2xp33_ASAP7_75t_SL g152 ( 
.A(n_136),
.B(n_95),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_136),
.A2(n_117),
.B(n_113),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_158),
.B(n_161),
.Y(n_168)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

NAND4xp25_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_119),
.C(n_107),
.D(n_112),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_112),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_128),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_166),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_148),
.A2(n_130),
.B1(n_127),
.B2(n_132),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_163),
.A2(n_152),
.B1(n_141),
.B2(n_155),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_173),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_169),
.C(n_172),
.Y(n_176)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_137),
.C(n_131),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_140),
.C(n_139),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_147),
.B1(n_158),
.B2(n_150),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_184),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_171),
.A3(n_168),
.B1(n_149),
.B2(n_165),
.C1(n_157),
.C2(n_161),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_121),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_133),
.B1(n_144),
.B2(n_107),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_162),
.B(n_156),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_180),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_147),
.C(n_156),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_169),
.C(n_160),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_186),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_141),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_111),
.C(n_121),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_189),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_190),
.B(n_179),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_179),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_194),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_188),
.B(n_182),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_195),
.A2(n_180),
.B(n_183),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_176),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_187),
.B(n_185),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_196),
.Y(n_201)
);

AOI31xp67_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_175),
.A3(n_178),
.B(n_186),
.Y(n_200)
);

OAI21x1_ASAP7_75t_L g203 ( 
.A1(n_200),
.A2(n_87),
.B(n_92),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_201),
.B(n_202),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_197),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_201),
.C(n_86),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_204),
.Y(n_207)
);


endmodule